
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule



module b15_ori ( clk, reset, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,  DATAI_9_,
DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
DATAI_1_, DATAI_0_, NA_N, BS16_N, READY_N, HOLD, BE_N_REG_3_,
BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
ADDRESS_REG_0_, W_R_N_REG, D_C_N_REG, M_IO_N_REG, ADS_N_REG,
DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
DATAO_REG_1_, DATAO_REG_0_ );
input clk, reset, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
DATAI_1_, DATAI_0_, NA_N, BS16_N, READY_N, HOLD;
output BE_N_REG_3_, BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
ADDRESS_REG_0_, W_R_N_REG, D_C_N_REG, M_IO_N_REG, ADS_N_REG,
DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_,
DATAO_REG_7_, DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_,
DATAO_REG_2_, DATAO_REG_1_, DATAO_REG_0_;
wire ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, ex_wire30, ex_wire31, ex_wire32, ex_wire33, ex_wire34, ex_wire35, ex_wire36, ex_wire37, ex_wire38, ex_wire39, ex_wire40, ex_wire41, ex_wire42, ex_wire43, ex_wire44, ex_wire45, ex_wire46, ex_wire47, ex_wire48, ex_wire49, ex_wire50, ex_wire51, ex_wire52, ex_wire53, ex_wire54, ex_wire55, ex_wire56, ex_wire57, ex_wire58, ex_wire59, ex_wire60, ex_wire61, ex_wire62, ex_wire63, ex_wire64, ex_wire65, ex_wire66, ex_wire67, ex_wire68, ex_wire69, ex_wire70, ex_wire71, ex_wire72, ex_wire73, ex_wire74, ex_wire75, ex_wire76, ex_wire77, ex_wire78, ex_wire79, ex_wire80, ex_wire81, ex_wire82, ex_wire83, ex_wire84, ex_wire85, ex_wire86, ex_wire87, ex_wire88, ex_wire89, ex_wire90, ex_wire91, ex_wire92, ex_wire93,n2384, n2375, n2370, n2362, n2352, n2342, n2328, n2318, n2313, n2308,
n2303, n2298, n2293, n2288, n2283, n2278, n2273, n2268, n2263, n2258,
n2253, n2248, n2243, n2238, n2233, n2228, n2223, n2218, n2213, n2208,
n2203, n2198, n2193, n2188, n2183, n2178, n2173, n2168, n2163, n2158,
n2153, n2148, n2143, n2138, n2133, n2128, n2123, n2118, n2113, n2108,
n2103, n2098, n2093, n2088, n2083, n2078, n2073, n2068, n2063, n2058,
n2053, n2048, n2043, n2038, n2033, n2028, n2023, n2018, n2013, n2008,
n2003, n1998, n1993, n1988, n1983, n1978, n1973, n1968, n1963, n1958,
n1953, n1948, n1943, n1938, n1933, n1928, n1923, n1918, n1913, n1908,
n1903, n1898, n1893, n1888, n1883, n1878, n1873, n1868, n1863, n1858,
n1853, n1848, n1843, n1838, n1834, n1830, n1826, n1822, n1818, n1814,
n1810, n1806, n1802, n1798, n1794, n1790, n1786, n1782, n1778, n1774,
n1770, n1766, n1762, n1758, n1754, n1750, n1746, n1742, n1738, n1734,
n1730, n1726, n1722, n1718, n1714, n1710, n1705, n1700, n1695, n1690,
n1685, n1680, n1675, n1670, n1665, n1660, n1655, n1650, n1645, n1640,
n1635, n1630, n1625, n1620, n1615, n1610, n1605, n1600, n1595, n1590,
n1585, n1580, n1575, n1570, n1565, n1560, n1555, n1550, n1545, n1540,
n1535, n1530, n1525, n1520, n1515, n1510, n1505, n1500, n1495, n1490,
n1485, n1480, n1475, n1470, n1465, n1460, n1455, n1450, n1445, n1440,
n1435, n1430, n1425, n1420, n1415, n1410, n1405, n1400, n1395, n1390,
n1385, n1380, n1375, n1370, n1365, n1360, n1355, n1350, n1345, n1340,
n1335, n1330, n1325, n1320, n1315, n1310, n1305, n1300, n1295, n1290,
n1285, n1280, n1275, n1270, n1265, n1260, n1255, n1250, n1245, n1240,
n1235, n1210, n1180, n1175, n1170, n1165, n1160, n1155, n1150, n1145,
n1140, n1135, n1130, n1125, n1120, n1115, n1110, n1105, n1100, n1095,
n1090, n1085, n1080, n1075, n1070, n1065, n1060, n1055, n1050, n1045,
n1040, n1035, n1030, n1025, n1020, n1015, n1010, n1005, n1000, n995,
n990, n985, n980, n975, n970, n965, n960, n955, n950, n945, n940,
n935, n930, n925, n920, n915, n910, n905, n900, n895, n890, n885,
n880, n875, n870, n865, n860, n855, n850, n845, n840, n835, n830,
n825, n820, n815, n810, n805, n800, n795, n790, n785, n780, n775,
n770, n765, n760, n755, n750, n745, n740, n735, n730, n725, n720,
n715, n710, n705, n700, n695, n690, n685, n680, n675, n670, n665,
n660, n655, n650, n645, n640, n635, n630, n625, n620, n615, n610,
n605, n600, n595, n590, n585, n580, n575, n570, n565, n560, n555,
n550, n545, n540, n535, n530, n520, n515, n510, n505, n500, n495,
n490, n485, n480, n475, n470, n465, n460, n455, n450, n445, n440,
n435, n430, n425, n420, n415, n410, n405, n400, n395, n390, n385,
n380, n375, n360, n355, n350, n346, n342, n338, n334, n330, n326,
n322, n318, n314, n310, n306, n302, n298, n294, n290, n286, n282,
n278, n274, n270, n266, n262, n258, n254, n250, n246, n242, n238,
n234, n230, n214, n218, n222, n226, n365, n370, n525, n1185, n1190,
n1195, n1200, n1205, n1215, n1220, n1225, n1230, n2323, n2333, n2338,
n2347, n2357, n2366, n2379, n7797, n7798, n7799, n7800, n7801, n7802,
n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
n15346, n15347, n15348, n15349, n15350, n15351, n15352;

dff REQUESTPENDING_REG_reg ( clk, reset, n8016, n2357 );
not U_inv0 ( n15352, n8016 );
dff STATE_REG_2__reg ( clk, reset, n7819, n350 );
not U_inv1 ( n15025, n7819 );
dff STATE_REG_1__reg ( clk, reset, n7802, n355 );
not U_inv2 ( n15026, n7802 );
dff STATE_REG_0__reg ( clk, reset, n7805, n360 );
not U_inv3 ( n15027, n7805 );
dff DATAWIDTH_REG_0__reg ( clk, reset, n7874, n365 );
not U_inv4 ( n15028, n7874 );
dff DATAWIDTH_REG_31__reg ( clk, reset, ex_wire0, n520 );
not U_inv5 ( n15059, ex_wire0 );
dff DATAWIDTH_REG_30__reg ( clk, reset, ex_wire1, n515 );
not U_inv6 ( n15058, ex_wire1 );
dff DATAWIDTH_REG_29__reg ( clk, reset, ex_wire2, n510 );
not U_inv7 ( n15057, ex_wire2 );
dff DATAWIDTH_REG_28__reg ( clk, reset, ex_wire3, n505 );
not U_inv8 ( n15056, ex_wire3 );
dff DATAWIDTH_REG_27__reg ( clk, reset, ex_wire4, n500 );
not U_inv9 ( n15055, ex_wire4 );
dff DATAWIDTH_REG_26__reg ( clk, reset, ex_wire5, n495 );
not U_inv10 ( n15054, ex_wire5 );
dff DATAWIDTH_REG_25__reg ( clk, reset, ex_wire6, n490 );
not U_inv11 ( n15053, ex_wire6 );
dff DATAWIDTH_REG_24__reg ( clk, reset, ex_wire7, n485 );
not U_inv12 ( n15052, ex_wire7 );
dff DATAWIDTH_REG_23__reg ( clk, reset, ex_wire8, n480 );
not U_inv13 ( n15051, ex_wire8 );
dff DATAWIDTH_REG_22__reg ( clk, reset, ex_wire9, n475 );
not U_inv14 ( n15050, ex_wire9 );
dff DATAWIDTH_REG_21__reg ( clk, reset, ex_wire10, n470 );
not U_inv15 ( n15049, ex_wire10 );
dff DATAWIDTH_REG_20__reg ( clk, reset, ex_wire11, n465 );
not U_inv16 ( n15048, ex_wire11 );
dff DATAWIDTH_REG_19__reg ( clk, reset, ex_wire12, n460 );
not U_inv17 ( n15047, ex_wire12 );
dff DATAWIDTH_REG_18__reg ( clk, reset, ex_wire13, n455 );
not U_inv18 ( n15046, ex_wire13 );
dff DATAWIDTH_REG_17__reg ( clk, reset, ex_wire14, n450 );
not U_inv19 ( n15045, ex_wire14 );
dff DATAWIDTH_REG_16__reg ( clk, reset, ex_wire15, n445 );
not U_inv20 ( n15044, ex_wire15 );
dff DATAWIDTH_REG_15__reg ( clk, reset, ex_wire16, n440 );
not U_inv21 ( n15043, ex_wire16 );
dff DATAWIDTH_REG_14__reg ( clk, reset, ex_wire17, n435 );
not U_inv22 ( n15042, ex_wire17 );
dff DATAWIDTH_REG_13__reg ( clk, reset, ex_wire18, n430 );
not U_inv23 ( n15041, ex_wire18 );
dff DATAWIDTH_REG_12__reg ( clk, reset, ex_wire19, n425 );
not U_inv24 ( n15040, ex_wire19 );
dff DATAWIDTH_REG_11__reg ( clk, reset, ex_wire20, n420 );
not U_inv25 ( n15039, ex_wire20 );
dff DATAWIDTH_REG_10__reg ( clk, reset, ex_wire21, n415 );
not U_inv26 ( n15038, ex_wire21 );
dff DATAWIDTH_REG_9__reg ( clk, reset, ex_wire22, n410 );
not U_inv27 ( n15037, ex_wire22 );
dff DATAWIDTH_REG_8__reg ( clk, reset, ex_wire23, n405 );
not U_inv28 ( n15036, ex_wire23 );
dff DATAWIDTH_REG_7__reg ( clk, reset, ex_wire24, n400 );
not U_inv29 ( n15035, ex_wire24 );
dff DATAWIDTH_REG_6__reg ( clk, reset, ex_wire25, n395 );
not U_inv30 ( n15034, ex_wire25 );
dff DATAWIDTH_REG_5__reg ( clk, reset, ex_wire26, n390 );
not U_inv31 ( n15033, ex_wire26 );
dff DATAWIDTH_REG_4__reg ( clk, reset, ex_wire27, n385 );
not U_inv32 ( n15032, ex_wire27 );
dff DATAWIDTH_REG_3__reg ( clk, reset, ex_wire28, n380 );
not U_inv33 ( n15031, ex_wire28 );
dff DATAWIDTH_REG_2__reg ( clk, reset, n8081, n375 );
not U_inv34 ( n15030, n8081 );
dff DATAWIDTH_REG_1__reg ( clk, reset, n7812, n370 );
not U_inv35 ( n15029, n7812 );
dff STATEBS16_REG_reg ( clk, reset, n7830, n2352 );
not U_inv36 ( n15351, n7830 );
dff INSTQUEUE_REG_4__4__reg ( clk, reset, ex_wire29, n1000 );
not U_inv37 ( n15155, ex_wire29 );
dff PHYADDRPOINTER_REG_20__reg ( clk, reset, n7849, n1495 );
not U_inv38 ( n15247, n7849 );
dff PHYADDRPOINTER_REG_21__reg ( clk, reset, ex_wire30, n1500 );
not U_inv39 ( n15248, ex_wire30 );
dff REIP_REG_21__reg ( clk, reset, ex_wire31, n2263 );
not U_inv40 ( n15340, ex_wire31 );
dff INSTADDRPOINTER_REG_21__reg ( clk, reset, n7833, n1340 );
not U_inv41 ( n15221, n7833 );
dff INSTADDRPOINTER_REG_22__reg ( clk, reset, n7862, n1345 );
not U_inv42 ( n15222, n7862 );
dff EBX_REG_22__reg ( clk, reset, n7883, n2108 );
dff REIP_REG_22__reg ( clk, reset, n8052, n2268 );
not U_inv43 ( n15341, n8052 );
dff ADDRESS_REG_20__reg ( clk, reset, ADDRESS_REG_20_, n266 );
dff PHYADDRPOINTER_REG_22__reg ( clk, reset, n7921, n1505 );
not U_inv44 ( n15249, n7921 );
dff PHYADDRPOINTER_REG_23__reg ( clk, reset, n8020, n1510 );
not U_inv45 ( n15250, n8020 );
dff REIP_REG_23__reg ( clk, reset, n7908, n2273 );
not U_inv46 ( n15342, n7908 );
dff ADDRESS_REG_21__reg ( clk, reset, ADDRESS_REG_21_, n262 );
dff REIP_REG_24__reg ( clk, reset, ex_wire32, n2278 );
not U_inv47 ( n15343, ex_wire32 );
dff ADDRESS_REG_22__reg ( clk, reset, ADDRESS_REG_22_, n258 );
dff INSTADDRPOINTER_REG_24__reg ( clk, reset, n7824, n1355 );
not U_inv48 ( n15224, n7824 );
dff PHYADDRPOINTER_REG_24__reg ( clk, reset, n7848, n1515 );
not U_inv49 ( n15015, n7848 );
dff EBX_REG_24__reg ( clk, reset, n7881, n2118 );
dff INSTADDRPOINTER_REG_25__reg ( clk, reset, n7807, n1360 );
not U_inv50 ( n15225, n7807 );
dff INSTADDRPOINTER_REG_26__reg ( clk, reset, n7841, n1365 );
not U_inv51 ( n15226, n7841 );
dff INSTADDRPOINTER_REG_27__reg ( clk, reset, n7801, n1370 );
not U_inv52 ( n15227, n7801 );
dff INSTADDRPOINTER_REG_28__reg ( clk, reset, n7860, n1375 );
not U_inv53 ( n15021, n7860 );
dff PHYADDRPOINTER_REG_28__reg ( clk, reset, n7847, n1535 );
not U_inv54 ( n15254, n7847 );
dff PHYADDRPOINTER_REG_29__reg ( clk, reset, ex_wire33, n1540 );
not U_inv55 ( n15255, ex_wire33 );
dff REIP_REG_29__reg ( clk, reset, n7915, n2303 );
not U_inv56 ( n15348, n7915 );
dff REIP_REG_30__reg ( clk, reset, ex_wire34, n2308 );
not U_inv57 ( n15349, ex_wire34 );
dff ADDRESS_REG_28__reg ( clk, reset, ADDRESS_REG_28_, n234 );
dff INSTADDRPOINTER_REG_30__reg ( clk, reset, n7845, n1385 );
not U_inv58 ( n15229, n7845 );
dff PHYADDRPOINTER_REG_30__reg ( clk, reset, n8017, n1545 );
not U_inv59 ( n15014, n8017 );
dff EBX_REG_30__reg ( clk, reset, n7875, n2148 );
dff INSTADDRPOINTER_REG_31__reg ( clk, reset, n7834, n1390 );
not U_inv60 ( n15230, n7834 );
dff PHYADDRPOINTER_REG_31__reg ( clk, reset, n7852, n1550 );
not U_inv61 ( n15256, n7852 );
dff REIP_REG_1__reg ( clk, reset, ex_wire35, n2163 );
not U_inv62 ( n15320, ex_wire35 );
dff INSTADDRPOINTER_REG_1__reg ( clk, reset, n7806, n1240 );
not U_inv63 ( n15203, n7806 );
dff INSTQUEUERD_ADDR_REG_1__reg ( clk, reset, n7821, n1200 );
not U_inv64 ( n15195, n7821 );
dff INSTQUEUE_REG_4__3__reg ( clk, reset, ex_wire36, n1005 );
not U_inv65 ( n15156, ex_wire36 );
dff INSTQUEUERD_ADDR_REG_3__reg ( clk, reset, n7816, n1190 );
not U_inv66 ( n15193, n7816 );
dff INSTADDRPOINTER_REG_0__reg ( clk, reset, n7817, n1235 );
not U_inv67 ( n15202, n7817 );
dff INSTQUEUERD_ADDR_REG_2__reg ( clk, reset, n7800, n1195 );
not U_inv68 ( n15194, n7800 );
dff INSTQUEUE_REG_15__7__reg ( clk, reset, n8067, n545 );
not U_inv69 ( n15064, n8067 );
dff INSTQUEUE_REG_2__6__reg ( clk, reset, n8008, n1070 );
not U_inv70 ( n15169, n8008 );
dff STATE2_REG_3__reg ( clk, reset, n7815, n525 );
not U_inv71 ( n15060, n7815 );
dff STATE2_REG_1__reg ( clk, reset, n7799, n535 );
not U_inv72 ( n15062, n7799 );
dff STATE2_REG_2__reg ( clk, reset, n7797, n530 );
not U_inv73 ( n15061, n7797 );
dff INSTQUEUE_REG_4__2__reg ( clk, reset, ex_wire37, n1010 );
not U_inv74 ( n15157, ex_wire37 );
dff INSTQUEUE_REG_3__1__reg ( clk, reset, n8010, n1055 );
not U_inv75 ( n15166, n8010 );
dff FLUSH_REG_reg ( clk, reset, n7813, n2342 );
not U_inv76 ( n15024, n7813 );
dff INSTQUEUERD_ADDR_REG_4__reg ( clk, reset, n7831, n1185 );
not U_inv77 ( n15192, n7831 );
dff INSTQUEUEWR_ADDR_REG_1__reg ( clk, reset, n7825, n1225 );
not U_inv78 ( n15200, n7825 );
dff INSTQUEUEWR_ADDR_REG_2__reg ( clk, reset, n7826, n1220 );
not U_inv79 ( n15199, n7826 );
dff INSTQUEUEWR_ADDR_REG_4__reg ( clk, reset, ex_wire38, n1210 );
not U_inv80 ( n15197, ex_wire38 );
dff INSTQUEUE_REG_4__0__reg ( clk, reset, ex_wire39, n1020 );
not U_inv81 ( n15159, ex_wire39 );
dff INSTQUEUEWR_ADDR_REG_0__reg ( clk, reset, n7803, n1230 );
not U_inv82 ( n15201, n7803 );
dff INSTQUEUEWR_ADDR_REG_3__reg ( clk, reset, n7804, n1215 );
not U_inv83 ( n15198, n7804 );
dff INSTQUEUE_REG_9__0__reg ( clk, reset, n7984, n820 );
not U_inv84 ( n15119, n7984 );
dff INSTQUEUE_REG_9__6__reg ( clk, reset, n7924, n790 );
not U_inv85 ( n15113, n7924 );
dff INSTQUEUE_REG_9__7__reg ( clk, reset, n8061, n785 );
not U_inv86 ( n15112, n8061 );
dff INSTQUEUE_REG_13__0__reg ( clk, reset, n7987, n660 );
not U_inv87 ( n15087, n7987 );
dff INSTQUEUE_REG_13__6__reg ( clk, reset, n7927, n630 );
not U_inv88 ( n15081, n7927 );
dff INSTQUEUE_REG_13__7__reg ( clk, reset, n8065, n625 );
not U_inv89 ( n15080, n8065 );
dff INSTQUEUE_REG_8__0__reg ( clk, reset, n7871, n860 );
not U_inv90 ( n15127, n7871 );
dff INSTQUEUE_REG_8__6__reg ( clk, reset, n7865, n830 );
not U_inv91 ( n15121, n7865 );
dff INSTQUEUE_REG_8__7__reg ( clk, reset, n7994, n825 );
not U_inv92 ( n15120, n7994 );
dff INSTQUEUE_REG_12__0__reg ( clk, reset, n7988, n700 );
not U_inv93 ( n15095, n7988 );
dff INSTQUEUE_REG_12__6__reg ( clk, reset, n7928, n670 );
not U_inv94 ( n15089, n7928 );
dff INSTQUEUE_REG_12__7__reg ( clk, reset, n8064, n665 );
not U_inv95 ( n15088, n8064 );
dff INSTQUEUE_REG_0__0__reg ( clk, reset, n7916, n1180 );
not U_inv96 ( n15191, n7916 );
dff INSTQUEUE_REG_0__6__reg ( clk, reset, n7858, n1150 );
not U_inv97 ( n15185, n7858 );
dff INSTQUEUE_REG_0__7__reg ( clk, reset, n7919, n1145 );
not U_inv98 ( n15184, n7919 );
dff INSTQUEUE_REG_4__6__reg ( clk, reset, ex_wire40, n990 );
not U_inv99 ( n15153, ex_wire40 );
dff INSTQUEUE_REG_4__7__reg ( clk, reset, ex_wire41, n985 );
not U_inv100 ( n15152, ex_wire41 );
dff INSTQUEUE_REG_6__0__reg ( clk, reset, n7992, n940 );
not U_inv101 ( n15143, n7992 );
dff INSTQUEUE_REG_6__6__reg ( clk, reset, n7932, n910 );
not U_inv102 ( n15137, n7932 );
dff INSTQUEUE_REG_6__7__reg ( clk, reset, n8059, n905 );
not U_inv103 ( n15136, n8059 );
dff INSTQUEUE_REG_10__0__reg ( clk, reset, n7985, n780 );
not U_inv104 ( n15111, n7985 );
dff INSTQUEUE_REG_10__6__reg ( clk, reset, n7925, n750 );
not U_inv105 ( n15105, n7925 );
dff INSTQUEUE_REG_10__7__reg ( clk, reset, n8062, n745 );
not U_inv106 ( n15104, n8062 );
dff INSTQUEUE_REG_14__0__reg ( clk, reset, n7989, n620 );
not U_inv107 ( n15079, n7989 );
dff INSTQUEUE_REG_14__6__reg ( clk, reset, n7929, n590 );
not U_inv108 ( n15073, n7929 );
dff INSTQUEUE_REG_14__7__reg ( clk, reset, n8066, n585 );
not U_inv109 ( n15072, n8066 );
dff INSTQUEUE_REG_2__0__reg ( clk, reset, n8002, n1100 );
not U_inv110 ( n15175, n8002 );
dff INSTQUEUE_REG_11__0__reg ( clk, reset, n7986, n740 );
not U_inv111 ( n15103, n7986 );
dff INSTQUEUE_REG_11__6__reg ( clk, reset, n7926, n710 );
not U_inv112 ( n15097, n7926 );
dff INSTQUEUE_REG_11__7__reg ( clk, reset, n8063, n705 );
not U_inv113 ( n15096, n8063 );
dff INSTQUEUE_REG_15__0__reg ( clk, reset, n7990, n580 );
not U_inv114 ( n15071, n7990 );
dff INSTQUEUE_REG_15__6__reg ( clk, reset, n7930, n550 );
not U_inv115 ( n15065, n7930 );
dff INSTQUEUE_REG_3__0__reg ( clk, reset, n8009, n1060 );
not U_inv116 ( n15167, n8009 );
dff INSTQUEUE_REG_3__6__reg ( clk, reset, ex_wire42, n1030 );
not U_inv117 ( n15161, ex_wire42 );
dff INSTQUEUE_REG_5__0__reg ( clk, reset, n7991, n980 );
not U_inv118 ( n15151, n7991 );
dff INSTQUEUE_REG_5__6__reg ( clk, reset, n7931, n950 );
not U_inv119 ( n15145, n7931 );
dff INSTQUEUE_REG_5__7__reg ( clk, reset, n8058, n945 );
not U_inv120 ( n15144, n8058 );
dff INSTQUEUE_REG_7__0__reg ( clk, reset, n7993, n900 );
not U_inv121 ( n15135, n7993 );
dff INSTQUEUE_REG_7__6__reg ( clk, reset, n7933, n870 );
not U_inv122 ( n15129, n7933 );
dff INSTQUEUE_REG_7__7__reg ( clk, reset, n8060, n865 );
not U_inv123 ( n15128, n8060 );
dff INSTQUEUE_REG_1__0__reg ( clk, reset, n7995, n1140 );
not U_inv124 ( n15183, n7995 );
dff INSTQUEUE_REG_1__5__reg ( clk, reset, n8000, n1115 );
not U_inv125 ( n15178, n8000 );
dff INSTQUEUE_REG_4__5__reg ( clk, reset, ex_wire43, n995 );
not U_inv126 ( n15154, ex_wire43 );
dff INSTQUEUE_REG_3__5__reg ( clk, reset, ex_wire44, n1035 );
not U_inv127 ( n15162, ex_wire44 );
dff INSTQUEUE_REG_5__5__reg ( clk, reset, n7941, n955 );
not U_inv128 ( n15146, n7941 );
dff INSTQUEUE_REG_6__5__reg ( clk, reset, n7942, n915 );
not U_inv129 ( n15138, n7942 );
dff INSTQUEUE_REG_7__5__reg ( clk, reset, n7943, n875 );
not U_inv130 ( n15130, n7943 );
dff INSTQUEUE_REG_8__5__reg ( clk, reset, n7866, n835 );
not U_inv131 ( n15122, n7866 );
dff INSTQUEUE_REG_9__5__reg ( clk, reset, n7934, n795 );
not U_inv132 ( n15114, n7934 );
dff INSTQUEUE_REG_10__5__reg ( clk, reset, n7935, n755 );
not U_inv133 ( n15106, n7935 );
dff INSTQUEUE_REG_11__5__reg ( clk, reset, n7936, n715 );
not U_inv134 ( n15098, n7936 );
dff INSTQUEUE_REG_12__5__reg ( clk, reset, n7938, n675 );
not U_inv135 ( n15090, n7938 );
dff INSTQUEUE_REG_13__5__reg ( clk, reset, n7937, n635 );
not U_inv136 ( n15082, n7937 );
dff INSTQUEUE_REG_14__5__reg ( clk, reset, n7939, n595 );
not U_inv137 ( n15074, n7939 );
dff INSTQUEUE_REG_15__5__reg ( clk, reset, n7940, n555 );
not U_inv138 ( n15066, n7940 );
dff INSTQUEUE_REG_0__5__reg ( clk, reset, n7857, n1155 );
not U_inv139 ( n15186, n7857 );
dff INSTQUEUE_REG_2__5__reg ( clk, reset, n8007, n1075 );
not U_inv140 ( n15170, n8007 );
dff INSTQUEUERD_ADDR_REG_0__reg ( clk, reset, n7798, n1205 );
not U_inv141 ( n15196, n7798 );
dff INSTQUEUE_REG_1__6__reg ( clk, reset, n8001, n1110 );
not U_inv142 ( n15177, n8001 );
dff INSTQUEUE_REG_1__7__reg ( clk, reset, n8068, n1105 );
not U_inv143 ( n15176, n8068 );
dff INSTQUEUE_REG_5__1__reg ( clk, reset, n7981, n975 );
not U_inv144 ( n15150, n7981 );
dff INSTQUEUE_REG_6__1__reg ( clk, reset, n7982, n935 );
not U_inv145 ( n15142, n7982 );
dff INSTQUEUE_REG_7__1__reg ( clk, reset, n7983, n895 );
not U_inv146 ( n15134, n7983 );
dff INSTQUEUE_REG_8__1__reg ( clk, reset, n7870, n855 );
not U_inv147 ( n15126, n7870 );
dff INSTQUEUE_REG_9__1__reg ( clk, reset, n7974, n815 );
not U_inv148 ( n15118, n7974 );
dff INSTQUEUE_REG_10__1__reg ( clk, reset, n7975, n775 );
not U_inv149 ( n15110, n7975 );
dff INSTQUEUE_REG_11__1__reg ( clk, reset, n7976, n735 );
not U_inv150 ( n15102, n7976 );
dff INSTQUEUE_REG_12__1__reg ( clk, reset, n7978, n695 );
not U_inv151 ( n15094, n7978 );
dff INSTQUEUE_REG_13__1__reg ( clk, reset, n7977, n655 );
not U_inv152 ( n15086, n7977 );
dff INSTQUEUE_REG_14__1__reg ( clk, reset, n7979, n615 );
not U_inv153 ( n15078, n7979 );
dff INSTQUEUE_REG_15__1__reg ( clk, reset, n7980, n575 );
not U_inv154 ( n15070, n7980 );
dff INSTQUEUE_REG_0__1__reg ( clk, reset, n7917, n1175 );
not U_inv155 ( n15190, n7917 );
dff INSTQUEUE_REG_1__1__reg ( clk, reset, n7996, n1135 );
not U_inv156 ( n15182, n7996 );
dff INSTQUEUE_REG_2__1__reg ( clk, reset, n8003, n1095 );
not U_inv157 ( n15174, n8003 );
dff INSTQUEUE_REG_4__1__reg ( clk, reset, ex_wire45, n1015 );
not U_inv158 ( n15158, ex_wire45 );
dff INSTQUEUE_REG_5__2__reg ( clk, reset, n7971, n970 );
not U_inv159 ( n15149, n7971 );
dff INSTQUEUE_REG_6__2__reg ( clk, reset, n7972, n930 );
not U_inv160 ( n15141, n7972 );
dff INSTQUEUE_REG_7__2__reg ( clk, reset, n7973, n890 );
not U_inv161 ( n15133, n7973 );
dff INSTQUEUE_REG_8__2__reg ( clk, reset, n7869, n850 );
not U_inv162 ( n15125, n7869 );
dff INSTQUEUE_REG_9__2__reg ( clk, reset, n7964, n810 );
not U_inv163 ( n15117, n7964 );
dff INSTQUEUE_REG_10__2__reg ( clk, reset, n7965, n770 );
not U_inv164 ( n15109, n7965 );
dff INSTQUEUE_REG_11__2__reg ( clk, reset, n7966, n730 );
not U_inv165 ( n15101, n7966 );
dff INSTQUEUE_REG_12__2__reg ( clk, reset, n7968, n690 );
not U_inv166 ( n15093, n7968 );
dff INSTQUEUE_REG_13__2__reg ( clk, reset, n7967, n650 );
not U_inv167 ( n15085, n7967 );
dff INSTQUEUE_REG_14__2__reg ( clk, reset, n7969, n610 );
not U_inv168 ( n15077, n7969 );
dff INSTQUEUE_REG_15__2__reg ( clk, reset, n7970, n570 );
not U_inv169 ( n15069, n7970 );
dff INSTQUEUE_REG_0__2__reg ( clk, reset, n7859, n1170 );
not U_inv170 ( n15189, n7859 );
dff INSTQUEUE_REG_1__2__reg ( clk, reset, n7997, n1130 );
not U_inv171 ( n15181, n7997 );
dff INSTQUEUE_REG_2__2__reg ( clk, reset, n8004, n1090 );
not U_inv172 ( n15173, n8004 );
dff MORE_REG_reg ( clk, reset, n8048, n2347 );
dff EBX_REG_31__reg ( clk, reset, n8022, n2153 );
not U_inv173 ( n15020, n8022 );
dff DATAO_REG_31__reg ( clk, reset, DATAO_REG_31_, n1834 );
not U_inv174 ( n15012, DATAO_REG_31_ );
dff INSTQUEUE_REG_3__2__reg ( clk, reset, n8011, n1050 );
not U_inv175 ( n15165, n8011 );
dff INSTQUEUE_REG_3__7__reg ( clk, reset, ex_wire46, n1025 );
not U_inv176 ( n15160, ex_wire46 );
dff INSTQUEUE_REG_5__3__reg ( clk, reset, n7961, n965 );
not U_inv177 ( n15148, n7961 );
dff INSTQUEUE_REG_6__3__reg ( clk, reset, n7962, n925 );
not U_inv178 ( n15140, n7962 );
dff INSTQUEUE_REG_7__3__reg ( clk, reset, n7963, n885 );
not U_inv179 ( n15132, n7963 );
dff INSTQUEUE_REG_8__3__reg ( clk, reset, n7868, n845 );
not U_inv180 ( n15124, n7868 );
dff INSTQUEUE_REG_9__3__reg ( clk, reset, n7954, n805 );
not U_inv181 ( n15116, n7954 );
dff INSTQUEUE_REG_10__3__reg ( clk, reset, n7955, n765 );
not U_inv182 ( n15108, n7955 );
dff INSTQUEUE_REG_11__3__reg ( clk, reset, n7956, n725 );
not U_inv183 ( n15100, n7956 );
dff INSTQUEUE_REG_12__3__reg ( clk, reset, n7958, n685 );
not U_inv184 ( n15092, n7958 );
dff INSTQUEUE_REG_13__3__reg ( clk, reset, n7957, n645 );
not U_inv185 ( n15084, n7957 );
dff INSTQUEUE_REG_14__3__reg ( clk, reset, n7959, n605 );
not U_inv186 ( n15076, n7959 );
dff INSTQUEUE_REG_15__3__reg ( clk, reset, n7960, n565 );
not U_inv187 ( n15068, n7960 );
dff INSTQUEUE_REG_0__3__reg ( clk, reset, n7918, n1165 );
not U_inv188 ( n15188, n7918 );
dff INSTQUEUE_REG_1__3__reg ( clk, reset, n7998, n1125 );
not U_inv189 ( n15180, n7998 );
dff INSTQUEUE_REG_2__3__reg ( clk, reset, n8005, n1085 );
not U_inv190 ( n15172, n8005 );
dff INSTQUEUE_REG_3__3__reg ( clk, reset, n8012, n1045 );
not U_inv191 ( n15164, n8012 );
dff INSTQUEUE_REG_5__4__reg ( clk, reset, n7951, n960 );
not U_inv192 ( n15147, n7951 );
dff INSTQUEUE_REG_6__4__reg ( clk, reset, n7952, n920 );
not U_inv193 ( n15139, n7952 );
dff INSTQUEUE_REG_7__4__reg ( clk, reset, n7953, n880 );
not U_inv194 ( n15131, n7953 );
dff INSTQUEUE_REG_8__4__reg ( clk, reset, n7867, n840 );
not U_inv195 ( n15123, n7867 );
dff INSTQUEUE_REG_9__4__reg ( clk, reset, n7944, n800 );
not U_inv196 ( n15115, n7944 );
dff INSTQUEUE_REG_10__4__reg ( clk, reset, n7945, n760 );
not U_inv197 ( n15107, n7945 );
dff INSTQUEUE_REG_11__4__reg ( clk, reset, n7946, n720 );
not U_inv198 ( n15099, n7946 );
dff INSTQUEUE_REG_12__4__reg ( clk, reset, n7948, n680 );
not U_inv199 ( n15091, n7948 );
dff INSTQUEUE_REG_13__4__reg ( clk, reset, n7947, n640 );
not U_inv200 ( n15083, n7947 );
dff INSTQUEUE_REG_14__4__reg ( clk, reset, n7949, n600 );
not U_inv201 ( n15075, n7949 );
dff INSTQUEUE_REG_15__4__reg ( clk, reset, n7950, n560 );
not U_inv202 ( n15067, n7950 );
dff INSTQUEUE_REG_0__4__reg ( clk, reset, n7856, n1160 );
not U_inv203 ( n15187, n7856 );
dff INSTQUEUE_REG_1__4__reg ( clk, reset, n7999, n1120 );
not U_inv204 ( n15179, n7999 );
dff INSTQUEUE_REG_2__4__reg ( clk, reset, n8006, n1080 );
not U_inv205 ( n15171, n8006 );
dff INSTQUEUE_REG_3__4__reg ( clk, reset, n8013, n1040 );
not U_inv206 ( n15163, n8013 );
dff EAX_REG_20__reg ( clk, reset, n8075, n1938 );
not U_inv207 ( n15308, n8075 );
dff EAX_REG_0__reg ( clk, reset, n7873, n1838 );
not U_inv208 ( n15288, n7873 );
dff EBX_REG_0__reg ( clk, reset, n7905, n1998 );
dff PHYADDRPOINTER_REG_0__reg ( clk, reset, n8043, n1395 );
not U_inv209 ( n15231, n8043 );
dff REIP_REG_0__reg ( clk, reset, n7855, n2158 );
not U_inv210 ( n15319, n7855 );
dff BYTEENABLE_REG_0__reg ( clk, reset, ex_wire47, n2333 );
not U_inv211 ( n15009, ex_wire47 );
dff BE_N_REG_0__reg ( clk, reset, BE_N_REG_0_, n226 );
dff BYTEENABLE_REG_2__reg ( clk, reset, ex_wire48, n2323 );
not U_inv212 ( n15010, ex_wire48 );
dff BE_N_REG_2__reg ( clk, reset, BE_N_REG_2_, n218 );
dff BYTEENABLE_REG_1__reg ( clk, reset, n8046, n2328 );
dff BE_N_REG_1__reg ( clk, reset, BE_N_REG_1_, n222 );
dff BYTEENABLE_REG_3__reg ( clk, reset, ex_wire49, n2318 );
not U_inv213 ( n15011, ex_wire49 );
dff BE_N_REG_3__reg ( clk, reset, BE_N_REG_3_, n214 );
dff UWORD_REG_4__reg ( clk, reset, ex_wire50, n1685 );
not U_inv214 ( n15283, ex_wire50 );
dff DATAO_REG_20__reg ( clk, reset, DATAO_REG_20_, n1790 );
dff LWORD_REG_0__reg ( clk, reset, ex_wire51, n1630 );
not U_inv215 ( n15272, ex_wire51 );
dff DATAO_REG_0__reg ( clk, reset, DATAO_REG_0_, n1710 );
dff INSTQUEUE_REG_2__7__reg ( clk, reset, n8069, n1065 );
not U_inv216 ( n15168, n8069 );
dff PHYADDRPOINTER_REG_1__reg ( clk, reset, n7850, n1400 );
not U_inv217 ( n15232, n7850 );
dff EBX_REG_1__reg ( clk, reset, n7904, n2003 );
dff EAX_REG_1__reg ( clk, reset, n8023, n1843 );
not U_inv218 ( n15289, n8023 );
dff LWORD_REG_1__reg ( clk, reset, ex_wire52, n1625 );
not U_inv219 ( n15271, ex_wire52 );
dff DATAO_REG_1__reg ( clk, reset, DATAO_REG_1_, n1714 );
dff INSTADDRPOINTER_REG_2__reg ( clk, reset, n7853, n1245 );
not U_inv220 ( n15204, n7853 );
dff EBX_REG_2__reg ( clk, reset, n7903, n2008 );
dff REIP_REG_2__reg ( clk, reset, ex_wire53, n2168 );
not U_inv221 ( n15321, ex_wire53 );
dff ADDRESS_REG_0__reg ( clk, reset, ADDRESS_REG_0_, n346 );
dff PHYADDRPOINTER_REG_2__reg ( clk, reset, ex_wire54, n1405 );
not U_inv222 ( n15233, ex_wire54 );
dff EAX_REG_2__reg ( clk, reset, n8024, n1848 );
not U_inv223 ( n15290, n8024 );
dff LWORD_REG_2__reg ( clk, reset, ex_wire55, n1620 );
not U_inv224 ( n15270, ex_wire55 );
dff DATAO_REG_2__reg ( clk, reset, DATAO_REG_2_, n1718 );
dff REIP_REG_3__reg ( clk, reset, n7846, n2173 );
not U_inv225 ( n15322, n7846 );
dff ADDRESS_REG_1__reg ( clk, reset, ADDRESS_REG_1_, n342 );
dff INSTADDRPOINTER_REG_3__reg ( clk, reset, n7808, n1250 );
not U_inv226 ( n15205, n7808 );
dff PHYADDRPOINTER_REG_3__reg ( clk, reset, n7851, n1410 );
not U_inv227 ( n15234, n7851 );
dff EAX_REG_3__reg ( clk, reset, n8025, n1853 );
not U_inv228 ( n15291, n8025 );
dff LWORD_REG_3__reg ( clk, reset, ex_wire56, n1615 );
not U_inv229 ( n15269, ex_wire56 );
dff DATAO_REG_3__reg ( clk, reset, DATAO_REG_3_, n1722 );
dff EBX_REG_3__reg ( clk, reset, n7902, n2013 );
dff REIP_REG_4__reg ( clk, reset, n8049, n2178 );
not U_inv230 ( n15323, n8049 );
dff ADDRESS_REG_2__reg ( clk, reset, ADDRESS_REG_2_, n338 );
dff INSTADDRPOINTER_REG_4__reg ( clk, reset, n7832, n1255 );
not U_inv231 ( n15023, n7832 );
dff PHYADDRPOINTER_REG_4__reg ( clk, reset, n7923, n1415 );
not U_inv232 ( n15235, n7923 );
dff EBX_REG_4__reg ( clk, reset, n7901, n2018 );
dff EAX_REG_4__reg ( clk, reset, n8026, n1858 );
not U_inv233 ( n15292, n8026 );
dff LWORD_REG_4__reg ( clk, reset, ex_wire57, n1610 );
not U_inv234 ( n15268, ex_wire57 );
dff DATAO_REG_4__reg ( clk, reset, DATAO_REG_4_, n1726 );
dff PHYADDRPOINTER_REG_5__reg ( clk, reset, n7811, n1420 );
not U_inv235 ( n15236, n7811 );
dff EBX_REG_5__reg ( clk, reset, n7900, n2023 );
dff REIP_REG_5__reg ( clk, reset, n7914, n2183 );
not U_inv236 ( n15324, n7914 );
dff ADDRESS_REG_3__reg ( clk, reset, ADDRESS_REG_3_, n334 );
dff INSTADDRPOINTER_REG_5__reg ( clk, reset, n7827, n1260 );
not U_inv237 ( n15206, n7827 );
dff EAX_REG_5__reg ( clk, reset, n8027, n1863 );
not U_inv238 ( n15293, n8027 );
dff LWORD_REG_5__reg ( clk, reset, ex_wire58, n1605 );
not U_inv239 ( n15267, ex_wire58 );
dff DATAO_REG_5__reg ( clk, reset, DATAO_REG_5_, n1730 );
dff EAX_REG_6__reg ( clk, reset, n8028, n1868 );
not U_inv240 ( n15294, n8028 );
dff LWORD_REG_6__reg ( clk, reset, ex_wire59, n1600 );
not U_inv241 ( n15266, ex_wire59 );
dff DATAO_REG_6__reg ( clk, reset, DATAO_REG_6_, n1734 );
dff PHYADDRPOINTER_REG_6__reg ( clk, reset, n7838, n1425 );
not U_inv242 ( n15019, n7838 );
dff REIP_REG_6__reg ( clk, reset, ex_wire60, n2188 );
not U_inv243 ( n15325, ex_wire60 );
dff ADDRESS_REG_4__reg ( clk, reset, ADDRESS_REG_4_, n330 );
dff INSTADDRPOINTER_REG_6__reg ( clk, reset, n7844, n1265 );
not U_inv244 ( n15207, n7844 );
dff EBX_REG_6__reg ( clk, reset, n7899, n2028 );
dff EBX_REG_7__reg ( clk, reset, n7898, n2033 );
dff INSTADDRPOINTER_REG_7__reg ( clk, reset, n7820, n1270 );
not U_inv245 ( n15208, n7820 );
dff PHYADDRPOINTER_REG_7__reg ( clk, reset, n8015, n1430 );
not U_inv246 ( n15237, n8015 );
dff REIP_REG_7__reg ( clk, reset, n8057, n2193 );
not U_inv247 ( n15326, n8057 );
dff ADDRESS_REG_5__reg ( clk, reset, ADDRESS_REG_5_, n326 );
dff EAX_REG_7__reg ( clk, reset, n8029, n1873 );
not U_inv248 ( n15295, n8029 );
dff LWORD_REG_7__reg ( clk, reset, ex_wire61, n1595 );
not U_inv249 ( n15265, ex_wire61 );
dff DATAO_REG_7__reg ( clk, reset, DATAO_REG_7_, n1738 );
dff EAX_REG_8__reg ( clk, reset, n8030, n1878 );
not U_inv250 ( n15296, n8030 );
dff LWORD_REG_8__reg ( clk, reset, ex_wire62, n1590 );
not U_inv251 ( n15264, ex_wire62 );
dff DATAO_REG_8__reg ( clk, reset, DATAO_REG_8_, n1742 );
dff PHYADDRPOINTER_REG_8__reg ( clk, reset, n7864, n1435 );
not U_inv252 ( n15018, n7864 );
dff REIP_REG_8__reg ( clk, reset, n7913, n2198 );
not U_inv253 ( n15327, n7913 );
dff ADDRESS_REG_6__reg ( clk, reset, ADDRESS_REG_6_, n322 );
dff INSTADDRPOINTER_REG_8__reg ( clk, reset, n7822, n1275 );
not U_inv254 ( n15209, n7822 );
dff EBX_REG_8__reg ( clk, reset, n7897, n2038 );
dff EAX_REG_9__reg ( clk, reset, n8031, n1883 );
not U_inv255 ( n15297, n8031 );
dff LWORD_REG_9__reg ( clk, reset, ex_wire63, n1585 );
not U_inv256 ( n15263, ex_wire63 );
dff DATAO_REG_9__reg ( clk, reset, DATAO_REG_9_, n1746 );
dff PHYADDRPOINTER_REG_9__reg ( clk, reset, n7810, n1440 );
not U_inv257 ( n15238, n7810 );
dff REIP_REG_9__reg ( clk, reset, ex_wire64, n2203 );
not U_inv258 ( n15328, ex_wire64 );
dff ADDRESS_REG_7__reg ( clk, reset, ADDRESS_REG_7_, n318 );
dff INSTADDRPOINTER_REG_9__reg ( clk, reset, n7872, n1280 );
not U_inv259 ( n15210, n7872 );
dff EBX_REG_9__reg ( clk, reset, n7896, n2043 );
dff EAX_REG_10__reg ( clk, reset, n8032, n1888 );
not U_inv260 ( n15298, n8032 );
dff LWORD_REG_10__reg ( clk, reset, ex_wire65, n1580 );
not U_inv261 ( n15262, ex_wire65 );
dff DATAO_REG_10__reg ( clk, reset, DATAO_REG_10_, n1750 );
dff PHYADDRPOINTER_REG_10__reg ( clk, reset, n7837, n1445 );
not U_inv262 ( n15017, n7837 );
dff REIP_REG_10__reg ( clk, reset, n8056, n2208 );
not U_inv263 ( n15329, n8056 );
dff ADDRESS_REG_8__reg ( clk, reset, ADDRESS_REG_8_, n314 );
dff INSTADDRPOINTER_REG_10__reg ( clk, reset, n7920, n1285 );
not U_inv264 ( n15022, n7920 );
dff EBX_REG_10__reg ( clk, reset, n7895, n2048 );
dff EBX_REG_11__reg ( clk, reset, n7894, n2053 );
dff INSTADDRPOINTER_REG_11__reg ( clk, reset, n7843, n1290 );
not U_inv265 ( n15211, n7843 );
dff PHYADDRPOINTER_REG_11__reg ( clk, reset, n8014, n1450 );
not U_inv266 ( n15239, n8014 );
dff REIP_REG_11__reg ( clk, reset, n7912, n2213 );
not U_inv267 ( n15330, n7912 );
dff ADDRESS_REG_9__reg ( clk, reset, ADDRESS_REG_9_, n310 );
dff EAX_REG_11__reg ( clk, reset, n8033, n1893 );
not U_inv268 ( n15299, n8033 );
dff LWORD_REG_11__reg ( clk, reset, ex_wire66, n1575 );
not U_inv269 ( n15261, ex_wire66 );
dff DATAO_REG_11__reg ( clk, reset, DATAO_REG_11_, n1754 );
dff EAX_REG_12__reg ( clk, reset, n8034, n1898 );
not U_inv270 ( n15300, n8034 );
dff LWORD_REG_12__reg ( clk, reset, ex_wire67, n1570 );
not U_inv271 ( n15260, ex_wire67 );
dff DATAO_REG_12__reg ( clk, reset, DATAO_REG_12_, n1758 );
dff PHYADDRPOINTER_REG_12__reg ( clk, reset, n7863, n1455 );
not U_inv272 ( n15016, n7863 );
dff REIP_REG_12__reg ( clk, reset, ex_wire68, n2218 );
not U_inv273 ( n15331, ex_wire68 );
dff ADDRESS_REG_10__reg ( clk, reset, ADDRESS_REG_10_, n306 );
dff INSTADDRPOINTER_REG_12__reg ( clk, reset, n7922, n1295 );
not U_inv274 ( n15212, n7922 );
dff EBX_REG_12__reg ( clk, reset, n7893, n2058 );
dff EAX_REG_13__reg ( clk, reset, n8035, n1903 );
not U_inv275 ( n15301, n8035 );
dff LWORD_REG_13__reg ( clk, reset, ex_wire69, n1565 );
not U_inv276 ( n15259, ex_wire69 );
dff DATAO_REG_13__reg ( clk, reset, DATAO_REG_13_, n1762 );
dff PHYADDRPOINTER_REG_13__reg ( clk, reset, n7809, n1460 );
not U_inv277 ( n15240, n7809 );
dff REIP_REG_13__reg ( clk, reset, n8055, n2223 );
not U_inv278 ( n15332, n8055 );
dff ADDRESS_REG_11__reg ( clk, reset, ADDRESS_REG_11_, n302 );
dff INSTADDRPOINTER_REG_13__reg ( clk, reset, n7840, n1300 );
not U_inv279 ( n15213, n7840 );
dff EBX_REG_13__reg ( clk, reset, n7892, n2063 );
dff EAX_REG_14__reg ( clk, reset, n8036, n1908 );
not U_inv280 ( n15302, n8036 );
dff LWORD_REG_14__reg ( clk, reset, ex_wire70, n1560 );
not U_inv281 ( n15258, ex_wire70 );
dff DATAO_REG_14__reg ( clk, reset, DATAO_REG_14_, n1766 );
dff PHYADDRPOINTER_REG_14__reg ( clk, reset, n7836, n1465 );
not U_inv282 ( n15241, n7836 );
dff REIP_REG_14__reg ( clk, reset, n7911, n2228 );
not U_inv283 ( n15333, n7911 );
dff ADDRESS_REG_12__reg ( clk, reset, ADDRESS_REG_12_, n298 );
dff INSTADDRPOINTER_REG_14__reg ( clk, reset, n7854, n1305 );
not U_inv284 ( n15214, n7854 );
dff EBX_REG_14__reg ( clk, reset, n7891, n2068 );
dff PHYADDRPOINTER_REG_15__reg ( clk, reset, n8021, n1470 );
not U_inv285 ( n15242, n8021 );
dff EAX_REG_15__reg ( clk, reset, n8037, n1913 );
not U_inv286 ( n15303, n8037 );
dff LWORD_REG_15__reg ( clk, reset, ex_wire71, n1555 );
not U_inv287 ( n15257, ex_wire71 );
dff DATAO_REG_15__reg ( clk, reset, DATAO_REG_15_, n1770 );
dff REIP_REG_15__reg ( clk, reset, ex_wire72, n2233 );
not U_inv288 ( n15334, ex_wire72 );
dff ADDRESS_REG_13__reg ( clk, reset, ADDRESS_REG_13_, n294 );
dff INSTADDRPOINTER_REG_15__reg ( clk, reset, n7906, n1310 );
not U_inv289 ( n15215, n7906 );
dff INSTADDRPOINTER_REG_16__reg ( clk, reset, n7842, n1315 );
not U_inv290 ( n15216, n7842 );
dff PHYADDRPOINTER_REG_16__reg ( clk, reset, ex_wire73, n1475 );
not U_inv291 ( n15243, ex_wire73 );
dff EBX_REG_16__reg ( clk, reset, n7889, n2078 );
dff EAX_REG_16__reg ( clk, reset, n8071, n1918 );
not U_inv292 ( n15304, n8071 );
dff UWORD_REG_0__reg ( clk, reset, ex_wire74, n1705 );
not U_inv293 ( n15287, ex_wire74 );
dff DATAO_REG_16__reg ( clk, reset, DATAO_REG_16_, n1774 );
dff REIP_REG_16__reg ( clk, reset, n8054, n2238 );
not U_inv294 ( n15335, n8054 );
dff ADDRESS_REG_14__reg ( clk, reset, ADDRESS_REG_14_, n290 );
dff INSTADDRPOINTER_REG_17__reg ( clk, reset, n7828, n1320 );
not U_inv295 ( n15217, n7828 );
dff PHYADDRPOINTER_REG_17__reg ( clk, reset, ex_wire75, n1480 );
not U_inv296 ( n15244, ex_wire75 );
dff EBX_REG_17__reg ( clk, reset, n7888, n2083 );
dff EAX_REG_17__reg ( clk, reset, n8072, n1923 );
not U_inv297 ( n15305, n8072 );
dff UWORD_REG_1__reg ( clk, reset, ex_wire76, n1700 );
not U_inv298 ( n15286, ex_wire76 );
dff DATAO_REG_17__reg ( clk, reset, DATAO_REG_17_, n1778 );
dff REIP_REG_17__reg ( clk, reset, n7910, n2243 );
not U_inv299 ( n15336, n7910 );
dff ADDRESS_REG_15__reg ( clk, reset, ADDRESS_REG_15_, n286 );
dff REIP_REG_18__reg ( clk, reset, ex_wire77, n2248 );
not U_inv300 ( n15337, ex_wire77 );
dff ADDRESS_REG_16__reg ( clk, reset, ADDRESS_REG_16_, n282 );
dff INSTADDRPOINTER_REG_18__reg ( clk, reset, n7835, n1325 );
not U_inv301 ( n15218, n7835 );
dff PHYADDRPOINTER_REG_18__reg ( clk, reset, n8044, n1485 );
not U_inv302 ( n15245, n8044 );
dff EAX_REG_18__reg ( clk, reset, n8073, n1928 );
not U_inv303 ( n15306, n8073 );
dff UWORD_REG_2__reg ( clk, reset, ex_wire78, n1695 );
not U_inv304 ( n15285, ex_wire78 );
dff DATAO_REG_18__reg ( clk, reset, DATAO_REG_18_, n1782 );
dff EBX_REG_18__reg ( clk, reset, n7887, n2088 );
dff EBX_REG_15__reg ( clk, reset, n7890, n2073 );
dff EAX_REG_21__reg ( clk, reset, n8076, n1943 );
not U_inv305 ( n15309, n8076 );
dff UWORD_REG_5__reg ( clk, reset, ex_wire79, n1680 );
not U_inv306 ( n15282, ex_wire79 );
dff DATAO_REG_21__reg ( clk, reset, DATAO_REG_21_, n1794 );
dff EAX_REG_22__reg ( clk, reset, n8077, n1948 );
not U_inv307 ( n15310, n8077 );
dff UWORD_REG_6__reg ( clk, reset, ex_wire80, n1675 );
not U_inv308 ( n15281, ex_wire80 );
dff DATAO_REG_22__reg ( clk, reset, DATAO_REG_22_, n1798 );
dff EAX_REG_23__reg ( clk, reset, n8042, n1953 );
not U_inv309 ( n15311, n8042 );
dff UWORD_REG_7__reg ( clk, reset, ex_wire81, n1670 );
not U_inv310 ( n15280, ex_wire81 );
dff DATAO_REG_23__reg ( clk, reset, DATAO_REG_23_, n1802 );
dff EAX_REG_19__reg ( clk, reset, n8074, n1933 );
not U_inv311 ( n15307, n8074 );
dff UWORD_REG_3__reg ( clk, reset, ex_wire82, n1690 );
not U_inv312 ( n15284, ex_wire82 );
dff DATAO_REG_19__reg ( clk, reset, DATAO_REG_19_, n1786 );
dff PHYADDRPOINTER_REG_19__reg ( clk, reset, ex_wire83, n1490 );
not U_inv313 ( n15246, ex_wire83 );
dff REIP_REG_19__reg ( clk, reset, n8053, n2253 );
not U_inv314 ( n15338, n8053 );
dff ADDRESS_REG_17__reg ( clk, reset, ADDRESS_REG_17_, n278 );
dff INSTADDRPOINTER_REG_19__reg ( clk, reset, n7829, n1330 );
not U_inv315 ( n15219, n7829 );
dff EBX_REG_20__reg ( clk, reset, n7885, n2098 );
dff REIP_REG_20__reg ( clk, reset, n7909, n2258 );
not U_inv316 ( n15339, n7909 );
dff ADDRESS_REG_18__reg ( clk, reset, ADDRESS_REG_18_, n274 );
dff ADDRESS_REG_19__reg ( clk, reset, ADDRESS_REG_19_, n270 );
dff INSTADDRPOINTER_REG_20__reg ( clk, reset, n7839, n1335 );
not U_inv317 ( n15220, n7839 );
dff EBX_REG_21__reg ( clk, reset, n7884, n2103 );
dff EBX_REG_23__reg ( clk, reset, n7882, n2113 );
dff INSTADDRPOINTER_REG_23__reg ( clk, reset, n7823, n1350 );
not U_inv318 ( n15223, n7823 );
dff PHYADDRPOINTER_REG_25__reg ( clk, reset, n8019, n1520 );
not U_inv319 ( n15251, n8019 );
dff EBX_REG_25__reg ( clk, reset, n7880, n2123 );
dff EAX_REG_25__reg ( clk, reset, n8041, n1963 );
not U_inv320 ( n15313, n8041 );
dff UWORD_REG_9__reg ( clk, reset, ex_wire84, n1660 );
not U_inv321 ( n15278, ex_wire84 );
dff DATAO_REG_25__reg ( clk, reset, DATAO_REG_25_, n1810 );
dff REIP_REG_25__reg ( clk, reset, n8051, n2283 );
not U_inv322 ( n15344, n8051 );
dff ADDRESS_REG_23__reg ( clk, reset, ADDRESS_REG_23_, n254 );
dff REIP_REG_26__reg ( clk, reset, n7907, n2288 );
not U_inv323 ( n15345, n7907 );
dff ADDRESS_REG_24__reg ( clk, reset, ADDRESS_REG_24_, n250 );
dff PHYADDRPOINTER_REG_26__reg ( clk, reset, n7861, n1525 );
not U_inv324 ( n15252, n7861 );
dff EBX_REG_26__reg ( clk, reset, n7879, n2128 );
dff EAX_REG_26__reg ( clk, reset, n8040, n1968 );
not U_inv325 ( n15314, n8040 );
dff UWORD_REG_10__reg ( clk, reset, ex_wire85, n1655 );
not U_inv326 ( n15277, ex_wire85 );
dff DATAO_REG_26__reg ( clk, reset, DATAO_REG_26_, n1814 );
dff REIP_REG_27__reg ( clk, reset, ex_wire86, n2293 );
not U_inv327 ( n15346, ex_wire86 );
dff ADDRESS_REG_25__reg ( clk, reset, ADDRESS_REG_25_, n246 );
dff PHYADDRPOINTER_REG_27__reg ( clk, reset, n8018, n1530 );
not U_inv328 ( n15253, n8018 );
dff EBX_REG_28__reg ( clk, reset, n7877, n2138 );
dff EAX_REG_28__reg ( clk, reset, n8079, n1978 );
not U_inv329 ( n15316, n8079 );
dff UWORD_REG_12__reg ( clk, reset, ex_wire87, n1645 );
not U_inv330 ( n15275, ex_wire87 );
dff DATAO_REG_28__reg ( clk, reset, DATAO_REG_28_, n1822 );
dff EBX_REG_29__reg ( clk, reset, n7876, n2143 );
dff INSTADDRPOINTER_REG_29__reg ( clk, reset, n7818, n1380 );
not U_inv331 ( n15228, n7818 );
dff EAX_REG_29__reg ( clk, reset, n8080, n1983 );
not U_inv332 ( n15317, n8080 );
dff UWORD_REG_13__reg ( clk, reset, ex_wire88, n1640 );
not U_inv333 ( n15274, ex_wire88 );
dff DATAO_REG_29__reg ( clk, reset, DATAO_REG_29_, n1826 );
dff EAX_REG_31__reg ( clk, reset, ex_wire89, n1993 );
not U_inv334 ( n15013, ex_wire89 );
dff REIP_REG_28__reg ( clk, reset, n8050, n2298 );
not U_inv335 ( n15347, n8050 );
dff ADDRESS_REG_26__reg ( clk, reset, ADDRESS_REG_26_, n242 );
dff ADDRESS_REG_27__reg ( clk, reset, ADDRESS_REG_27_, n238 );
dff REIP_REG_31__reg ( clk, reset, n8070, n2313 );
not U_inv336 ( n15350, n8070 );
dff ADDRESS_REG_29__reg ( clk, reset, ADDRESS_REG_29_, n230 );
dff EBX_REG_27__reg ( clk, reset, n7878, n2133 );
dff EAX_REG_27__reg ( clk, reset, n8039, n1973 );
not U_inv337 ( n15315, n8039 );
dff UWORD_REG_11__reg ( clk, reset, ex_wire90, n1650 );
not U_inv338 ( n15276, ex_wire90 );
dff DATAO_REG_27__reg ( clk, reset, DATAO_REG_27_, n1818 );
dff EBX_REG_19__reg ( clk, reset, n7886, n2093 );
dff EAX_REG_30__reg ( clk, reset, n8038, n1988 );
not U_inv339 ( n15318, n8038 );
dff UWORD_REG_14__reg ( clk, reset, ex_wire91, n1635 );
not U_inv340 ( n15273, ex_wire91 );
dff DATAO_REG_30__reg ( clk, reset, DATAO_REG_30_, n1830 );
dff EAX_REG_24__reg ( clk, reset, n8078, n1958 );
not U_inv341 ( n15312, n8078 );
dff UWORD_REG_8__reg ( clk, reset, ex_wire92, n1665 );
not U_inv342 ( n15279, ex_wire92 );
dff DATAO_REG_24__reg ( clk, reset, DATAO_REG_24_, n1806 );
dff CODEFETCH_REG_reg ( clk, reset, n8047, n2370 );
dff D_C_N_REG_reg ( clk, reset, D_C_N_REG, n2362 );
not U_inv343 ( n15007, D_C_N_REG );
dff ADS_N_REG_reg ( clk, reset, ADS_N_REG, n2375 );
dff READREQUEST_REG_reg ( clk, reset, ex_wire93, n2379 );
not U_inv344 ( n15008, ex_wire93 );
dff W_R_N_REG_reg ( clk, reset, W_R_N_REG, n2338 );
dff MEMORYFETCH_REG_reg ( clk, reset, n8045, n2384 );
dff M_IO_N_REG_reg ( clk, reset, M_IO_N_REG, n2366 );
dff STATE2_REG_0__reg ( clk, reset, n7814, n540 );
not U_inv345 ( n15063, n7814 );
nand U7799 ( n9226, n9196, n7819 );
nand U7800 ( n9530, n10167, n10168 );
nand U7801 ( n10843, n10361, n7797 );
nand U7802 ( n8235, n15063, n14353 );
not U7803 ( n10579, n10576 );
nand U7804 ( n9217, n9196, n15025 );
nand U7805 ( n12196, n9363, n13712 );
nand U7806 ( n9174, n9401, n9402 );
nor U7807 ( n8184, n10452, n8235 );
nor U7808 ( n8172, n10459, n8235 );
nor U7809 ( n8106, n10438, n8235 );
nor U7810 ( n8160, n10466, n8235 );
nor U7811 ( n8148, n10473, n8235 );
nor U7812 ( n8131, n10481, n8235 );
nor U7813 ( n8089, n10445, n8235 );
nor U7814 ( n8118, n10431, n8235 );
and U7815 ( n10841, n15351, n15061 );
not U7816 ( n8082, n10841 );
not U7817 ( n10188, n8082 );
not U7818 ( n10847, n11209 );
nor U7819 ( n14267, n13789, n8235 );
not U7820 ( n10835, n12106 );
nand U7821 ( n10851, n7814, n10854 );
not U7822 ( n10210, n10202 );
not U7823 ( n9517, n9545 );
not U7824 ( n9536, n9509 );
and U7825 ( n10714, n10717, n10822 );
not U7826 ( n12220, n12188 );
or U7827 ( n10209, n10203, n10361 );
nand U7828 ( n10582, n15063, n10576 );
nand U7829 ( n10384, n10375, n10554 );
nand U7830 ( n10855, n9095, n10854 );
nand U7831 ( n12207, n15061, n12409 );
and U7832 ( n12176, n13720, n13721 );
and U7833 ( n10717, n10826, n10827 );
nand U7834 ( n10203, n9098, n10362 );
nand U7835 ( n10854, n12146, n12147 );
not U7836 ( n10822, n10825 );
not U7837 ( n12254, n9363 );
nand U7838 ( n9216, n15027, n7802 );
nor U7839 ( n9528, n10164, n10165 );
nand U7840 ( n995, n8083, n8084 );
nor U7841 ( n8084, n8085, n8086 );
nand U7842 ( n8086, n8087, n8088 );
nand U7843 ( n8088, n8089, n8090 );
nand U7844 ( n8087, n8091, n8092 );
nor U7845 ( n8085, n8093, n8094 );
nor U7846 ( n8083, n8095, n8096 );
nor U7847 ( n8096, n15154, n8097 );
nor U7848 ( n8095, n8098, n8099 );
nand U7849 ( n990, n8100, n8101 );
nor U7850 ( n8101, n8102, n8103 );
nand U7851 ( n8103, n8104, n8105 );
nand U7852 ( n8105, n8106, n8090 );
nand U7853 ( n8104, n8107, n8091 );
nor U7854 ( n8102, n8094, n8108 );
nor U7855 ( n8100, n8109, n8110 );
nor U7856 ( n8110, n15153, n8097 );
nor U7857 ( n8109, n8099, n8111 );
nand U7858 ( n985, n8112, n8113 );
nor U7859 ( n8113, n8114, n8115 );
nand U7860 ( n8115, n8116, n8117 );
nand U7861 ( n8117, n8118, n8090 );
or U7862 ( n8116, n8119, n8120 );
nor U7863 ( n8114, n8099, n8121 );
nor U7864 ( n8112, n8122, n8123 );
nor U7865 ( n8123, n15152, n8097 );
nor U7866 ( n8122, n8094, n8124 );
nand U7867 ( n980, n8125, n8126 );
nor U7868 ( n8126, n8127, n8128 );
nand U7869 ( n8128, n8129, n8130 );
nand U7870 ( n8130, n8131, n8132 );
nand U7871 ( n8129, n8133, n7991 );
nor U7872 ( n8127, n8134, n8135 );
nor U7873 ( n8125, n8136, n8137 );
nor U7874 ( n8137, n8138, n8139 );
nor U7875 ( n8136, n8140, n8141 );
nand U7876 ( n975, n8142, n8143 );
nor U7877 ( n8143, n8144, n8145 );
nand U7878 ( n8145, n8146, n8147 );
nand U7879 ( n8147, n8148, n8132 );
nand U7880 ( n8146, n8133, n7981 );
nor U7881 ( n8144, n8134, n8149 );
nor U7882 ( n8142, n8150, n8151 );
nor U7883 ( n8151, n8138, n8152 );
nor U7884 ( n8150, n8140, n8153 );
nand U7885 ( n970, n8154, n8155 );
nor U7886 ( n8155, n8156, n8157 );
nand U7887 ( n8157, n8158, n8159 );
nand U7888 ( n8159, n8160, n8132 );
nand U7889 ( n8158, n8133, n7971 );
nor U7890 ( n8156, n8134, n8161 );
nor U7891 ( n8154, n8162, n8163 );
nor U7892 ( n8163, n8138, n8164 );
nor U7893 ( n8162, n8140, n8165 );
nand U7894 ( n965, n8166, n8167 );
nor U7895 ( n8167, n8168, n8169 );
nand U7896 ( n8169, n8170, n8171 );
nand U7897 ( n8171, n8172, n8132 );
nand U7898 ( n8170, n8133, n7961 );
nor U7899 ( n8168, n8134, n8173 );
nor U7900 ( n8166, n8174, n8175 );
nor U7901 ( n8175, n8138, n8176 );
nor U7902 ( n8174, n8140, n8177 );
nand U7903 ( n960, n8178, n8179 );
nor U7904 ( n8179, n8180, n8181 );
nand U7905 ( n8181, n8182, n8183 );
nand U7906 ( n8183, n8184, n8132 );
nand U7907 ( n8182, n8133, n7951 );
nor U7908 ( n8180, n8134, n8185 );
nor U7909 ( n8178, n8186, n8187 );
nor U7910 ( n8187, n8138, n8188 );
nor U7911 ( n8186, n8140, n8189 );
nand U7912 ( n955, n8190, n8191 );
nor U7913 ( n8191, n8192, n8193 );
nand U7914 ( n8193, n8194, n8195 );
nand U7915 ( n8195, n8089, n8132 );
nand U7916 ( n8194, n8133, n7941 );
nor U7917 ( n8192, n8196, n8134 );
nor U7918 ( n8190, n8197, n8198 );
nor U7919 ( n8198, n8093, n8138 );
nor U7920 ( n8197, n8098, n8140 );
nand U7921 ( n950, n8199, n8200 );
nor U7922 ( n8200, n8201, n8202 );
nand U7923 ( n8202, n8203, n8204 );
nand U7924 ( n8204, n8106, n8132 );
nand U7925 ( n8203, n8133, n7931 );
nor U7926 ( n8201, n8205, n8134 );
nor U7927 ( n8199, n8206, n8207 );
nor U7928 ( n8207, n8108, n8138 );
nor U7929 ( n8206, n8111, n8140 );
nand U7930 ( n945, n8208, n8209 );
nor U7931 ( n8209, n8210, n8211 );
nand U7932 ( n8211, n8212, n8213 );
nand U7933 ( n8213, n8118, n8132 );
nand U7934 ( n8132, n8214, n8215 );
nand U7935 ( n8215, n8216, n7797 );
nand U7936 ( n8214, n8217, n8218 );
nand U7937 ( n8212, n8133, n8058 );
nand U7938 ( n8133, n8219, n8220 );
nor U7939 ( n8220, n8221, n8222 );
nor U7940 ( n8222, n15061, n8216 );
nand U7941 ( n8216, n8134, n8223 );
nand U7942 ( n8223, n8224, n8225 );
nor U7943 ( n8221, n8226, n8217 );
nand U7944 ( n8217, n8134, n8227 );
nand U7945 ( n8227, n8228, n8229 );
nor U7946 ( n8226, n8230, n8231 );
nor U7947 ( n8230, n8232, n8233 );
nand U7948 ( n8233, n8140, n8138 );
nor U7949 ( n8219, n8234, n8235 );
and U7950 ( n8234, n7815, n8134 );
nor U7951 ( n8210, n8119, n8134 );
nand U7952 ( n8134, n8236, n8237 );
nor U7953 ( n8208, n8238, n8239 );
nor U7954 ( n8239, n8124, n8138 );
nand U7955 ( n8138, n8240, n8241 );
nor U7956 ( n8238, n8121, n8140 );
nand U7957 ( n8140, n8242, n8243 );
nand U7958 ( n940, n8244, n8245 );
nor U7959 ( n8245, n8246, n8247 );
nand U7960 ( n8247, n8248, n8249 );
nand U7961 ( n8249, n8131, n8250 );
nand U7962 ( n8248, n8251, n7992 );
nor U7963 ( n8246, n8135, n8252 );
nor U7964 ( n8244, n8253, n8254 );
nor U7965 ( n8254, n8139, n8255 );
nor U7966 ( n8253, n8141, n8256 );
nand U7967 ( n935, n8257, n8258 );
nor U7968 ( n8258, n8259, n8260 );
nand U7969 ( n8260, n8261, n8262 );
nand U7970 ( n8262, n8148, n8250 );
nand U7971 ( n8261, n8251, n7982 );
nor U7972 ( n8259, n8149, n8252 );
nor U7973 ( n8257, n8263, n8264 );
nor U7974 ( n8264, n8152, n8255 );
nor U7975 ( n8263, n8153, n8256 );
nand U7976 ( n930, n8265, n8266 );
nor U7977 ( n8266, n8267, n8268 );
nand U7978 ( n8268, n8269, n8270 );
nand U7979 ( n8270, n8160, n8250 );
nand U7980 ( n8269, n8251, n7972 );
nor U7981 ( n8267, n8161, n8252 );
nor U7982 ( n8265, n8271, n8272 );
nor U7983 ( n8272, n8164, n8255 );
nor U7984 ( n8271, n8165, n8256 );
nand U7985 ( n925, n8273, n8274 );
nor U7986 ( n8274, n8275, n8276 );
nand U7987 ( n8276, n8277, n8278 );
nand U7988 ( n8278, n8172, n8250 );
nand U7989 ( n8277, n8251, n7962 );
nor U7990 ( n8275, n8173, n8252 );
nor U7991 ( n8273, n8279, n8280 );
nor U7992 ( n8280, n8176, n8255 );
nor U7993 ( n8279, n8177, n8256 );
nand U7994 ( n920, n8281, n8282 );
nor U7995 ( n8282, n8283, n8284 );
nand U7996 ( n8284, n8285, n8286 );
nand U7997 ( n8286, n8184, n8250 );
nand U7998 ( n8285, n8251, n7952 );
nor U7999 ( n8283, n8185, n8252 );
nor U8000 ( n8281, n8287, n8288 );
nor U8001 ( n8288, n8188, n8255 );
nor U8002 ( n8287, n8189, n8256 );
nand U8003 ( n915, n8289, n8290 );
nor U8004 ( n8290, n8291, n8292 );
nand U8005 ( n8292, n8293, n8294 );
nand U8006 ( n8294, n8089, n8250 );
nand U8007 ( n8293, n8251, n7942 );
nor U8008 ( n8291, n8196, n8252 );
nor U8009 ( n8289, n8295, n8296 );
nor U8010 ( n8296, n8093, n8255 );
nor U8011 ( n8295, n8098, n8256 );
nand U8012 ( n910, n8297, n8298 );
nor U8013 ( n8298, n8299, n8300 );
nand U8014 ( n8300, n8301, n8302 );
nand U8015 ( n8302, n8106, n8250 );
nand U8016 ( n8301, n8251, n7932 );
nor U8017 ( n8299, n8205, n8252 );
nor U8018 ( n8297, n8303, n8304 );
nor U8019 ( n8304, n8108, n8255 );
nor U8020 ( n8303, n8111, n8256 );
nand U8021 ( n905, n8305, n8306 );
nor U8022 ( n8306, n8307, n8308 );
nand U8023 ( n8308, n8309, n8310 );
nand U8024 ( n8310, n8118, n8250 );
nand U8025 ( n8250, n8311, n8312 );
nand U8026 ( n8312, n8313, n8229 );
nand U8027 ( n8311, n8314, n8225 );
nand U8028 ( n8309, n8251, n8059 );
nand U8029 ( n8251, n8315, n8316 );
not U8030 ( n8316, n8317 );
nor U8031 ( n8315, n8318, n8319 );
and U8032 ( n8318, n7815, n8252 );
nor U8033 ( n8307, n8119, n8252 );
nand U8034 ( n8252, n8320, n8237 );
nor U8035 ( n8305, n8321, n8322 );
nor U8036 ( n8322, n8124, n8255 );
nand U8037 ( n8255, n8323, n8241 );
nor U8038 ( n8321, n8121, n8256 );
nand U8039 ( n8256, n8324, n8243 );
nand U8040 ( n900, n8325, n8326 );
nor U8041 ( n8326, n8327, n8328 );
nand U8042 ( n8328, n8329, n8330 );
nand U8043 ( n8330, n8131, n8331 );
nand U8044 ( n8329, n8332, n7993 );
nor U8045 ( n8327, n8141, n8333 );
nor U8046 ( n8325, n8334, n8335 );
nor U8047 ( n8335, n8139, n8336 );
nor U8048 ( n8334, n8135, n8337 );
nand U8049 ( n895, n8338, n8339 );
nor U8050 ( n8339, n8340, n8341 );
nand U8051 ( n8341, n8342, n8343 );
nand U8052 ( n8343, n8148, n8331 );
nand U8053 ( n8342, n8332, n7983 );
nor U8054 ( n8340, n8153, n8333 );
nor U8055 ( n8338, n8344, n8345 );
nor U8056 ( n8345, n8152, n8336 );
nor U8057 ( n8344, n8149, n8337 );
nand U8058 ( n890, n8346, n8347 );
nor U8059 ( n8347, n8348, n8349 );
nand U8060 ( n8349, n8350, n8351 );
nand U8061 ( n8351, n8160, n8331 );
nand U8062 ( n8350, n8332, n7973 );
nor U8063 ( n8348, n8165, n8333 );
nor U8064 ( n8346, n8352, n8353 );
nor U8065 ( n8353, n8164, n8336 );
nor U8066 ( n8352, n8161, n8337 );
nand U8067 ( n885, n8354, n8355 );
nor U8068 ( n8355, n8356, n8357 );
nand U8069 ( n8357, n8358, n8359 );
nand U8070 ( n8359, n8172, n8331 );
nand U8071 ( n8358, n8332, n7963 );
nor U8072 ( n8356, n8177, n8333 );
nor U8073 ( n8354, n8360, n8361 );
nor U8074 ( n8361, n8176, n8336 );
nor U8075 ( n8360, n8173, n8337 );
nand U8076 ( n880, n8362, n8363 );
nor U8077 ( n8363, n8364, n8365 );
nand U8078 ( n8365, n8366, n8367 );
nand U8079 ( n8367, n8184, n8331 );
nand U8080 ( n8366, n8332, n7953 );
nor U8081 ( n8364, n8189, n8333 );
nor U8082 ( n8362, n8368, n8369 );
nor U8083 ( n8369, n8188, n8336 );
nor U8084 ( n8368, n8185, n8337 );
nand U8085 ( n875, n8370, n8371 );
nor U8086 ( n8371, n8372, n8373 );
nand U8087 ( n8373, n8374, n8375 );
nand U8088 ( n8375, n8089, n8331 );
nand U8089 ( n8374, n8332, n7943 );
nor U8090 ( n8372, n8098, n8333 );
nor U8091 ( n8370, n8376, n8377 );
nor U8092 ( n8377, n8093, n8336 );
nor U8093 ( n8376, n8196, n8337 );
nand U8094 ( n870, n8378, n8379 );
nor U8095 ( n8379, n8380, n8381 );
nand U8096 ( n8381, n8382, n8383 );
nand U8097 ( n8383, n8106, n8331 );
nand U8098 ( n8382, n8332, n7933 );
nor U8099 ( n8380, n8111, n8333 );
nor U8100 ( n8378, n8384, n8385 );
nor U8101 ( n8385, n8108, n8336 );
nor U8102 ( n8384, n8205, n8337 );
nand U8103 ( n865, n8386, n8387 );
nor U8104 ( n8387, n8388, n8389 );
nand U8105 ( n8389, n8390, n8391 );
nand U8106 ( n8391, n8118, n8331 );
nand U8107 ( n8331, n8392, n8393 );
nand U8108 ( n8393, n8394, n7797 );
nand U8109 ( n8392, n8395, n8218 );
nand U8110 ( n8390, n8332, n8060 );
nand U8111 ( n8332, n8396, n8397 );
nor U8112 ( n8397, n8398, n8399 );
nor U8113 ( n8399, n15061, n8394 );
nand U8114 ( n8394, n8337, n8400 );
nand U8115 ( n8400, n8401, n8225 );
nor U8116 ( n8398, n8402, n8395 );
nand U8117 ( n8395, n8337, n8403 );
nand U8118 ( n8403, n8404, n8229 );
nor U8119 ( n8402, n8405, n8231 );
nor U8120 ( n8405, n8232, n8406 );
nand U8121 ( n8406, n8333, n8336 );
nor U8122 ( n8396, n8407, n8235 );
nor U8123 ( n8407, n15060, n8408 );
nor U8124 ( n8388, n8121, n8333 );
nor U8125 ( n8386, n8409, n8410 );
nor U8126 ( n8410, n8124, n8336 );
nor U8127 ( n8409, n8119, n8337 );
nand U8128 ( n860, n8411, n8412 );
nor U8129 ( n8412, n8413, n8414 );
nand U8130 ( n8414, n8415, n8416 );
nand U8131 ( n8416, n8131, n8417 );
nand U8132 ( n8415, n8418, n7871 );
nor U8133 ( n8413, n8135, n8419 );
nor U8134 ( n8411, n8420, n8421 );
nor U8135 ( n8421, n8139, n8422 );
nor U8136 ( n8420, n8141, n8423 );
nand U8137 ( n855, n8424, n8425 );
nor U8138 ( n8425, n8426, n8427 );
nand U8139 ( n8427, n8428, n8429 );
nand U8140 ( n8429, n8148, n8417 );
nand U8141 ( n8428, n8418, n7870 );
nor U8142 ( n8426, n8149, n8419 );
nor U8143 ( n8424, n8430, n8431 );
nor U8144 ( n8431, n8152, n8422 );
nor U8145 ( n8430, n8153, n8423 );
nand U8146 ( n850, n8432, n8433 );
nor U8147 ( n8433, n8434, n8435 );
nand U8148 ( n8435, n8436, n8437 );
nand U8149 ( n8437, n8160, n8417 );
nand U8150 ( n8436, n8418, n7869 );
nor U8151 ( n8434, n8161, n8419 );
nor U8152 ( n8432, n8438, n8439 );
nor U8153 ( n8439, n8164, n8422 );
nor U8154 ( n8438, n8165, n8423 );
nand U8155 ( n845, n8440, n8441 );
nor U8156 ( n8441, n8442, n8443 );
nand U8157 ( n8443, n8444, n8445 );
nand U8158 ( n8445, n8172, n8417 );
nand U8159 ( n8444, n8418, n7868 );
nor U8160 ( n8442, n8173, n8419 );
nor U8161 ( n8440, n8446, n8447 );
nor U8162 ( n8447, n8176, n8422 );
nor U8163 ( n8446, n8177, n8423 );
nand U8164 ( n840, n8448, n8449 );
nor U8165 ( n8449, n8450, n8451 );
nand U8166 ( n8451, n8452, n8453 );
nand U8167 ( n8453, n8184, n8417 );
nand U8168 ( n8452, n8418, n7867 );
nor U8169 ( n8450, n8185, n8419 );
nor U8170 ( n8448, n8454, n8455 );
nor U8171 ( n8455, n8188, n8422 );
nor U8172 ( n8454, n8189, n8423 );
nand U8173 ( n835, n8456, n8457 );
nor U8174 ( n8457, n8458, n8459 );
nand U8175 ( n8459, n8460, n8461 );
nand U8176 ( n8461, n8089, n8417 );
nand U8177 ( n8460, n8418, n7866 );
nor U8178 ( n8458, n8196, n8419 );
nor U8179 ( n8456, n8462, n8463 );
nor U8180 ( n8463, n8093, n8422 );
nor U8181 ( n8462, n8098, n8423 );
nand U8182 ( n830, n8464, n8465 );
nor U8183 ( n8465, n8466, n8467 );
nand U8184 ( n8467, n8468, n8469 );
nand U8185 ( n8469, n8106, n8417 );
nand U8186 ( n8468, n8418, n7865 );
nor U8187 ( n8466, n8205, n8419 );
nor U8188 ( n8464, n8470, n8471 );
nor U8189 ( n8471, n8108, n8422 );
nor U8190 ( n8470, n8111, n8423 );
nand U8191 ( n825, n8472, n8473 );
nor U8192 ( n8473, n8474, n8475 );
nand U8193 ( n8475, n8476, n8477 );
nand U8194 ( n8477, n8118, n8417 );
nand U8195 ( n8417, n8478, n8479 );
nand U8196 ( n8479, n8480, n8218 );
nand U8197 ( n8478, n8481, n8482 );
nand U8198 ( n8476, n8418, n7994 );
nand U8199 ( n8418, n8483, n8484 );
nor U8200 ( n8484, n8485, n8486 );
and U8201 ( n8486, n7815, n8419 );
nor U8202 ( n8485, n8487, n8480 );
nand U8203 ( n8480, n8419, n8488 );
nand U8204 ( n8488, n8489, n8490 );
nor U8205 ( n8487, n8491, n8231 );
and U8206 ( n8491, n8422, n8423 );
nor U8207 ( n8483, n8492, n8235 );
nor U8208 ( n8492, n15061, n8481 );
nor U8209 ( n8474, n8119, n8419 );
nand U8210 ( n8419, n8493, n8494 );
nor U8211 ( n8472, n8495, n8496 );
nor U8212 ( n8496, n8124, n8422 );
nand U8213 ( n8422, n8497, n8498 );
nor U8214 ( n8495, n8121, n8423 );
nand U8215 ( n8423, n8499, n8500 );
nand U8216 ( n820, n8501, n8502 );
nor U8217 ( n8502, n8503, n8504 );
nand U8218 ( n8504, n8505, n8506 );
nand U8219 ( n8506, n8131, n8507 );
nand U8220 ( n8505, n8508, n7984 );
nor U8221 ( n8503, n8135, n8509 );
nor U8222 ( n8501, n8510, n8511 );
nor U8223 ( n8511, n8139, n8512 );
nor U8224 ( n8510, n8141, n8513 );
nand U8225 ( n815, n8514, n8515 );
nor U8226 ( n8515, n8516, n8517 );
nand U8227 ( n8517, n8518, n8519 );
nand U8228 ( n8519, n8148, n8507 );
nand U8229 ( n8518, n8508, n7974 );
nor U8230 ( n8516, n8149, n8509 );
nor U8231 ( n8514, n8520, n8521 );
nor U8232 ( n8521, n8152, n8512 );
nor U8233 ( n8520, n8153, n8513 );
nand U8234 ( n810, n8522, n8523 );
nor U8235 ( n8523, n8524, n8525 );
nand U8236 ( n8525, n8526, n8527 );
nand U8237 ( n8527, n8160, n8507 );
nand U8238 ( n8526, n8508, n7964 );
nor U8239 ( n8524, n8161, n8509 );
nor U8240 ( n8522, n8528, n8529 );
nor U8241 ( n8529, n8164, n8512 );
nor U8242 ( n8528, n8165, n8513 );
nand U8243 ( n805, n8530, n8531 );
nor U8244 ( n8531, n8532, n8533 );
nand U8245 ( n8533, n8534, n8535 );
nand U8246 ( n8535, n8172, n8507 );
nand U8247 ( n8534, n8508, n7954 );
nor U8248 ( n8532, n8173, n8509 );
nor U8249 ( n8530, n8536, n8537 );
nor U8250 ( n8537, n8176, n8512 );
nor U8251 ( n8536, n8177, n8513 );
nand U8252 ( n800, n8538, n8539 );
nor U8253 ( n8539, n8540, n8541 );
nand U8254 ( n8541, n8542, n8543 );
nand U8255 ( n8543, n8184, n8507 );
nand U8256 ( n8542, n8508, n7944 );
nor U8257 ( n8540, n8185, n8509 );
nor U8258 ( n8538, n8544, n8545 );
nor U8259 ( n8545, n8188, n8512 );
nor U8260 ( n8544, n8189, n8513 );
nand U8261 ( n795, n8546, n8547 );
nor U8262 ( n8547, n8548, n8549 );
nand U8263 ( n8549, n8550, n8551 );
nand U8264 ( n8551, n8089, n8507 );
nand U8265 ( n8550, n8508, n7934 );
nor U8266 ( n8548, n8196, n8509 );
nor U8267 ( n8546, n8552, n8553 );
nor U8268 ( n8553, n8093, n8512 );
nor U8269 ( n8552, n8098, n8513 );
nand U8270 ( n790, n8554, n8555 );
nor U8271 ( n8555, n8556, n8557 );
nand U8272 ( n8557, n8558, n8559 );
nand U8273 ( n8559, n8106, n8507 );
nand U8274 ( n8558, n8508, n7924 );
nor U8275 ( n8556, n8205, n8509 );
nor U8276 ( n8554, n8560, n8561 );
nor U8277 ( n8561, n8108, n8512 );
nor U8278 ( n8560, n8111, n8513 );
nand U8279 ( n785, n8562, n8563 );
nor U8280 ( n8563, n8564, n8565 );
nand U8281 ( n8565, n8566, n8567 );
nand U8282 ( n8567, n8118, n8507 );
nand U8283 ( n8507, n8568, n8569 );
nand U8284 ( n8569, n8570, n7797 );
nand U8285 ( n8568, n8571, n8218 );
nand U8286 ( n8566, n8508, n8061 );
nand U8287 ( n8508, n8572, n8573 );
nor U8288 ( n8573, n8574, n8575 );
nor U8289 ( n8575, n15061, n8570 );
nand U8290 ( n8570, n8509, n8576 );
nand U8291 ( n8576, n8481, n8224 );
nor U8292 ( n8574, n8577, n8571 );
nand U8293 ( n8571, n8509, n8578 );
nand U8294 ( n8578, n8489, n8228 );
nor U8295 ( n8577, n8579, n8231 );
nor U8296 ( n8579, n8232, n8580 );
nand U8297 ( n8580, n8513, n8512 );
nor U8298 ( n8572, n8581, n8235 );
and U8299 ( n8581, n7815, n8509 );
nor U8300 ( n8564, n8119, n8509 );
nand U8301 ( n8509, n8493, n8236 );
nor U8302 ( n8562, n8582, n8583 );
nor U8303 ( n8583, n8124, n8512 );
nand U8304 ( n8512, n8497, n8240 );
nor U8305 ( n8582, n8121, n8513 );
nand U8306 ( n8513, n8499, n8242 );
nand U8307 ( n780, n8584, n8585 );
nor U8308 ( n8585, n8586, n8587 );
nand U8309 ( n8587, n8588, n8589 );
nand U8310 ( n8589, n8131, n8590 );
nand U8311 ( n8588, n8591, n7985 );
nor U8312 ( n8586, n8135, n8592 );
nor U8313 ( n8584, n8593, n8594 );
nor U8314 ( n8594, n8139, n8595 );
nor U8315 ( n8593, n8141, n8596 );
nand U8316 ( n775, n8597, n8598 );
nor U8317 ( n8598, n8599, n8600 );
nand U8318 ( n8600, n8601, n8602 );
nand U8319 ( n8602, n8148, n8590 );
nand U8320 ( n8601, n8591, n7975 );
nor U8321 ( n8599, n8149, n8592 );
nor U8322 ( n8597, n8603, n8604 );
nor U8323 ( n8604, n8152, n8595 );
nor U8324 ( n8603, n8153, n8596 );
nand U8325 ( n770, n8605, n8606 );
nor U8326 ( n8606, n8607, n8608 );
nand U8327 ( n8608, n8609, n8610 );
nand U8328 ( n8610, n8160, n8590 );
nand U8329 ( n8609, n8591, n7965 );
nor U8330 ( n8607, n8161, n8592 );
nor U8331 ( n8605, n8611, n8612 );
nor U8332 ( n8612, n8164, n8595 );
nor U8333 ( n8611, n8165, n8596 );
nand U8334 ( n765, n8613, n8614 );
nor U8335 ( n8614, n8615, n8616 );
nand U8336 ( n8616, n8617, n8618 );
nand U8337 ( n8618, n8172, n8590 );
nand U8338 ( n8617, n8591, n7955 );
nor U8339 ( n8615, n8173, n8592 );
nor U8340 ( n8613, n8619, n8620 );
nor U8341 ( n8620, n8176, n8595 );
nor U8342 ( n8619, n8177, n8596 );
nand U8343 ( n760, n8621, n8622 );
nor U8344 ( n8622, n8623, n8624 );
nand U8345 ( n8624, n8625, n8626 );
nand U8346 ( n8626, n8184, n8590 );
nand U8347 ( n8625, n8591, n7945 );
nor U8348 ( n8623, n8185, n8592 );
nor U8349 ( n8621, n8627, n8628 );
nor U8350 ( n8628, n8188, n8595 );
nor U8351 ( n8627, n8189, n8596 );
nand U8352 ( n755, n8629, n8630 );
nor U8353 ( n8630, n8631, n8632 );
nand U8354 ( n8632, n8633, n8634 );
nand U8355 ( n8634, n8089, n8590 );
nand U8356 ( n8633, n8591, n7935 );
nor U8357 ( n8631, n8196, n8592 );
nor U8358 ( n8629, n8635, n8636 );
nor U8359 ( n8636, n8093, n8595 );
nor U8360 ( n8635, n8098, n8596 );
nand U8361 ( n750, n8637, n8638 );
nor U8362 ( n8638, n8639, n8640 );
nand U8363 ( n8640, n8641, n8642 );
nand U8364 ( n8642, n8106, n8590 );
nand U8365 ( n8641, n8591, n7925 );
nor U8366 ( n8639, n8205, n8592 );
nor U8367 ( n8637, n8643, n8644 );
nor U8368 ( n8644, n8108, n8595 );
nor U8369 ( n8643, n8111, n8596 );
nand U8370 ( n745, n8645, n8646 );
nor U8371 ( n8646, n8647, n8648 );
nand U8372 ( n8648, n8649, n8650 );
nand U8373 ( n8650, n8118, n8590 );
nand U8374 ( n8590, n8651, n8652 );
nand U8375 ( n8652, n8489, n8313 );
nand U8376 ( n8651, n8481, n8314 );
nand U8377 ( n8649, n8591, n8062 );
nand U8378 ( n8591, n8653, n8481 );
nor U8379 ( n8653, n8654, n8317 );
and U8380 ( n8654, n7815, n8592 );
nor U8381 ( n8647, n8119, n8592 );
nand U8382 ( n8592, n8493, n8320 );
nor U8383 ( n8645, n8655, n8656 );
nor U8384 ( n8656, n8124, n8595 );
nand U8385 ( n8595, n8497, n8323 );
nor U8386 ( n8655, n8121, n8596 );
nand U8387 ( n8596, n8499, n8324 );
nand U8388 ( n740, n8657, n8658 );
nor U8389 ( n8658, n8659, n8660 );
nand U8390 ( n8660, n8661, n8662 );
nand U8391 ( n8662, n8131, n8663 );
nand U8392 ( n8661, n8664, n7986 );
nor U8393 ( n8659, n8135, n8665 );
nor U8394 ( n8657, n8666, n8667 );
nor U8395 ( n8667, n8139, n8668 );
nor U8396 ( n8666, n8141, n8669 );
nand U8397 ( n735, n8670, n8671 );
nor U8398 ( n8671, n8672, n8673 );
nand U8399 ( n8673, n8674, n8675 );
nand U8400 ( n8675, n8148, n8663 );
nand U8401 ( n8674, n8664, n7976 );
nor U8402 ( n8672, n8149, n8665 );
nor U8403 ( n8670, n8676, n8677 );
nor U8404 ( n8677, n8152, n8668 );
nor U8405 ( n8676, n8153, n8669 );
nand U8406 ( n730, n8678, n8679 );
nor U8407 ( n8679, n8680, n8681 );
nand U8408 ( n8681, n8682, n8683 );
nand U8409 ( n8683, n8160, n8663 );
nand U8410 ( n8682, n8664, n7966 );
nor U8411 ( n8680, n8161, n8665 );
nor U8412 ( n8678, n8684, n8685 );
nor U8413 ( n8685, n8164, n8668 );
nor U8414 ( n8684, n8165, n8669 );
nand U8415 ( n725, n8686, n8687 );
nor U8416 ( n8687, n8688, n8689 );
nand U8417 ( n8689, n8690, n8691 );
nand U8418 ( n8691, n8172, n8663 );
nand U8419 ( n8690, n8664, n7956 );
nor U8420 ( n8688, n8173, n8665 );
nor U8421 ( n8686, n8692, n8693 );
nor U8422 ( n8693, n8176, n8668 );
nor U8423 ( n8692, n8177, n8669 );
nand U8424 ( n720, n8694, n8695 );
nor U8425 ( n8695, n8696, n8697 );
nand U8426 ( n8697, n8698, n8699 );
nand U8427 ( n8699, n8184, n8663 );
nand U8428 ( n8698, n8664, n7946 );
nor U8429 ( n8696, n8185, n8665 );
nor U8430 ( n8694, n8700, n8701 );
nor U8431 ( n8701, n8188, n8668 );
nor U8432 ( n8700, n8189, n8669 );
nand U8433 ( n715, n8702, n8703 );
nor U8434 ( n8703, n8704, n8705 );
nand U8435 ( n8705, n8706, n8707 );
nand U8436 ( n8707, n8089, n8663 );
nand U8437 ( n8706, n8664, n7936 );
nor U8438 ( n8704, n8196, n8665 );
nor U8439 ( n8702, n8708, n8709 );
nor U8440 ( n8709, n8093, n8668 );
nor U8441 ( n8708, n8098, n8669 );
nand U8442 ( n710, n8710, n8711 );
nor U8443 ( n8711, n8712, n8713 );
nand U8444 ( n8713, n8714, n8715 );
nand U8445 ( n8715, n8106, n8663 );
nand U8446 ( n8714, n8664, n7926 );
nor U8447 ( n8712, n8205, n8665 );
nor U8448 ( n8710, n8716, n8717 );
nor U8449 ( n8717, n8108, n8668 );
nor U8450 ( n8716, n8111, n8669 );
nand U8451 ( n705, n8718, n8719 );
nor U8452 ( n8719, n8720, n8721 );
nand U8453 ( n8721, n8722, n8723 );
nand U8454 ( n8723, n8118, n8663 );
nand U8455 ( n8663, n8724, n8725 );
nand U8456 ( n8725, n8726, n7797 );
nand U8457 ( n8724, n8727, n8218 );
nand U8458 ( n8722, n8664, n8063 );
nand U8459 ( n8664, n8728, n8729 );
nor U8460 ( n8729, n8730, n8731 );
nor U8461 ( n8731, n15061, n8726 );
nand U8462 ( n8726, n8665, n8732 );
nand U8463 ( n8732, n8481, n8401 );
nor U8464 ( n8481, n8733, n8734 );
nor U8465 ( n8730, n8735, n8727 );
nand U8466 ( n8727, n8665, n8736 );
nand U8467 ( n8736, n8489, n8404 );
nor U8468 ( n8489, n8737, n8738 );
nor U8469 ( n8735, n8739, n8231 );
nor U8470 ( n8739, n8232, n8740 );
nand U8471 ( n8740, n8669, n8668 );
nor U8472 ( n8728, n8741, n8235 );
and U8473 ( n8741, n7815, n8665 );
nor U8474 ( n8720, n8119, n8665 );
nand U8475 ( n8665, n8493, n8742 );
nor U8476 ( n8718, n8743, n8744 );
nor U8477 ( n8744, n8124, n8668 );
nand U8478 ( n8668, n8497, n8745 );
nor U8479 ( n8743, n8121, n8669 );
nand U8480 ( n8669, n8499, n8746 );
nor U8481 ( n8499, n8747, n8748 );
nand U8482 ( n700, n8749, n8750 );
nor U8483 ( n8750, n8751, n8752 );
nand U8484 ( n8752, n8753, n8754 );
nand U8485 ( n8754, n8131, n8755 );
nand U8486 ( n8753, n8756, n7988 );
nor U8487 ( n8751, n8135, n8757 );
nor U8488 ( n8749, n8758, n8759 );
nor U8489 ( n8759, n8139, n8760 );
nor U8490 ( n8758, n8141, n8761 );
nand U8491 ( n695, n8762, n8763 );
nor U8492 ( n8763, n8764, n8765 );
nand U8493 ( n8765, n8766, n8767 );
nand U8494 ( n8767, n8148, n8755 );
nand U8495 ( n8766, n8756, n7978 );
nor U8496 ( n8764, n8149, n8757 );
nor U8497 ( n8762, n8768, n8769 );
nor U8498 ( n8769, n8152, n8760 );
nor U8499 ( n8768, n8153, n8761 );
nand U8500 ( n690, n8770, n8771 );
nor U8501 ( n8771, n8772, n8773 );
nand U8502 ( n8773, n8774, n8775 );
nand U8503 ( n8775, n8160, n8755 );
nand U8504 ( n8774, n8756, n7968 );
nor U8505 ( n8772, n8161, n8757 );
nor U8506 ( n8770, n8776, n8777 );
nor U8507 ( n8777, n8164, n8760 );
nor U8508 ( n8776, n8165, n8761 );
nand U8509 ( n685, n8778, n8779 );
nor U8510 ( n8779, n8780, n8781 );
nand U8511 ( n8781, n8782, n8783 );
nand U8512 ( n8783, n8172, n8755 );
nand U8513 ( n8782, n8756, n7958 );
nor U8514 ( n8780, n8173, n8757 );
nor U8515 ( n8778, n8784, n8785 );
nor U8516 ( n8785, n8176, n8760 );
nor U8517 ( n8784, n8177, n8761 );
nand U8518 ( n680, n8786, n8787 );
nor U8519 ( n8787, n8788, n8789 );
nand U8520 ( n8789, n8790, n8791 );
nand U8521 ( n8791, n8184, n8755 );
nand U8522 ( n8790, n8756, n7948 );
nor U8523 ( n8788, n8185, n8757 );
nor U8524 ( n8786, n8792, n8793 );
nor U8525 ( n8793, n8188, n8760 );
nor U8526 ( n8792, n8189, n8761 );
nand U8527 ( n675, n8794, n8795 );
nor U8528 ( n8795, n8796, n8797 );
nand U8529 ( n8797, n8798, n8799 );
nand U8530 ( n8799, n8089, n8755 );
nand U8531 ( n8798, n8756, n7938 );
nor U8532 ( n8796, n8196, n8757 );
nor U8533 ( n8794, n8800, n8801 );
nor U8534 ( n8801, n8093, n8760 );
nor U8535 ( n8800, n8098, n8761 );
nand U8536 ( n670, n8802, n8803 );
nor U8537 ( n8803, n8804, n8805 );
nand U8538 ( n8805, n8806, n8807 );
nand U8539 ( n8807, n8106, n8755 );
nand U8540 ( n8806, n8756, n7928 );
nor U8541 ( n8804, n8205, n8757 );
nor U8542 ( n8802, n8808, n8809 );
nor U8543 ( n8809, n8108, n8760 );
nor U8544 ( n8808, n8111, n8761 );
nand U8545 ( n665, n8810, n8811 );
nor U8546 ( n8811, n8812, n8813 );
nand U8547 ( n8813, n8814, n8815 );
nand U8548 ( n8815, n8118, n8755 );
nand U8549 ( n8755, n8816, n8817 );
nand U8550 ( n8817, n8818, n8218 );
nand U8551 ( n8816, n8819, n8482 );
nand U8552 ( n8814, n8756, n8064 );
nand U8553 ( n8756, n8820, n8821 );
nor U8554 ( n8821, n8822, n8823 );
and U8555 ( n8823, n7815, n8757 );
nor U8556 ( n8822, n8824, n8818 );
nand U8557 ( n8818, n8757, n8825 );
nand U8558 ( n8825, n8826, n8490 );
nor U8559 ( n8824, n8827, n8231 );
and U8560 ( n8827, n8760, n8761 );
nor U8561 ( n8820, n8828, n8235 );
nor U8562 ( n8828, n15061, n8819 );
nor U8563 ( n8812, n8119, n8757 );
nand U8564 ( n8757, n8829, n8494 );
nor U8565 ( n8810, n8830, n8831 );
nor U8566 ( n8831, n8124, n8760 );
nand U8567 ( n8760, n8832, n8498 );
nor U8568 ( n8830, n8121, n8761 );
nand U8569 ( n8761, n8833, n8500 );
nand U8570 ( n660, n8834, n8835 );
nor U8571 ( n8835, n8836, n8837 );
nand U8572 ( n8837, n8838, n8839 );
nand U8573 ( n8839, n8131, n8840 );
nand U8574 ( n8838, n8841, n7987 );
nor U8575 ( n8836, n8135, n8842 );
nor U8576 ( n8834, n8843, n8844 );
nor U8577 ( n8844, n8139, n8845 );
nor U8578 ( n8843, n8141, n8846 );
nand U8579 ( n655, n8847, n8848 );
nor U8580 ( n8848, n8849, n8850 );
nand U8581 ( n8850, n8851, n8852 );
nand U8582 ( n8852, n8148, n8840 );
nand U8583 ( n8851, n8841, n7977 );
nor U8584 ( n8849, n8149, n8842 );
nor U8585 ( n8847, n8853, n8854 );
nor U8586 ( n8854, n8152, n8845 );
nor U8587 ( n8853, n8153, n8846 );
nand U8588 ( n650, n8855, n8856 );
nor U8589 ( n8856, n8857, n8858 );
nand U8590 ( n8858, n8859, n8860 );
nand U8591 ( n8860, n8160, n8840 );
nand U8592 ( n8859, n8841, n7967 );
nor U8593 ( n8857, n8161, n8842 );
nor U8594 ( n8855, n8861, n8862 );
nor U8595 ( n8862, n8164, n8845 );
nor U8596 ( n8861, n8165, n8846 );
nand U8597 ( n645, n8863, n8864 );
nor U8598 ( n8864, n8865, n8866 );
nand U8599 ( n8866, n8867, n8868 );
nand U8600 ( n8868, n8172, n8840 );
nand U8601 ( n8867, n8841, n7957 );
nor U8602 ( n8865, n8173, n8842 );
nor U8603 ( n8863, n8869, n8870 );
nor U8604 ( n8870, n8176, n8845 );
nor U8605 ( n8869, n8177, n8846 );
nand U8606 ( n640, n8871, n8872 );
nor U8607 ( n8872, n8873, n8874 );
nand U8608 ( n8874, n8875, n8876 );
nand U8609 ( n8876, n8184, n8840 );
nand U8610 ( n8875, n8841, n7947 );
nor U8611 ( n8873, n8185, n8842 );
nor U8612 ( n8871, n8877, n8878 );
nor U8613 ( n8878, n8188, n8845 );
nor U8614 ( n8877, n8189, n8846 );
nand U8615 ( n635, n8879, n8880 );
nor U8616 ( n8880, n8881, n8882 );
nand U8617 ( n8882, n8883, n8884 );
nand U8618 ( n8884, n8089, n8840 );
nand U8619 ( n8883, n8841, n7937 );
nor U8620 ( n8881, n8196, n8842 );
nor U8621 ( n8879, n8885, n8886 );
nor U8622 ( n8886, n8093, n8845 );
nor U8623 ( n8885, n8098, n8846 );
nand U8624 ( n630, n8887, n8888 );
nor U8625 ( n8888, n8889, n8890 );
nand U8626 ( n8890, n8891, n8892 );
nand U8627 ( n8892, n8106, n8840 );
nand U8628 ( n8891, n8841, n7927 );
nor U8629 ( n8889, n8205, n8842 );
nor U8630 ( n8887, n8893, n8894 );
nor U8631 ( n8894, n8108, n8845 );
nor U8632 ( n8893, n8111, n8846 );
nand U8633 ( n625, n8895, n8896 );
nor U8634 ( n8896, n8897, n8898 );
nand U8635 ( n8898, n8899, n8900 );
nand U8636 ( n8900, n8118, n8840 );
nand U8637 ( n8840, n8901, n8902 );
nand U8638 ( n8902, n8903, n7797 );
nand U8639 ( n8901, n8904, n8218 );
nand U8640 ( n8899, n8841, n8065 );
nand U8641 ( n8841, n8905, n8906 );
nor U8642 ( n8906, n8907, n8908 );
nor U8643 ( n8908, n15061, n8903 );
nand U8644 ( n8903, n8842, n8909 );
nand U8645 ( n8909, n8819, n8224 );
nor U8646 ( n8907, n8910, n8904 );
nand U8647 ( n8904, n8842, n8911 );
nand U8648 ( n8911, n8826, n8228 );
nor U8649 ( n8910, n8912, n8231 );
nor U8650 ( n8912, n8232, n8913 );
nand U8651 ( n8913, n8846, n8845 );
nor U8652 ( n8905, n8914, n8235 );
and U8653 ( n8914, n7815, n8842 );
nor U8654 ( n8897, n8119, n8842 );
nand U8655 ( n8842, n8829, n8236 );
nor U8656 ( n8895, n8915, n8916 );
nor U8657 ( n8916, n8124, n8845 );
nand U8658 ( n8845, n8832, n8240 );
nor U8659 ( n8915, n8121, n8846 );
nand U8660 ( n8846, n8833, n8242 );
nand U8661 ( n620, n8917, n8918 );
nor U8662 ( n8918, n8919, n8920 );
nand U8663 ( n8920, n8921, n8922 );
nand U8664 ( n8922, n8131, n8923 );
nand U8665 ( n8921, n8924, n7989 );
nor U8666 ( n8919, n8135, n8925 );
nor U8667 ( n8917, n8926, n8927 );
nor U8668 ( n8927, n8139, n8928 );
nor U8669 ( n8926, n8141, n8929 );
nand U8670 ( n615, n8930, n8931 );
nor U8671 ( n8931, n8932, n8933 );
nand U8672 ( n8933, n8934, n8935 );
nand U8673 ( n8935, n8148, n8923 );
nand U8674 ( n8934, n8924, n7979 );
nor U8675 ( n8932, n8149, n8925 );
nor U8676 ( n8930, n8936, n8937 );
nor U8677 ( n8937, n8152, n8928 );
nor U8678 ( n8936, n8153, n8929 );
nand U8679 ( n610, n8938, n8939 );
nor U8680 ( n8939, n8940, n8941 );
nand U8681 ( n8941, n8942, n8943 );
nand U8682 ( n8943, n8160, n8923 );
nand U8683 ( n8942, n8924, n7969 );
nor U8684 ( n8940, n8161, n8925 );
nor U8685 ( n8938, n8944, n8945 );
nor U8686 ( n8945, n8164, n8928 );
nor U8687 ( n8944, n8165, n8929 );
nand U8688 ( n605, n8946, n8947 );
nor U8689 ( n8947, n8948, n8949 );
nand U8690 ( n8949, n8950, n8951 );
nand U8691 ( n8951, n8172, n8923 );
nand U8692 ( n8950, n8924, n7959 );
nor U8693 ( n8948, n8173, n8925 );
nor U8694 ( n8946, n8952, n8953 );
nor U8695 ( n8953, n8176, n8928 );
nor U8696 ( n8952, n8177, n8929 );
nand U8697 ( n600, n8954, n8955 );
nor U8698 ( n8955, n8956, n8957 );
nand U8699 ( n8957, n8958, n8959 );
nand U8700 ( n8959, n8184, n8923 );
nand U8701 ( n8958, n8924, n7949 );
nor U8702 ( n8956, n8185, n8925 );
nor U8703 ( n8954, n8960, n8961 );
nor U8704 ( n8961, n8188, n8928 );
nor U8705 ( n8960, n8189, n8929 );
nand U8706 ( n595, n8962, n8963 );
nor U8707 ( n8963, n8964, n8965 );
nand U8708 ( n8965, n8966, n8967 );
nand U8709 ( n8967, n8089, n8923 );
nand U8710 ( n8966, n8924, n7939 );
nor U8711 ( n8964, n8196, n8925 );
nor U8712 ( n8962, n8968, n8969 );
nor U8713 ( n8969, n8093, n8928 );
nor U8714 ( n8968, n8098, n8929 );
nand U8715 ( n590, n8970, n8971 );
nor U8716 ( n8971, n8972, n8973 );
nand U8717 ( n8973, n8974, n8975 );
nand U8718 ( n8975, n8106, n8923 );
nand U8719 ( n8974, n8924, n7929 );
nor U8720 ( n8972, n8205, n8925 );
nor U8721 ( n8970, n8976, n8977 );
nor U8722 ( n8977, n8108, n8928 );
nor U8723 ( n8976, n8111, n8929 );
nand U8724 ( n585, n8978, n8979 );
nor U8725 ( n8979, n8980, n8981 );
nand U8726 ( n8981, n8982, n8983 );
nand U8727 ( n8983, n8118, n8923 );
nand U8728 ( n8923, n8984, n8985 );
nand U8729 ( n8985, n8826, n8313 );
nand U8730 ( n8984, n8819, n8314 );
nand U8731 ( n8982, n8924, n8066 );
nand U8732 ( n8924, n8986, n8819 );
nor U8733 ( n8986, n8987, n8317 );
and U8734 ( n8987, n7815, n8925 );
nor U8735 ( n8980, n8119, n8925 );
nand U8736 ( n8925, n8829, n8320 );
nor U8737 ( n8978, n8988, n8989 );
nor U8738 ( n8989, n8124, n8928 );
nand U8739 ( n8928, n8832, n8323 );
nor U8740 ( n8988, n8121, n8929 );
nand U8741 ( n8929, n8833, n8324 );
nor U8742 ( n8833, n8990, n8748 );
nand U8743 ( n580, n8991, n8992 );
nor U8744 ( n8992, n8993, n8994 );
nand U8745 ( n8994, n8995, n8996 );
nand U8746 ( n8996, n8131, n8997 );
nand U8747 ( n8995, n8998, n7990 );
nor U8748 ( n8993, n8135, n8999 );
nor U8749 ( n8991, n9000, n9001 );
nor U8750 ( n9001, n8139, n9002 );
nor U8751 ( n9000, n8141, n9003 );
nand U8752 ( n575, n9004, n9005 );
nor U8753 ( n9005, n9006, n9007 );
nand U8754 ( n9007, n9008, n9009 );
nand U8755 ( n9009, n8148, n8997 );
nand U8756 ( n9008, n8998, n7980 );
nor U8757 ( n9006, n8149, n8999 );
nor U8758 ( n9004, n9010, n9011 );
nor U8759 ( n9011, n8152, n9002 );
nor U8760 ( n9010, n8153, n9003 );
nand U8761 ( n570, n9012, n9013 );
nor U8762 ( n9013, n9014, n9015 );
nand U8763 ( n9015, n9016, n9017 );
nand U8764 ( n9017, n8160, n8997 );
nand U8765 ( n9016, n8998, n7970 );
nor U8766 ( n9014, n8161, n8999 );
nor U8767 ( n9012, n9018, n9019 );
nor U8768 ( n9019, n8164, n9002 );
nor U8769 ( n9018, n8165, n9003 );
nand U8770 ( n565, n9020, n9021 );
nor U8771 ( n9021, n9022, n9023 );
nand U8772 ( n9023, n9024, n9025 );
nand U8773 ( n9025, n8172, n8997 );
nand U8774 ( n9024, n8998, n7960 );
nor U8775 ( n9022, n8173, n8999 );
nor U8776 ( n9020, n9026, n9027 );
nor U8777 ( n9027, n8176, n9002 );
nor U8778 ( n9026, n8177, n9003 );
nand U8779 ( n560, n9028, n9029 );
nor U8780 ( n9029, n9030, n9031 );
nand U8781 ( n9031, n9032, n9033 );
nand U8782 ( n9033, n8184, n8997 );
nand U8783 ( n9032, n8998, n7950 );
nor U8784 ( n9030, n8185, n8999 );
nor U8785 ( n9028, n9034, n9035 );
nor U8786 ( n9035, n8188, n9002 );
nor U8787 ( n9034, n8189, n9003 );
nand U8788 ( n555, n9036, n9037 );
nor U8789 ( n9037, n9038, n9039 );
nand U8790 ( n9039, n9040, n9041 );
nand U8791 ( n9041, n8089, n8997 );
nand U8792 ( n9040, n8998, n7940 );
nor U8793 ( n9038, n8196, n8999 );
nor U8794 ( n9036, n9042, n9043 );
nor U8795 ( n9043, n8093, n9002 );
nor U8796 ( n9042, n8098, n9003 );
nand U8797 ( n550, n9044, n9045 );
nor U8798 ( n9045, n9046, n9047 );
nand U8799 ( n9047, n9048, n9049 );
nand U8800 ( n9049, n8106, n8997 );
nand U8801 ( n9048, n8998, n7930 );
nor U8802 ( n9046, n8205, n8999 );
nor U8803 ( n9044, n9050, n9051 );
nor U8804 ( n9051, n8108, n9002 );
nor U8805 ( n9050, n8111, n9003 );
nand U8806 ( n545, n9052, n9053 );
nor U8807 ( n9053, n9054, n9055 );
nand U8808 ( n9055, n9056, n9057 );
nand U8809 ( n9057, n8118, n8997 );
nand U8810 ( n8997, n9058, n9059 );
nand U8811 ( n9059, n9060, n7797 );
nand U8812 ( n9058, n9061, n8218 );
nand U8813 ( n9056, n8998, n8067 );
nand U8814 ( n8998, n9062, n9063 );
nor U8815 ( n9063, n9064, n9065 );
nor U8816 ( n9065, n15061, n9060 );
nand U8817 ( n9060, n8999, n9066 );
nand U8818 ( n9066, n8819, n8401 );
nor U8819 ( n8819, n9067, n8734 );
nor U8820 ( n9064, n9068, n9061 );
nand U8821 ( n9061, n8999, n9069 );
nand U8822 ( n9069, n8826, n8404 );
nor U8823 ( n8826, n8737, n9070 );
nor U8824 ( n9068, n9071, n8231 );
nor U8825 ( n9071, n8232, n9072 );
nand U8826 ( n9072, n9003, n9002 );
nor U8827 ( n9062, n9073, n8235 );
and U8828 ( n9073, n7815, n8999 );
nor U8829 ( n9054, n8119, n8999 );
nand U8830 ( n8999, n8829, n8742 );
nor U8831 ( n8829, n15198, n15199 );
nor U8832 ( n9052, n9074, n9075 );
nor U8833 ( n9075, n8124, n9002 );
nand U8834 ( n9002, n8832, n8745 );
nor U8835 ( n8832, n9076, n9077 );
nor U8836 ( n9074, n8121, n9003 );
nand U8837 ( n9003, n9078, n9079 );
nand U8838 ( n540, n9080, n9081 );
nor U8839 ( n9081, n9082, n9083 );
nand U8840 ( n9083, n9084, n9085 );
nor U8841 ( n9082, n9086, n9087 );
nor U8842 ( n9080, n9088, n9089 );
nand U8843 ( n9089, n9090, n9091 );
nand U8844 ( n9091, n9092, n7814 );
nand U8845 ( n9090, n9093, n15063 );
nor U8846 ( n9093, n9092, n9094 );
and U8847 ( n9094, n9095, n9096 );
and U8848 ( n9088, n9097, n9098 );
nand U8849 ( n535, n9099, n9100 );
nor U8850 ( n9100, n9101, n9102 );
nor U8851 ( n9102, n9103, n9104 );
nand U8852 ( n9104, n9105, n9106 );
nor U8853 ( n9099, n9107, n9108 );
nor U8854 ( n9108, n9092, n9109 );
not U8855 ( n9092, n9110 );
nor U8856 ( n9107, n15062, n9111 );
and U8857 ( n9111, n9084, n9110 );
nand U8858 ( n9084, n9112, READY_N );
nor U8859 ( n9112, n15063, n7797 );
nand U8860 ( n530, n9113, n9114 );
nor U8861 ( n9114, n9115, n9116 );
nor U8862 ( n9116, n7814, n9117 );
nand U8863 ( n9117, n7830, n7799 );
nor U8864 ( n9115, n15063, n9118 );
or U8865 ( n9118, n9119, READY_N );
nor U8866 ( n9113, n9120, n9121 );
nor U8867 ( n9121, n15061, n9122 );
nand U8868 ( n525, n9123, n9124 );
nand U8869 ( n9124, n9122, n9125 );
not U8870 ( n9122, n9103 );
nand U8871 ( n9123, n9103, n7815 );
nand U8872 ( n9103, n7814, n9110 );
nand U8873 ( n9110, n9126, n9127 );
nor U8874 ( n9127, n9128, n9129 );
nor U8875 ( n9129, n15063, n9130 );
nor U8876 ( n9130, n7799, n9097 );
nand U8877 ( n9097, n9131, n9132 );
nor U8878 ( n9132, n9133, n9134 );
nand U8879 ( n9134, n9135, n9136 );
nand U8880 ( n9135, n9137, n9138 );
nor U8881 ( n9137, n9139, n9140 );
nor U8882 ( n9133, n9141, n9142 );
nor U8883 ( n9141, n7813, n8048 );
nor U8884 ( n9131, n9143, n9144 );
nand U8885 ( n9144, n9145, n9146 );
nand U8886 ( n9146, n15197, n9147 );
nand U8887 ( n9147, n9148, n9149 );
nand U8888 ( n9149, n15198, n9150 );
or U8889 ( n9150, n9151, n9152 );
nand U8890 ( n9148, n9152, n9151 );
nand U8891 ( n9151, n9153, n9154 );
nand U8892 ( n9154, n15199, n9155 );
or U8893 ( n9155, n9156, n9157 );
nand U8894 ( n9153, n9157, n9156 );
nand U8895 ( n9156, n9158, n9159 );
nand U8896 ( n9159, n9160, n9161 );
nand U8897 ( n9160, n7825, n9162 );
nand U8898 ( n9158, n9163, n9164 );
nand U8899 ( n9163, n9162, n9165 );
nand U8900 ( n9162, n9166, n9167 );
nand U8901 ( n9145, n9168, n9169 );
nor U8902 ( n9128, n9170, n7814 );
nor U8903 ( n9170, n15062, n9106 );
nor U8904 ( n9126, n15061, n9171 );
nor U8905 ( n9171, n9172, n9173 );
nor U8906 ( n520, n15059, n9174 );
nor U8907 ( n515, n15058, n9174 );
nor U8908 ( n510, n15057, n9174 );
nor U8909 ( n505, n15056, n9174 );
nor U8910 ( n500, n15055, n9174 );
nor U8911 ( n495, n15054, n9174 );
nor U8912 ( n490, n15053, n9174 );
nor U8913 ( n485, n15052, n9174 );
nor U8914 ( n480, n15051, n9174 );
nor U8915 ( n475, n15050, n9174 );
nor U8916 ( n470, n15049, n9174 );
nor U8917 ( n465, n15048, n9174 );
nor U8918 ( n460, n15047, n9174 );
nor U8919 ( n455, n15046, n9174 );
nor U8920 ( n450, n15045, n9174 );
nor U8921 ( n445, n15044, n9174 );
nor U8922 ( n440, n15043, n9174 );
nor U8923 ( n435, n15042, n9174 );
nor U8924 ( n430, n15041, n9174 );
nor U8925 ( n425, n15040, n9174 );
nor U8926 ( n420, n15039, n9174 );
nor U8927 ( n415, n15038, n9174 );
nor U8928 ( n410, n15037, n9174 );
nor U8929 ( n405, n15036, n9174 );
nor U8930 ( n400, n15035, n9174 );
nor U8931 ( n395, n15034, n9174 );
nor U8932 ( n390, n15033, n9174 );
nor U8933 ( n385, n15032, n9174 );
nor U8934 ( n380, n15031, n9174 );
nor U8935 ( n375, n15030, n9174 );
nand U8936 ( n370, n9175, n9176 );
nand U8937 ( n9176, n9174, n9177 );
nand U8938 ( n9177, n9178, n9179 );
nand U8939 ( n9175, n9180, n7812 );
nand U8940 ( n365, n9181, n9182 );
nand U8941 ( n9182, n9180, n7874 );
nand U8942 ( n9181, n9183, n9174 );
nor U8943 ( n9183, BS16_N, n9184 );
nand U8944 ( n360, n9185, n9186 );
nor U8945 ( n9186, n9187, n9188 );
nor U8946 ( n9188, n15026, n9189 );
nand U8947 ( n9189, HOLD, n7805 );
nor U8948 ( n9187, n9190, n7802 );
nor U8949 ( n9190, n9191, n9192 );
nor U8950 ( n9191, n7805, n9193 );
nor U8951 ( n9185, n9194, n9195 );
nor U8952 ( n9195, n9196, n8016 );
nor U8953 ( n9194, n9197, n7819 );
nor U8954 ( n9197, n9198, n15027 );
nor U8955 ( n9198, n15026, n9106 );
nand U8956 ( n355, n9199, n9200 );
nor U8957 ( n9200, n9201, n9202 );
nor U8958 ( n9202, n15026, n9203 );
nand U8959 ( n9203, n9204, n9205 );
nand U8960 ( n9204, n9206, n9106 );
nand U8961 ( n9206, n9207, n9208 );
nand U8962 ( n9208, n15352, n9209 );
nor U8963 ( n9201, n9210, n7802 );
nor U8964 ( n9210, n9211, n9212 );
not U8965 ( n9212, n9205 );
nor U8966 ( n9211, n9192, n9213 );
nand U8967 ( n9213, n8016, n7805 );
not U8968 ( n9192, n9207 );
nand U8969 ( n9207, HOLD, n7819 );
nor U8970 ( n9199, n9214, n9215 );
nor U8971 ( n9215, n9106, n9216 );
not U8972 ( n9214, n9217 );
nand U8973 ( n350, n9218, n9219 );
nor U8974 ( n9219, n9220, n9221 );
nor U8975 ( n9221, n9106, n9222 );
nand U8976 ( n9222, n9223, n7802 );
nand U8977 ( n9223, n15025, n9224 );
nand U8978 ( n9224, n9225, n9193 );
nor U8979 ( n9225, n15027, n15352 );
not U8980 ( n9220, n9226 );
nor U8981 ( n9218, n9227, n9228 );
nor U8982 ( n9228, NA_N, n9205 );
nand U8983 ( n9205, n15027, n7819 );
nor U8984 ( n9227, n9209, n9229 );
nand U8985 ( n9229, n9230, n7805 );
nand U8986 ( n9230, n15025, n9231 );
nand U8987 ( n9231, n15352, n9232 );
nand U8988 ( n9232, n7802, n9233 );
nand U8989 ( n9233, READY_N, n9193 );
not U8990 ( n9193, NA_N );
not U8991 ( n9209, HOLD );
nand U8992 ( n346, n9234, n9235 );
nand U8993 ( n9235, n9216, ADDRESS_REG_0_ );
nor U8994 ( n9234, n9236, n9237 );
nor U8995 ( n9237, n15321, n9217 );
nor U8996 ( n9236, n15320, n9226 );
nand U8997 ( n342, n9238, n9239 );
nand U8998 ( n9239, n9216, ADDRESS_REG_1_ );
nor U8999 ( n9238, n9240, n9241 );
nor U9000 ( n9241, n15322, n9217 );
nor U9001 ( n9240, n15321, n9226 );
nand U9002 ( n338, n9242, n9243 );
nand U9003 ( n9243, n9216, ADDRESS_REG_2_ );
nor U9004 ( n9242, n9244, n9245 );
nor U9005 ( n9245, n15323, n9217 );
nor U9006 ( n9244, n15322, n9226 );
nand U9007 ( n334, n9246, n9247 );
nand U9008 ( n9247, n9216, ADDRESS_REG_3_ );
nor U9009 ( n9246, n9248, n9249 );
nor U9010 ( n9249, n15324, n9217 );
nor U9011 ( n9248, n15323, n9226 );
nand U9012 ( n330, n9250, n9251 );
nand U9013 ( n9251, n9216, ADDRESS_REG_4_ );
nor U9014 ( n9250, n9252, n9253 );
nor U9015 ( n9253, n15325, n9217 );
nor U9016 ( n9252, n15324, n9226 );
nand U9017 ( n326, n9254, n9255 );
nand U9018 ( n9255, n9216, ADDRESS_REG_5_ );
nor U9019 ( n9254, n9256, n9257 );
nor U9020 ( n9257, n15326, n9217 );
nor U9021 ( n9256, n15325, n9226 );
nand U9022 ( n322, n9258, n9259 );
nand U9023 ( n9259, n9216, ADDRESS_REG_6_ );
nor U9024 ( n9258, n9260, n9261 );
nor U9025 ( n9261, n15327, n9217 );
nor U9026 ( n9260, n15326, n9226 );
nand U9027 ( n318, n9262, n9263 );
nand U9028 ( n9263, n9216, ADDRESS_REG_7_ );
nor U9029 ( n9262, n9264, n9265 );
nor U9030 ( n9265, n15328, n9217 );
nor U9031 ( n9264, n15327, n9226 );
nand U9032 ( n314, n9266, n9267 );
nand U9033 ( n9267, n9216, ADDRESS_REG_8_ );
nor U9034 ( n9266, n9268, n9269 );
nor U9035 ( n9269, n15329, n9217 );
nor U9036 ( n9268, n15328, n9226 );
nand U9037 ( n310, n9270, n9271 );
nand U9038 ( n9271, n9216, ADDRESS_REG_9_ );
nor U9039 ( n9270, n9272, n9273 );
nor U9040 ( n9273, n15330, n9217 );
nor U9041 ( n9272, n15329, n9226 );
nand U9042 ( n306, n9274, n9275 );
nand U9043 ( n9275, n9216, ADDRESS_REG_10_ );
nor U9044 ( n9274, n9276, n9277 );
nor U9045 ( n9277, n15331, n9217 );
nor U9046 ( n9276, n15330, n9226 );
nand U9047 ( n302, n9278, n9279 );
nand U9048 ( n9279, n9216, ADDRESS_REG_11_ );
nor U9049 ( n9278, n9280, n9281 );
nor U9050 ( n9281, n15332, n9217 );
nor U9051 ( n9280, n15331, n9226 );
nand U9052 ( n298, n9282, n9283 );
nand U9053 ( n9283, n9216, ADDRESS_REG_12_ );
nor U9054 ( n9282, n9284, n9285 );
nor U9055 ( n9285, n15333, n9217 );
nor U9056 ( n9284, n15332, n9226 );
nand U9057 ( n294, n9286, n9287 );
nand U9058 ( n9287, n9216, ADDRESS_REG_13_ );
nor U9059 ( n9286, n9288, n9289 );
nor U9060 ( n9289, n15334, n9217 );
nor U9061 ( n9288, n15333, n9226 );
nand U9062 ( n290, n9290, n9291 );
nand U9063 ( n9291, n9216, ADDRESS_REG_14_ );
nor U9064 ( n9290, n9292, n9293 );
nor U9065 ( n9293, n15335, n9217 );
nor U9066 ( n9292, n15334, n9226 );
nand U9067 ( n286, n9294, n9295 );
nand U9068 ( n9295, n9216, ADDRESS_REG_15_ );
nor U9069 ( n9294, n9296, n9297 );
nor U9070 ( n9297, n15336, n9217 );
nor U9071 ( n9296, n15335, n9226 );
nand U9072 ( n282, n9298, n9299 );
nand U9073 ( n9299, n9216, ADDRESS_REG_16_ );
nor U9074 ( n9298, n9300, n9301 );
nor U9075 ( n9301, n15337, n9217 );
nor U9076 ( n9300, n15336, n9226 );
nand U9077 ( n278, n9302, n9303 );
nand U9078 ( n9303, n9216, ADDRESS_REG_17_ );
nor U9079 ( n9302, n9304, n9305 );
nor U9080 ( n9305, n15338, n9217 );
nor U9081 ( n9304, n15337, n9226 );
nand U9082 ( n274, n9306, n9307 );
nand U9083 ( n9307, n9216, ADDRESS_REG_18_ );
nor U9084 ( n9306, n9308, n9309 );
nor U9085 ( n9309, n15339, n9217 );
nor U9086 ( n9308, n15338, n9226 );
nand U9087 ( n270, n9310, n9311 );
nand U9088 ( n9311, n9216, ADDRESS_REG_19_ );
nor U9089 ( n9310, n9312, n9313 );
nor U9090 ( n9313, n15340, n9217 );
nor U9091 ( n9312, n15339, n9226 );
nand U9092 ( n266, n9314, n9315 );
nand U9093 ( n9315, n9216, ADDRESS_REG_20_ );
nor U9094 ( n9314, n9316, n9317 );
nor U9095 ( n9317, n15341, n9217 );
nor U9096 ( n9316, n15340, n9226 );
nand U9097 ( n262, n9318, n9319 );
nand U9098 ( n9319, n9216, ADDRESS_REG_21_ );
nor U9099 ( n9318, n9320, n9321 );
nor U9100 ( n9321, n15342, n9217 );
nor U9101 ( n9320, n15341, n9226 );
nand U9102 ( n258, n9322, n9323 );
nand U9103 ( n9323, n9216, ADDRESS_REG_22_ );
nor U9104 ( n9322, n9324, n9325 );
nor U9105 ( n9325, n15343, n9217 );
nor U9106 ( n9324, n15342, n9226 );
nand U9107 ( n254, n9326, n9327 );
nand U9108 ( n9327, n9216, ADDRESS_REG_23_ );
nor U9109 ( n9326, n9328, n9329 );
nor U9110 ( n9329, n15344, n9217 );
nor U9111 ( n9328, n15343, n9226 );
nand U9112 ( n250, n9330, n9331 );
nand U9113 ( n9331, n9216, ADDRESS_REG_24_ );
nor U9114 ( n9330, n9332, n9333 );
nor U9115 ( n9333, n15345, n9217 );
nor U9116 ( n9332, n15344, n9226 );
nand U9117 ( n246, n9334, n9335 );
nand U9118 ( n9335, n9216, ADDRESS_REG_25_ );
nor U9119 ( n9334, n9336, n9337 );
nor U9120 ( n9337, n15346, n9217 );
nor U9121 ( n9336, n15345, n9226 );
nand U9122 ( n242, n9338, n9339 );
nand U9123 ( n9339, n9216, ADDRESS_REG_26_ );
nor U9124 ( n9338, n9340, n9341 );
nor U9125 ( n9341, n15347, n9217 );
nor U9126 ( n9340, n15346, n9226 );
nand U9127 ( n2384, n9342, n9343 );
nand U9128 ( n9343, n9344, n8045 );
nand U9129 ( n9344, n9345, n9346 );
and U9130 ( n9346, n9347, n9348 );
nor U9131 ( n9345, n9349, n9350 );
and U9132 ( n9342, n9351, n9352 );
nand U9133 ( n238, n9353, n9354 );
nand U9134 ( n9354, n9216, ADDRESS_REG_27_ );
nor U9135 ( n9353, n9355, n9356 );
nor U9136 ( n9356, n15348, n9217 );
nor U9137 ( n9355, n15347, n9226 );
nand U9138 ( n2379, n9357, n9358 );
or U9139 ( n9358, n9359, n15008 );
nand U9140 ( n9357, n9360, n9361 );
nand U9141 ( n9361, n9362, n9363 );
nor U9142 ( n9362, n15061, n9364 );
or U9143 ( n9360, n9359, n9365 );
nand U9144 ( n2375, n9180, n9366 );
nand U9145 ( n9366, n7805, ADS_N_REG );
nand U9146 ( n2370, n9367, n9368 );
nand U9147 ( n9368, n9369, n8047 );
nand U9148 ( n9369, n9098, n9370 );
nand U9149 ( n9367, n9365, n7814 );
nand U9150 ( n2366, n9371, n9372 );
nand U9151 ( n9372, n9196, n8045 );
nand U9152 ( n9371, n9216, M_IO_N_REG );
nand U9153 ( n2362, n9373, n9374 );
nor U9154 ( n9373, n9375, n9376 );
nor U9155 ( n9376, n15007, n9196 );
nor U9156 ( n9375, n9216, n8047 );
nand U9157 ( n2357, n9377, n9378 );
or U9158 ( n9378, n9379, n15352 );
nand U9159 ( n9377, n9380, n9379 );
nand U9160 ( n9379, n9381, n9382 );
nor U9161 ( n9382, n9383, n9384 );
nor U9162 ( n9381, n9385, n9359 );
nor U9163 ( n9385, n9386, n9387 );
nand U9164 ( n9387, n15063, n9106 );
nand U9165 ( n9380, n9388, n9389 );
nand U9166 ( n9389, n9390, n7814 );
nand U9167 ( n9390, n9391, n9392 );
nand U9168 ( n9392, n9393, n9394 );
nand U9169 ( n9394, n9395, n7830 );
nor U9170 ( n9391, n15061, READY_N );
nor U9171 ( n9388, n9095, n9396 );
nor U9172 ( n9396, n9395, n9397 );
nand U9173 ( n2352, n9398, n9374 );
nand U9174 ( n9374, n9184, n15027 );
not U9175 ( n9184, n9179 );
nor U9176 ( n9398, n9399, n9400 );
nor U9177 ( n9400, n15351, n9174 );
nor U9178 ( n9399, n9180, n9178 );
not U9179 ( n9178, BS16_N );
not U9180 ( n9180, n9174 );
nand U9181 ( n9402, n9403, n7802 );
nor U9182 ( n9403, n15027, n7819 );
nand U9183 ( n9401, n15027, n15026 );
nand U9184 ( n2347, n9404, n9405 );
or U9185 ( n9405, n9136, n9406 );
nand U9186 ( n9136, n9407, n9408 );
nand U9187 ( n9408, n9409, n9410 );
nand U9188 ( n9410, n9411, n9349 );
nor U9189 ( n9409, n9412, n9413 );
nor U9190 ( n9413, n9414, n9415 );
nor U9191 ( n9414, n9416, n9417 );
nand U9192 ( n9417, n9418, n9419 );
nor U9193 ( n9416, n9420, n9421 );
nand U9194 ( n9421, n9138, n9422 );
nand U9195 ( n9420, n9423, n9424 );
nand U9196 ( n9423, n9140, n9425 );
nand U9197 ( n9425, n9426, n9427 );
nor U9198 ( n9412, n9428, n9429 );
nand U9199 ( n9404, n9406, n8048 );
nand U9200 ( n2342, n9430, n9431 );
nand U9201 ( n9431, n9406, n7813 );
nand U9202 ( n9406, n9098, n9142 );
nand U9203 ( n9142, n9370, n9432 );
nand U9204 ( n9432, n9433, n9106 );
nand U9205 ( n9433, n9434, n9435 );
and U9206 ( n9370, n9436, n9437 );
nor U9207 ( n9436, n9438, n9439 );
nor U9208 ( n9439, n9139, n9440 );
nor U9209 ( n9438, n9348, n9424 );
nand U9210 ( n234, n9441, n9442 );
nand U9211 ( n9442, n9216, ADDRESS_REG_28_ );
nor U9212 ( n9441, n9443, n9444 );
nor U9213 ( n9444, n15349, n9217 );
nor U9214 ( n9443, n15348, n9226 );
nand U9215 ( n2338, n9445, n9446 );
nand U9216 ( n9446, n15008, n9196 );
nand U9217 ( n9445, n9216, W_R_N_REG );
nand U9218 ( n2333, n9447, n9448 );
nor U9219 ( n9447, n9449, n9450 );
nor U9220 ( n9450, n15009, n9451 );
nor U9221 ( n9449, n15319, n9452 );
nand U9222 ( n2328, n9453, n9454 );
nand U9223 ( n9454, n9452, n8046 );
and U9224 ( n9453, n9455, n9448 );
not U9225 ( n9448, n9456 );
nand U9226 ( n2323, n9457, n9458 );
nand U9227 ( n9458, n9456, n7855 );
nor U9228 ( n9456, n9452, n15320 );
nor U9229 ( n9457, n9459, n9460 );
nor U9230 ( n9460, n9452, n9461 );
nand U9231 ( n9461, n9462, n15320 );
nor U9232 ( n9462, n9463, n7812 );
nor U9233 ( n9463, n15028, n15319 );
nor U9234 ( n9459, n15010, n9451 );
nand U9235 ( n2318, n9464, n9455 );
nand U9236 ( n9455, n9465, n9466 );
nor U9237 ( n9466, n9452, n7855 );
nor U9238 ( n9465, n7812, n7874 );
nor U9239 ( n9464, n9467, n9468 );
nor U9240 ( n9468, n9452, n9469 );
nand U9241 ( n9469, n15320, n15029 );
nor U9242 ( n9467, n15011, n9451 );
not U9243 ( n9451, n9452 );
nand U9244 ( n9452, n9470, n9471 );
nor U9245 ( n9471, n9472, n9473 );
nand U9246 ( n9473, n9474, n9475 );
nor U9247 ( n9475, n9476, n9477 );
nand U9248 ( n9477, n15049, n15050 );
nand U9249 ( n9476, n15051, n15052 );
nor U9250 ( n9474, n9478, n9479 );
nand U9251 ( n9479, n15045, n15046 );
nand U9252 ( n9478, n15047, n15048 );
nand U9253 ( n9472, n9480, n9481 );
nor U9254 ( n9481, n9482, n9483 );
nand U9255 ( n9483, n15057, n15058 );
nand U9256 ( n9482, n15059, n9484 );
nand U9257 ( n9484, n7812, n7874 );
nor U9258 ( n9480, n9485, n9486 );
nand U9259 ( n9486, n15053, n15054 );
nand U9260 ( n9485, n15055, n15056 );
nor U9261 ( n9470, n9487, n9488 );
nand U9262 ( n9488, n9489, n9490 );
nor U9263 ( n9490, n9491, n9492 );
nand U9264 ( n9492, n15033, n15034 );
nand U9265 ( n9491, n15035, n15036 );
nor U9266 ( n9489, n8081, n9493 );
nand U9267 ( n9493, n15031, n15032 );
nand U9268 ( n9487, n9494, n9495 );
nor U9269 ( n9495, n9496, n9497 );
nand U9270 ( n9497, n15041, n15042 );
nand U9271 ( n9496, n15043, n15044 );
nor U9272 ( n9494, n9498, n9499 );
nand U9273 ( n9499, n15037, n15038 );
nand U9274 ( n9498, n15039, n15040 );
nand U9275 ( n2313, n9500, n9501 );
nor U9276 ( n9501, n9502, n9503 );
nand U9277 ( n9503, n9504, n9505 );
nand U9278 ( n9505, n9506, n7852 );
nand U9279 ( n9504, n9507, n9508 );
nor U9280 ( n9502, n15020, n9509 );
nor U9281 ( n9500, n9510, n9511 );
nand U9282 ( n9511, n9512, n9513 );
nand U9283 ( n9513, n9514, n8070 );
nand U9284 ( n9514, n9515, n9516 );
nand U9285 ( n9516, n15349, n9517 );
nand U9286 ( n9512, n9518, n15350 );
nor U9287 ( n9518, n15349, n9519 );
and U9288 ( n9510, n9520, n9521 );
nand U9289 ( n2308, n9522, n9523 );
nor U9290 ( n9523, n9524, n9525 );
nand U9291 ( n9525, n9526, n9527 );
nand U9292 ( n9527, n9506, n8017 );
nand U9293 ( n9526, n9528, n9529 );
nor U9294 ( n9524, n9530, n9531 );
nor U9295 ( n9522, n9532, n9533 );
nand U9296 ( n9533, n9534, n9535 );
nand U9297 ( n9535, n9536, n7875 );
nand U9298 ( n9534, n9537, n9521 );
nand U9299 ( n9532, n9538, n9539 );
nand U9300 ( n9539, n15349, n9540 );
not U9301 ( n9540, n9519 );
nand U9302 ( n9519, n9541, n9517 );
nor U9303 ( n9541, n15348, n9542 );
or U9304 ( n9538, n9515, n15349 );
nor U9305 ( n9515, n9543, n9544 );
nor U9306 ( n9544, n7915, n9545 );
nand U9307 ( n2303, n9546, n9547 );
nor U9308 ( n9547, n9548, n9549 );
nand U9309 ( n9549, n9550, n9551 );
or U9310 ( n9551, n9552, n15255 );
nand U9311 ( n9550, n9528, n9553 );
nor U9312 ( n9548, n9530, n9554 );
nor U9313 ( n9546, n9555, n9556 );
nand U9314 ( n9556, n9557, n9558 );
nand U9315 ( n9558, n9536, n7876 );
nand U9316 ( n9557, n9559, n9521 );
nand U9317 ( n9555, n9560, n9561 );
nand U9318 ( n9561, n9543, n7915 );
nand U9319 ( n9543, n9562, n9563 );
nand U9320 ( n9563, n9517, n9542 );
nand U9321 ( n9560, n9564, n15348 );
nor U9322 ( n9564, n9542, n9545 );
nand U9323 ( n9542, n9565, n9566 );
nor U9324 ( n9566, n15345, n15346 );
nor U9325 ( n9565, n15347, n9567 );
nand U9326 ( n230, n9568, n9569 );
nand U9327 ( n9569, n9216, ADDRESS_REG_29_ );
nor U9328 ( n9568, n9570, n9571 );
nor U9329 ( n9571, n15350, n9217 );
nor U9330 ( n9570, n15349, n9226 );
nand U9331 ( n2298, n9572, n9573 );
nor U9332 ( n9573, n9574, n9575 );
nand U9333 ( n9575, n9576, n9577 );
nand U9334 ( n9577, n9506, n7847 );
nand U9335 ( n9576, n9528, n9578 );
nor U9336 ( n9574, n9530, n9579 );
nor U9337 ( n9572, n9580, n9581 );
nand U9338 ( n9581, n9582, n9583 );
nand U9339 ( n9583, n9536, n7877 );
nand U9340 ( n9582, n9584, n9521 );
nand U9341 ( n9580, n9585, n9586 );
nand U9342 ( n9586, n9587, n8050 );
nand U9343 ( n9587, n9588, n9589 );
nand U9344 ( n9589, n15346, n9517 );
nand U9345 ( n9585, n9590, n15347 );
nor U9346 ( n9590, n15346, n9591 );
nand U9347 ( n2293, n9592, n9593 );
nor U9348 ( n9593, n9594, n9595 );
nand U9349 ( n9595, n9596, n9597 );
nand U9350 ( n9597, n9506, n8018 );
nand U9351 ( n9596, n9528, n9598 );
nor U9352 ( n9594, n9530, n9599 );
nor U9353 ( n9592, n9600, n9601 );
nand U9354 ( n9601, n9602, n9603 );
nand U9355 ( n9603, n9536, n7878 );
nand U9356 ( n9602, n9604, n9521 );
nand U9357 ( n9600, n9605, n9606 );
nand U9358 ( n9606, n15346, n9607 );
not U9359 ( n9607, n9591 );
nand U9360 ( n9591, n9608, n9517 );
nor U9361 ( n9608, n15345, n9567 );
or U9362 ( n9605, n9588, n15346 );
nor U9363 ( n9588, n9609, n9610 );
nor U9364 ( n9610, n7907, n9545 );
nand U9365 ( n2288, n9611, n9612 );
nor U9366 ( n9612, n9613, n9614 );
nand U9367 ( n9614, n9615, n9616 );
nand U9368 ( n9616, n9506, n7861 );
nand U9369 ( n9615, n9528, n9617 );
nor U9370 ( n9613, n9530, n9618 );
nor U9371 ( n9611, n9619, n9620 );
nand U9372 ( n9620, n9621, n9622 );
nand U9373 ( n9622, n9536, n7879 );
nand U9374 ( n9621, n9623, n9521 );
nand U9375 ( n9619, n9624, n9625 );
nand U9376 ( n9625, n9609, n7907 );
nand U9377 ( n9609, n9562, n9626 );
nand U9378 ( n9626, n9517, n9567 );
nand U9379 ( n9624, n9627, n15345 );
nor U9380 ( n9627, n9567, n9545 );
nand U9381 ( n9567, n9628, n9629 );
nor U9382 ( n9629, n15342, n15343 );
nor U9383 ( n9628, n15344, n9630 );
nand U9384 ( n2283, n9631, n9632 );
nor U9385 ( n9632, n9633, n9634 );
nand U9386 ( n9634, n9635, n9636 );
nand U9387 ( n9636, n9506, n8019 );
nand U9388 ( n9635, n9528, n9637 );
nor U9389 ( n9633, n9530, n9638 );
nor U9390 ( n9631, n9639, n9640 );
nand U9391 ( n9640, n9641, n9642 );
nand U9392 ( n9642, n9536, n7880 );
nand U9393 ( n9641, n9643, n9521 );
nand U9394 ( n9639, n9644, n9645 );
nand U9395 ( n9645, n9646, n8051 );
nand U9396 ( n9646, n9647, n9648 );
nand U9397 ( n9648, n15343, n9517 );
nand U9398 ( n9644, n9649, n15344 );
nor U9399 ( n9649, n15343, n9650 );
nand U9400 ( n2278, n9651, n9652 );
nor U9401 ( n9652, n9653, n9654 );
nand U9402 ( n9654, n9655, n9656 );
nand U9403 ( n9656, n9506, n7848 );
nand U9404 ( n9655, n9528, n9657 );
nor U9405 ( n9653, n9530, n9658 );
nor U9406 ( n9651, n9659, n9660 );
nand U9407 ( n9660, n9661, n9662 );
nand U9408 ( n9662, n9536, n7881 );
nand U9409 ( n9661, n9663, n9521 );
nand U9410 ( n9659, n9664, n9665 );
nand U9411 ( n9665, n15343, n9666 );
not U9412 ( n9666, n9650 );
nand U9413 ( n9650, n9667, n9517 );
nor U9414 ( n9667, n15342, n9630 );
or U9415 ( n9664, n9647, n15343 );
nor U9416 ( n9647, n9668, n9669 );
nor U9417 ( n9669, n7908, n9545 );
nand U9418 ( n2273, n9670, n9671 );
nor U9419 ( n9671, n9672, n9673 );
nand U9420 ( n9673, n9674, n9675 );
nand U9421 ( n9675, n9506, n8020 );
nand U9422 ( n9674, n9528, n9676 );
nor U9423 ( n9672, n9530, n9677 );
nor U9424 ( n9670, n9678, n9679 );
nand U9425 ( n9679, n9680, n9681 );
nand U9426 ( n9681, n9536, n7882 );
nand U9427 ( n9680, n9682, n9521 );
nand U9428 ( n9678, n9683, n9684 );
nand U9429 ( n9684, n9668, n7908 );
nand U9430 ( n9668, n9562, n9685 );
nand U9431 ( n9685, n9517, n9630 );
nand U9432 ( n9683, n9686, n15342 );
nor U9433 ( n9686, n9630, n9545 );
nand U9434 ( n9630, n9687, n9688 );
nor U9435 ( n9688, n15339, n15340 );
nor U9436 ( n9687, n15341, n9689 );
nand U9437 ( n2268, n9690, n9691 );
nor U9438 ( n9691, n9692, n9693 );
nand U9439 ( n9693, n9694, n9695 );
nand U9440 ( n9695, n9506, n7921 );
nand U9441 ( n9694, n9528, n9696 );
nor U9442 ( n9692, n9530, n9697 );
nor U9443 ( n9690, n9698, n9699 );
nand U9444 ( n9699, n9700, n9701 );
nand U9445 ( n9701, n9536, n7883 );
nand U9446 ( n9700, n9702, n9521 );
nand U9447 ( n9698, n9703, n9704 );
nand U9448 ( n9704, n9705, n8052 );
nand U9449 ( n9705, n9706, n9707 );
nand U9450 ( n9707, n15340, n9517 );
nand U9451 ( n9703, n9708, n15341 );
nor U9452 ( n9708, n15340, n9709 );
nand U9453 ( n2263, n9710, n9711 );
nor U9454 ( n9711, n9712, n9713 );
nand U9455 ( n9713, n9714, n9715 );
or U9456 ( n9715, n9552, n15248 );
nand U9457 ( n9714, n9528, n9716 );
nor U9458 ( n9712, n9530, n9717 );
nor U9459 ( n9710, n9718, n9719 );
nand U9460 ( n9719, n9720, n9721 );
nand U9461 ( n9721, n9536, n7884 );
nand U9462 ( n9720, n9722, n9521 );
nand U9463 ( n9718, n9723, n9724 );
nand U9464 ( n9724, n15340, n9725 );
not U9465 ( n9725, n9709 );
nand U9466 ( n9709, n9726, n9517 );
nor U9467 ( n9726, n15339, n9689 );
or U9468 ( n9723, n9706, n15340 );
nor U9469 ( n9706, n9727, n9728 );
nor U9470 ( n9728, n7909, n9545 );
nand U9471 ( n226, n9729, n9730 );
or U9472 ( n9730, n9216, n15009 );
nand U9473 ( n9729, n9216, BE_N_REG_0_ );
nand U9474 ( n2258, n9731, n9732 );
nor U9475 ( n9732, n9733, n9734 );
nand U9476 ( n9734, n9735, n9736 );
nand U9477 ( n9736, n9506, n7849 );
nand U9478 ( n9735, n9528, n9737 );
nor U9479 ( n9733, n9530, n9738 );
nor U9480 ( n9731, n9739, n9740 );
nand U9481 ( n9740, n9741, n9742 );
nand U9482 ( n9742, n9536, n7885 );
nand U9483 ( n9741, n9743, n9521 );
nand U9484 ( n9739, n9744, n9745 );
nand U9485 ( n9745, n9727, n7909 );
nand U9486 ( n9727, n9562, n9746 );
nand U9487 ( n9746, n9517, n9689 );
nand U9488 ( n9744, n9747, n15339 );
nor U9489 ( n9747, n9689, n9545 );
nand U9490 ( n9689, n9748, n9749 );
nor U9491 ( n9749, n15336, n15337 );
nor U9492 ( n9748, n15338, n9750 );
nand U9493 ( n2253, n9751, n9752 );
nor U9494 ( n9752, n9753, n9754 );
nand U9495 ( n9754, n9755, n9756 );
nand U9496 ( n9756, n9528, n9757 );
or U9497 ( n9755, n9758, n9530 );
nand U9498 ( n9753, n9759, n9760 );
or U9499 ( n9759, n9552, n15246 );
nor U9500 ( n9751, n9761, n9762 );
nand U9501 ( n9762, n9763, n9764 );
nand U9502 ( n9764, n9536, n7886 );
nand U9503 ( n9763, n9765, n9521 );
nand U9504 ( n9761, n9766, n9767 );
nand U9505 ( n9767, n9768, n8053 );
nand U9506 ( n9768, n9769, n9770 );
nand U9507 ( n9770, n15337, n9517 );
nand U9508 ( n9766, n9771, n15338 );
nor U9509 ( n9771, n15337, n9772 );
nand U9510 ( n2248, n9773, n9774 );
nor U9511 ( n9774, n9775, n9776 );
nand U9512 ( n9776, n9777, n9778 );
nand U9513 ( n9778, n9528, n9779 );
or U9514 ( n9777, n9780, n9530 );
nand U9515 ( n9775, n9781, n9760 );
nand U9516 ( n9781, n9506, n8044 );
nor U9517 ( n9773, n9782, n9783 );
nand U9518 ( n9783, n9784, n9785 );
nand U9519 ( n9785, n9536, n7887 );
nand U9520 ( n9784, n9786, n9521 );
nand U9521 ( n9782, n9787, n9788 );
nand U9522 ( n9788, n15337, n9789 );
not U9523 ( n9789, n9772 );
nand U9524 ( n9772, n9790, n9517 );
nor U9525 ( n9790, n15336, n9750 );
or U9526 ( n9787, n9769, n15337 );
nor U9527 ( n9769, n9791, n9792 );
nor U9528 ( n9792, n7910, n9545 );
nand U9529 ( n2243, n9793, n9794 );
nor U9530 ( n9794, n9795, n9796 );
nand U9531 ( n9796, n9797, n9798 );
nand U9532 ( n9798, n9528, n9799 );
or U9533 ( n9797, n9800, n9530 );
nand U9534 ( n9795, n9801, n9760 );
or U9535 ( n9801, n9552, n15244 );
nor U9536 ( n9793, n9802, n9803 );
nand U9537 ( n9803, n9804, n9805 );
nand U9538 ( n9805, n9536, n7888 );
nand U9539 ( n9804, n9806, n9521 );
nand U9540 ( n9802, n9807, n9808 );
nand U9541 ( n9808, n9791, n7910 );
nand U9542 ( n9791, n9562, n9809 );
nand U9543 ( n9809, n9517, n9750 );
nand U9544 ( n9807, n9810, n15336 );
nor U9545 ( n9810, n9750, n9545 );
nand U9546 ( n9750, n9811, n9812 );
nor U9547 ( n9812, n15333, n15334 );
nor U9548 ( n9811, n15335, n9813 );
nand U9549 ( n2238, n9814, n9815 );
nor U9550 ( n9815, n9816, n9817 );
nand U9551 ( n9817, n9818, n9819 );
or U9552 ( n9819, n9820, n9821 );
or U9553 ( n9818, n9822, n9530 );
nand U9554 ( n9816, n9823, n9760 );
or U9555 ( n9823, n9552, n15243 );
nor U9556 ( n9814, n9824, n9825 );
nand U9557 ( n9825, n9826, n9827 );
nand U9558 ( n9827, n9536, n7889 );
nand U9559 ( n9826, n9828, n9521 );
nand U9560 ( n9824, n9829, n9830 );
nand U9561 ( n9830, n9831, n8054 );
nand U9562 ( n9831, n9832, n9833 );
nand U9563 ( n9833, n15334, n9517 );
nand U9564 ( n9829, n9834, n15335 );
nor U9565 ( n9834, n15334, n9835 );
nand U9566 ( n2233, n9836, n9837 );
nor U9567 ( n9837, n9838, n9839 );
nand U9568 ( n9839, n9840, n9841 );
nand U9569 ( n9841, n9528, n9842 );
or U9570 ( n9840, n9843, n9530 );
nand U9571 ( n9838, n9844, n9760 );
nand U9572 ( n9844, n9506, n8021 );
nor U9573 ( n9836, n9845, n9846 );
nand U9574 ( n9846, n9847, n9848 );
nand U9575 ( n9848, n9536, n7890 );
nand U9576 ( n9847, n9849, n9521 );
nand U9577 ( n9845, n9850, n9851 );
nand U9578 ( n9851, n15334, n9852 );
not U9579 ( n9852, n9835 );
nand U9580 ( n9835, n9853, n9517 );
nor U9581 ( n9853, n15333, n9813 );
or U9582 ( n9850, n9832, n15334 );
nor U9583 ( n9832, n9854, n9855 );
nor U9584 ( n9855, n7911, n9545 );
nand U9585 ( n2228, n9856, n9857 );
nor U9586 ( n9857, n9858, n9859 );
nand U9587 ( n9859, n9860, n9861 );
nand U9588 ( n9861, n9528, n9862 );
or U9589 ( n9860, n9863, n9530 );
nand U9590 ( n9858, n9864, n9760 );
nand U9591 ( n9864, n9506, n7836 );
nor U9592 ( n9856, n9865, n9866 );
nand U9593 ( n9866, n9867, n9868 );
nand U9594 ( n9868, n9536, n7891 );
nand U9595 ( n9867, n9521, n9869 );
nand U9596 ( n9865, n9870, n9871 );
nand U9597 ( n9871, n9854, n7911 );
nand U9598 ( n9854, n9562, n9872 );
nand U9599 ( n9872, n9517, n9813 );
nand U9600 ( n9870, n9873, n15333 );
nor U9601 ( n9873, n9813, n9545 );
nand U9602 ( n9813, n9874, n9875 );
nor U9603 ( n9875, n15330, n15331 );
nor U9604 ( n9874, n15332, n9876 );
nand U9605 ( n2223, n9877, n9878 );
nor U9606 ( n9878, n9879, n9880 );
nand U9607 ( n9880, n9881, n9882 );
nand U9608 ( n9882, n9528, n9883 );
or U9609 ( n9881, n9884, n9530 );
nand U9610 ( n9879, n9885, n9760 );
nand U9611 ( n9885, n9506, n7809 );
nor U9612 ( n9877, n9886, n9887 );
nand U9613 ( n9887, n9888, n9889 );
nand U9614 ( n9889, n9536, n7892 );
nand U9615 ( n9888, n9890, n9521 );
nand U9616 ( n9886, n9891, n9892 );
nand U9617 ( n9892, n9893, n8055 );
nand U9618 ( n9893, n9894, n9895 );
nand U9619 ( n9895, n15331, n9517 );
nand U9620 ( n9891, n9896, n15332 );
nor U9621 ( n9896, n15331, n9897 );
nand U9622 ( n222, n9898, n9899 );
nand U9623 ( n9899, n9196, n8046 );
not U9624 ( n9196, n9216 );
nand U9625 ( n9898, n9216, BE_N_REG_1_ );
nand U9626 ( n2218, n9900, n9901 );
nor U9627 ( n9901, n9902, n9903 );
nand U9628 ( n9903, n9904, n9905 );
nand U9629 ( n9905, n9528, n9906 );
or U9630 ( n9904, n9907, n9530 );
nand U9631 ( n9902, n9908, n9760 );
nand U9632 ( n9908, n9506, n7863 );
nor U9633 ( n9900, n9909, n9910 );
nand U9634 ( n9910, n9911, n9912 );
nand U9635 ( n9912, n9536, n7893 );
nand U9636 ( n9911, n9913, n9521 );
nand U9637 ( n9909, n9914, n9915 );
nand U9638 ( n9915, n15331, n9916 );
not U9639 ( n9916, n9897 );
nand U9640 ( n9897, n9917, n9517 );
nor U9641 ( n9917, n15330, n9876 );
or U9642 ( n9914, n9894, n15331 );
nor U9643 ( n9894, n9918, n9919 );
nor U9644 ( n9919, n7912, n9545 );
nand U9645 ( n2213, n9920, n9921 );
nor U9646 ( n9921, n9922, n9923 );
nand U9647 ( n9923, n9924, n9925 );
nand U9648 ( n9925, n9528, n9926 );
or U9649 ( n9924, n9927, n9530 );
nand U9650 ( n9922, n9928, n9760 );
nand U9651 ( n9928, n9506, n8014 );
nor U9652 ( n9920, n9929, n9930 );
nand U9653 ( n9930, n9931, n9932 );
nand U9654 ( n9932, n9536, n7894 );
nand U9655 ( n9931, n9933, n9521 );
nand U9656 ( n9929, n9934, n9935 );
nand U9657 ( n9935, n9918, n7912 );
nand U9658 ( n9918, n9562, n9936 );
nand U9659 ( n9936, n9517, n9876 );
nand U9660 ( n9934, n9937, n15330 );
nor U9661 ( n9937, n9876, n9545 );
nand U9662 ( n9876, n9938, n9939 );
nor U9663 ( n9939, n15327, n15328 );
nor U9664 ( n9938, n15329, n9940 );
nand U9665 ( n2208, n9941, n9942 );
nor U9666 ( n9942, n9943, n9944 );
nand U9667 ( n9944, n9945, n9946 );
nand U9668 ( n9946, n9528, n9947 );
or U9669 ( n9945, n9948, n9530 );
nand U9670 ( n9943, n9949, n9760 );
nand U9671 ( n9949, n9506, n7837 );
nor U9672 ( n9941, n9950, n9951 );
nand U9673 ( n9951, n9952, n9953 );
nand U9674 ( n9953, n9536, n7895 );
nand U9675 ( n9952, n9954, n9521 );
nand U9676 ( n9950, n9955, n9956 );
nand U9677 ( n9956, n9957, n8056 );
nand U9678 ( n9957, n9958, n9959 );
nand U9679 ( n9959, n15328, n9517 );
nand U9680 ( n9955, n9960, n15329 );
nor U9681 ( n9960, n15328, n9961 );
nand U9682 ( n2203, n9962, n9963 );
nor U9683 ( n9963, n9964, n9965 );
nand U9684 ( n9965, n9966, n9967 );
nand U9685 ( n9967, n9528, n9968 );
or U9686 ( n9966, n9969, n9530 );
nand U9687 ( n9964, n9970, n9760 );
nand U9688 ( n9970, n9506, n7810 );
nor U9689 ( n9962, n9971, n9972 );
nand U9690 ( n9972, n9973, n9974 );
nand U9691 ( n9974, n9536, n7896 );
nand U9692 ( n9973, n9975, n9521 );
nand U9693 ( n9971, n9976, n9977 );
nand U9694 ( n9977, n15328, n9978 );
not U9695 ( n9978, n9961 );
nand U9696 ( n9961, n9979, n9517 );
nor U9697 ( n9979, n15327, n9940 );
or U9698 ( n9976, n9958, n15328 );
nor U9699 ( n9958, n9980, n9981 );
nor U9700 ( n9981, n7913, n9545 );
nand U9701 ( n2198, n9982, n9983 );
nor U9702 ( n9983, n9984, n9985 );
nand U9703 ( n9985, n9986, n9987 );
nand U9704 ( n9987, n9528, n9988 );
or U9705 ( n9986, n9989, n9530 );
nand U9706 ( n9984, n9990, n9760 );
nand U9707 ( n9990, n9506, n7864 );
nor U9708 ( n9982, n9991, n9992 );
nand U9709 ( n9992, n9993, n9994 );
nand U9710 ( n9994, n9536, n7897 );
nand U9711 ( n9993, n9995, n9521 );
nand U9712 ( n9991, n9996, n9997 );
nand U9713 ( n9997, n9980, n7913 );
nand U9714 ( n9980, n9562, n9998 );
nand U9715 ( n9998, n9517, n9940 );
nand U9716 ( n9996, n9999, n15327 );
nor U9717 ( n9999, n9940, n9545 );
nand U9718 ( n9940, n10000, n10001 );
nor U9719 ( n10001, n15324, n15325 );
nor U9720 ( n10000, n15326, n10002 );
nand U9721 ( n2193, n10003, n10004 );
nor U9722 ( n10004, n10005, n10006 );
nand U9723 ( n10006, n10007, n10008 );
nand U9724 ( n10008, n9528, n10009 );
or U9725 ( n10007, n10010, n9530 );
nand U9726 ( n10005, n10011, n9760 );
nand U9727 ( n10011, n9506, n8015 );
nor U9728 ( n10003, n10012, n10013 );
nand U9729 ( n10013, n10014, n10015 );
nand U9730 ( n10015, n9536, n7898 );
nand U9731 ( n10014, n10016, n9521 );
nand U9732 ( n10012, n10017, n10018 );
nand U9733 ( n10018, n10019, n8057 );
nand U9734 ( n10019, n10020, n10021 );
nand U9735 ( n10021, n15325, n9517 );
nand U9736 ( n10017, n10022, n15326 );
nor U9737 ( n10022, n15325, n10023 );
nand U9738 ( n2188, n10024, n10025 );
nor U9739 ( n10025, n10026, n10027 );
nand U9740 ( n10027, n10028, n10029 );
nand U9741 ( n10029, n9528, n10030 );
or U9742 ( n10028, n10031, n9530 );
nand U9743 ( n10026, n10032, n9760 );
nand U9744 ( n10032, n9506, n7838 );
nor U9745 ( n10024, n10033, n10034 );
nand U9746 ( n10034, n10035, n10036 );
nand U9747 ( n10036, n9536, n7899 );
nand U9748 ( n10035, n10037, n9521 );
not U9749 ( n9521, n10038 );
nand U9750 ( n10033, n10039, n10040 );
nand U9751 ( n10040, n15325, n10041 );
not U9752 ( n10041, n10023 );
nand U9753 ( n10023, n10042, n9517 );
nor U9754 ( n10042, n15324, n10002 );
or U9755 ( n10039, n10020, n15325 );
nor U9756 ( n10020, n10043, n10044 );
nor U9757 ( n10044, n7914, n9545 );
nand U9758 ( n2183, n10045, n10046 );
nor U9759 ( n10046, n10047, n10048 );
nand U9760 ( n10048, n10049, n10050 );
nand U9761 ( n10050, n9528, n10051 );
or U9762 ( n10049, n10052, n9530 );
nand U9763 ( n10047, n10053, n9760 );
nand U9764 ( n10053, n9506, n7811 );
nor U9765 ( n10045, n10054, n10055 );
nand U9766 ( n10055, n10056, n10057 );
nand U9767 ( n10057, n9536, n7900 );
nand U9768 ( n10056, n10058, n10059 );
nand U9769 ( n10054, n10060, n10061 );
nand U9770 ( n10061, n10043, n7914 );
nand U9771 ( n10043, n9562, n10062 );
nand U9772 ( n10062, n9517, n10002 );
nand U9773 ( n10060, n10063, n15324 );
nor U9774 ( n10063, n10002, n9545 );
nand U9775 ( n10002, n10064, n10065 );
nor U9776 ( n10064, n15322, n15323 );
nand U9777 ( n218, n10066, n10067 );
or U9778 ( n10067, n9216, n15010 );
nand U9779 ( n10066, n9216, BE_N_REG_2_ );
nand U9780 ( n2178, n10068, n10069 );
nor U9781 ( n10069, n10070, n10071 );
nand U9782 ( n10071, n10072, n10073 );
nand U9783 ( n10073, n9528, n10074 );
or U9784 ( n10072, n10075, n9530 );
nand U9785 ( n10070, n10076, n9760 );
nand U9786 ( n9760, n9365, n9562 );
not U9787 ( n9365, n9351 );
nand U9788 ( n9351, n9383, n15062 );
nand U9789 ( n10076, n9506, n7923 );
nor U9790 ( n10068, n10077, n10078 );
nand U9791 ( n10078, n10079, n10080 );
nand U9792 ( n10080, n10081, n10059 );
nor U9793 ( n10079, n10082, n10083 );
nor U9794 ( n10083, n8049, n10084 );
nand U9795 ( n10084, n10085, n7846 );
nor U9796 ( n10082, n15323, n10086 );
nor U9797 ( n10086, n10087, n10088 );
nor U9798 ( n10087, n9545, n7846 );
nand U9799 ( n10077, n10089, n10090 );
nand U9800 ( n10090, n9536, n7901 );
nand U9801 ( n10089, n10091, n10092 );
nand U9802 ( n2173, n10093, n10094 );
nor U9803 ( n10094, n10095, n10096 );
nand U9804 ( n10096, n10097, n10098 );
or U9805 ( n10098, n10099, n9530 );
nand U9806 ( n10097, n9536, n7902 );
nand U9807 ( n10095, n10100, n10101 );
nand U9808 ( n10101, n9506, n7851 );
nand U9809 ( n10100, n9528, n10102 );
nor U9810 ( n10093, n10103, n10104 );
nand U9811 ( n10104, n10105, n10106 );
nand U9812 ( n10106, n10091, n10107 );
nand U9813 ( n10105, n10108, n10059 );
nand U9814 ( n10103, n10109, n10110 );
nand U9815 ( n10110, n15322, n10085 );
and U9816 ( n10085, n10065, n9517 );
nor U9817 ( n10065, n15320, n15321 );
nand U9818 ( n10109, n10088, n7846 );
nand U9819 ( n10088, n10111, n10112 );
nand U9820 ( n10112, n15321, n9517 );
nand U9821 ( n2168, n10113, n10114 );
nor U9822 ( n10114, n10115, n10116 );
nand U9823 ( n10116, n10117, n10118 );
nand U9824 ( n10118, n10119, n9507 );
not U9825 ( n9507, n9530 );
nand U9826 ( n10117, n9536, n7903 );
nand U9827 ( n10115, n10120, n10121 );
or U9828 ( n10121, n9552, n15233 );
nand U9829 ( n10120, n9528, n10122 );
nor U9830 ( n10113, n10123, n10124 );
nand U9831 ( n10124, n10125, n10126 );
nand U9832 ( n10126, n10091, n8738 );
nand U9833 ( n10125, n10127, n10059 );
nand U9834 ( n10123, n10128, n10129 );
or U9835 ( n10129, n10111, n15321 );
and U9836 ( n10111, n9562, n10130 );
nand U9837 ( n10130, n9517, n15320 );
nand U9838 ( n10128, n10131, n15321 );
nor U9839 ( n10131, n15320, n9545 );
nand U9840 ( n2163, n10132, n10133 );
nor U9841 ( n10133, n10134, n10135 );
nand U9842 ( n10135, n10136, n10137 );
or U9843 ( n10137, n10138, n9530 );
nand U9844 ( n10136, n9536, n7904 );
nor U9845 ( n10134, n8490, n10139 );
nor U9846 ( n10132, n10140, n10141 );
nand U9847 ( n10141, n10142, n10143 );
or U9848 ( n10143, n10144, n10145 );
nor U9849 ( n10142, n10146, n10147 );
and U9850 ( n10147, n15320, n9517 );
nor U9851 ( n10146, n15320, n9562 );
nand U9852 ( n10140, n10148, n10149 );
nand U9853 ( n10149, n9506, n7850 );
not U9854 ( n9506, n9552 );
nand U9855 ( n10148, n15232, n9528 );
nand U9856 ( n2158, n10150, n10151 );
nor U9857 ( n10151, n10152, n10153 );
nand U9858 ( n10153, n10154, n10155 );
nand U9859 ( n10155, n10156, n7855 );
nand U9860 ( n10156, n9562, n9545 );
nand U9861 ( n9545, n10157, n10158 );
nor U9862 ( n10158, n9434, n10159 );
nor U9863 ( n10159, n9393, n10160 );
and U9864 ( n10157, n10161, n10162 );
nand U9865 ( n10154, n10163, n8043 );
nand U9866 ( n10163, n9820, n9552 );
nand U9867 ( n9552, n7815, n9562 );
not U9868 ( n9820, n9528 );
nand U9869 ( n10164, n7799, n9562 );
nor U9870 ( n10152, n10166, n9530 );
nor U9871 ( n10168, n15020, n10161 );
and U9872 ( n10167, n10160, n10162 );
nor U9873 ( n10150, n10169, n10170 );
nand U9874 ( n10170, n10171, n10172 );
nand U9875 ( n10172, n9536, n7905 );
nand U9876 ( n9509, n10162, n10173 );
nand U9877 ( n10173, n10174, n10175 );
nand U9878 ( n10175, n10176, n15020 );
nor U9879 ( n10176, n10161, n10177 );
nand U9880 ( n10174, n9393, n9172 );
nand U9881 ( n9172, n10161, n9395 );
nor U9882 ( n10161, n7830, READY_N );
nand U9883 ( n10171, n10091, n10178 );
not U9884 ( n10091, n10139 );
nand U9885 ( n10139, n10179, n10162 );
nor U9886 ( n10169, n10145, n10180 );
not U9887 ( n10145, n10059 );
nand U9888 ( n10059, n10038, n10181 );
nand U9889 ( n10181, n10162, n9364 );
nor U9890 ( n10162, n10182, n15061 );
nand U9891 ( n10038, n10183, n10165 );
nor U9892 ( n10183, n15062, n10182 );
not U9893 ( n10182, n9562 );
nand U9894 ( n9562, n10184, n10185 );
nor U9895 ( n10185, n10186, n9101 );
and U9896 ( n9101, n10187, n10188 );
nor U9897 ( n10187, n15062, n7814 );
not U9898 ( n10186, n9085 );
nand U9899 ( n9085, n10189, n9095 );
nor U9900 ( n10189, n15060, n15063 );
nor U9901 ( n10184, n10190, n9359 );
nand U9902 ( n9359, n10191, n10192 );
nand U9903 ( n10192, n9120, n10193 );
nand U9904 ( n10193, n9352, n10194 );
nand U9905 ( n10194, n10195, n9437 );
not U9906 ( n9437, n9349 );
nand U9907 ( n9352, n10196, n10197 );
nor U9908 ( n10196, n9139, n10198 );
nand U9909 ( n10191, n10197, n10199 );
nand U9910 ( n2153, n10200, n10201 );
nand U9911 ( n10201, n10202, n9508 );
nand U9912 ( n10200, n10203, n8022 );
nand U9913 ( n2148, n10204, n10205 );
nand U9914 ( n10205, n10203, n7875 );
nor U9915 ( n10204, n10206, n10207 );
nor U9916 ( n10207, n10208, n10209 );
nor U9917 ( n10206, n9531, n10210 );
nand U9918 ( n2143, n10211, n10212 );
nand U9919 ( n10212, n10203, n7876 );
nor U9920 ( n10211, n10213, n10214 );
nor U9921 ( n10214, n10215, n10209 );
nor U9922 ( n10213, n9554, n10210 );
nand U9923 ( n214, n10216, n10217 );
or U9924 ( n10217, n9216, n15011 );
nand U9925 ( n10216, n9216, BE_N_REG_3_ );
nand U9926 ( n2138, n10218, n10219 );
nand U9927 ( n10219, n10203, n7877 );
nor U9928 ( n10218, n10220, n10221 );
nor U9929 ( n10221, n10222, n10209 );
nor U9930 ( n10220, n9579, n10210 );
nand U9931 ( n2133, n10223, n10224 );
nand U9932 ( n10224, n10203, n7878 );
nor U9933 ( n10223, n10225, n10226 );
nor U9934 ( n10226, n10227, n10209 );
nor U9935 ( n10225, n9599, n10210 );
nand U9936 ( n2128, n10228, n10229 );
nand U9937 ( n10229, n10203, n7879 );
nor U9938 ( n10228, n10230, n10231 );
nor U9939 ( n10231, n10232, n10209 );
nor U9940 ( n10230, n9618, n10210 );
nand U9941 ( n2123, n10233, n10234 );
nand U9942 ( n10234, n10203, n7880 );
nor U9943 ( n10233, n10235, n10236 );
nor U9944 ( n10236, n10237, n10209 );
nor U9945 ( n10235, n9638, n10210 );
nand U9946 ( n2118, n10238, n10239 );
nand U9947 ( n10239, n10203, n7881 );
nor U9948 ( n10238, n10240, n10241 );
nor U9949 ( n10241, n10242, n10209 );
nor U9950 ( n10240, n9658, n10210 );
nand U9951 ( n2113, n10243, n10244 );
nand U9952 ( n10244, n10203, n7882 );
nor U9953 ( n10243, n10245, n10246 );
nor U9954 ( n10246, n10247, n10209 );
nor U9955 ( n10245, n9677, n10210 );
nand U9956 ( n2108, n10248, n10249 );
nand U9957 ( n10249, n10203, n7883 );
nor U9958 ( n10248, n10250, n10251 );
nor U9959 ( n10251, n10252, n10209 );
nor U9960 ( n10250, n9697, n10210 );
nand U9961 ( n2103, n10253, n10254 );
nand U9962 ( n10254, n10203, n7884 );
nor U9963 ( n10253, n10255, n10256 );
nor U9964 ( n10256, n10257, n10209 );
nor U9965 ( n10255, n9717, n10210 );
nand U9966 ( n2098, n10258, n10259 );
nand U9967 ( n10259, n10203, n7885 );
nor U9968 ( n10258, n10260, n10261 );
nor U9969 ( n10261, n10262, n10209 );
nor U9970 ( n10260, n9738, n10210 );
nand U9971 ( n2093, n10263, n10264 );
nand U9972 ( n10264, n10203, n7886 );
nor U9973 ( n10263, n10265, n10266 );
nor U9974 ( n10266, n10267, n10209 );
nor U9975 ( n10265, n9758, n10210 );
nand U9976 ( n2088, n10268, n10269 );
nand U9977 ( n10269, n10203, n7887 );
nor U9978 ( n10268, n10270, n10271 );
nor U9979 ( n10271, n10272, n10209 );
nor U9980 ( n10270, n9780, n10210 );
nand U9981 ( n2083, n10273, n10274 );
nand U9982 ( n10274, n10203, n7888 );
nor U9983 ( n10273, n10275, n10276 );
nor U9984 ( n10276, n10277, n10209 );
nor U9985 ( n10275, n9800, n10210 );
nand U9986 ( n2078, n10278, n10279 );
nand U9987 ( n10279, n10203, n7889 );
nor U9988 ( n10278, n10280, n10281 );
nor U9989 ( n10281, n10282, n10209 );
nor U9990 ( n10280, n9822, n10210 );
nand U9991 ( n2073, n10283, n10284 );
nand U9992 ( n10284, n10203, n7890 );
nor U9993 ( n10283, n10285, n10286 );
nor U9994 ( n10286, n10287, n10209 );
nor U9995 ( n10285, n9843, n10210 );
nand U9996 ( n2068, n10288, n10289 );
nand U9997 ( n10289, n10203, n7891 );
nor U9998 ( n10288, n10290, n10291 );
nor U9999 ( n10291, n10292, n10209 );
nor U10000 ( n10290, n9863, n10210 );
nand U10001 ( n2063, n10293, n10294 );
nand U10002 ( n10294, n10203, n7892 );
nor U10003 ( n10293, n10295, n10296 );
nor U10004 ( n10296, n10297, n10209 );
nor U10005 ( n10295, n9884, n10210 );
nand U10006 ( n2058, n10298, n10299 );
nand U10007 ( n10299, n10203, n7893 );
nor U10008 ( n10298, n10300, n10301 );
nor U10009 ( n10301, n10302, n10209 );
nor U10010 ( n10300, n9907, n10210 );
nand U10011 ( n2053, n10303, n10304 );
nand U10012 ( n10304, n10203, n7894 );
nor U10013 ( n10303, n10305, n10306 );
nor U10014 ( n10306, n10307, n10209 );
nor U10015 ( n10305, n9927, n10210 );
nand U10016 ( n2048, n10308, n10309 );
nand U10017 ( n10309, n10203, n7895 );
nor U10018 ( n10308, n10310, n10311 );
nor U10019 ( n10311, n10312, n10209 );
nor U10020 ( n10310, n9948, n10210 );
nand U10021 ( n2043, n10313, n10314 );
nand U10022 ( n10314, n10203, n7896 );
nor U10023 ( n10313, n10315, n10316 );
nor U10024 ( n10316, n10317, n10209 );
nor U10025 ( n10315, n9969, n10210 );
nand U10026 ( n2038, n10318, n10319 );
nand U10027 ( n10319, n10203, n7897 );
nor U10028 ( n10318, n10320, n10321 );
nor U10029 ( n10321, n10322, n10209 );
nor U10030 ( n10320, n9989, n10210 );
nand U10031 ( n2033, n10323, n10324 );
nand U10032 ( n10324, n10203, n7898 );
nor U10033 ( n10323, n10325, n10326 );
nor U10034 ( n10326, n10327, n10209 );
nor U10035 ( n10325, n10010, n10210 );
nand U10036 ( n2028, n10328, n10329 );
nand U10037 ( n10329, n10203, n7899 );
nor U10038 ( n10328, n10330, n10331 );
nor U10039 ( n10331, n10332, n10209 );
nor U10040 ( n10330, n10031, n10210 );
nand U10041 ( n2023, n10333, n10334 );
nand U10042 ( n10334, n10203, n7900 );
nor U10043 ( n10333, n10335, n10336 );
nor U10044 ( n10336, n10337, n10209 );
nor U10045 ( n10335, n10052, n10210 );
nand U10046 ( n2018, n10338, n10339 );
nand U10047 ( n10339, n10203, n7901 );
nor U10048 ( n10338, n10340, n10341 );
nor U10049 ( n10341, n10342, n10209 );
nor U10050 ( n10340, n10075, n10210 );
nand U10051 ( n2013, n10343, n10344 );
nand U10052 ( n10344, n10203, n7902 );
nor U10053 ( n10343, n10345, n10346 );
nor U10054 ( n10346, n10347, n10209 );
nor U10055 ( n10345, n10099, n10210 );
nand U10056 ( n2008, n10348, n10349 );
nand U10057 ( n10349, n10203, n7903 );
nor U10058 ( n10348, n10350, n10351 );
nor U10059 ( n10351, n10352, n10209 );
and U10060 ( n10350, n10119, n10202 );
nand U10061 ( n2003, n10353, n10354 );
nand U10062 ( n10354, n10203, n7904 );
nor U10063 ( n10353, n10355, n10356 );
nor U10064 ( n10356, n10144, n10209 );
nor U10065 ( n10355, n10138, n10210 );
nand U10066 ( n1998, n10357, n10358 );
nand U10067 ( n10358, n10203, n7905 );
nor U10068 ( n10357, n10359, n10360 );
nor U10069 ( n10360, n10180, n10209 );
nor U10070 ( n10359, n10166, n10210 );
nor U10071 ( n10202, n10203, n9407 );
nand U10072 ( n10362, n10363, n10364 );
nand U10073 ( n10364, n10365, n10366 );
and U10074 ( n10365, n10160, n10367 );
nand U10075 ( n1993, n10368, n10369 );
nand U10076 ( n10369, n10370, DATAI_31_ );
nor U10077 ( n10368, n10371, n10372 );
nor U10078 ( n10372, n10373, n10374 );
nand U10079 ( n10374, n10361, n9520 );
nor U10080 ( n10371, n15013, n10375 );
nand U10081 ( n1988, n10376, n10377 );
nor U10082 ( n10377, n10378, n10379 );
and U10083 ( n10379, DATAI_30_, n10370 );
nor U10084 ( n10378, n10380, n10381 );
nor U10085 ( n10376, n10382, n10383 );
nor U10086 ( n10383, n15318, n10375 );
nor U10087 ( n10382, n10208, n10384 );
not U10088 ( n10208, n9537 );
nand U10089 ( n1983, n10385, n10386 );
nor U10090 ( n10386, n10387, n10388 );
and U10091 ( n10388, DATAI_29_, n10370 );
nor U10092 ( n10387, n10380, n10389 );
nor U10093 ( n10385, n10390, n10391 );
nor U10094 ( n10391, n15317, n10375 );
nor U10095 ( n10390, n10215, n10384 );
not U10096 ( n10215, n9559 );
nand U10097 ( n1978, n10392, n10393 );
nor U10098 ( n10393, n10394, n10395 );
and U10099 ( n10395, DATAI_28_, n10370 );
nor U10100 ( n10394, n10380, n10396 );
nor U10101 ( n10392, n10397, n10398 );
nor U10102 ( n10398, n15316, n10375 );
nor U10103 ( n10397, n10222, n10384 );
not U10104 ( n10222, n9584 );
nand U10105 ( n1973, n10399, n10400 );
nor U10106 ( n10400, n10401, n10402 );
and U10107 ( n10402, DATAI_27_, n10370 );
nor U10108 ( n10401, n10380, n10403 );
nor U10109 ( n10399, n10404, n10405 );
nor U10110 ( n10405, n15315, n10375 );
nor U10111 ( n10404, n10227, n10384 );
not U10112 ( n10227, n9604 );
nand U10113 ( n1968, n10406, n10407 );
nor U10114 ( n10407, n10408, n10409 );
and U10115 ( n10409, DATAI_26_, n10370 );
nor U10116 ( n10408, n10380, n10410 );
nor U10117 ( n10406, n10411, n10412 );
nor U10118 ( n10412, n15314, n10375 );
nor U10119 ( n10411, n10232, n10384 );
not U10120 ( n10232, n9623 );
nand U10121 ( n1963, n10413, n10414 );
nor U10122 ( n10414, n10415, n10416 );
and U10123 ( n10416, DATAI_25_, n10370 );
nor U10124 ( n10415, n10380, n10417 );
nor U10125 ( n10413, n10418, n10419 );
nor U10126 ( n10419, n15313, n10375 );
nor U10127 ( n10418, n10237, n10384 );
not U10128 ( n10237, n9643 );
nand U10129 ( n1958, n10420, n10421 );
nor U10130 ( n10421, n10422, n10423 );
and U10131 ( n10423, DATAI_24_, n10370 );
nor U10132 ( n10422, n10380, n10424 );
nor U10133 ( n10420, n10425, n10426 );
nor U10134 ( n10426, n15312, n10375 );
nor U10135 ( n10425, n10242, n10384 );
not U10136 ( n10242, n9663 );
nand U10137 ( n1953, n10427, n10428 );
nor U10138 ( n10428, n10429, n10430 );
and U10139 ( n10430, DATAI_23_, n10370 );
nor U10140 ( n10429, n10431, n10380 );
nor U10141 ( n10427, n10432, n10433 );
nor U10142 ( n10433, n15311, n10375 );
nor U10143 ( n10432, n10247, n10384 );
not U10144 ( n10247, n9682 );
nand U10145 ( n1948, n10434, n10435 );
nor U10146 ( n10435, n10436, n10437 );
and U10147 ( n10437, DATAI_22_, n10370 );
nor U10148 ( n10436, n10438, n10380 );
nor U10149 ( n10434, n10439, n10440 );
nor U10150 ( n10440, n15310, n10375 );
nor U10151 ( n10439, n10252, n10384 );
not U10152 ( n10252, n9702 );
nand U10153 ( n1943, n10441, n10442 );
nor U10154 ( n10442, n10443, n10444 );
and U10155 ( n10444, DATAI_21_, n10370 );
nor U10156 ( n10443, n10445, n10380 );
nor U10157 ( n10441, n10446, n10447 );
nor U10158 ( n10447, n15309, n10375 );
nor U10159 ( n10446, n10257, n10384 );
nand U10160 ( n1938, n10448, n10449 );
nor U10161 ( n10449, n10450, n10451 );
and U10162 ( n10451, DATAI_20_, n10370 );
nor U10163 ( n10450, n10452, n10380 );
nor U10164 ( n10448, n10453, n10454 );
nor U10165 ( n10454, n15308, n10375 );
nor U10166 ( n10453, n10262, n10384 );
not U10167 ( n10262, n9743 );
nand U10168 ( n1933, n10455, n10456 );
nor U10169 ( n10456, n10457, n10458 );
and U10170 ( n10458, DATAI_19_, n10370 );
nor U10171 ( n10457, n10459, n10380 );
nor U10172 ( n10455, n10460, n10461 );
nor U10173 ( n10461, n15307, n10375 );
nor U10174 ( n10460, n10267, n10384 );
not U10175 ( n10267, n9765 );
nand U10176 ( n1928, n10462, n10463 );
nor U10177 ( n10463, n10464, n10465 );
and U10178 ( n10465, DATAI_18_, n10370 );
nor U10179 ( n10464, n10466, n10380 );
nor U10180 ( n10462, n10467, n10468 );
nor U10181 ( n10468, n15306, n10375 );
nor U10182 ( n10467, n10272, n10384 );
not U10183 ( n10272, n9786 );
nand U10184 ( n1923, n10469, n10470 );
nor U10185 ( n10470, n10471, n10472 );
and U10186 ( n10472, DATAI_17_, n10370 );
nor U10187 ( n10471, n10473, n10380 );
nor U10188 ( n10469, n10474, n10475 );
nor U10189 ( n10475, n15305, n10375 );
nor U10190 ( n10474, n10277, n10384 );
not U10191 ( n10277, n9806 );
nand U10192 ( n1918, n10476, n10477 );
nor U10193 ( n10477, n10478, n10479 );
and U10194 ( n10479, DATAI_16_, n10370 );
nor U10195 ( n10370, n10373, n10480 );
nor U10196 ( n10478, n10481, n10380 );
nand U10197 ( n10380, n10482, n10375 );
nor U10198 ( n10482, n10361, n10483 );
nor U10199 ( n10476, n10484, n10485 );
nor U10200 ( n10485, n15304, n10375 );
nor U10201 ( n10484, n10282, n10384 );
nand U10202 ( n1913, n10486, n10487 );
nand U10203 ( n10487, n10373, n8037 );
nor U10204 ( n10486, n10488, n10489 );
nor U10205 ( n10489, n10490, n10491 );
nor U10206 ( n10488, n10287, n10384 );
nand U10207 ( n1908, n10492, n10493 );
nand U10208 ( n10493, n10373, n8036 );
nor U10209 ( n10492, n10494, n10495 );
nor U10210 ( n10495, n10381, n10490 );
nor U10211 ( n10494, n10292, n10384 );
nand U10212 ( n1903, n10496, n10497 );
nand U10213 ( n10497, n10373, n8035 );
nor U10214 ( n10496, n10498, n10499 );
nor U10215 ( n10499, n10389, n10490 );
nor U10216 ( n10498, n10297, n10384 );
not U10217 ( n10297, n9890 );
nand U10218 ( n1898, n10500, n10501 );
nand U10219 ( n10501, n10373, n8034 );
nor U10220 ( n10500, n10502, n10503 );
nor U10221 ( n10503, n10396, n10490 );
nor U10222 ( n10502, n10302, n10384 );
nand U10223 ( n1893, n10504, n10505 );
nand U10224 ( n10505, n10373, n8033 );
nor U10225 ( n10504, n10506, n10507 );
nor U10226 ( n10507, n10403, n10490 );
nor U10227 ( n10506, n10307, n10384 );
not U10228 ( n10307, n9933 );
nand U10229 ( n1888, n10508, n10509 );
nand U10230 ( n10509, n10373, n8032 );
nor U10231 ( n10508, n10510, n10511 );
nor U10232 ( n10511, n10410, n10490 );
nor U10233 ( n10510, n10312, n10384 );
nand U10234 ( n1883, n10512, n10513 );
nand U10235 ( n10513, n10373, n8031 );
nor U10236 ( n10512, n10514, n10515 );
nor U10237 ( n10515, n10417, n10490 );
nor U10238 ( n10514, n10317, n10384 );
not U10239 ( n10317, n9975 );
nand U10240 ( n1878, n10516, n10517 );
nand U10241 ( n10517, n10373, n8030 );
nor U10242 ( n10516, n10518, n10519 );
nor U10243 ( n10519, n10424, n10490 );
nor U10244 ( n10518, n10322, n10384 );
nand U10245 ( n1873, n10520, n10521 );
nand U10246 ( n10521, n10373, n8029 );
nor U10247 ( n10520, n10522, n10523 );
nor U10248 ( n10523, n10431, n10490 );
nor U10249 ( n10522, n10327, n10384 );
not U10250 ( n10327, n10016 );
nand U10251 ( n1868, n10524, n10525 );
nand U10252 ( n10525, n10373, n8028 );
nor U10253 ( n10524, n10526, n10527 );
nor U10254 ( n10527, n10438, n10490 );
nor U10255 ( n10526, n10332, n10384 );
not U10256 ( n10332, n10037 );
nand U10257 ( n1863, n10528, n10529 );
nand U10258 ( n10529, n10373, n8027 );
nor U10259 ( n10528, n10530, n10531 );
nor U10260 ( n10531, n10445, n10490 );
nor U10261 ( n10530, n10337, n10384 );
not U10262 ( n10337, n10058 );
nand U10263 ( n1858, n10532, n10533 );
nand U10264 ( n10533, n10373, n8026 );
nor U10265 ( n10532, n10534, n10535 );
nor U10266 ( n10535, n10452, n10490 );
nor U10267 ( n10534, n10342, n10384 );
not U10268 ( n10342, n10081 );
nand U10269 ( n1853, n10536, n10537 );
nand U10270 ( n10537, n10373, n8025 );
nor U10271 ( n10536, n10538, n10539 );
nor U10272 ( n10539, n10459, n10490 );
nor U10273 ( n10538, n10347, n10384 );
nand U10274 ( n1848, n10540, n10541 );
nand U10275 ( n10541, n10373, n8024 );
nor U10276 ( n10540, n10542, n10543 );
nor U10277 ( n10543, n10466, n10490 );
nor U10278 ( n10542, n10352, n10384 );
nand U10279 ( n1843, n10544, n10545 );
nand U10280 ( n10545, n10373, n8023 );
nor U10281 ( n10544, n10546, n10547 );
nor U10282 ( n10547, n10473, n10490 );
nor U10283 ( n10546, n10144, n10384 );
nand U10284 ( n1838, n10548, n10549 );
nand U10285 ( n10549, n10373, n7873 );
nor U10286 ( n10548, n10550, n10551 );
nor U10287 ( n10551, n10481, n10490 );
nand U10288 ( n10490, n10552, n10375 );
nor U10289 ( n10552, n10361, n10553 );
nor U10290 ( n10550, n10180, n10384 );
nand U10291 ( n10554, n10555, n9407 );
not U10292 ( n10375, n10373 );
nand U10293 ( n10373, n9120, n10556 );
nand U10294 ( n10556, n10557, n10558 );
nand U10295 ( n10558, n10559, n10560 );
nor U10296 ( n10560, n9428, n10561 );
nand U10297 ( n10561, n9106, n7814 );
nand U10298 ( n10557, n10562, n10563 );
nand U10299 ( n10563, n10564, n10565 );
nand U10300 ( n10565, n10366, n10367 );
and U10301 ( n10366, n10566, n10567 );
nor U10302 ( n10567, n10568, n10569 );
nor U10303 ( n10566, n10570, n9407 );
nor U10304 ( n10564, n10571, n10572 );
nor U10305 ( n10572, n10573, n10574 );
nand U10306 ( n10574, n9415, n10569 );
nor U10307 ( n10571, n9349, n10575 );
nand U10308 ( n10575, n9348, n9106 );
nor U10309 ( n1834, n15012, n10576 );
nand U10310 ( n1830, n10577, n10578 );
nand U10311 ( n10578, n10579, DATAO_REG_30_ );
nor U10312 ( n10577, n10580, n10581 );
nor U10313 ( n10581, n15273, n10582 );
nor U10314 ( n10580, n15318, n10583 );
nand U10315 ( n1826, n10584, n10585 );
nand U10316 ( n10585, n10579, DATAO_REG_29_ );
nor U10317 ( n10584, n10586, n10587 );
nor U10318 ( n10587, n15274, n10582 );
nor U10319 ( n10586, n15317, n10583 );
nand U10320 ( n1822, n10588, n10589 );
nand U10321 ( n10589, n10579, DATAO_REG_28_ );
nor U10322 ( n10588, n10590, n10591 );
nor U10323 ( n10591, n15275, n10582 );
nor U10324 ( n10590, n15316, n10583 );
nand U10325 ( n1818, n10592, n10593 );
nand U10326 ( n10593, n10579, DATAO_REG_27_ );
nor U10327 ( n10592, n10594, n10595 );
nor U10328 ( n10595, n15276, n10582 );
nor U10329 ( n10594, n15315, n10583 );
nand U10330 ( n1814, n10596, n10597 );
nand U10331 ( n10597, n10579, DATAO_REG_26_ );
nor U10332 ( n10596, n10598, n10599 );
nor U10333 ( n10599, n15277, n10582 );
nor U10334 ( n10598, n15314, n10583 );
nand U10335 ( n1810, n10600, n10601 );
nand U10336 ( n10601, n10579, DATAO_REG_25_ );
nor U10337 ( n10600, n10602, n10603 );
nor U10338 ( n10603, n15278, n10582 );
nor U10339 ( n10602, n15313, n10583 );
nand U10340 ( n1806, n10604, n10605 );
nand U10341 ( n10605, n10579, DATAO_REG_24_ );
nor U10342 ( n10604, n10606, n10607 );
nor U10343 ( n10607, n15279, n10582 );
nor U10344 ( n10606, n15312, n10583 );
nand U10345 ( n1802, n10608, n10609 );
nand U10346 ( n10609, n10579, DATAO_REG_23_ );
nor U10347 ( n10608, n10610, n10611 );
nor U10348 ( n10611, n15280, n10582 );
nor U10349 ( n10610, n15311, n10583 );
nand U10350 ( n1798, n10612, n10613 );
nand U10351 ( n10613, n10579, DATAO_REG_22_ );
nor U10352 ( n10612, n10614, n10615 );
nor U10353 ( n10615, n15281, n10582 );
nor U10354 ( n10614, n15310, n10583 );
nand U10355 ( n1794, n10616, n10617 );
nand U10356 ( n10617, n10579, DATAO_REG_21_ );
nor U10357 ( n10616, n10618, n10619 );
nor U10358 ( n10619, n15282, n10582 );
nor U10359 ( n10618, n15309, n10583 );
nand U10360 ( n1790, n10620, n10621 );
nand U10361 ( n10621, n10579, DATAO_REG_20_ );
nor U10362 ( n10620, n10622, n10623 );
nor U10363 ( n10623, n15283, n10582 );
nor U10364 ( n10622, n15308, n10583 );
nand U10365 ( n1786, n10624, n10625 );
nand U10366 ( n10625, n10579, DATAO_REG_19_ );
nor U10367 ( n10624, n10626, n10627 );
nor U10368 ( n10627, n15284, n10582 );
nor U10369 ( n10626, n15307, n10583 );
nand U10370 ( n1782, n10628, n10629 );
nand U10371 ( n10629, n10579, DATAO_REG_18_ );
nor U10372 ( n10628, n10630, n10631 );
nor U10373 ( n10631, n15285, n10582 );
nor U10374 ( n10630, n15306, n10583 );
nand U10375 ( n1778, n10632, n10633 );
nand U10376 ( n10633, n10579, DATAO_REG_17_ );
nor U10377 ( n10632, n10634, n10635 );
nor U10378 ( n10635, n15286, n10582 );
nor U10379 ( n10634, n15305, n10583 );
nand U10380 ( n1774, n10636, n10637 );
nand U10381 ( n10637, n10579, DATAO_REG_16_ );
nor U10382 ( n10636, n10638, n10639 );
nor U10383 ( n10639, n15287, n10582 );
nor U10384 ( n10638, n15304, n10583 );
or U10385 ( n10583, n10640, n9139 );
nand U10386 ( n1770, n10641, n10642 );
nand U10387 ( n10642, n10579, DATAO_REG_15_ );
nor U10388 ( n10641, n10643, n10644 );
nor U10389 ( n10644, n15257, n10582 );
nor U10390 ( n10643, n15303, n10640 );
nand U10391 ( n1766, n10645, n10646 );
nand U10392 ( n10646, n10579, DATAO_REG_14_ );
nor U10393 ( n10645, n10647, n10648 );
nor U10394 ( n10648, n15258, n10582 );
nor U10395 ( n10647, n15302, n10640 );
nand U10396 ( n1762, n10649, n10650 );
nand U10397 ( n10650, n10579, DATAO_REG_13_ );
nor U10398 ( n10649, n10651, n10652 );
nor U10399 ( n10652, n15259, n10582 );
nor U10400 ( n10651, n15301, n10640 );
nand U10401 ( n1758, n10653, n10654 );
nand U10402 ( n10654, n10579, DATAO_REG_12_ );
nor U10403 ( n10653, n10655, n10656 );
nor U10404 ( n10656, n15260, n10582 );
nor U10405 ( n10655, n15300, n10640 );
nand U10406 ( n1754, n10657, n10658 );
nand U10407 ( n10658, n10579, DATAO_REG_11_ );
nor U10408 ( n10657, n10659, n10660 );
nor U10409 ( n10660, n15261, n10582 );
nor U10410 ( n10659, n15299, n10640 );
nand U10411 ( n1750, n10661, n10662 );
nand U10412 ( n10662, n10579, DATAO_REG_10_ );
nor U10413 ( n10661, n10663, n10664 );
nor U10414 ( n10664, n15262, n10582 );
nor U10415 ( n10663, n15298, n10640 );
nand U10416 ( n1746, n10665, n10666 );
nand U10417 ( n10666, n10579, DATAO_REG_9_ );
nor U10418 ( n10665, n10667, n10668 );
nor U10419 ( n10668, n15263, n10582 );
nor U10420 ( n10667, n15297, n10640 );
nand U10421 ( n1742, n10669, n10670 );
nand U10422 ( n10670, n10579, DATAO_REG_8_ );
nor U10423 ( n10669, n10671, n10672 );
nor U10424 ( n10672, n15264, n10582 );
nor U10425 ( n10671, n15296, n10640 );
nand U10426 ( n1738, n10673, n10674 );
nand U10427 ( n10674, n10579, DATAO_REG_7_ );
nor U10428 ( n10673, n10675, n10676 );
nor U10429 ( n10676, n15265, n10582 );
nor U10430 ( n10675, n15295, n10640 );
nand U10431 ( n1734, n10677, n10678 );
nand U10432 ( n10678, n10579, DATAO_REG_6_ );
nor U10433 ( n10677, n10679, n10680 );
nor U10434 ( n10680, n15266, n10582 );
nor U10435 ( n10679, n15294, n10640 );
nand U10436 ( n1730, n10681, n10682 );
nand U10437 ( n10682, n10579, DATAO_REG_5_ );
nor U10438 ( n10681, n10683, n10684 );
nor U10439 ( n10684, n15267, n10582 );
nor U10440 ( n10683, n15293, n10640 );
nand U10441 ( n1726, n10685, n10686 );
nand U10442 ( n10686, n10579, DATAO_REG_4_ );
nor U10443 ( n10685, n10687, n10688 );
nor U10444 ( n10688, n15268, n10582 );
nor U10445 ( n10687, n15292, n10640 );
nand U10446 ( n1722, n10689, n10690 );
nand U10447 ( n10690, n10579, DATAO_REG_3_ );
nor U10448 ( n10689, n10691, n10692 );
nor U10449 ( n10692, n15269, n10582 );
nor U10450 ( n10691, n15291, n10640 );
nand U10451 ( n1718, n10693, n10694 );
nand U10452 ( n10694, n10579, DATAO_REG_2_ );
nor U10453 ( n10693, n10695, n10696 );
nor U10454 ( n10696, n15270, n10582 );
nor U10455 ( n10695, n15290, n10640 );
nand U10456 ( n1714, n10697, n10698 );
nand U10457 ( n10698, n10579, DATAO_REG_1_ );
nor U10458 ( n10697, n10699, n10700 );
nor U10459 ( n10700, n15271, n10582 );
nor U10460 ( n10699, n15289, n10640 );
nand U10461 ( n1710, n10701, n10702 );
nand U10462 ( n10702, n10579, DATAO_REG_0_ );
nor U10463 ( n10701, n10703, n10704 );
nor U10464 ( n10704, n15272, n10582 );
nor U10465 ( n10703, n15288, n10640 );
nand U10466 ( n10640, n7814, n10576 );
nand U10467 ( n10576, n10705, n10706 );
nand U10468 ( n10706, n10707, n10197 );
not U10469 ( n10197, n10708 );
nor U10470 ( n10707, n10709, n10710 );
nor U10471 ( n10709, n10711, n10199 );
nand U10472 ( n10705, n9125, n15063 );
nand U10473 ( n1705, n10712, n10713 );
nand U10474 ( n10713, n10714, n8071 );
nor U10475 ( n10712, n10715, n10716 );
nor U10476 ( n10715, n15287, n10717 );
nand U10477 ( n1700, n10718, n10719 );
nand U10478 ( n10719, n10714, n8072 );
nor U10479 ( n10718, n10720, n10721 );
nor U10480 ( n10720, n15286, n10717 );
nand U10481 ( n1695, n10722, n10723 );
nand U10482 ( n10723, n10714, n8073 );
nor U10483 ( n10722, n10724, n10725 );
nor U10484 ( n10724, n15285, n10717 );
nand U10485 ( n1690, n10726, n10727 );
nand U10486 ( n10727, n10714, n8074 );
nor U10487 ( n10726, n10728, n10729 );
nor U10488 ( n10728, n15284, n10717 );
nand U10489 ( n1685, n10730, n10731 );
nand U10490 ( n10731, n10714, n8075 );
nor U10491 ( n10730, n10732, n10733 );
nor U10492 ( n10732, n15283, n10717 );
nand U10493 ( n1680, n10734, n10735 );
nand U10494 ( n10735, n10714, n8076 );
nor U10495 ( n10734, n10736, n10737 );
nor U10496 ( n10736, n15282, n10717 );
nand U10497 ( n1675, n10738, n10739 );
nand U10498 ( n10739, n10714, n8077 );
nor U10499 ( n10738, n10740, n10741 );
nor U10500 ( n10740, n15281, n10717 );
nand U10501 ( n1670, n10742, n10743 );
nand U10502 ( n10743, n10714, n8042 );
nor U10503 ( n10742, n10744, n10745 );
nor U10504 ( n10744, n15280, n10717 );
nand U10505 ( n1665, n10746, n10747 );
nand U10506 ( n10747, n10714, n8078 );
nor U10507 ( n10746, n10748, n10749 );
nor U10508 ( n10748, n15279, n10717 );
nand U10509 ( n1660, n10750, n10751 );
nand U10510 ( n10751, n10714, n8041 );
nor U10511 ( n10750, n10752, n10753 );
nor U10512 ( n10752, n15278, n10717 );
nand U10513 ( n1655, n10754, n10755 );
nand U10514 ( n10755, n10714, n8040 );
nor U10515 ( n10754, n10756, n10757 );
nor U10516 ( n10756, n15277, n10717 );
nand U10517 ( n1650, n10758, n10759 );
nand U10518 ( n10759, n10714, n8039 );
nor U10519 ( n10758, n10760, n10761 );
nor U10520 ( n10760, n15276, n10717 );
nand U10521 ( n1645, n10762, n10763 );
nand U10522 ( n10763, n10714, n8079 );
nor U10523 ( n10762, n10764, n10765 );
nor U10524 ( n10764, n15275, n10717 );
nand U10525 ( n1640, n10766, n10767 );
nand U10526 ( n10767, n10714, n8080 );
nor U10527 ( n10766, n10768, n10769 );
nor U10528 ( n10768, n15274, n10717 );
nand U10529 ( n1635, n10770, n10771 );
nand U10530 ( n10771, n10714, n8038 );
nor U10531 ( n10770, n10772, n10773 );
nor U10532 ( n10772, n15273, n10717 );
nand U10533 ( n1630, n10774, n10775 );
nand U10534 ( n10775, n10714, n7873 );
nor U10535 ( n10774, n10776, n10716 );
nor U10536 ( n10716, n10481, n10777 );
nor U10537 ( n10776, n15272, n10717 );
nand U10538 ( n1625, n10778, n10779 );
nand U10539 ( n10779, n10714, n8023 );
nor U10540 ( n10778, n10780, n10721 );
nor U10541 ( n10721, n10473, n10777 );
nor U10542 ( n10780, n15271, n10717 );
nand U10543 ( n1620, n10781, n10782 );
nand U10544 ( n10782, n10714, n8024 );
nor U10545 ( n10781, n10783, n10725 );
nor U10546 ( n10725, n10466, n10777 );
nor U10547 ( n10783, n15270, n10717 );
nand U10548 ( n1615, n10784, n10785 );
nand U10549 ( n10785, n10714, n8025 );
nor U10550 ( n10784, n10786, n10729 );
nor U10551 ( n10729, n10459, n10777 );
nor U10552 ( n10786, n15269, n10717 );
nand U10553 ( n1610, n10787, n10788 );
nand U10554 ( n10788, n10714, n8026 );
nor U10555 ( n10787, n10789, n10733 );
nor U10556 ( n10733, n10452, n10777 );
nor U10557 ( n10789, n15268, n10717 );
nand U10558 ( n1605, n10790, n10791 );
nand U10559 ( n10791, n10714, n8027 );
nor U10560 ( n10790, n10792, n10737 );
nor U10561 ( n10737, n10445, n10777 );
nor U10562 ( n10792, n15267, n10717 );
nand U10563 ( n1600, n10793, n10794 );
nand U10564 ( n10794, n10714, n8028 );
nor U10565 ( n10793, n10795, n10741 );
nor U10566 ( n10741, n10438, n10777 );
nor U10567 ( n10795, n15266, n10717 );
nand U10568 ( n1595, n10796, n10797 );
nand U10569 ( n10797, n10714, n8029 );
nor U10570 ( n10796, n10798, n10745 );
nor U10571 ( n10745, n10431, n10777 );
nor U10572 ( n10798, n15265, n10717 );
nand U10573 ( n1590, n10799, n10800 );
nand U10574 ( n10800, n10714, n8030 );
nor U10575 ( n10799, n10801, n10749 );
nor U10576 ( n10749, n10424, n10777 );
not U10577 ( n10424, DATAI_8_ );
nor U10578 ( n10801, n15264, n10717 );
nand U10579 ( n1585, n10802, n10803 );
nand U10580 ( n10803, n10714, n8031 );
nor U10581 ( n10802, n10804, n10753 );
nor U10582 ( n10753, n10417, n10777 );
not U10583 ( n10417, DATAI_9_ );
nor U10584 ( n10804, n15263, n10717 );
nand U10585 ( n1580, n10805, n10806 );
nand U10586 ( n10806, n10714, n8032 );
nor U10587 ( n10805, n10807, n10757 );
nor U10588 ( n10757, n10410, n10777 );
not U10589 ( n10410, DATAI_10_ );
nor U10590 ( n10807, n15262, n10717 );
nand U10591 ( n1575, n10808, n10809 );
nand U10592 ( n10809, n10714, n8033 );
nor U10593 ( n10808, n10810, n10761 );
nor U10594 ( n10761, n10403, n10777 );
not U10595 ( n10403, DATAI_11_ );
nor U10596 ( n10810, n15261, n10717 );
nand U10597 ( n1570, n10811, n10812 );
nand U10598 ( n10812, n10714, n8034 );
nor U10599 ( n10811, n10813, n10765 );
nor U10600 ( n10765, n10396, n10777 );
not U10601 ( n10396, DATAI_12_ );
nor U10602 ( n10813, n15260, n10717 );
nand U10603 ( n1565, n10814, n10815 );
nand U10604 ( n10815, n10714, n8035 );
nor U10605 ( n10814, n10816, n10769 );
nor U10606 ( n10769, n10389, n10777 );
not U10607 ( n10389, DATAI_13_ );
nor U10608 ( n10816, n15259, n10717 );
nand U10609 ( n1560, n10817, n10818 );
nand U10610 ( n10818, n10714, n8036 );
nor U10611 ( n10817, n10819, n10773 );
nor U10612 ( n10773, n10381, n10777 );
not U10613 ( n10381, DATAI_14_ );
nor U10614 ( n10819, n15258, n10717 );
nand U10615 ( n1555, n10820, n10821 );
nand U10616 ( n10821, n10714, n8037 );
nor U10617 ( n10820, n10823, n10824 );
nor U10618 ( n10824, n10491, n10777 );
nand U10619 ( n10777, n10717, n10825 );
not U10620 ( n10491, DATAI_15_ );
nor U10621 ( n10823, n15257, n10717 );
nor U10622 ( n10827, n9139, n10828 );
nor U10623 ( n10828, n9393, n9106 );
nor U10624 ( n10826, n10198, n10708 );
nand U10625 ( n1550, n10829, n10830 );
nor U10626 ( n10830, n10831, n10832 );
nand U10627 ( n10832, n10833, n10834 );
nand U10628 ( n10834, n10835, n9520 );
xor U10629 ( n9520, n10836, n10837 );
nor U10630 ( n10837, n10838, n10839 );
nand U10631 ( n10839, n10840, n8082 );
nand U10632 ( n10840, n10842, n7852 );
nor U10633 ( n10838, n15013, n10843 );
xor U10634 ( n10836, n8082, n10844 );
nor U10635 ( n10844, n10845, n10846 );
nand U10636 ( n10833, n10847, n10165 );
xor U10637 ( n10165, n7852, n10848 );
nor U10638 ( n10848, n15014, n10849 );
nor U10639 ( n10831, n10850, n10851 );
nor U10640 ( n10829, n10852, n10853 );
nor U10641 ( n10853, n15256, n10854 );
nor U10642 ( n10852, n15350, n10855 );
nand U10643 ( n1545, n10856, n10857 );
nor U10644 ( n10857, n10858, n10859 );
nand U10645 ( n10859, n10860, n10861 );
nand U10646 ( n10861, n10835, n9537 );
xor U10647 ( n9537, n10846, n10845 );
xor U10648 ( n10845, n10188, n10862 );
nor U10649 ( n10862, n10863, n10864 );
nand U10650 ( n10864, n10865, n10866 );
nand U10651 ( n10866, n10842, n8017 );
nand U10652 ( n10865, n10867, n8038 );
nand U10653 ( n10863, n10868, n10869 );
nand U10654 ( n10869, n10870, n10871 );
xor U10655 ( n10870, n10872, n10873 );
nor U10656 ( n10873, n10874, n10875 );
nand U10657 ( n10872, n10876, n10877 );
nor U10658 ( n10877, n10878, n10879 );
nand U10659 ( n10879, n10880, n10881 );
nor U10660 ( n10881, n10882, n10883 );
nor U10661 ( n10883, n15168, n10884 );
nor U10662 ( n10882, n15160, n10885 );
nor U10663 ( n10880, n10886, n10887 );
nor U10664 ( n10887, n15176, n10888 );
nor U10665 ( n10886, n15184, n10889 );
nand U10666 ( n10878, n10890, n10891 );
nor U10667 ( n10891, n10892, n10893 );
nor U10668 ( n10893, n15136, n10894 );
nor U10669 ( n10892, n15128, n10895 );
nor U10670 ( n10890, n10896, n10897 );
nor U10671 ( n10897, n15144, n10898 );
nor U10672 ( n10896, n15152, n10899 );
nor U10673 ( n10876, n10900, n10901 );
nand U10674 ( n10901, n10902, n10903 );
nor U10675 ( n10903, n10904, n10905 );
nor U10676 ( n10905, n15072, n10906 );
nor U10677 ( n10904, n15064, n10907 );
nor U10678 ( n10902, n10908, n10909 );
nor U10679 ( n10909, n15080, n10910 );
nor U10680 ( n10908, n15088, n10911 );
nand U10681 ( n10900, n10912, n10913 );
nor U10682 ( n10913, n10914, n10915 );
nor U10683 ( n10915, n15104, n10916 );
nor U10684 ( n10914, n15096, n10917 );
nor U10685 ( n10912, n10918, n10919 );
nor U10686 ( n10919, n15112, n10920 );
nor U10687 ( n10918, n15120, n10921 );
nand U10688 ( n10868, n9529, n10188 );
or U10689 ( n10846, n10922, n10923 );
nand U10690 ( n10860, n10847, n9529 );
xor U10691 ( n9529, n10849, n15014 );
nor U10692 ( n10858, n10924, n10851 );
nor U10693 ( n10856, n10925, n10926 );
nor U10694 ( n10926, n15014, n10854 );
nor U10695 ( n10925, n15349, n10855 );
nand U10696 ( n1540, n10927, n10928 );
nor U10697 ( n10928, n10929, n10930 );
nand U10698 ( n10930, n10931, n10932 );
nand U10699 ( n10932, n10835, n9559 );
xor U10700 ( n9559, n10922, n10923 );
xnor U10701 ( n10923, n10933, n10188 );
nand U10702 ( n10933, n10934, n10935 );
nor U10703 ( n10935, n10936, n10937 );
nor U10704 ( n10937, n8082, n10938 );
nor U10705 ( n10936, n10939, n10940 );
xnor U10706 ( n10940, n10875, n10874 );
and U10707 ( n10874, n10941, n10942 );
nor U10708 ( n10942, n10943, n10944 );
nand U10709 ( n10944, n10945, n10946 );
nor U10710 ( n10946, n10947, n10948 );
nor U10711 ( n10948, n15169, n10884 );
nor U10712 ( n10947, n15161, n10885 );
nor U10713 ( n10945, n10949, n10950 );
nor U10714 ( n10950, n15177, n10888 );
nor U10715 ( n10949, n15185, n10889 );
nand U10716 ( n10943, n10951, n10952 );
nor U10717 ( n10952, n10953, n10954 );
nor U10718 ( n10954, n15137, n10894 );
nor U10719 ( n10953, n15129, n10895 );
nor U10720 ( n10951, n10955, n10956 );
nor U10721 ( n10956, n15145, n10898 );
nor U10722 ( n10955, n15153, n10899 );
nor U10723 ( n10941, n10957, n10958 );
nand U10724 ( n10958, n10959, n10960 );
nor U10725 ( n10960, n10961, n10962 );
nor U10726 ( n10962, n15073, n10906 );
nor U10727 ( n10961, n15065, n10907 );
nor U10728 ( n10959, n10963, n10964 );
nor U10729 ( n10964, n15081, n10910 );
nor U10730 ( n10963, n15089, n10911 );
nand U10731 ( n10957, n10965, n10966 );
nor U10732 ( n10966, n10967, n10968 );
nor U10733 ( n10968, n15105, n10916 );
nor U10734 ( n10967, n15097, n10917 );
nor U10735 ( n10965, n10969, n10970 );
nor U10736 ( n10970, n15113, n10920 );
nor U10737 ( n10969, n15121, n10921 );
nand U10738 ( n10875, n10971, n10972 );
nor U10739 ( n10934, n10973, n10974 );
nor U10740 ( n10974, n15317, n10843 );
nor U10741 ( n10973, n15255, n10975 );
nand U10742 ( n10922, n10976, n10977 );
nand U10743 ( n10931, n10847, n9553 );
not U10744 ( n9553, n10938 );
nand U10745 ( n10938, n10849, n10978 );
nand U10746 ( n10978, n15255, n10979 );
nand U10747 ( n10979, n10980, n7847 );
nand U10748 ( n10849, n10981, n10980 );
nor U10749 ( n10981, n15254, n15255 );
nor U10750 ( n10929, n10851, n10982 );
nor U10751 ( n10927, n10983, n10984 );
nor U10752 ( n10984, n15255, n10854 );
nor U10753 ( n10983, n15348, n10855 );
nand U10754 ( n1535, n10985, n10986 );
nor U10755 ( n10986, n10987, n10988 );
nand U10756 ( n10988, n10989, n10990 );
nand U10757 ( n10990, n10835, n9584 );
xor U10758 ( n9584, n10976, n10977 );
xnor U10759 ( n10977, n10991, n8082 );
nand U10760 ( n10991, n10992, n10993 );
nor U10761 ( n10993, n10994, n10995 );
nor U10762 ( n10995, n15254, n10975 );
nor U10763 ( n10994, n8082, n10996 );
nor U10764 ( n10992, n10997, n10998 );
nand U10765 ( n10998, n10999, n11000 );
nand U10766 ( n11000, n11001, n10972 );
nor U10767 ( n11001, n10939, n10971 );
nand U10768 ( n10999, n11002, n10971 );
nor U10769 ( n10971, n11003, n11004 );
not U10770 ( n11002, n10972 );
nand U10771 ( n10972, n11005, n11006 );
nor U10772 ( n11006, n11007, n11008 );
nand U10773 ( n11008, n11009, n11010 );
nor U10774 ( n11010, n11011, n11012 );
nor U10775 ( n11012, n15106, n10916 );
nor U10776 ( n11011, n15098, n10917 );
nor U10777 ( n11009, n11013, n11014 );
nor U10778 ( n11014, n15114, n10920 );
nor U10779 ( n11013, n15122, n10921 );
nand U10780 ( n11007, n11015, n11016 );
nor U10781 ( n11016, n11017, n11018 );
nor U10782 ( n11018, n15074, n10906 );
nor U10783 ( n11017, n15066, n10907 );
nor U10784 ( n11015, n11019, n11020 );
nor U10785 ( n11020, n15082, n10910 );
nor U10786 ( n11019, n15090, n10911 );
nor U10787 ( n11005, n11021, n11022 );
nand U10788 ( n11022, n11023, n11024 );
nor U10789 ( n11024, n11025, n11026 );
nor U10790 ( n11026, n15138, n10894 );
nor U10791 ( n11025, n15130, n10895 );
nor U10792 ( n11023, n11027, n11028 );
nor U10793 ( n11028, n15146, n10898 );
nor U10794 ( n11027, n15154, n10899 );
nand U10795 ( n11021, n11029, n11030 );
nor U10796 ( n11030, n11031, n11032 );
nor U10797 ( n11032, n15170, n10884 );
nor U10798 ( n11031, n15162, n10885 );
nor U10799 ( n11029, n11033, n11034 );
nor U10800 ( n11034, n15178, n10888 );
nor U10801 ( n11033, n15186, n10889 );
nor U10802 ( n10997, n15316, n10843 );
nor U10803 ( n10976, n11035, n11036 );
nand U10804 ( n10989, n10847, n9578 );
not U10805 ( n9578, n10996 );
xnor U10806 ( n10996, n7847, n10980 );
not U10807 ( n10980, n11037 );
nor U10808 ( n10987, n11038, n10851 );
nor U10809 ( n10985, n11039, n11040 );
nor U10810 ( n11040, n15254, n10854 );
nor U10811 ( n11039, n15347, n10855 );
nand U10812 ( n1530, n11041, n11042 );
nor U10813 ( n11042, n11043, n11044 );
nand U10814 ( n11044, n11045, n11046 );
nand U10815 ( n11046, n10835, n9604 );
xor U10816 ( n9604, n11035, n11036 );
xnor U10817 ( n11036, n8082, n11047 );
nor U10818 ( n11047, n11048, n11049 );
nand U10819 ( n11049, n11050, n11051 );
nand U10820 ( n11051, n10842, n8018 );
nand U10821 ( n11050, n10867, n8039 );
nand U10822 ( n11048, n11052, n11053 );
nand U10823 ( n11053, n11054, n10871 );
xor U10824 ( n11054, n11003, n11004 );
and U10825 ( n11004, n11055, n11056 );
nor U10826 ( n11056, n11057, n11058 );
nand U10827 ( n11058, n11059, n11060 );
nor U10828 ( n11060, n11061, n11062 );
nor U10829 ( n11062, n15171, n10884 );
nor U10830 ( n11061, n15163, n10885 );
nor U10831 ( n11059, n11063, n11064 );
nor U10832 ( n11064, n15179, n10888 );
nor U10833 ( n11063, n15187, n10889 );
nand U10834 ( n11057, n11065, n11066 );
nor U10835 ( n11066, n11067, n11068 );
nor U10836 ( n11068, n15139, n10894 );
nor U10837 ( n11067, n15131, n10895 );
nor U10838 ( n11065, n11069, n11070 );
nor U10839 ( n11070, n15147, n10898 );
nor U10840 ( n11069, n15155, n10899 );
nor U10841 ( n11055, n11071, n11072 );
nand U10842 ( n11072, n11073, n11074 );
nor U10843 ( n11074, n11075, n11076 );
nor U10844 ( n11076, n15075, n10906 );
nor U10845 ( n11075, n15067, n10907 );
nor U10846 ( n11073, n11077, n11078 );
nor U10847 ( n11078, n15083, n10910 );
nor U10848 ( n11077, n15091, n10911 );
nand U10849 ( n11071, n11079, n11080 );
nor U10850 ( n11080, n11081, n11082 );
nor U10851 ( n11082, n15107, n10916 );
nor U10852 ( n11081, n15099, n10917 );
nor U10853 ( n11079, n11083, n11084 );
nor U10854 ( n11084, n15115, n10920 );
nor U10855 ( n11083, n15123, n10921 );
nand U10856 ( n11003, n11085, n11086 );
nand U10857 ( n11052, n9598, n10188 );
nand U10858 ( n11035, n11087, n11088 );
nand U10859 ( n11045, n10847, n9598 );
and U10860 ( n9598, n11037, n11089 );
nand U10861 ( n11089, n15253, n11090 );
nand U10862 ( n11090, n11091, n7861 );
nand U10863 ( n11037, n11092, n11091 );
not U10864 ( n11091, n11093 );
nor U10865 ( n11092, n15252, n15253 );
nor U10866 ( n11043, n10851, n11094 );
nor U10867 ( n11041, n11095, n11096 );
nor U10868 ( n11096, n15253, n10854 );
nor U10869 ( n11095, n15346, n10855 );
nand U10870 ( n1525, n11097, n11098 );
nor U10871 ( n11098, n11099, n11100 );
nand U10872 ( n11100, n11101, n11102 );
nand U10873 ( n11102, n10835, n9623 );
xor U10874 ( n9623, n11087, n11088 );
xnor U10875 ( n11088, n10188, n11103 );
nor U10876 ( n11103, n11104, n11105 );
nand U10877 ( n11105, n11106, n11107 );
nand U10878 ( n11107, n10867, n8040 );
nor U10879 ( n11106, n11108, n11109 );
nor U10880 ( n11109, n11110, n11086 );
nor U10881 ( n11108, n11085, n11111 );
nand U10882 ( n11111, n11086, n10871 );
nand U10883 ( n11086, n11112, n11113 );
nor U10884 ( n11113, n11114, n11115 );
nand U10885 ( n11115, n11116, n11117 );
nor U10886 ( n11117, n11118, n11119 );
nor U10887 ( n11119, n15172, n10884 );
nor U10888 ( n11118, n15164, n10885 );
nor U10889 ( n11116, n11120, n11121 );
nor U10890 ( n11121, n15180, n10888 );
nor U10891 ( n11120, n15188, n10889 );
nand U10892 ( n11114, n11122, n11123 );
nor U10893 ( n11123, n11124, n11125 );
nor U10894 ( n11125, n15140, n10894 );
nor U10895 ( n11124, n15132, n10895 );
nor U10896 ( n11122, n11126, n11127 );
nor U10897 ( n11127, n15148, n10898 );
nor U10898 ( n11126, n15156, n10899 );
nor U10899 ( n11112, n11128, n11129 );
nand U10900 ( n11129, n11130, n11131 );
nor U10901 ( n11131, n11132, n11133 );
nor U10902 ( n11133, n15076, n10906 );
nor U10903 ( n11132, n15068, n10907 );
nor U10904 ( n11130, n11134, n11135 );
nor U10905 ( n11135, n15084, n10910 );
nor U10906 ( n11134, n15092, n10911 );
nand U10907 ( n11128, n11136, n11137 );
nor U10908 ( n11137, n11138, n11139 );
nor U10909 ( n11139, n15108, n10916 );
nor U10910 ( n11138, n15100, n10917 );
nor U10911 ( n11136, n11140, n11141 );
nor U10912 ( n11141, n15116, n10920 );
nor U10913 ( n11140, n15124, n10921 );
not U10914 ( n11085, n11110 );
nand U10915 ( n11110, n11142, n11143 );
nor U10916 ( n11142, n11144, n11145 );
nand U10917 ( n11104, n11146, n11147 );
nand U10918 ( n11147, n9617, n10188 );
nand U10919 ( n11146, n10842, n7861 );
nor U10920 ( n11087, n11148, n11149 );
nand U10921 ( n11101, n10847, n9617 );
xor U10922 ( n9617, n11093, n15252 );
nor U10923 ( n11099, n10851, n11150 );
nor U10924 ( n11097, n11151, n11152 );
nor U10925 ( n11152, n15252, n10854 );
nor U10926 ( n11151, n15345, n10855 );
nand U10927 ( n1520, n11153, n11154 );
nor U10928 ( n11154, n11155, n11156 );
nand U10929 ( n11156, n11157, n11158 );
nand U10930 ( n11158, n11159, n11160 );
and U10931 ( n11159, n11161, n11162 );
nand U10932 ( n11157, n10835, n9643 );
xor U10933 ( n9643, n11148, n11149 );
xnor U10934 ( n11149, n8082, n11163 );
nor U10935 ( n11163, n11164, n11165 );
nand U10936 ( n11165, n11166, n11167 );
nand U10937 ( n11167, n10842, n8019 );
nand U10938 ( n11166, n10867, n8041 );
nand U10939 ( n11164, n11168, n11169 );
nand U10940 ( n11169, n11170, n10871 );
xnor U10941 ( n11170, n11145, n11171 );
nor U10942 ( n11171, n11144, n11172 );
and U10943 ( n11145, n11173, n11174 );
nor U10944 ( n11174, n11175, n11176 );
nand U10945 ( n11176, n11177, n11178 );
nor U10946 ( n11178, n11179, n11180 );
nor U10947 ( n11180, n15173, n10884 );
nor U10948 ( n11179, n15165, n10885 );
nor U10949 ( n11177, n11181, n11182 );
nor U10950 ( n11182, n15181, n10888 );
nor U10951 ( n11181, n15189, n10889 );
nand U10952 ( n11175, n11183, n11184 );
nor U10953 ( n11184, n11185, n11186 );
nor U10954 ( n11186, n15141, n10894 );
nor U10955 ( n11185, n15133, n10895 );
nor U10956 ( n11183, n11187, n11188 );
nor U10957 ( n11188, n15149, n10898 );
nor U10958 ( n11187, n15157, n10899 );
nor U10959 ( n11173, n11189, n11190 );
nand U10960 ( n11190, n11191, n11192 );
nor U10961 ( n11192, n11193, n11194 );
nor U10962 ( n11194, n15077, n10906 );
nor U10963 ( n11193, n15069, n10907 );
nor U10964 ( n11191, n11195, n11196 );
nor U10965 ( n11196, n15085, n10910 );
nor U10966 ( n11195, n15093, n10911 );
nand U10967 ( n11189, n11197, n11198 );
nor U10968 ( n11198, n11199, n11200 );
nor U10969 ( n11200, n15109, n10916 );
nor U10970 ( n11199, n15101, n10917 );
nor U10971 ( n11197, n11201, n11202 );
nor U10972 ( n11202, n15117, n10920 );
nor U10973 ( n11201, n15125, n10921 );
nand U10974 ( n11168, n9637, n10188 );
not U10975 ( n9637, n11203 );
nand U10976 ( n11148, n11204, n11205 );
nor U10977 ( n11204, n11206, n11207 );
not U10978 ( n11206, n11208 );
nor U10979 ( n11155, n11203, n11209 );
nand U10980 ( n11203, n11093, n11210 );
nand U10981 ( n11210, n15251, n11211 );
nand U10982 ( n11211, n11212, n7848 );
nand U10983 ( n11093, n11213, n11212 );
nor U10984 ( n11213, n15015, n15251 );
nor U10985 ( n11153, n11214, n11215 );
nor U10986 ( n11215, n15251, n10854 );
nor U10987 ( n11214, n15344, n10855 );
nand U10988 ( n1515, n11216, n11217 );
nor U10989 ( n11217, n11218, n11219 );
nand U10990 ( n11219, n11220, n11221 );
nand U10991 ( n11221, n10835, n9663 );
xor U10992 ( n9663, n11222, n11207 );
xor U10993 ( n11207, n11223, n8082 );
nand U10994 ( n11223, n11224, n11225 );
nor U10995 ( n11225, n11226, n11227 );
nor U10996 ( n11227, n15015, n10975 );
nor U10997 ( n11226, n8082, n11228 );
nor U10998 ( n11224, n11229, n11230 );
nand U10999 ( n11230, n11231, n11232 );
nand U11000 ( n11232, n11233, n11172 );
nor U11001 ( n11233, n10939, n11144 );
nand U11002 ( n11231, n11144, n11143 );
not U11003 ( n11143, n11172 );
and U11004 ( n11144, n11234, n11235 );
nor U11005 ( n11235, n11236, n11237 );
nand U11006 ( n11237, n11238, n11239 );
nor U11007 ( n11239, n11240, n11241 );
nor U11008 ( n11241, n15174, n10884 );
nor U11009 ( n11240, n15166, n10885 );
nor U11010 ( n11238, n11242, n11243 );
nor U11011 ( n11243, n15182, n10888 );
nor U11012 ( n11242, n15190, n10889 );
nand U11013 ( n11236, n11244, n11245 );
nor U11014 ( n11245, n11246, n11247 );
nor U11015 ( n11247, n15142, n10894 );
nor U11016 ( n11246, n15134, n10895 );
nor U11017 ( n11244, n11248, n11249 );
nor U11018 ( n11249, n15150, n10898 );
nor U11019 ( n11248, n15158, n10899 );
nor U11020 ( n11234, n11250, n11251 );
nand U11021 ( n11251, n11252, n11253 );
nor U11022 ( n11253, n11254, n11255 );
nor U11023 ( n11255, n15078, n10906 );
nor U11024 ( n11254, n15070, n10907 );
nor U11025 ( n11252, n11256, n11257 );
nor U11026 ( n11257, n15086, n10910 );
nor U11027 ( n11256, n15094, n10911 );
nand U11028 ( n11250, n11258, n11259 );
nor U11029 ( n11259, n11260, n11261 );
nor U11030 ( n11261, n15110, n10916 );
nor U11031 ( n11260, n15102, n10917 );
nor U11032 ( n11258, n11262, n11263 );
nor U11033 ( n11263, n15118, n10920 );
nor U11034 ( n11262, n15126, n10921 );
nor U11035 ( n11229, n15312, n10843 );
nand U11036 ( n11222, n11205, n11208 );
nand U11037 ( n11220, n10847, n9657 );
not U11038 ( n9657, n11228 );
xnor U11039 ( n11228, n7848, n11212 );
not U11040 ( n11212, n11264 );
nor U11041 ( n11218, n10851, n11265 );
nor U11042 ( n11216, n11266, n11267 );
nor U11043 ( n11267, n15015, n10854 );
nor U11044 ( n11266, n15343, n10855 );
nand U11045 ( n1510, n11268, n11269 );
nor U11046 ( n11269, n11270, n11271 );
nand U11047 ( n11271, n11272, n11273 );
nand U11048 ( n11273, n11274, n11160 );
and U11049 ( n11274, n11275, n11276 );
nand U11050 ( n11272, n10835, n9682 );
xor U11051 ( n9682, n11205, n11208 );
xor U11052 ( n11208, n8082, n11277 );
nor U11053 ( n11277, n11278, n11279 );
nand U11054 ( n11279, n11280, n11281 );
nand U11055 ( n11281, n10842, n8020 );
nand U11056 ( n11280, n10867, n8042 );
nand U11057 ( n11278, n11282, n11283 );
nand U11058 ( n11283, n11284, n11172 );
nand U11059 ( n11172, n11285, n11286 );
and U11060 ( n11285, n10871, n11287 );
nor U11061 ( n11284, n11288, n10939 );
nor U11062 ( n11288, n11286, n11287 );
nand U11063 ( n11287, n11289, n11290 );
nor U11064 ( n11290, n11291, n11292 );
nand U11065 ( n11292, n11293, n11294 );
nor U11066 ( n11294, n11295, n11296 );
nor U11067 ( n11296, n15120, n11297 );
nor U11068 ( n11295, n15112, n11298 );
nor U11069 ( n11293, n11299, n11300 );
nor U11070 ( n11300, n15096, n11301 );
nor U11071 ( n11299, n15104, n11302 );
nand U11072 ( n11291, n11303, n11304 );
nor U11073 ( n11304, n11305, n11306 );
nor U11074 ( n11306, n15088, n11307 );
nor U11075 ( n11305, n15080, n11308 );
nor U11076 ( n11303, n11309, n11310 );
nor U11077 ( n11310, n15064, n11311 );
nor U11078 ( n11309, n15072, n11312 );
nor U11079 ( n11289, n11313, n11314 );
nand U11080 ( n11314, n11315, n11316 );
nor U11081 ( n11316, n11317, n11318 );
nor U11082 ( n11318, n15152, n11319 );
nor U11083 ( n11317, n15144, n11320 );
nor U11084 ( n11315, n11321, n11322 );
nor U11085 ( n11322, n15128, n11323 );
nor U11086 ( n11321, n15136, n11324 );
nand U11087 ( n11313, n11325, n11326 );
nor U11088 ( n11326, n11327, n11328 );
nor U11089 ( n11328, n15184, n11329 );
nor U11090 ( n11327, n15176, n11330 );
nor U11091 ( n11325, n11331, n11332 );
nor U11092 ( n11332, n15160, n11333 );
nor U11093 ( n11331, n15168, n11334 );
nand U11094 ( n11286, n11335, n11336 );
nor U11095 ( n11336, n11337, n11338 );
nand U11096 ( n11338, n11339, n11340 );
nor U11097 ( n11340, n11341, n11342 );
nor U11098 ( n11342, n15111, n10916 );
nand U11099 ( n10916, n11343, n11344 );
nor U11100 ( n11341, n15103, n10917 );
nand U11101 ( n10917, n11343, n11345 );
nor U11102 ( n11339, n11346, n11347 );
nor U11103 ( n11347, n15119, n10920 );
nand U11104 ( n10920, n11343, n11348 );
nor U11105 ( n11346, n15127, n10921 );
nand U11106 ( n10921, n11343, n11349 );
nor U11107 ( n11343, n15194, n11350 );
nand U11108 ( n11337, n11351, n11352 );
nor U11109 ( n11352, n11353, n11354 );
nor U11110 ( n11354, n15079, n10906 );
nand U11111 ( n10906, n11355, n11344 );
nor U11112 ( n11353, n15071, n10907 );
nand U11113 ( n10907, n11355, n11345 );
nor U11114 ( n11351, n11356, n11357 );
nor U11115 ( n11357, n15087, n10910 );
nand U11116 ( n10910, n11355, n11348 );
nor U11117 ( n11355, n7800, n11350 );
nor U11118 ( n11356, n15095, n10911 );
nand U11119 ( n10911, n11358, n11359 );
nor U11120 ( n11335, n11360, n11361 );
nand U11121 ( n11361, n11362, n11363 );
nor U11122 ( n11363, n11364, n11365 );
nor U11123 ( n11365, n15143, n10894 );
nand U11124 ( n10894, n11366, n11344 );
nor U11125 ( n11364, n15135, n10895 );
nand U11126 ( n10895, n11366, n11345 );
nor U11127 ( n11362, n11367, n11368 );
nor U11128 ( n11368, n15151, n10898 );
nand U11129 ( n10898, n11366, n11348 );
nor U11130 ( n11366, n11359, n7800 );
nor U11131 ( n11367, n15159, n10899 );
nand U11132 ( n10899, n11350, n11358 );
not U11133 ( n11350, n11359 );
nand U11134 ( n11360, n11369, n11370 );
nor U11135 ( n11370, n11371, n11372 );
nor U11136 ( n11372, n15175, n10884 );
nand U11137 ( n10884, n11373, n11344 );
nor U11138 ( n11371, n15167, n10885 );
nand U11139 ( n10885, n11373, n11345 );
nor U11140 ( n11369, n11374, n11375 );
nor U11141 ( n11375, n15183, n10888 );
nand U11142 ( n10888, n11373, n11348 );
nor U11143 ( n11374, n15191, n10889 );
nand U11144 ( n10889, n11373, n11349 );
nor U11145 ( n11373, n11359, n15194 );
nand U11146 ( n11359, n11376, n11377 );
nand U11147 ( n11282, n9676, n10188 );
not U11148 ( n9676, n11378 );
nor U11149 ( n11205, n11379, n11380 );
nor U11150 ( n11270, n11378, n11209 );
nand U11151 ( n11378, n11264, n11381 );
nand U11152 ( n11381, n15250, n11382 );
nand U11153 ( n11382, n11383, n7921 );
nand U11154 ( n11264, n11384, n11383 );
not U11155 ( n11383, n11385 );
nor U11156 ( n11384, n15249, n15250 );
nor U11157 ( n11268, n11386, n11387 );
nor U11158 ( n11387, n15250, n10854 );
nor U11159 ( n11386, n15342, n10855 );
nand U11160 ( n1505, n11388, n11389 );
nor U11161 ( n11389, n11390, n11391 );
nand U11162 ( n11391, n11392, n11393 );
nand U11163 ( n11393, n10835, n9702 );
xor U11164 ( n9702, n11379, n11380 );
xnor U11165 ( n11380, n11394, n10188 );
nand U11166 ( n11394, n11395, n11396 );
nor U11167 ( n11396, n11397, n11398 );
nor U11168 ( n11398, n8082, n11399 );
nor U11169 ( n11397, n11400, n10939 );
nor U11170 ( n11400, n11401, n11402 );
nand U11171 ( n11402, n11403, n11404 );
nor U11172 ( n11404, n11405, n11406 );
nand U11173 ( n11406, n11407, n11408 );
nand U11174 ( n11408, n11409, n7924 );
nand U11175 ( n11407, n11410, n7865 );
nand U11176 ( n11405, n11411, n11412 );
nand U11177 ( n11412, n11413, n7925 );
nand U11178 ( n11411, n11414, n7926 );
nor U11179 ( n11403, n11415, n11416 );
nand U11180 ( n11416, n11417, n11418 );
nand U11181 ( n11418, n11419, n7927 );
nand U11182 ( n11417, n11420, n7928 );
nand U11183 ( n11415, n11421, n11422 );
nand U11184 ( n11422, n11423, n7929 );
nand U11185 ( n11421, n11424, n7930 );
nand U11186 ( n11401, n11425, n11426 );
nor U11187 ( n11426, n11427, n11428 );
nand U11188 ( n11428, n11429, n11430 );
nand U11189 ( n11430, n11431, n7931 );
or U11190 ( n11429, n11319, n15153 );
nand U11191 ( n11427, n11432, n11433 );
nand U11192 ( n11433, n11434, n7932 );
nand U11193 ( n11432, n11435, n7933 );
nor U11194 ( n11425, n11436, n11437 );
nand U11195 ( n11437, n11438, n11439 );
nand U11196 ( n11439, n11440, n8001 );
nand U11197 ( n11438, n11441, n7858 );
nand U11198 ( n11436, n11442, n11443 );
nand U11199 ( n11443, n11444, n8008 );
or U11200 ( n11442, n11333, n15161 );
nor U11201 ( n11395, n11445, n11446 );
nor U11202 ( n11446, n15310, n10843 );
nor U11203 ( n11445, n15249, n10975 );
nand U11204 ( n11392, n10847, n9696 );
not U11205 ( n9696, n11399 );
xnor U11206 ( n11399, n11385, n15249 );
nor U11207 ( n11390, n10851, n11447 );
nor U11208 ( n11388, n11448, n11449 );
nor U11209 ( n11449, n15249, n10854 );
nor U11210 ( n11448, n15341, n10855 );
nand U11211 ( n1500, n11450, n11451 );
nor U11212 ( n11451, n11452, n11453 );
nand U11213 ( n11453, n11454, n11455 );
nand U11214 ( n11455, n10835, n9722 );
not U11215 ( n9722, n10257 );
nand U11216 ( n10257, n11379, n11456 );
nand U11217 ( n11456, n11457, n11458 );
or U11218 ( n11379, n11458, n11457 );
xnor U11219 ( n11457, n11459, n10188 );
nand U11220 ( n11459, n11460, n11461 );
nor U11221 ( n11461, n11462, n11463 );
nor U11222 ( n11463, n8082, n11464 );
nor U11223 ( n11462, n11465, n10939 );
nor U11224 ( n11465, n11466, n11467 );
nand U11225 ( n11467, n11468, n11469 );
nor U11226 ( n11469, n11470, n11471 );
nand U11227 ( n11471, n11472, n11473 );
nand U11228 ( n11473, n11409, n7934 );
nand U11229 ( n11472, n11410, n7866 );
nand U11230 ( n11470, n11474, n11475 );
nand U11231 ( n11475, n11413, n7935 );
nand U11232 ( n11474, n11414, n7936 );
nor U11233 ( n11468, n11476, n11477 );
nand U11234 ( n11477, n11478, n11479 );
nand U11235 ( n11479, n11419, n7937 );
nand U11236 ( n11478, n11420, n7938 );
nand U11237 ( n11476, n11480, n11481 );
nand U11238 ( n11481, n11423, n7939 );
nand U11239 ( n11480, n11424, n7940 );
nand U11240 ( n11466, n11482, n11483 );
nor U11241 ( n11483, n11484, n11485 );
nand U11242 ( n11485, n11486, n11487 );
nand U11243 ( n11487, n11431, n7941 );
or U11244 ( n11486, n11319, n15154 );
nand U11245 ( n11484, n11488, n11489 );
nand U11246 ( n11489, n11434, n7942 );
nand U11247 ( n11488, n11435, n7943 );
nor U11248 ( n11482, n11490, n11491 );
nand U11249 ( n11491, n11492, n11493 );
nand U11250 ( n11493, n11440, n8000 );
nand U11251 ( n11492, n11441, n7857 );
nand U11252 ( n11490, n11494, n11495 );
nand U11253 ( n11495, n11444, n8007 );
or U11254 ( n11494, n11333, n15162 );
nor U11255 ( n11460, n11496, n11497 );
nor U11256 ( n11497, n15309, n10843 );
nor U11257 ( n11496, n15248, n10975 );
nand U11258 ( n11458, n11498, n11499 );
nand U11259 ( n11454, n10847, n9716 );
not U11260 ( n9716, n11464 );
nand U11261 ( n11464, n11385, n11500 );
nand U11262 ( n11500, n15248, n11501 );
nand U11263 ( n11501, n11502, n7849 );
nand U11264 ( n11385, n11503, n11502 );
nor U11265 ( n11503, n15247, n15248 );
nor U11266 ( n11452, n10851, n11504 );
nor U11267 ( n11450, n11505, n11506 );
nor U11268 ( n11506, n15248, n10854 );
nor U11269 ( n11505, n15340, n10855 );
nand U11270 ( n1495, n11507, n11508 );
nor U11271 ( n11508, n11509, n11510 );
nand U11272 ( n11510, n11511, n11512 );
nand U11273 ( n11512, n10835, n9743 );
xor U11274 ( n9743, n11498, n11499 );
xnor U11275 ( n11499, n11513, n8082 );
nand U11276 ( n11513, n11514, n11515 );
nor U11277 ( n11515, n11516, n11517 );
and U11278 ( n11517, n10188, n9737 );
nor U11279 ( n11516, n11518, n10939 );
nor U11280 ( n11518, n11519, n11520 );
nand U11281 ( n11520, n11521, n11522 );
nor U11282 ( n11522, n11523, n11524 );
nand U11283 ( n11524, n11525, n11526 );
nand U11284 ( n11526, n11409, n7944 );
nand U11285 ( n11525, n11410, n7867 );
nand U11286 ( n11523, n11527, n11528 );
nand U11287 ( n11528, n11413, n7945 );
nand U11288 ( n11527, n11414, n7946 );
nor U11289 ( n11521, n11529, n11530 );
nand U11290 ( n11530, n11531, n11532 );
nand U11291 ( n11532, n11419, n7947 );
nand U11292 ( n11531, n11420, n7948 );
nand U11293 ( n11529, n11533, n11534 );
nand U11294 ( n11534, n11423, n7949 );
nand U11295 ( n11533, n11424, n7950 );
nand U11296 ( n11519, n11535, n11536 );
nor U11297 ( n11536, n11537, n11538 );
nand U11298 ( n11538, n11539, n11540 );
nand U11299 ( n11540, n11431, n7951 );
or U11300 ( n11539, n11319, n15155 );
nand U11301 ( n11537, n11541, n11542 );
nand U11302 ( n11542, n11434, n7952 );
nand U11303 ( n11541, n11435, n7953 );
nor U11304 ( n11535, n11543, n11544 );
nand U11305 ( n11544, n11545, n11546 );
nand U11306 ( n11546, n11440, n7999 );
nand U11307 ( n11545, n11441, n7856 );
nand U11308 ( n11543, n11547, n11548 );
nand U11309 ( n11548, n11444, n8006 );
nand U11310 ( n11547, n11549, n8013 );
nor U11311 ( n11514, n11550, n11551 );
nor U11312 ( n11551, n15308, n10843 );
nor U11313 ( n11550, n15247, n10975 );
nor U11314 ( n11498, n11552, n11553 );
nand U11315 ( n11511, n10847, n9737 );
xor U11316 ( n9737, n7849, n11502 );
and U11317 ( n11502, n11554, n11555 );
nor U11318 ( n11554, n15245, n15246 );
nor U11319 ( n11509, n10851, n11556 );
nor U11320 ( n11507, n11557, n11558 );
nor U11321 ( n11558, n15247, n10854 );
nor U11322 ( n11557, n15339, n10855 );
nand U11323 ( n1490, n11559, n11560 );
nor U11324 ( n11560, n11561, n11562 );
nand U11325 ( n11562, n11563, n11564 );
nand U11326 ( n11564, n10835, n9765 );
xor U11327 ( n9765, n11552, n11553 );
xnor U11328 ( n11553, n11565, n10188 );
nand U11329 ( n11565, n11566, n11567 );
nor U11330 ( n11567, n11568, n11569 );
and U11331 ( n11569, n10188, n9757 );
nor U11332 ( n11568, n11570, n10939 );
nor U11333 ( n11570, n11571, n11572 );
nand U11334 ( n11572, n11573, n11574 );
nor U11335 ( n11574, n11575, n11576 );
nand U11336 ( n11576, n11577, n11578 );
nand U11337 ( n11578, n11409, n7954 );
nand U11338 ( n11577, n11410, n7868 );
nand U11339 ( n11575, n11579, n11580 );
nand U11340 ( n11580, n11413, n7955 );
nand U11341 ( n11579, n11414, n7956 );
nor U11342 ( n11573, n11581, n11582 );
nand U11343 ( n11582, n11583, n11584 );
nand U11344 ( n11584, n11419, n7957 );
nand U11345 ( n11583, n11420, n7958 );
nand U11346 ( n11581, n11585, n11586 );
nand U11347 ( n11586, n11423, n7959 );
nand U11348 ( n11585, n11424, n7960 );
nand U11349 ( n11571, n11587, n11588 );
nor U11350 ( n11588, n11589, n11590 );
nand U11351 ( n11590, n11591, n11592 );
nand U11352 ( n11592, n11431, n7961 );
or U11353 ( n11591, n11319, n15156 );
nand U11354 ( n11589, n11593, n11594 );
nand U11355 ( n11594, n11434, n7962 );
nand U11356 ( n11593, n11435, n7963 );
nor U11357 ( n11587, n11595, n11596 );
nand U11358 ( n11596, n11597, n11598 );
nand U11359 ( n11598, n11440, n7998 );
nand U11360 ( n11597, n11441, n7918 );
nand U11361 ( n11595, n11599, n11600 );
nand U11362 ( n11600, n11444, n8005 );
nand U11363 ( n11599, n11549, n8012 );
nor U11364 ( n11566, n11601, n11602 );
nor U11365 ( n11602, n15307, n10843 );
nor U11366 ( n11601, n15246, n10975 );
nand U11367 ( n11552, n11603, n11604 );
nand U11368 ( n11563, n10847, n9757 );
xnor U11369 ( n9757, n15246, n11605 );
and U11370 ( n11605, n8044, n11555 );
nor U11371 ( n11561, n11606, n10851 );
nor U11372 ( n11559, n11607, n11608 );
nor U11373 ( n11608, n15246, n10854 );
nor U11374 ( n11607, n15338, n10855 );
nand U11375 ( n1485, n11609, n11610 );
nor U11376 ( n11610, n11611, n11612 );
nand U11377 ( n11612, n11613, n11614 );
nand U11378 ( n11614, n10835, n9786 );
xor U11379 ( n9786, n11603, n11604 );
xnor U11380 ( n11604, n11615, n8082 );
nand U11381 ( n11615, n11616, n11617 );
nor U11382 ( n11617, n11618, n11619 );
and U11383 ( n11619, n10188, n9779 );
nor U11384 ( n11618, n11620, n10939 );
nor U11385 ( n11620, n11621, n11622 );
nand U11386 ( n11622, n11623, n11624 );
nor U11387 ( n11624, n11625, n11626 );
nand U11388 ( n11626, n11627, n11628 );
nand U11389 ( n11628, n11409, n7964 );
nand U11390 ( n11627, n11410, n7869 );
nand U11391 ( n11625, n11629, n11630 );
nand U11392 ( n11630, n11413, n7965 );
nand U11393 ( n11629, n11414, n7966 );
nor U11394 ( n11623, n11631, n11632 );
nand U11395 ( n11632, n11633, n11634 );
nand U11396 ( n11634, n11419, n7967 );
nand U11397 ( n11633, n11420, n7968 );
nand U11398 ( n11631, n11635, n11636 );
nand U11399 ( n11636, n11423, n7969 );
nand U11400 ( n11635, n11424, n7970 );
nand U11401 ( n11621, n11637, n11638 );
nor U11402 ( n11638, n11639, n11640 );
nand U11403 ( n11640, n11641, n11642 );
nand U11404 ( n11642, n11431, n7971 );
or U11405 ( n11641, n11319, n15157 );
nand U11406 ( n11639, n11643, n11644 );
nand U11407 ( n11644, n11434, n7972 );
nand U11408 ( n11643, n11435, n7973 );
nor U11409 ( n11637, n11645, n11646 );
nand U11410 ( n11646, n11647, n11648 );
nand U11411 ( n11648, n11440, n7997 );
nand U11412 ( n11647, n11441, n7859 );
nand U11413 ( n11645, n11649, n11650 );
nand U11414 ( n11650, n11444, n8004 );
nand U11415 ( n11649, n11549, n8011 );
nor U11416 ( n11616, n11651, n11652 );
nor U11417 ( n11652, n15306, n10843 );
nor U11418 ( n11651, n15245, n10975 );
nor U11419 ( n11603, n11653, n11654 );
nand U11420 ( n11613, n10847, n9779 );
xnor U11421 ( n9779, n11555, n15245 );
nor U11422 ( n11555, n11655, n15244 );
nor U11423 ( n11611, n11656, n10851 );
nor U11424 ( n11609, n11657, n11658 );
nor U11425 ( n11658, n15245, n10854 );
nor U11426 ( n11657, n15337, n10855 );
nand U11427 ( n1480, n11659, n11660 );
nor U11428 ( n11660, n11661, n11662 );
nand U11429 ( n11662, n11663, n11664 );
nand U11430 ( n11664, n10835, n9806 );
xor U11431 ( n9806, n11653, n11654 );
xnor U11432 ( n11654, n11665, n10188 );
nand U11433 ( n11665, n11666, n11667 );
nor U11434 ( n11667, n11668, n11669 );
and U11435 ( n11669, n10188, n9799 );
nor U11436 ( n11668, n11670, n10939 );
nor U11437 ( n11670, n11671, n11672 );
nand U11438 ( n11672, n11673, n11674 );
nor U11439 ( n11674, n11675, n11676 );
nand U11440 ( n11676, n11677, n11678 );
nand U11441 ( n11678, n11409, n7974 );
nand U11442 ( n11677, n11410, n7870 );
nand U11443 ( n11675, n11679, n11680 );
nand U11444 ( n11680, n11413, n7975 );
nand U11445 ( n11679, n11414, n7976 );
nor U11446 ( n11673, n11681, n11682 );
nand U11447 ( n11682, n11683, n11684 );
nand U11448 ( n11684, n11419, n7977 );
nand U11449 ( n11683, n11420, n7978 );
nand U11450 ( n11681, n11685, n11686 );
nand U11451 ( n11686, n11423, n7979 );
nand U11452 ( n11685, n11424, n7980 );
nand U11453 ( n11671, n11687, n11688 );
nor U11454 ( n11688, n11689, n11690 );
nand U11455 ( n11690, n11691, n11692 );
nand U11456 ( n11692, n11431, n7981 );
or U11457 ( n11691, n11319, n15158 );
nand U11458 ( n11689, n11693, n11694 );
nand U11459 ( n11694, n11434, n7982 );
nand U11460 ( n11693, n11435, n7983 );
nor U11461 ( n11687, n11695, n11696 );
nand U11462 ( n11696, n11697, n11698 );
nand U11463 ( n11698, n11440, n7996 );
nand U11464 ( n11697, n11441, n7917 );
nand U11465 ( n11695, n11699, n11700 );
nand U11466 ( n11700, n11444, n8003 );
nand U11467 ( n11699, n11549, n8010 );
nor U11468 ( n11666, n11701, n11702 );
nor U11469 ( n11702, n15305, n10843 );
nor U11470 ( n11701, n15244, n10975 );
nand U11471 ( n11663, n10847, n9799 );
xor U11472 ( n9799, n15244, n11655 );
nor U11473 ( n11661, n11703, n10851 );
nor U11474 ( n11659, n11704, n11705 );
nor U11475 ( n11705, n15244, n10854 );
nor U11476 ( n11704, n15336, n10855 );
nand U11477 ( n1475, n11706, n11707 );
nor U11478 ( n11707, n11708, n11709 );
nand U11479 ( n11709, n11710, n11711 );
nand U11480 ( n11711, n11712, n11160 );
and U11481 ( n11712, n11713, n11714 );
nand U11482 ( n11710, n10835, n9828 );
not U11483 ( n9828, n10282 );
nand U11484 ( n10282, n11653, n11715 );
nand U11485 ( n11715, n11716, n11717 );
or U11486 ( n11653, n11717, n11716 );
xnor U11487 ( n11716, n11718, n10188 );
nand U11488 ( n11718, n11719, n11720 );
nor U11489 ( n11720, n11721, n11722 );
nor U11490 ( n11722, n8082, n9821 );
nor U11491 ( n11721, n11723, n10939 );
not U11492 ( n10939, n10871 );
nand U11493 ( n10871, n11724, n11725 );
nand U11494 ( n11725, n11726, n7814 );
nand U11495 ( n11724, n11727, n10562 );
nor U11496 ( n11723, n11728, n11729 );
nand U11497 ( n11729, n11730, n11731 );
nor U11498 ( n11731, n11732, n11733 );
nand U11499 ( n11733, n11734, n11735 );
nand U11500 ( n11735, n11409, n7984 );
not U11501 ( n11409, n11298 );
nand U11502 ( n11298, n11736, n11737 );
nand U11503 ( n11734, n11410, n7871 );
not U11504 ( n11410, n11297 );
nand U11505 ( n11297, n11736, n11738 );
nand U11506 ( n11732, n11739, n11740 );
nand U11507 ( n11740, n11413, n7985 );
not U11508 ( n11413, n11302 );
nand U11509 ( n11302, n11736, n11741 );
nand U11510 ( n11739, n11414, n7986 );
not U11511 ( n11414, n11301 );
nand U11512 ( n11301, n11736, n11742 );
and U11513 ( n11736, n11743, n11744 );
nor U11514 ( n11730, n11745, n11746 );
nand U11515 ( n11746, n11747, n11748 );
nand U11516 ( n11748, n11419, n7987 );
not U11517 ( n11419, n11308 );
nand U11518 ( n11308, n11749, n11737 );
nand U11519 ( n11747, n11420, n7988 );
not U11520 ( n11420, n11307 );
nand U11521 ( n11307, n11749, n11738 );
nand U11522 ( n11745, n11750, n11751 );
nand U11523 ( n11751, n11423, n7989 );
not U11524 ( n11423, n11312 );
nand U11525 ( n11312, n11749, n11741 );
nand U11526 ( n11750, n11424, n7990 );
not U11527 ( n11424, n11311 );
nand U11528 ( n11311, n11749, n11742 );
and U11529 ( n11749, n11752, n11744 );
nand U11530 ( n11728, n11753, n11754 );
nor U11531 ( n11754, n11755, n11756 );
nand U11532 ( n11756, n11757, n11758 );
nand U11533 ( n11758, n11431, n7991 );
not U11534 ( n11431, n11320 );
nand U11535 ( n11320, n11759, n11737 );
or U11536 ( n11757, n11319, n15159 );
nand U11537 ( n11319, n11759, n11738 );
nand U11538 ( n11755, n11760, n11761 );
nand U11539 ( n11761, n11434, n7992 );
not U11540 ( n11434, n11324 );
nand U11541 ( n11324, n11759, n11741 );
nand U11542 ( n11760, n11435, n7993 );
not U11543 ( n11435, n11323 );
nand U11544 ( n11323, n11759, n11742 );
nor U11545 ( n11759, n11743, n11744 );
not U11546 ( n11743, n11752 );
nor U11547 ( n11753, n11762, n11763 );
nand U11548 ( n11763, n11764, n11765 );
nand U11549 ( n11765, n11440, n7995 );
not U11550 ( n11440, n11330 );
nand U11551 ( n11330, n11766, n11737 );
nand U11552 ( n11764, n11441, n7916 );
not U11553 ( n11441, n11329 );
nand U11554 ( n11329, n11766, n11738 );
nand U11555 ( n11762, n11767, n11768 );
nand U11556 ( n11768, n11444, n8002 );
not U11557 ( n11444, n11334 );
nand U11558 ( n11334, n11766, n11741 );
nand U11559 ( n11767, n11549, n8009 );
not U11560 ( n11549, n11333 );
nand U11561 ( n11333, n11766, n11742 );
nor U11562 ( n11766, n11744, n11752 );
nor U11563 ( n11752, n11769, n11358 );
nor U11564 ( n11769, n15194, n11349 );
nand U11565 ( n11744, n11770, n11377 );
nor U11566 ( n11770, n11771, n11772 );
nor U11567 ( n11772, n11349, n11376 );
nor U11568 ( n11771, n15193, n11773 );
nor U11569 ( n11719, n11774, n11775 );
nor U11570 ( n11775, n15304, n10843 );
nor U11571 ( n11774, n15243, n10975 );
nor U11572 ( n11708, n9821, n11209 );
nand U11573 ( n9821, n11655, n11776 );
nand U11574 ( n11776, n15243, n11777 );
or U11575 ( n11655, n11777, n15243 );
nor U11576 ( n11706, n11778, n11779 );
nor U11577 ( n11779, n15243, n10854 );
nor U11578 ( n11778, n15335, n10855 );
nand U11579 ( n1470, n11780, n11781 );
nor U11580 ( n11781, n11782, n11783 );
nand U11581 ( n11783, n11784, n11785 );
nand U11582 ( n11785, n10835, n9849 );
not U11583 ( n9849, n10287 );
nand U11584 ( n10287, n11717, n11786 );
nand U11585 ( n11786, n11787, n11788 );
nand U11586 ( n11788, n11789, n11790 );
not U11587 ( n11787, n11791 );
nand U11588 ( n11717, n11792, n11791 );
nand U11589 ( n11791, n11793, n11794 );
nand U11590 ( n11794, n11795, n11796 );
xor U11591 ( n11793, n10188, n11797 );
nor U11592 ( n11797, n11798, n11799 );
nand U11593 ( n11799, n11800, n11801 );
nand U11594 ( n11801, n9842, n10188 );
nand U11595 ( n11800, n10842, n8021 );
nor U11596 ( n11798, n15303, n10843 );
and U11597 ( n11792, n11789, n11790 );
nand U11598 ( n11784, n10847, n9842 );
and U11599 ( n9842, n11777, n11802 );
nand U11600 ( n11802, n15242, n11803 );
nand U11601 ( n11803, n11804, n7836 );
nand U11602 ( n11777, n11805, n11804 );
nor U11603 ( n11805, n15241, n15242 );
nor U11604 ( n11782, n10851, n11806 );
nor U11605 ( n11780, n11807, n11808 );
nor U11606 ( n11808, n15242, n10854 );
nor U11607 ( n11807, n15334, n10855 );
nand U11608 ( n1465, n11809, n11810 );
nor U11609 ( n11810, n11811, n11812 );
nand U11610 ( n11812, n11813, n11814 );
nand U11611 ( n11814, n10835, n9869 );
not U11612 ( n9869, n10292 );
xnor U11613 ( n10292, n11789, n11790 );
nand U11614 ( n11790, n11815, n11816 );
nand U11615 ( n11816, n11817, n11818 );
nand U11616 ( n11789, n11819, n11820 );
nand U11617 ( n11820, n11821, n11796 );
xor U11618 ( n11819, n10188, n11822 );
nor U11619 ( n11822, n11823, n11824 );
nand U11620 ( n11824, n11825, n11826 );
nand U11621 ( n11826, n9862, n10188 );
nand U11622 ( n11825, n10842, n7836 );
nor U11623 ( n11823, n15302, n10843 );
nand U11624 ( n11813, n10847, n9862 );
xor U11625 ( n9862, n7836, n11804 );
nor U11626 ( n11804, n11827, n11828 );
nand U11627 ( n11827, n7863, n7809 );
nor U11628 ( n11811, n10851, n11829 );
nor U11629 ( n11809, n11830, n11831 );
nor U11630 ( n11831, n15241, n10854 );
nor U11631 ( n11830, n15333, n10855 );
nand U11632 ( n1460, n11832, n11833 );
nor U11633 ( n11833, n11834, n11835 );
nand U11634 ( n11835, n11836, n11837 );
nand U11635 ( n11837, n10835, n9890 );
xor U11636 ( n9890, n11818, n11838 );
nor U11637 ( n11838, n11839, n11840 );
not U11638 ( n11840, n11815 );
nand U11639 ( n11815, n11841, n11842 );
and U11640 ( n11841, n11796, n11817 );
nor U11641 ( n11839, n11817, n11843 );
nor U11642 ( n11843, n11844, n11845 );
and U11643 ( n11817, n11846, n11847 );
xor U11644 ( n11818, n8082, n11848 );
nor U11645 ( n11848, n11849, n11850 );
nand U11646 ( n11850, n11851, n11852 );
nand U11647 ( n11852, n9883, n10188 );
nand U11648 ( n11851, n10842, n7809 );
nor U11649 ( n11849, n15301, n10843 );
nand U11650 ( n11836, n10847, n9883 );
xor U11651 ( n9883, n7809, n11853 );
nor U11652 ( n11853, n15016, n11828 );
nor U11653 ( n11834, n10851, n11854 );
nor U11654 ( n11832, n11855, n11856 );
nor U11655 ( n11856, n15240, n10854 );
nor U11656 ( n11855, n15332, n10855 );
nand U11657 ( n1455, n11857, n11858 );
nor U11658 ( n11858, n11859, n11860 );
nand U11659 ( n11860, n11861, n11862 );
nand U11660 ( n11862, n10835, n9913 );
not U11661 ( n9913, n10302 );
xnor U11662 ( n10302, n11846, n11847 );
nand U11663 ( n11847, n11863, n11864 );
nand U11664 ( n11864, n11865, n11796 );
xor U11665 ( n11863, n10188, n11866 );
nor U11666 ( n11866, n11867, n11868 );
nand U11667 ( n11868, n11869, n11870 );
nand U11668 ( n11870, n9906, n10188 );
nand U11669 ( n11869, n10842, n7863 );
nor U11670 ( n11867, n15300, n10843 );
nand U11671 ( n11861, n10847, n9906 );
xor U11672 ( n9906, n11828, n15016 );
nand U11673 ( n11828, n11871, n11872 );
nor U11674 ( n11871, n15017, n15239 );
nor U11675 ( n11859, n10851, n11873 );
nor U11676 ( n11857, n11874, n11875 );
nor U11677 ( n11875, n15016, n10854 );
nor U11678 ( n11874, n15331, n10855 );
nand U11679 ( n1450, n11876, n11877 );
nor U11680 ( n11877, n11878, n11879 );
nand U11681 ( n11879, n11880, n11881 );
nand U11682 ( n11881, n10835, n9933 );
nor U11683 ( n9933, n11846, n11882 );
and U11684 ( n11882, n11883, n11884 );
nor U11685 ( n11846, n11884, n11883 );
and U11686 ( n11883, n11885, n11886 );
nand U11687 ( n11886, n11887, n11796 );
xor U11688 ( n11885, n10188, n11888 );
nor U11689 ( n11888, n11889, n11890 );
nand U11690 ( n11890, n11891, n11892 );
nand U11691 ( n11892, n9926, n10188 );
nand U11692 ( n11891, n10842, n8014 );
nor U11693 ( n11889, n15299, n10843 );
nand U11694 ( n11880, n10847, n9926 );
xor U11695 ( n9926, n11893, n15239 );
nand U11696 ( n11893, n11872, n7837 );
nor U11697 ( n11878, n10851, n11894 );
nor U11698 ( n11876, n11895, n11896 );
nor U11699 ( n11896, n15239, n10854 );
nor U11700 ( n11895, n15330, n10855 );
nand U11701 ( n1445, n11897, n11898 );
nor U11702 ( n11898, n11899, n11900 );
nand U11703 ( n11900, n11901, n11902 );
nand U11704 ( n11902, n10835, n9954 );
not U11705 ( n9954, n10312 );
nand U11706 ( n10312, n11903, n11884 );
nand U11707 ( n11884, n11904, n11905 );
nor U11708 ( n11904, n11906, n11907 );
not U11709 ( n11907, n11908 );
nand U11710 ( n11903, n11906, n11909 );
nand U11711 ( n11909, n11905, n11908 );
nand U11712 ( n11908, n11910, n11911 );
nand U11713 ( n11911, n11912, n11796 );
and U11714 ( n11906, n11913, n11914 );
nand U11715 ( n11914, n11915, n11796 );
xor U11716 ( n11913, n10188, n11916 );
nor U11717 ( n11916, n11917, n11918 );
nand U11718 ( n11918, n11919, n11920 );
nand U11719 ( n11920, n9947, n10188 );
nand U11720 ( n11919, n10842, n7837 );
nor U11721 ( n11917, n15298, n10843 );
nand U11722 ( n11901, n10847, n9947 );
xor U11723 ( n9947, n7837, n11872 );
nor U11724 ( n11872, n11921, n11922 );
nand U11725 ( n11921, n7864, n7810 );
nor U11726 ( n11899, n10851, n11923 );
nor U11727 ( n11897, n11924, n11925 );
nor U11728 ( n11925, n15017, n10854 );
nor U11729 ( n11924, n15329, n10855 );
nand U11730 ( n1440, n11926, n11927 );
nor U11731 ( n11927, n11928, n11929 );
nand U11732 ( n11929, n11930, n11931 );
nand U11733 ( n11931, n10835, n9975 );
xor U11734 ( n9975, n11932, n11910 );
xor U11735 ( n11910, n10188, n11933 );
nor U11736 ( n11933, n11934, n11935 );
nand U11737 ( n11935, n11936, n11937 );
nand U11738 ( n11937, n9968, n10188 );
nand U11739 ( n11936, n10842, n7810 );
nor U11740 ( n11934, n15297, n10843 );
xnor U11741 ( n11932, n11905, n11938 );
nor U11742 ( n11938, n11844, n11939 );
and U11743 ( n11905, n11940, n11941 );
nand U11744 ( n11930, n10847, n9968 );
xor U11745 ( n9968, n7810, n11942 );
nor U11746 ( n11942, n15018, n11922 );
nor U11747 ( n11928, n10851, n11943 );
nor U11748 ( n11926, n11944, n11945 );
nor U11749 ( n11945, n15238, n10854 );
nor U11750 ( n11944, n15328, n10855 );
nand U11751 ( n1435, n11946, n11947 );
nor U11752 ( n11947, n11948, n11949 );
nand U11753 ( n11949, n11950, n11951 );
nand U11754 ( n11951, n10835, n9995 );
not U11755 ( n9995, n10322 );
xnor U11756 ( n10322, n11940, n11941 );
nand U11757 ( n11941, n11952, n11953 );
nand U11758 ( n11953, n11954, n11796 );
xor U11759 ( n11952, n10188, n11955 );
nor U11760 ( n11955, n11956, n11957 );
nand U11761 ( n11957, n11958, n11959 );
nand U11762 ( n11959, n9988, n10188 );
nand U11763 ( n11958, n10842, n7864 );
nor U11764 ( n11956, n15296, n10843 );
nand U11765 ( n11950, n10847, n9988 );
xor U11766 ( n9988, n11922, n15018 );
nand U11767 ( n11922, n11960, n11961 );
nor U11768 ( n11960, n15019, n15237 );
nor U11769 ( n11948, n10851, n11962 );
nor U11770 ( n11946, n11963, n11964 );
nor U11771 ( n11964, n15018, n10854 );
nor U11772 ( n11963, n15327, n10855 );
nand U11773 ( n1430, n11965, n11966 );
nor U11774 ( n11966, n11967, n11968 );
nand U11775 ( n11968, n11969, n11970 );
nand U11776 ( n11970, n11971, n11160 );
not U11777 ( n11160, n10851 );
and U11778 ( n11971, n11972, n11973 );
nand U11779 ( n11969, n10835, n10016 );
nor U11780 ( n10016, n11940, n11974 );
and U11781 ( n11974, n11975, n11976 );
nor U11782 ( n11940, n11976, n11975 );
and U11783 ( n11975, n11977, n11978 );
nand U11784 ( n11978, n11979, n11796 );
xor U11785 ( n11977, n10188, n11980 );
nor U11786 ( n11980, n11981, n11982 );
nand U11787 ( n11982, n11983, n11984 );
nand U11788 ( n11984, n10009, n10188 );
nand U11789 ( n11983, n10842, n8015 );
nor U11790 ( n11981, n15295, n10843 );
nand U11791 ( n11976, n11985, n11986 );
nand U11792 ( n11986, n11987, n11988 );
and U11793 ( n11967, n10009, n10847 );
xor U11794 ( n10009, n11989, n15237 );
nand U11795 ( n11989, n11961, n7838 );
nor U11796 ( n11965, n11990, n11991 );
nor U11797 ( n11991, n15237, n10854 );
nor U11798 ( n11990, n15326, n10855 );
nand U11799 ( n1425, n11992, n11993 );
nor U11800 ( n11993, n11994, n11995 );
nand U11801 ( n11995, n11996, n11997 );
nand U11802 ( n11997, n10835, n10037 );
xor U11803 ( n10037, n11998, n11987 );
xor U11804 ( n11987, n10188, n11999 );
nor U11805 ( n11999, n12000, n12001 );
nand U11806 ( n12001, n12002, n12003 );
nand U11807 ( n12003, n10030, n10188 );
nand U11808 ( n12002, n10842, n7838 );
nor U11809 ( n12000, n15294, n10843 );
xor U11810 ( n11998, n11985, n11988 );
or U11811 ( n11988, n11844, n12004 );
nand U11812 ( n11996, n10847, n10030 );
xor U11813 ( n10030, n7838, n11961 );
nor U11814 ( n11961, n12005, n12006 );
nand U11815 ( n12005, n7923, n7811 );
nor U11816 ( n11994, n10851, n12007 );
nor U11817 ( n11992, n12008, n12009 );
nor U11818 ( n12009, n15019, n10854 );
nor U11819 ( n12008, n15325, n10855 );
nand U11820 ( n1420, n12010, n12011 );
nor U11821 ( n12011, n12012, n12013 );
nand U11822 ( n12013, n12014, n12015 );
nand U11823 ( n12015, n10835, n10058 );
nor U11824 ( n10058, n11985, n12016 );
and U11825 ( n12016, n12017, n12018 );
nor U11826 ( n11985, n12018, n12017 );
and U11827 ( n12017, n12019, n12020 );
nand U11828 ( n12020, n12021, n11796 );
xor U11829 ( n12019, n10188, n12022 );
nor U11830 ( n12022, n12023, n12024 );
nand U11831 ( n12024, n12025, n12026 );
nand U11832 ( n12026, n10051, n10188 );
nand U11833 ( n12025, n10842, n7811 );
nor U11834 ( n12023, n15293, n10843 );
nand U11835 ( n12018, n12027, n12028 );
nand U11836 ( n12014, n10847, n10051 );
xor U11837 ( n10051, n7811, n12029 );
nor U11838 ( n12029, n15235, n12006 );
nor U11839 ( n12012, n10851, n12030 );
nor U11840 ( n12010, n12031, n12032 );
nor U11841 ( n12032, n15236, n10854 );
nor U11842 ( n12031, n15324, n10855 );
nand U11843 ( n1415, n12033, n12034 );
nor U11844 ( n12034, n12035, n12036 );
nand U11845 ( n12036, n12037, n12038 );
nand U11846 ( n12038, n10835, n10081 );
xor U11847 ( n10081, n12027, n12028 );
nand U11848 ( n12028, n12039, n12040 );
nand U11849 ( n12040, n12041, n11796 );
xor U11850 ( n12039, n8082, n12042 );
nand U11851 ( n12042, n12043, n12044 );
nor U11852 ( n12044, n12045, n12046 );
nor U11853 ( n12046, n15235, n10975 );
and U11854 ( n12045, n10188, n10074 );
nor U11855 ( n12043, n12047, n12048 );
nor U11856 ( n12048, n15192, n12049 );
nor U11857 ( n12047, n15292, n10843 );
and U11858 ( n12027, n12050, n12051 );
nand U11859 ( n12051, n12052, n12053 );
nand U11860 ( n12052, n12054, n12055 );
nand U11861 ( n12055, n12056, n8082 );
nor U11862 ( n12054, n12057, n12058 );
and U11863 ( n12050, n12059, n12060 );
nand U11864 ( n12037, n10847, n10074 );
xor U11865 ( n10074, n12006, n15235 );
nand U11866 ( n12006, n12061, n7851 );
nor U11867 ( n12035, n10851, n12062 );
nor U11868 ( n12033, n12063, n12064 );
nor U11869 ( n12064, n15235, n10854 );
nor U11870 ( n12063, n15323, n10855 );
nand U11871 ( n1410, n12065, n12066 );
nor U11872 ( n12066, n12067, n12068 );
nand U11873 ( n12068, n12069, n12070 );
nand U11874 ( n12070, n10835, n10108 );
not U11875 ( n10108, n10347 );
xor U11876 ( n10347, n12060, n12071 );
and U11877 ( n12071, n12072, n12053 );
nand U11878 ( n12060, n12073, n12074 );
nand U11879 ( n12074, n11796, n12075 );
xor U11880 ( n12073, n8082, n12076 );
nand U11881 ( n12076, n12077, n12078 );
nor U11882 ( n12078, n12079, n12080 );
nor U11883 ( n12080, n15234, n10975 );
and U11884 ( n12079, n10188, n10102 );
nor U11885 ( n12077, n12081, n12082 );
nor U11886 ( n12082, n15193, n12049 );
nor U11887 ( n12081, n15291, n10843 );
nand U11888 ( n12069, n10847, n10102 );
xor U11889 ( n10102, n7851, n12061 );
nor U11890 ( n12061, n15233, n15232 );
nor U11891 ( n12067, n12083, n10851 );
nor U11892 ( n12065, n12084, n12085 );
nor U11893 ( n12085, n15234, n10854 );
nor U11894 ( n12084, n15322, n10855 );
nand U11895 ( n1405, n12086, n12087 );
nor U11896 ( n12087, n12088, n12089 );
nand U11897 ( n12089, n12090, n12091 );
nand U11898 ( n12091, n10835, n10127 );
not U11899 ( n10127, n10352 );
nand U11900 ( n10352, n12072, n12092 );
nand U11901 ( n12092, n12093, n12094 );
nand U11902 ( n12093, n12053, n12059 );
nand U11903 ( n12053, n10842, n12095 );
nand U11904 ( n12072, n12096, n12059 );
nand U11905 ( n12059, n12097, n12098 );
xor U11906 ( n12098, n8082, n12095 );
nand U11907 ( n12095, n12099, n12100 );
nor U11908 ( n12100, n12101, n12102 );
nor U11909 ( n12102, n15233, n10975 );
and U11910 ( n12101, n10122, n10188 );
nor U11911 ( n12099, n12103, n12104 );
nor U11912 ( n12104, n15194, n12049 );
nor U11913 ( n12103, n15290, n10843 );
nor U11914 ( n12097, n10842, n12105 );
nor U11915 ( n12105, n9077, n11844 );
nand U11916 ( n12090, n10847, n10122 );
xor U11917 ( n10122, n15233, n15232 );
nor U11918 ( n12088, n10851, n12107 );
nor U11919 ( n12086, n12108, n12109 );
nor U11920 ( n12109, n15233, n10854 );
nor U11921 ( n12108, n15321, n10855 );
nand U11922 ( n1400, n12110, n12111 );
nor U11923 ( n12111, n12112, n12113 );
nor U11924 ( n12113, n12114, n10851 );
nor U11925 ( n12112, n10144, n12106 );
nand U11926 ( n10144, n12094, n12115 );
nand U11927 ( n12115, n12058, n12116 );
not U11928 ( n12094, n12096 );
nor U11929 ( n12096, n12116, n12058 );
and U11930 ( n12058, n12117, n12118 );
nand U11931 ( n12118, n11796, n12119 );
xor U11932 ( n12117, n8082, n12120 );
nand U11933 ( n12120, n12121, n12122 );
nor U11934 ( n12122, n12123, n12124 );
nor U11935 ( n12124, n8082, n7850 );
nor U11936 ( n12123, n15232, n10975 );
nor U11937 ( n12121, n12125, n12126 );
nor U11938 ( n12126, n15195, n12049 );
nor U11939 ( n12125, n15289, n10843 );
and U11940 ( n12116, n12056, n12127 );
nand U11941 ( n12127, n10188, n12128 );
not U11942 ( n12056, n12129 );
nor U11943 ( n12110, n12130, n12131 );
nand U11944 ( n12131, n12132, n12133 );
nand U11945 ( n12133, n12134, n7850 );
nand U11946 ( n12132, n15232, n10847 );
nor U11947 ( n12130, n15320, n10855 );
nand U11948 ( n1395, n12135, n12136 );
nor U11949 ( n12136, n12137, n12138 );
nor U11950 ( n12138, n12139, n10851 );
nor U11951 ( n12137, n15231, n12140 );
nor U11952 ( n12140, n10847, n12134 );
nand U11953 ( n11209, n12141, n12142 );
nor U11954 ( n12142, n9095, n10842 );
not U11955 ( n10842, n10975 );
nor U11956 ( n12141, n12134, n7814 );
not U11957 ( n12134, n10854 );
nor U11958 ( n12135, n12143, n12144 );
nor U11959 ( n12144, n15319, n10855 );
nor U11960 ( n9095, n7797, n7799 );
nor U11961 ( n12143, n10180, n12106 );
nand U11962 ( n12106, n12145, n10854 );
nand U11963 ( n12147, n9383, n15063 );
and U11964 ( n12146, n12148, n9430 );
nand U11965 ( n9430, n12149, n12150 );
nor U11966 ( n12150, n12151, n12152 );
nand U11967 ( n12152, n12153, n9415 );
nand U11968 ( n12151, n9424, n7814 );
nor U11969 ( n12149, n12049, n12154 );
nand U11970 ( n12154, n9138, n15062 );
not U11971 ( n9138, n12155 );
nor U11972 ( n12145, n15062, n15351 );
and U11973 ( n10180, n12156, n12157 );
nand U11974 ( n12157, n12158, n12128 );
nor U11975 ( n12158, n10188, n12129 );
nor U11976 ( n12129, n12159, n12160 );
nand U11977 ( n12156, n12057, n10188 );
not U11978 ( n12057, n12128 );
nand U11979 ( n12128, n12160, n12159 );
nand U11980 ( n12159, n12161, n7797 );
nand U11981 ( n12161, n12162, n9426 );
xor U11982 ( n12160, n10188, n12163 );
nor U11983 ( n12163, n12164, n12165 );
nand U11984 ( n12165, n12166, n12167 );
nand U11985 ( n12167, n10867, n7873 );
not U11986 ( n10867, n10843 );
nand U11987 ( n12166, n12168, n7798 );
nand U11988 ( n12164, n12169, n12170 );
nand U11989 ( n12170, n12171, n8043 );
nand U11990 ( n12171, n8082, n10975 );
nand U11991 ( n10975, n15061, n7830 );
nand U11992 ( n12169, n11796, n10178 );
not U11993 ( n11796, n11844 );
nand U11994 ( n11844, n9426, n7797 );
nand U11995 ( n1390, n12172, n12173 );
nor U11996 ( n12173, n12174, n12175 );
nor U11997 ( n12175, n12176, n10850 );
xor U11998 ( n10850, n12177, n12178 );
xor U11999 ( n12178, n7834, n12179 );
nand U12000 ( n12177, n12180, n12181 );
nand U12001 ( n12181, n12182, n12183 );
nand U12002 ( n12183, n12184, n12185 );
nor U12003 ( n12185, n12186, n7818 );
nor U12004 ( n12184, n12187, n7845 );
nand U12005 ( n12180, n12186, n7845 );
and U12006 ( n12174, n12188, n9508 );
xnor U12007 ( n9508, n12189, n12190 );
nor U12008 ( n12190, n12191, n12192 );
nand U12009 ( n12189, n9363, n12193 );
nand U12010 ( n12193, n12194, n12195 );
nand U12011 ( n12195, n10822, n7834 );
nand U12012 ( n12194, n8022, n12196 );
nor U12013 ( n12172, n12197, n12198 );
nand U12014 ( n12198, n12199, n12200 );
nand U12015 ( n12200, n12201, n7834 );
nand U12016 ( n12201, n12202, n12203 );
nand U12017 ( n12203, n15229, n12204 );
nand U12018 ( n12199, n12205, n15230 );
nor U12019 ( n12205, n15229, n12206 );
nor U12020 ( n12197, n15350, n12207 );
nand U12021 ( n1385, n12208, n12209 );
nor U12022 ( n12209, n12210, n12211 );
nor U12023 ( n12211, n12176, n10924 );
xor U12024 ( n10924, n12179, n12212 );
xor U12025 ( n12212, n15229, n12213 );
nor U12026 ( n12213, n12186, n12214 );
nor U12027 ( n12214, n12215, n12179 );
nor U12028 ( n12215, n7818, n12187 );
and U12029 ( n12186, n12216, n12217 );
nor U12030 ( n12216, n12218, n12219 );
nor U12031 ( n12210, n12220, n9531 );
xnor U12032 ( n9531, n12192, n12191 );
xor U12033 ( n12191, n12221, n9363 );
nand U12034 ( n12221, n12222, n12223 );
nand U12035 ( n12223, n12196, n7875 );
nand U12036 ( n12222, n10822, n7845 );
nor U12037 ( n12208, n12224, n12225 );
nand U12038 ( n12225, n12226, n12227 );
or U12039 ( n12227, n12206, n7845 );
nand U12040 ( n12206, n12228, n7818 );
or U12041 ( n12226, n12202, n15229 );
nor U12042 ( n12202, n12229, n12230 );
and U12043 ( n12230, n15228, n12204 );
nor U12044 ( n12224, n15349, n12207 );
nand U12045 ( n1380, n12231, n12232 );
nor U12046 ( n12232, n12233, n12234 );
nor U12047 ( n12234, n12176, n10982 );
nand U12048 ( n10982, n12235, n12236 );
nand U12049 ( n12236, n12219, n12237 );
not U12050 ( n12237, n12238 );
nor U12051 ( n12219, n7818, n12182 );
nor U12052 ( n12235, n12239, n12240 );
nor U12053 ( n12240, n15228, n12241 );
xor U12054 ( n12241, n12179, n12238 );
nor U12055 ( n12239, n7818, n12242 );
nand U12056 ( n12242, n12182, n12238 );
nand U12057 ( n12238, n12243, n12244 );
nand U12058 ( n12244, n12182, n12187 );
nand U12059 ( n12187, n12245, n15021 );
nor U12060 ( n12245, n7841, n7801 );
nand U12061 ( n12243, n12217, n12246 );
and U12062 ( n12217, n12247, n12248 );
nand U12063 ( n12247, n12179, n12249 );
nor U12064 ( n12233, n12220, n9554 );
nand U12065 ( n9554, n12192, n12250 );
nand U12066 ( n12250, n12251, n12252 );
or U12067 ( n12192, n12252, n12251 );
xnor U12068 ( n12251, n12253, n12254 );
nand U12069 ( n12253, n12255, n12256 );
nand U12070 ( n12256, n12196, n7876 );
nand U12071 ( n12255, n10822, n7818 );
nor U12072 ( n12231, n12257, n12258 );
nand U12073 ( n12258, n12259, n12260 );
nand U12074 ( n12260, n15228, n12228 );
nand U12075 ( n12228, n12261, n12262 );
nand U12076 ( n12262, n12263, n12264 );
nand U12077 ( n12261, n12265, n12266 );
nand U12078 ( n12259, n12229, n7818 );
nand U12079 ( n12229, n12267, n12268 );
nor U12080 ( n12267, n12269, n12270 );
nor U12081 ( n12270, n12265, n12271 );
and U12082 ( n12265, n12272, n12273 );
nor U12083 ( n12272, n12274, n12249 );
nor U12084 ( n12269, n12263, n12275 );
not U12085 ( n12263, n12249 );
nand U12086 ( n12249, n7801, n7860 );
nor U12087 ( n12257, n15348, n12207 );
nand U12088 ( n1375, n12276, n12277 );
nor U12089 ( n12277, n12278, n12279 );
nor U12090 ( n12279, n12176, n11038 );
xor U12091 ( n11038, n12280, n12182 );
xor U12092 ( n12280, n12281, n15021 );
nand U12093 ( n12281, n12282, n12283 );
nand U12094 ( n12283, n12182, n7801 );
nor U12095 ( n12282, n12284, n12285 );
nor U12096 ( n12285, n12286, n12287 );
nand U12097 ( n12287, n12248, n12246 );
nor U12098 ( n12278, n12220, n9579 );
nand U12099 ( n9579, n12252, n12288 );
nand U12100 ( n12288, n12289, n12290 );
or U12101 ( n12252, n12290, n12289 );
xnor U12102 ( n12289, n12291, n12254 );
nand U12103 ( n12291, n12292, n12293 );
nand U12104 ( n12293, n12196, n7877 );
nand U12105 ( n12292, n10822, n7860 );
nor U12106 ( n12276, n12294, n12295 );
nand U12107 ( n12295, n12296, n12297 );
nand U12108 ( n12297, n12298, n7860 );
nand U12109 ( n12298, n12299, n12300 );
nand U12110 ( n12300, n15227, n12204 );
not U12111 ( n12299, n12301 );
nand U12112 ( n12296, n12302, n15021 );
nor U12113 ( n12302, n15227, n12303 );
nor U12114 ( n12294, n15347, n12207 );
nand U12115 ( n1370, n12304, n12305 );
nor U12116 ( n12305, n12306, n12307 );
nor U12117 ( n12307, n12176, n11094 );
nand U12118 ( n11094, n12308, n12309 );
nand U12119 ( n12309, n12286, n12310 );
nor U12120 ( n12286, n7801, n12182 );
nor U12121 ( n12308, n12311, n12312 );
nor U12122 ( n12312, n15227, n12313 );
xor U12123 ( n12313, n12179, n12314 );
nor U12124 ( n12311, n7801, n12315 );
nand U12125 ( n12315, n12182, n12314 );
not U12126 ( n12314, n12310 );
nor U12127 ( n12310, n12284, n12316 );
nor U12128 ( n12316, n12317, n12218 );
nor U12129 ( n12306, n12220, n9599 );
nand U12130 ( n9599, n12290, n12318 );
nand U12131 ( n12318, n12319, n12320 );
or U12132 ( n12290, n12320, n12319 );
xnor U12133 ( n12319, n12321, n12254 );
nand U12134 ( n12321, n12322, n12323 );
nand U12135 ( n12323, n12196, n7878 );
nand U12136 ( n12322, n10822, n7801 );
nor U12137 ( n12304, n12324, n12325 );
nand U12138 ( n12325, n12326, n12327 );
or U12139 ( n12327, n7801, n12303 );
nor U12140 ( n12303, n12264, n12328 );
and U12141 ( n12328, n12329, n12266 );
nor U12142 ( n12329, n12274, n12330 );
nand U12143 ( n12264, n12331, n12332 );
nand U12144 ( n12332, n12333, n12334 );
or U12145 ( n12331, n12335, n12336 );
nand U12146 ( n12326, n12301, n7801 );
nand U12147 ( n12301, n12268, n12337 );
nand U12148 ( n12337, n12266, n12338 );
nand U12149 ( n12338, n12273, n12339 );
and U12150 ( n12268, n12340, n12341 );
nand U12151 ( n12341, n12342, n12335 );
nand U12152 ( n12335, n12343, n12344 );
nor U12153 ( n12343, n15224, n12274 );
nor U12154 ( n12340, n12345, n12346 );
nor U12155 ( n12346, n12334, n12347 );
and U12156 ( n12334, n12348, n12339 );
not U12157 ( n12339, n12274 );
nand U12158 ( n12274, n7807, n7841 );
nor U12159 ( n12348, n15224, n12349 );
nor U12160 ( n12324, n15346, n12207 );
nand U12161 ( n1365, n12350, n12351 );
nor U12162 ( n12351, n12352, n12353 );
nor U12163 ( n12353, n12220, n9618 );
nand U12164 ( n9618, n12320, n12354 );
nand U12165 ( n12354, n12355, n12356 );
or U12166 ( n12320, n12356, n12355 );
xnor U12167 ( n12355, n12357, n12254 );
nand U12168 ( n12357, n12358, n12359 );
nand U12169 ( n12359, n12196, n7879 );
nand U12170 ( n12358, n10822, n7841 );
nor U12171 ( n12352, n12176, n11150 );
xor U12172 ( n11150, n12218, n12360 );
nor U12173 ( n12360, n12284, n12317 );
not U12174 ( n12317, n12248 );
nand U12175 ( n12248, n15226, n12179 );
nor U12176 ( n12284, n12179, n15226 );
not U12177 ( n12218, n12246 );
nand U12178 ( n12246, n12361, n12362 );
nand U12179 ( n12362, n12182, n12363 );
nand U12180 ( n12363, n12364, n12365 );
not U12181 ( n12364, n12366 );
nand U12182 ( n12361, n12367, n7807 );
nand U12183 ( n12367, n12368, n12179 );
nand U12184 ( n12368, n12366, n7824 );
nor U12185 ( n12350, n12369, n12370 );
nand U12186 ( n12370, n12371, n12372 );
nand U12187 ( n12372, n12373, n7841 );
nand U12188 ( n12373, n12374, n12375 );
nand U12189 ( n12375, n15225, n12204 );
not U12190 ( n12374, n12376 );
nand U12191 ( n12371, n12377, n15226 );
and U12192 ( n12377, n7807, n12378 );
nor U12193 ( n12369, n15345, n12207 );
nand U12194 ( n1360, n12379, n12380 );
nor U12195 ( n12380, n12381, n12382 );
nor U12196 ( n12382, n12220, n9638 );
nand U12197 ( n9638, n12356, n12383 );
nand U12198 ( n12383, n12384, n12385 );
or U12199 ( n12356, n12385, n12384 );
xnor U12200 ( n12384, n12386, n12254 );
nand U12201 ( n12386, n12387, n12388 );
nand U12202 ( n12388, n12196, n7880 );
nand U12203 ( n12387, n10822, n7807 );
nor U12204 ( n12381, n12176, n12389 );
nand U12205 ( n12389, n11162, n11161 );
or U12206 ( n11161, n12390, n12391 );
nand U12207 ( n11162, n12391, n12390 );
xor U12208 ( n12390, n12179, n7807 );
and U12209 ( n12391, n12392, n12365 );
nand U12210 ( n12392, n12366, n12393 );
nor U12211 ( n12379, n12394, n12395 );
nand U12212 ( n12395, n12396, n12397 );
nand U12213 ( n12397, n15225, n12378 );
nand U12214 ( n12378, n12398, n12399 );
nand U12215 ( n12399, n12400, n7824 );
nand U12216 ( n12400, n12401, n12402 );
nand U12217 ( n12402, n12333, n12403 );
nand U12218 ( n12398, n12266, n12273 );
nand U12219 ( n12396, n12376, n7807 );
nand U12220 ( n12376, n12404, n12405 );
nor U12221 ( n12405, n12406, n12407 );
nand U12222 ( n12407, n12408, n12409 );
nand U12223 ( n12408, n12333, n12349 );
not U12224 ( n12349, n12403 );
nor U12225 ( n12403, n12410, n15223 );
nor U12226 ( n12406, n12273, n12271 );
not U12227 ( n12273, n12330 );
nand U12228 ( n12330, n12411, n12412 );
nor U12229 ( n12411, n15223, n15224 );
nor U12230 ( n12404, n12413, n12414 );
nor U12231 ( n12414, n12275, n7824 );
nor U12232 ( n12394, n15344, n12207 );
nand U12233 ( n1355, n12415, n12416 );
nor U12234 ( n12416, n12417, n12418 );
nor U12235 ( n12418, n12176, n11265 );
xor U12236 ( n11265, n12419, n12366 );
nand U12237 ( n12366, n12420, n12421 );
nor U12238 ( n12420, n12422, n12423 );
nor U12239 ( n12422, n12424, n12425 );
nand U12240 ( n12419, n12365, n12393 );
nand U12241 ( n12393, n15224, n12179 );
nand U12242 ( n12365, n12182, n7824 );
nor U12243 ( n12417, n12220, n9658 );
nand U12244 ( n9658, n12385, n12426 );
nand U12245 ( n12426, n12427, n12428 );
or U12246 ( n12385, n12428, n12427 );
xnor U12247 ( n12427, n12429, n12254 );
nand U12248 ( n12429, n12430, n12431 );
nand U12249 ( n12431, n12196, n7881 );
nand U12250 ( n12430, n10822, n7824 );
nor U12251 ( n12415, n12432, n12433 );
nand U12252 ( n12433, n12434, n12435 );
nand U12253 ( n12435, n12436, n7824 );
nand U12254 ( n12436, n12437, n12438 );
nor U12255 ( n12437, n12413, n12439 );
nor U12256 ( n12439, n12440, n7823 );
nor U12257 ( n12413, n12344, n12336 );
nand U12258 ( n12434, n15224, n12441 );
nand U12259 ( n12441, n12442, n12401 );
nand U12260 ( n12401, n12342, n12344 );
nor U12261 ( n12344, n12443, n15223 );
nand U12262 ( n12442, n12444, n7823 );
nor U12263 ( n12432, n15343, n12207 );
nand U12264 ( n1350, n12445, n12446 );
nor U12265 ( n12446, n12447, n12448 );
nor U12266 ( n12448, n12220, n9677 );
nand U12267 ( n9677, n12428, n12449 );
nand U12268 ( n12449, n12450, n12451 );
or U12269 ( n12428, n12451, n12450 );
xnor U12270 ( n12450, n12452, n12254 );
nand U12271 ( n12452, n12453, n12454 );
nand U12272 ( n12454, n12196, n7882 );
nand U12273 ( n12453, n10822, n7823 );
nor U12274 ( n12447, n12176, n12455 );
nand U12275 ( n12455, n11276, n11275 );
nand U12276 ( n11275, n12456, n12457 );
nand U12277 ( n12457, n12182, n7823 );
nor U12278 ( n12456, n12424, n12458 );
and U12279 ( n12458, n12425, n12421 );
nand U12280 ( n11276, n12459, n12421 );
nor U12281 ( n12421, n12460, n12461 );
and U12282 ( n12460, n12182, n12462 );
nand U12283 ( n12462, n15220, n15221 );
nor U12284 ( n12459, n12463, n12464 );
nor U12285 ( n12464, n12424, n12423 );
nor U12286 ( n12423, n15223, n12179 );
nor U12287 ( n12424, n7823, n12182 );
not U12288 ( n12463, n12425 );
nand U12289 ( n12425, n12465, n12466 );
nor U12290 ( n12465, n12467, n12468 );
nor U12291 ( n12445, n12469, n12470 );
nand U12292 ( n12470, n12471, n12472 );
nand U12293 ( n12472, n15223, n12473 );
nand U12294 ( n12473, n12474, n12475 );
or U12295 ( n12475, n12336, n12443 );
not U12296 ( n12474, n12444 );
nand U12297 ( n12444, n12476, n12477 );
nand U12298 ( n12477, n12266, n12412 );
or U12299 ( n12476, n12347, n12410 );
nand U12300 ( n12471, n12478, n7823 );
nand U12301 ( n12478, n12438, n12479 );
nand U12302 ( n12479, n12342, n12443 );
nand U12303 ( n12443, n12480, n12481 );
and U12304 ( n12438, n12482, n12483 );
nand U12305 ( n12483, n12333, n12410 );
nand U12306 ( n12410, n12480, n12484 );
nor U12307 ( n12482, n12345, n12485 );
nor U12308 ( n12485, n12412, n12271 );
and U12309 ( n12412, n12480, n12486 );
nor U12310 ( n12480, n15221, n15222 );
nor U12311 ( n12469, n15342, n12207 );
nand U12312 ( n1345, n12487, n12488 );
nor U12313 ( n12488, n12489, n12490 );
nor U12314 ( n12490, n12176, n11447 );
xnor U12315 ( n11447, n12491, n12492 );
nor U12316 ( n12492, n12468, n12461 );
nor U12317 ( n12461, n12179, n15222 );
nor U12318 ( n12468, n7862, n12182 );
nand U12319 ( n12491, n12493, n12494 );
nand U12320 ( n12494, n12182, n7833 );
nor U12321 ( n12493, n12495, n12496 );
nor U12322 ( n12496, n12467, n12497 );
not U12323 ( n12495, n12498 );
nor U12324 ( n12489, n12220, n9697 );
nand U12325 ( n9697, n12451, n12499 );
nand U12326 ( n12499, n12500, n12501 );
or U12327 ( n12451, n12501, n12500 );
xnor U12328 ( n12500, n12502, n12254 );
nand U12329 ( n12502, n12503, n12504 );
nand U12330 ( n12504, n12196, n7883 );
nand U12331 ( n12503, n10822, n7862 );
nor U12332 ( n12487, n12505, n12506 );
nand U12333 ( n12506, n12507, n12508 );
nand U12334 ( n12508, n12509, n7862 );
nand U12335 ( n12509, n12510, n12511 );
nand U12336 ( n12511, n15221, n12204 );
not U12337 ( n12510, n12512 );
nand U12338 ( n12507, n12513, n15222 );
and U12339 ( n12513, n7833, n12514 );
nor U12340 ( n12505, n15341, n12207 );
nand U12341 ( n1340, n12515, n12516 );
nor U12342 ( n12516, n12517, n12518 );
nor U12343 ( n12518, n12176, n11504 );
xnor U12344 ( n11504, n12519, n12520 );
nor U12345 ( n12520, n12467, n12521 );
nor U12346 ( n12521, n15221, n12179 );
nor U12347 ( n12467, n7833, n12182 );
nand U12348 ( n12519, n12498, n12497 );
nor U12349 ( n12517, n12220, n9717 );
nand U12350 ( n9717, n12501, n12522 );
nand U12351 ( n12522, n12523, n12524 );
or U12352 ( n12501, n12524, n12523 );
xnor U12353 ( n12523, n12525, n12254 );
nand U12354 ( n12525, n12526, n12527 );
nand U12355 ( n12527, n12196, n7884 );
nand U12356 ( n12526, n10822, n7833 );
nor U12357 ( n12515, n12528, n12529 );
nand U12358 ( n12529, n12530, n12531 );
nand U12359 ( n12531, n15221, n12514 );
nand U12360 ( n12514, n12532, n12533 );
nand U12361 ( n12533, n12342, n12481 );
nor U12362 ( n12532, n12534, n12535 );
nor U12363 ( n12535, n12536, n12347 );
nor U12364 ( n12534, n12537, n12271 );
nand U12365 ( n12530, n12512, n7833 );
nand U12366 ( n12512, n12538, n12539 );
nor U12367 ( n12539, n12345, n12540 );
nor U12368 ( n12540, n12486, n12271 );
not U12369 ( n12486, n12537 );
nand U12370 ( n12537, n12541, n7839 );
nor U12371 ( n12538, n12542, n12543 );
nor U12372 ( n12543, n12481, n12336 );
and U12373 ( n12481, n12544, n12545 );
nor U12374 ( n12545, n15218, n15219 );
nor U12375 ( n12544, n15220, n12546 );
nor U12376 ( n12542, n12484, n12347 );
not U12377 ( n12484, n12536 );
nand U12378 ( n12536, n12547, n12548 );
nor U12379 ( n12547, n15219, n15220 );
nor U12380 ( n12528, n15340, n12207 );
nand U12381 ( n1335, n12549, n12550 );
nor U12382 ( n12550, n12551, n12552 );
nor U12383 ( n12552, n12220, n9738 );
nand U12384 ( n9738, n12524, n12553 );
nand U12385 ( n12553, n12554, n12555 );
or U12386 ( n12524, n12555, n12554 );
xnor U12387 ( n12554, n12556, n12254 );
nand U12388 ( n12556, n12557, n12558 );
nand U12389 ( n12558, n12196, n7885 );
nand U12390 ( n12557, n10822, n7839 );
nor U12391 ( n12551, n12176, n11556 );
nand U12392 ( n11556, n12559, n12560 );
nand U12393 ( n12560, n12561, n12562 );
nand U12394 ( n12562, n12498, n12563 );
not U12395 ( n12561, n12564 );
nand U12396 ( n12559, n12466, n12498 );
nand U12397 ( n12498, n12182, n7839 );
not U12398 ( n12466, n12497 );
nand U12399 ( n12497, n12564, n12563 );
nand U12400 ( n12563, n15220, n12179 );
nand U12401 ( n12564, n12565, n12566 );
nand U12402 ( n12566, n12567, n7829 );
or U12403 ( n12567, n12568, n12182 );
nand U12404 ( n12565, n12182, n12568 );
nor U12405 ( n12549, n12569, n12570 );
nand U12406 ( n12570, n12571, n12572 );
nand U12407 ( n12572, n12573, n7839 );
nand U12408 ( n12573, n12574, n12575 );
nor U12409 ( n12574, n12576, n12577 );
nor U12410 ( n12577, n12275, n7829 );
nor U12411 ( n12576, n12541, n12271 );
nand U12412 ( n12571, n15220, n12578 );
nand U12413 ( n12578, n12579, n12580 );
nand U12414 ( n12580, n12266, n12541 );
nor U12415 ( n12541, n12581, n15219 );
nand U12416 ( n12579, n12582, n7829 );
nor U12417 ( n12569, n15339, n12207 );
nand U12418 ( n1330, n12583, n12584 );
nor U12419 ( n12584, n12585, n12586 );
nor U12420 ( n12586, n12176, n11606 );
xnor U12421 ( n11606, n12587, n12568 );
nand U12422 ( n12568, n12588, n12589 );
nand U12423 ( n12589, n12182, n12590 );
nand U12424 ( n12590, n12591, n15218 );
nor U12425 ( n12591, n12592, n12593 );
or U12426 ( n12588, n12594, n15218 );
xor U12427 ( n12587, n12179, n15219 );
nor U12428 ( n12585, n12220, n9758 );
nand U12429 ( n9758, n12555, n12595 );
nand U12430 ( n12595, n12596, n12597 );
or U12431 ( n12555, n12597, n12596 );
xnor U12432 ( n12596, n12598, n12254 );
nand U12433 ( n12598, n12599, n12600 );
nand U12434 ( n12600, n12196, n7886 );
nand U12435 ( n12599, n10822, n7829 );
nor U12436 ( n12583, n12601, n12602 );
nand U12437 ( n12602, n12603, n12604 );
nand U12438 ( n12604, n15219, n12605 );
nand U12439 ( n12605, n12606, n12607 );
or U12440 ( n12607, n12271, n12581 );
not U12441 ( n12606, n12582 );
nand U12442 ( n12582, n12608, n12609 );
nand U12443 ( n12609, n12610, n12342 );
nor U12444 ( n12610, n15218, n12546 );
not U12445 ( n12546, n12611 );
nand U12446 ( n12608, n12333, n12548 );
and U12447 ( n12548, n12612, n12613 );
nand U12448 ( n12603, n12614, n7829 );
nand U12449 ( n12614, n12575, n12615 );
nand U12450 ( n12615, n12266, n12581 );
nand U12451 ( n12581, n12612, n12616 );
nor U12452 ( n12612, n15217, n15218 );
and U12453 ( n12575, n12617, n12618 );
nor U12454 ( n12618, n12619, n12620 );
nor U12455 ( n12620, n12275, n7835 );
nor U12456 ( n12617, n12621, n12622 );
nor U12457 ( n12621, n7828, n12347 );
nor U12458 ( n12601, n15338, n12207 );
nand U12459 ( n1325, n12623, n12624 );
nor U12460 ( n12624, n12625, n12626 );
nor U12461 ( n12626, n12176, n11656 );
xor U12462 ( n11656, n12627, n12628 );
xor U12463 ( n12628, n7835, n12179 );
nand U12464 ( n12627, n12594, n12629 );
nand U12465 ( n12629, n12182, n12592 );
nand U12466 ( n12592, n15217, n12630 );
nand U12467 ( n12594, n12631, n12632 );
nand U12468 ( n12632, n15217, n12179 );
nor U12469 ( n12625, n12220, n9780 );
nand U12470 ( n9780, n12597, n12633 );
nand U12471 ( n12633, n12634, n12635 );
or U12472 ( n12597, n12635, n12634 );
xnor U12473 ( n12634, n12636, n12254 );
nand U12474 ( n12636, n12637, n12638 );
nand U12475 ( n12638, n12196, n7887 );
nand U12476 ( n12637, n10822, n7835 );
nor U12477 ( n12623, n12639, n12640 );
nand U12478 ( n12640, n12641, n12642 );
nand U12479 ( n12642, n12643, n7835 );
nand U12480 ( n12643, n12644, n12645 );
nor U12481 ( n12644, n12619, n12646 );
nor U12482 ( n12646, n12440, n7828 );
nor U12483 ( n12619, n12611, n12336 );
nand U12484 ( n12641, n15218, n12647 );
nand U12485 ( n12647, n12648, n12649 );
nand U12486 ( n12649, n12342, n12611 );
nor U12487 ( n12611, n12650, n15217 );
nand U12488 ( n12648, n12651, n7828 );
nor U12489 ( n12639, n15337, n12207 );
nand U12490 ( n1320, n12652, n12653 );
nor U12491 ( n12653, n12654, n12655 );
nor U12492 ( n12655, n12176, n11703 );
xor U12493 ( n11703, n12656, n12657 );
nor U12494 ( n12657, n12631, n12658 );
xor U12495 ( n12656, n12179, n15217 );
nor U12496 ( n12654, n12220, n9800 );
nand U12497 ( n9800, n12635, n12659 );
nand U12498 ( n12659, n12660, n12661 );
or U12499 ( n12635, n12661, n12660 );
xnor U12500 ( n12660, n12662, n12254 );
nand U12501 ( n12662, n12663, n12664 );
nand U12502 ( n12664, n12196, n7888 );
nand U12503 ( n12663, n10822, n7828 );
nor U12504 ( n12652, n12665, n12666 );
nand U12505 ( n12666, n12667, n12668 );
nand U12506 ( n12668, n15217, n12669 );
nand U12507 ( n12669, n12670, n12671 );
or U12508 ( n12671, n12336, n12650 );
not U12509 ( n12670, n12651 );
nand U12510 ( n12651, n12672, n12673 );
nand U12511 ( n12673, n12266, n12616 );
nand U12512 ( n12672, n12333, n12613 );
not U12513 ( n12613, n12674 );
nand U12514 ( n12667, n12675, n7828 );
nand U12515 ( n12675, n12645, n12676 );
nand U12516 ( n12676, n12342, n12650 );
nand U12517 ( n12650, n12677, n12678 );
nor U12518 ( n12645, n12622, n12679 );
nor U12519 ( n12679, n12271, n12616 );
and U12520 ( n12616, n12677, n12680 );
nand U12521 ( n12622, n12409, n12681 );
nand U12522 ( n12681, n12333, n12674 );
nand U12523 ( n12674, n12677, n12682 );
nor U12524 ( n12677, n15215, n15216 );
nor U12525 ( n12665, n15336, n12207 );
nand U12526 ( n1315, n12683, n12684 );
nor U12527 ( n12684, n12685, n12686 );
nor U12528 ( n12686, n12220, n9822 );
nand U12529 ( n9822, n12661, n12687 );
nand U12530 ( n12687, n12688, n12689 );
or U12531 ( n12661, n12689, n12688 );
xnor U12532 ( n12688, n12690, n12254 );
nand U12533 ( n12690, n12691, n12692 );
nand U12534 ( n12692, n12196, n7889 );
nand U12535 ( n12691, n10822, n7842 );
nor U12536 ( n12685, n12176, n12693 );
nand U12537 ( n12693, n11714, n11713 );
nand U12538 ( n11713, n12631, n12630 );
nor U12539 ( n12631, n12694, n12695 );
nand U12540 ( n11714, n12694, n12696 );
or U12541 ( n12696, n12658, n12695 );
nor U12542 ( n12695, n7842, n12182 );
not U12543 ( n12658, n12630 );
nand U12544 ( n12630, n12182, n7842 );
not U12545 ( n12182, n12179 );
nand U12546 ( n12179, n12697, n12698 );
nor U12547 ( n12697, n12699, n12700 );
not U12548 ( n12694, n12593 );
nand U12549 ( n12593, n12701, n12702 );
nand U12550 ( n12702, n12703, n12704 );
nand U12551 ( n12703, n12705, n12706 );
and U12552 ( n12706, n12707, n12708 );
nor U12553 ( n12705, n12709, n12710 );
nor U12554 ( n12710, n12711, n12712 );
nand U12555 ( n12712, n12713, n12714 );
nor U12556 ( n12683, n12715, n12716 );
nand U12557 ( n12716, n12717, n12718 );
nand U12558 ( n12718, n12719, n7842 );
nand U12559 ( n12719, n12720, n12721 );
nand U12560 ( n12721, n15215, n12204 );
not U12561 ( n12720, n12722 );
nand U12562 ( n12717, n12723, n15216 );
and U12563 ( n12723, n7906, n12724 );
nor U12564 ( n12715, n15335, n12207 );
nand U12565 ( n1310, n12725, n12726 );
nor U12566 ( n12726, n12727, n12728 );
nor U12567 ( n12728, n12220, n9843 );
nand U12568 ( n9843, n12689, n12729 );
nand U12569 ( n12729, n12730, n12731 );
or U12570 ( n12689, n12731, n12730 );
xnor U12571 ( n12730, n12732, n12254 );
nand U12572 ( n12732, n12733, n12734 );
nand U12573 ( n12734, n12196, n7890 );
nand U12574 ( n12733, n10822, n7906 );
nor U12575 ( n12727, n12176, n11806 );
xnor U12576 ( n11806, n12735, n12736 );
nor U12577 ( n12736, n12737, n12709 );
not U12578 ( n12709, n12738 );
nor U12579 ( n12737, n12739, n12740 );
not U12580 ( n12739, n12713 );
nand U12581 ( n12735, n12701, n12704 );
nand U12582 ( n12704, n15215, n12741 );
nand U12583 ( n12741, n11795, n12742 );
nand U12584 ( n12701, n12743, n11795 );
and U12585 ( n11795, n12744, n12745 );
nand U12586 ( n12745, n12746, n12747 );
nor U12587 ( n12747, n12748, n12749 );
nand U12588 ( n12749, n12750, n12751 );
nor U12589 ( n12751, n12752, n12753 );
nor U12590 ( n12753, n15080, n12754 );
nor U12591 ( n12752, n15088, n12755 );
nor U12592 ( n12750, n12756, n12757 );
nor U12593 ( n12757, n15072, n12758 );
nor U12594 ( n12756, n15064, n12759 );
nand U12595 ( n12748, n12760, n12761 );
nor U12596 ( n12761, n12762, n12763 );
nand U12597 ( n12763, n12764, n12765 );
nand U12598 ( n12764, n12766, n7994 );
nor U12599 ( n12762, n15112, n12767 );
nor U12600 ( n12760, n12768, n12769 );
nor U12601 ( n12769, n15104, n12770 );
nor U12602 ( n12768, n15096, n12771 );
nor U12603 ( n12746, n12772, n12773 );
nand U12604 ( n12773, n12774, n12775 );
nor U12605 ( n12775, n12776, n12777 );
nor U12606 ( n12777, n15176, n12778 );
nor U12607 ( n12776, n15184, n12779 );
nor U12608 ( n12774, n12780, n12781 );
nor U12609 ( n12781, n15168, n12782 );
nor U12610 ( n12780, n15160, n12783 );
nand U12611 ( n12772, n12784, n12785 );
nor U12612 ( n12785, n12786, n12787 );
nor U12613 ( n12787, n15144, n12788 );
nor U12614 ( n12786, n15152, n12789 );
nor U12615 ( n12784, n12790, n12791 );
nor U12616 ( n12791, n15136, n12792 );
nor U12617 ( n12790, n15128, n12793 );
nor U12618 ( n12743, n15215, n12700 );
nor U12619 ( n12725, n12794, n12795 );
nand U12620 ( n12795, n12796, n12797 );
nand U12621 ( n12797, n15215, n12724 );
nand U12622 ( n12724, n12798, n12799 );
nand U12623 ( n12799, n12342, n12678 );
nor U12624 ( n12798, n12800, n12801 );
nor U12625 ( n12801, n12802, n12347 );
nor U12626 ( n12800, n12803, n12271 );
nand U12627 ( n12796, n12722, n7906 );
nand U12628 ( n12722, n12804, n12805 );
nor U12629 ( n12805, n12345, n12806 );
nor U12630 ( n12806, n12680, n12271 );
not U12631 ( n12680, n12803 );
nand U12632 ( n12803, n12807, n7854 );
nor U12633 ( n12804, n12808, n12809 );
nor U12634 ( n12809, n12678, n12336 );
and U12635 ( n12678, n12810, n12811 );
nor U12636 ( n12808, n12682, n12347 );
not U12637 ( n12682, n12802 );
nand U12638 ( n12802, n12810, n12812 );
nor U12639 ( n12810, n15213, n15214 );
nor U12640 ( n12794, n15334, n12207 );
nand U12641 ( n1305, n12813, n12814 );
nor U12642 ( n12814, n12815, n12816 );
nor U12643 ( n12816, n12176, n11829 );
xnor U12644 ( n11829, n12817, n12740 );
and U12645 ( n12740, n12708, n12818 );
nand U12646 ( n12818, n12819, n12714 );
nand U12647 ( n12817, n12713, n12738 );
nand U12648 ( n12738, n12820, n11821 );
nor U12649 ( n12820, n15214, n12700 );
nand U12650 ( n12713, n15214, n12821 );
nand U12651 ( n12821, n11821, n12742 );
and U12652 ( n11821, n12744, n12822 );
nand U12653 ( n12822, n12823, n12824 );
nor U12654 ( n12824, n12825, n12826 );
nand U12655 ( n12826, n12827, n12828 );
nor U12656 ( n12828, n12829, n12830 );
nor U12657 ( n12830, n15081, n12754 );
nor U12658 ( n12829, n15089, n12755 );
nor U12659 ( n12827, n12831, n12832 );
nor U12660 ( n12832, n15073, n12758 );
nor U12661 ( n12831, n15065, n12759 );
nand U12662 ( n12825, n12833, n12834 );
nor U12663 ( n12834, n12835, n12836 );
nand U12664 ( n12836, n12837, n12765 );
nand U12665 ( n12837, n12766, n7865 );
nor U12666 ( n12835, n15113, n12767 );
nor U12667 ( n12833, n12838, n12839 );
nor U12668 ( n12839, n15105, n12770 );
nor U12669 ( n12838, n15097, n12771 );
nor U12670 ( n12823, n12840, n12841 );
nand U12671 ( n12841, n12842, n12843 );
nor U12672 ( n12843, n12844, n12845 );
nor U12673 ( n12845, n15177, n12778 );
nor U12674 ( n12844, n15185, n12779 );
nor U12675 ( n12842, n12846, n12847 );
nor U12676 ( n12847, n15169, n12782 );
nor U12677 ( n12846, n15161, n12783 );
nand U12678 ( n12840, n12848, n12849 );
nor U12679 ( n12849, n12850, n12851 );
nor U12680 ( n12851, n15145, n12788 );
nor U12681 ( n12850, n15153, n12789 );
nor U12682 ( n12848, n12852, n12853 );
nor U12683 ( n12853, n15137, n12792 );
nor U12684 ( n12852, n15129, n12793 );
nor U12685 ( n12815, n12220, n9863 );
nand U12686 ( n9863, n12731, n12854 );
nand U12687 ( n12854, n12855, n12856 );
or U12688 ( n12731, n12856, n12855 );
xnor U12689 ( n12855, n12857, n12254 );
nand U12690 ( n12857, n12858, n12859 );
nand U12691 ( n12859, n12196, n7891 );
nand U12692 ( n12858, n10822, n7854 );
nor U12693 ( n12813, n12860, n12861 );
nand U12694 ( n12861, n12862, n12863 );
nand U12695 ( n12863, n12864, n7854 );
nand U12696 ( n12864, n12865, n12866 );
nor U12697 ( n12865, n12867, n12868 );
nor U12698 ( n12868, n12275, n7840 );
nor U12699 ( n12867, n12807, n12271 );
nand U12700 ( n12862, n15214, n12869 );
nand U12701 ( n12869, n12870, n12871 );
nand U12702 ( n12871, n12266, n12807 );
nor U12703 ( n12807, n12872, n15213 );
nand U12704 ( n12870, n12873, n7840 );
nor U12705 ( n12860, n15333, n12207 );
nand U12706 ( n1300, n12874, n12875 );
nor U12707 ( n12875, n12876, n12877 );
nor U12708 ( n12877, n12176, n11854 );
xor U12709 ( n11854, n12878, n12819 );
nand U12710 ( n12819, n12711, n12707 );
nand U12711 ( n12878, n12714, n12708 );
nand U12712 ( n12708, n12879, n11842 );
nor U12713 ( n12879, n15213, n12700 );
nand U12714 ( n12714, n15213, n12880 );
nand U12715 ( n12880, n11842, n12742 );
not U12716 ( n11842, n11845 );
nand U12717 ( n11845, n12744, n12881 );
nand U12718 ( n12881, n12882, n12883 );
nor U12719 ( n12883, n12884, n12885 );
nand U12720 ( n12885, n12886, n12887 );
nor U12721 ( n12887, n12888, n12889 );
nor U12722 ( n12889, n15082, n12754 );
nor U12723 ( n12888, n15090, n12755 );
nor U12724 ( n12886, n12890, n12891 );
nor U12725 ( n12891, n15074, n12758 );
nor U12726 ( n12890, n15066, n12759 );
nand U12727 ( n12884, n12892, n12893 );
nor U12728 ( n12893, n12894, n12895 );
nand U12729 ( n12895, n12896, n12765 );
nand U12730 ( n12896, n12766, n7866 );
nor U12731 ( n12894, n15114, n12767 );
nor U12732 ( n12892, n12897, n12898 );
nor U12733 ( n12898, n15106, n12770 );
nor U12734 ( n12897, n15098, n12771 );
nor U12735 ( n12882, n12899, n12900 );
nand U12736 ( n12900, n12901, n12902 );
nor U12737 ( n12902, n12903, n12904 );
nor U12738 ( n12904, n15178, n12778 );
nor U12739 ( n12903, n15186, n12779 );
nor U12740 ( n12901, n12905, n12906 );
nor U12741 ( n12906, n15170, n12782 );
nor U12742 ( n12905, n15162, n12783 );
nand U12743 ( n12899, n12907, n12908 );
nor U12744 ( n12908, n12909, n12910 );
nor U12745 ( n12910, n15146, n12788 );
nor U12746 ( n12909, n15154, n12789 );
nor U12747 ( n12907, n12911, n12912 );
nor U12748 ( n12912, n15138, n12792 );
nor U12749 ( n12911, n15130, n12793 );
nor U12750 ( n12876, n12220, n9884 );
nand U12751 ( n9884, n12856, n12913 );
nand U12752 ( n12913, n12914, n12915 );
or U12753 ( n12856, n12915, n12914 );
xnor U12754 ( n12914, n12916, n12254 );
nand U12755 ( n12916, n12917, n12918 );
nand U12756 ( n12918, n12196, n7892 );
nand U12757 ( n12917, n10822, n7840 );
nor U12758 ( n12874, n12919, n12920 );
nand U12759 ( n12920, n12921, n12922 );
nand U12760 ( n12922, n15213, n12923 );
nand U12761 ( n12923, n12924, n12925 );
or U12762 ( n12925, n12271, n12872 );
not U12763 ( n12924, n12873 );
nand U12764 ( n12873, n12926, n12927 );
nand U12765 ( n12927, n12333, n12812 );
nand U12766 ( n12926, n12342, n12811 );
not U12767 ( n12811, n12928 );
nand U12768 ( n12921, n12929, n7840 );
nand U12769 ( n12929, n12866, n12930 );
nand U12770 ( n12930, n12266, n12872 );
nand U12771 ( n12872, n12931, n12932 );
and U12772 ( n12866, n12933, n12934 );
nand U12773 ( n12934, n12342, n12928 );
nand U12774 ( n12928, n12931, n12935 );
nor U12775 ( n12933, n12345, n12936 );
nor U12776 ( n12936, n12812, n12347 );
and U12777 ( n12812, n12931, n12937 );
nor U12778 ( n12931, n15211, n15212 );
nor U12779 ( n12919, n15332, n12207 );
nand U12780 ( n1295, n12938, n12939 );
nor U12781 ( n12939, n12940, n12941 );
nor U12782 ( n12941, n12176, n11873 );
nand U12783 ( n11873, n12942, n12943 );
nand U12784 ( n12943, n12944, n12945 );
nand U12785 ( n12945, n12707, n12946 );
not U12786 ( n12707, n12947 );
not U12787 ( n12944, n12948 );
or U12788 ( n12942, n12711, n12947 );
nor U12789 ( n12947, n12949, n15212 );
nand U12790 ( n12711, n12948, n12946 );
nand U12791 ( n12946, n15212, n12949 );
nand U12792 ( n12949, n11865, n12742 );
and U12793 ( n11865, n12744, n12950 );
nand U12794 ( n12950, n12951, n12952 );
nor U12795 ( n12952, n12953, n12954 );
nand U12796 ( n12954, n12955, n12956 );
nor U12797 ( n12956, n12957, n12958 );
nor U12798 ( n12958, n15083, n12754 );
nor U12799 ( n12957, n15091, n12755 );
nor U12800 ( n12955, n12959, n12960 );
nor U12801 ( n12960, n15075, n12758 );
nor U12802 ( n12959, n15067, n12759 );
nand U12803 ( n12953, n12961, n12962 );
nor U12804 ( n12962, n12963, n12964 );
nand U12805 ( n12964, n12965, n12765 );
nand U12806 ( n12965, n12766, n7867 );
nor U12807 ( n12963, n15115, n12767 );
nor U12808 ( n12961, n12966, n12967 );
nor U12809 ( n12967, n15107, n12770 );
nor U12810 ( n12966, n15099, n12771 );
nor U12811 ( n12951, n12968, n12969 );
nand U12812 ( n12969, n12970, n12971 );
nor U12813 ( n12971, n12972, n12973 );
nor U12814 ( n12973, n15179, n12778 );
nor U12815 ( n12972, n15187, n12779 );
nor U12816 ( n12970, n12974, n12975 );
nor U12817 ( n12975, n15171, n12782 );
nor U12818 ( n12974, n15163, n12783 );
nand U12819 ( n12968, n12976, n12977 );
nor U12820 ( n12977, n12978, n12979 );
nor U12821 ( n12979, n15147, n12788 );
nor U12822 ( n12978, n15155, n12789 );
nor U12823 ( n12976, n12980, n12981 );
nor U12824 ( n12981, n15139, n12792 );
nor U12825 ( n12980, n15131, n12793 );
nand U12826 ( n12948, n12982, n12983 );
nand U12827 ( n12983, n12984, n12985 );
and U12828 ( n12985, n12986, n12987 );
nor U12829 ( n12984, n12988, n12989 );
nor U12830 ( n12988, n12990, n7822 );
nor U12831 ( n12982, n12991, n12992 );
nor U12832 ( n12992, n12993, n12989 );
nand U12833 ( n12989, n12994, n12995 );
nand U12834 ( n12995, n15211, n12996 );
nand U12835 ( n12996, n11887, n12742 );
nor U12836 ( n12993, n12997, n12998 );
nand U12837 ( n12998, n12999, n13000 );
nor U12838 ( n12997, n13001, n13002 );
nand U12839 ( n13002, n12987, n7822 );
not U12840 ( n13001, n12990 );
nor U12841 ( n12940, n12220, n9907 );
nand U12842 ( n9907, n12915, n13003 );
nand U12843 ( n13003, n13004, n13005 );
or U12844 ( n12915, n13005, n13004 );
xnor U12845 ( n13004, n13006, n12254 );
nand U12846 ( n13006, n13007, n13008 );
nand U12847 ( n13008, n12196, n7893 );
nand U12848 ( n13007, n10822, n7922 );
nor U12849 ( n12938, n13009, n13010 );
nand U12850 ( n13010, n13011, n13012 );
nand U12851 ( n13012, n13013, n7922 );
nand U12852 ( n13013, n13014, n13015 );
nand U12853 ( n13015, n15211, n13016 );
nand U12854 ( n13016, n12440, n12336 );
not U12855 ( n13014, n13017 );
nand U12856 ( n13011, n13018, n15212 );
and U12857 ( n13018, n7843, n13019 );
nor U12858 ( n13009, n15331, n12207 );
nand U12859 ( n1290, n13020, n13021 );
nor U12860 ( n13021, n13022, n13023 );
nor U12861 ( n13023, n12220, n9927 );
nand U12862 ( n9927, n13005, n13024 );
nand U12863 ( n13024, n13025, n13026 );
or U12864 ( n13005, n13026, n13025 );
xnor U12865 ( n13025, n13027, n12254 );
nand U12866 ( n13027, n13028, n13029 );
nand U12867 ( n13029, n12196, n7894 );
nand U12868 ( n13028, n10822, n7843 );
nor U12869 ( n13022, n12176, n11894 );
xnor U12870 ( n11894, n13030, n13031 );
nor U12871 ( n13031, n12991, n13032 );
nor U12872 ( n13032, n13033, n7843 );
nor U12873 ( n13033, n12700, n13034 );
and U12874 ( n12991, n13035, n11887 );
not U12875 ( n11887, n13034 );
nand U12876 ( n13034, n12744, n13036 );
nand U12877 ( n13036, n13037, n13038 );
nor U12878 ( n13038, n13039, n13040 );
nand U12879 ( n13040, n13041, n13042 );
nor U12880 ( n13042, n13043, n13044 );
nor U12881 ( n13044, n15084, n12754 );
nor U12882 ( n13043, n15092, n12755 );
nor U12883 ( n13041, n13045, n13046 );
nor U12884 ( n13046, n15076, n12758 );
nor U12885 ( n13045, n15068, n12759 );
nand U12886 ( n13039, n13047, n13048 );
nor U12887 ( n13048, n13049, n13050 );
nand U12888 ( n13050, n13051, n12765 );
nand U12889 ( n13051, n12766, n7868 );
nor U12890 ( n13049, n15116, n12767 );
nor U12891 ( n13047, n13052, n13053 );
nor U12892 ( n13053, n15108, n12770 );
nor U12893 ( n13052, n15100, n12771 );
nor U12894 ( n13037, n13054, n13055 );
nand U12895 ( n13055, n13056, n13057 );
nor U12896 ( n13057, n13058, n13059 );
nor U12897 ( n13059, n15180, n12778 );
nor U12898 ( n13058, n15188, n12779 );
nor U12899 ( n13056, n13060, n13061 );
nor U12900 ( n13061, n15172, n12782 );
nor U12901 ( n13060, n15164, n12783 );
nand U12902 ( n13054, n13062, n13063 );
nor U12903 ( n13063, n13064, n13065 );
nor U12904 ( n13065, n15148, n12788 );
nor U12905 ( n13064, n15156, n12789 );
nor U12906 ( n13062, n13066, n13067 );
nor U12907 ( n13067, n15140, n12792 );
nor U12908 ( n13066, n15132, n12793 );
nor U12909 ( n13035, n15211, n12700 );
nand U12910 ( n13030, n12999, n13068 );
nand U12911 ( n13068, n13069, n12994 );
nor U12912 ( n13020, n13070, n13071 );
nand U12913 ( n13071, n13072, n13073 );
nand U12914 ( n13073, n15211, n13019 );
nand U12915 ( n13019, n13074, n13075 );
nand U12916 ( n13075, n12342, n12935 );
nor U12917 ( n13074, n13076, n13077 );
nor U12918 ( n13077, n13078, n12271 );
nor U12919 ( n13076, n13079, n12347 );
nand U12920 ( n13072, n13017, n7843 );
nand U12921 ( n13017, n13080, n13081 );
nor U12922 ( n13081, n12345, n13082 );
nor U12923 ( n13082, n12937, n12347 );
not U12924 ( n12937, n13079 );
nand U12925 ( n13079, n13083, n13084 );
nor U12926 ( n13080, n13085, n13086 );
nor U12927 ( n13086, n12935, n12336 );
and U12928 ( n12935, n13083, n13087 );
nor U12929 ( n13083, n15022, n15210 );
nor U12930 ( n13085, n12932, n12271 );
not U12931 ( n12932, n13078 );
nand U12932 ( n13078, n13088, n13089 );
nor U12933 ( n13089, n15022, n15209 );
nor U12934 ( n13088, n15210, n13090 );
nor U12935 ( n13070, n15330, n12207 );
nand U12936 ( n1285, n13091, n13092 );
nor U12937 ( n13092, n13093, n13094 );
nor U12938 ( n13094, n12176, n11923 );
xnor U12939 ( n11923, n13069, n13095 );
and U12940 ( n13095, n12994, n12999 );
or U12941 ( n12999, n13096, n15022 );
nand U12942 ( n12994, n15022, n13096 );
nand U12943 ( n13096, n11915, n12742 );
and U12944 ( n11915, n12744, n13097 );
nand U12945 ( n13097, n13098, n13099 );
nor U12946 ( n13099, n13100, n13101 );
nand U12947 ( n13101, n13102, n13103 );
nor U12948 ( n13103, n13104, n13105 );
nor U12949 ( n13105, n15085, n12754 );
nor U12950 ( n13104, n15093, n12755 );
nor U12951 ( n13102, n13106, n13107 );
nor U12952 ( n13107, n15077, n12758 );
nor U12953 ( n13106, n15069, n12759 );
nand U12954 ( n13100, n13108, n13109 );
nor U12955 ( n13109, n13110, n13111 );
nand U12956 ( n13111, n13112, n12765 );
nand U12957 ( n13112, n12766, n7869 );
nor U12958 ( n13110, n15117, n12767 );
nor U12959 ( n13108, n13113, n13114 );
nor U12960 ( n13114, n15109, n12770 );
nor U12961 ( n13113, n15101, n12771 );
nor U12962 ( n13098, n13115, n13116 );
nand U12963 ( n13116, n13117, n13118 );
nor U12964 ( n13118, n13119, n13120 );
nor U12965 ( n13120, n15181, n12778 );
nor U12966 ( n13119, n15189, n12779 );
nor U12967 ( n13117, n13121, n13122 );
nor U12968 ( n13122, n15173, n12782 );
nor U12969 ( n13121, n15165, n12783 );
nand U12970 ( n13115, n13123, n13124 );
nor U12971 ( n13124, n13125, n13126 );
nor U12972 ( n13126, n15149, n12788 );
nor U12973 ( n13125, n15157, n12789 );
nor U12974 ( n13123, n13127, n13128 );
nor U12975 ( n13128, n15141, n12792 );
nor U12976 ( n13127, n15133, n12793 );
nand U12977 ( n13069, n13000, n13129 );
nand U12978 ( n13129, n13130, n12987 );
nor U12979 ( n13093, n12220, n9948 );
nand U12980 ( n9948, n13026, n13131 );
nand U12981 ( n13131, n13132, n13133 );
or U12982 ( n13026, n13133, n13132 );
xnor U12983 ( n13132, n13134, n12254 );
nand U12984 ( n13134, n13135, n13136 );
nand U12985 ( n13136, n12196, n7895 );
nand U12986 ( n13135, n10822, n7920 );
nor U12987 ( n13091, n13137, n13138 );
nand U12988 ( n13138, n13139, n13140 );
nand U12989 ( n13140, n13141, n7920 );
nand U12990 ( n13141, n13142, n13143 );
nand U12991 ( n13143, n15210, n12204 );
not U12992 ( n13142, n13144 );
nand U12993 ( n13139, n13145, n15022 );
and U12994 ( n13145, n7872, n13146 );
nor U12995 ( n13137, n15329, n12207 );
nand U12996 ( n1280, n13147, n13148 );
nor U12997 ( n13148, n13149, n13150 );
nor U12998 ( n13150, n12176, n11943 );
xnor U12999 ( n11943, n13130, n13151 );
and U13000 ( n13151, n12987, n13000 );
nand U13001 ( n13000, n13152, n11912 );
nor U13002 ( n13152, n15210, n12700 );
nand U13003 ( n12987, n15210, n13153 );
nand U13004 ( n13153, n11912, n12742 );
not U13005 ( n11912, n11939 );
nand U13006 ( n11939, n12744, n13154 );
nand U13007 ( n13154, n13155, n13156 );
nor U13008 ( n13156, n13157, n13158 );
nand U13009 ( n13158, n13159, n13160 );
nor U13010 ( n13160, n13161, n13162 );
nor U13011 ( n13162, n15086, n12754 );
nor U13012 ( n13161, n15094, n12755 );
nor U13013 ( n13159, n13163, n13164 );
nor U13014 ( n13164, n15078, n12758 );
nor U13015 ( n13163, n15070, n12759 );
nand U13016 ( n13157, n13165, n13166 );
nor U13017 ( n13166, n13167, n13168 );
nand U13018 ( n13168, n13169, n12765 );
nand U13019 ( n13169, n12766, n7870 );
nor U13020 ( n13167, n15118, n12767 );
nor U13021 ( n13165, n13170, n13171 );
nor U13022 ( n13171, n15110, n12770 );
nor U13023 ( n13170, n15102, n12771 );
nor U13024 ( n13155, n13172, n13173 );
nand U13025 ( n13173, n13174, n13175 );
nor U13026 ( n13175, n13176, n13177 );
nor U13027 ( n13177, n15182, n12778 );
nor U13028 ( n13176, n15190, n12779 );
nor U13029 ( n13174, n13178, n13179 );
nor U13030 ( n13179, n15174, n12782 );
nor U13031 ( n13178, n15166, n12783 );
nand U13032 ( n13172, n13180, n13181 );
nor U13033 ( n13181, n13182, n13183 );
nor U13034 ( n13183, n15150, n12788 );
nor U13035 ( n13182, n15158, n12789 );
nor U13036 ( n13180, n13184, n13185 );
nor U13037 ( n13185, n15142, n12792 );
nor U13038 ( n13184, n15134, n12793 );
nand U13039 ( n13130, n13186, n13187 );
nand U13040 ( n13187, n13188, n7822 );
or U13041 ( n13188, n12986, n12990 );
nand U13042 ( n13186, n12990, n12986 );
nor U13043 ( n13149, n12220, n9969 );
nand U13044 ( n9969, n13133, n13189 );
nand U13045 ( n13189, n13190, n13191 );
or U13046 ( n13133, n13191, n13190 );
xnor U13047 ( n13190, n13192, n12254 );
nand U13048 ( n13192, n13193, n13194 );
nand U13049 ( n13194, n12196, n7896 );
nand U13050 ( n13193, n10822, n7872 );
nor U13051 ( n13147, n13195, n13196 );
nand U13052 ( n13196, n13197, n13198 );
nand U13053 ( n13198, n15210, n13146 );
nand U13054 ( n13146, n13199, n13200 );
nand U13055 ( n13200, n12333, n13084 );
nor U13056 ( n13199, n13201, n13202 );
nor U13057 ( n13202, n13203, n12336 );
nor U13058 ( n13201, n12271, n13204 );
nand U13059 ( n13204, n13205, n7822 );
nand U13060 ( n13197, n13144, n7872 );
nand U13061 ( n13144, n13206, n13207 );
nor U13062 ( n13207, n12345, n13208 );
nor U13063 ( n13208, n13209, n12271 );
nor U13064 ( n13209, n15209, n13090 );
not U13065 ( n13090, n13205 );
nor U13066 ( n13206, n13210, n13211 );
nor U13067 ( n13211, n13084, n12347 );
and U13068 ( n13084, n13212, n13213 );
nor U13069 ( n13212, n15208, n15209 );
nor U13070 ( n13210, n13087, n12336 );
not U13071 ( n13087, n13203 );
nand U13072 ( n13203, n13214, n13215 );
nor U13073 ( n13215, n15207, n15208 );
nor U13074 ( n13214, n15209, n13216 );
nor U13075 ( n13195, n15328, n12207 );
nand U13076 ( n1275, n13217, n13218 );
nor U13077 ( n13218, n13219, n13220 );
nor U13078 ( n13220, n12176, n11962 );
xor U13079 ( n11962, n13221, n12990 );
nand U13080 ( n12990, n13222, n13223 );
nand U13081 ( n13223, n13224, n13225 );
nor U13082 ( n13224, n13226, n13227 );
nand U13083 ( n13222, n11954, n12742 );
and U13084 ( n11954, n12744, n13228 );
nand U13085 ( n13228, n13229, n13230 );
nor U13086 ( n13230, n13231, n13232 );
nand U13087 ( n13232, n13233, n13234 );
nor U13088 ( n13234, n13235, n13236 );
nor U13089 ( n13236, n15087, n12754 );
nand U13090 ( n12754, n13237, n11345 );
nor U13091 ( n13235, n15095, n12755 );
nand U13092 ( n12755, n13237, n11344 );
nor U13093 ( n13233, n13238, n13239 );
nor U13094 ( n13239, n15079, n12758 );
nand U13095 ( n12758, n13237, n11349 );
nor U13096 ( n13238, n15071, n12759 );
nand U13097 ( n12759, n13237, n11348 );
nor U13098 ( n13237, n13240, n13241 );
nand U13099 ( n13231, n13242, n13243 );
nor U13100 ( n13243, n13244, n13245 );
nand U13101 ( n13245, n13246, n12765 );
nand U13102 ( n13246, n12766, n7871 );
and U13103 ( n12766, n13247, n11344 );
nor U13104 ( n13244, n15119, n12767 );
nand U13105 ( n12767, n13247, n11345 );
nor U13106 ( n13242, n13248, n13249 );
nor U13107 ( n13249, n15111, n12770 );
nand U13108 ( n12770, n13247, n11349 );
nor U13109 ( n13248, n15103, n12771 );
nand U13110 ( n12771, n13247, n11348 );
nor U13111 ( n13247, n13250, n13241 );
nor U13112 ( n13229, n13251, n13252 );
nand U13113 ( n13252, n13253, n13254 );
nor U13114 ( n13254, n13255, n13256 );
nor U13115 ( n13256, n15183, n12778 );
nand U13116 ( n12778, n13257, n11345 );
nor U13117 ( n13255, n15191, n12779 );
nand U13118 ( n12779, n13257, n11344 );
nor U13119 ( n13253, n13258, n13259 );
nor U13120 ( n13259, n15175, n12782 );
nand U13121 ( n12782, n13257, n11349 );
nor U13122 ( n13258, n15167, n12783 );
nand U13123 ( n12783, n13257, n11348 );
nor U13124 ( n13257, n13260, n13250 );
nand U13125 ( n13251, n13261, n13262 );
nor U13126 ( n13262, n13263, n13264 );
nor U13127 ( n13264, n15151, n12788 );
nand U13128 ( n12788, n13265, n11345 );
nor U13129 ( n13263, n15159, n12789 );
nand U13130 ( n12789, n13265, n11344 );
nor U13131 ( n13261, n13266, n13267 );
nor U13132 ( n13267, n15143, n12792 );
nand U13133 ( n12792, n13265, n11349 );
nor U13134 ( n13266, n15135, n12793 );
nand U13135 ( n12793, n13265, n11348 );
nor U13136 ( n13265, n13260, n13240 );
and U13137 ( n12744, n13268, n13269 );
nand U13138 ( n13269, n13270, n13271 );
nor U13139 ( n13270, n12698, n9347 );
xor U13140 ( n13221, n12986, n15209 );
nand U13141 ( n12986, n13272, n13273 );
or U13142 ( n13273, n13274, n13275 );
nor U13143 ( n13219, n12220, n9989 );
nand U13144 ( n9989, n13191, n13276 );
nand U13145 ( n13276, n13277, n13278 );
or U13146 ( n13191, n13278, n13277 );
xnor U13147 ( n13277, n13279, n12254 );
nand U13148 ( n13279, n13280, n13281 );
nand U13149 ( n13281, n12196, n7897 );
nand U13150 ( n13280, n10822, n7822 );
nor U13151 ( n13217, n13282, n13283 );
nand U13152 ( n13283, n13284, n13285 );
nand U13153 ( n13285, n13286, n7822 );
nand U13154 ( n13286, n13287, n13288 );
nor U13155 ( n13287, n13289, n13290 );
nor U13156 ( n13290, n12275, n7820 );
nor U13157 ( n13289, n13205, n12271 );
nand U13158 ( n13284, n15209, n13291 );
nand U13159 ( n13291, n13292, n13293 );
nand U13160 ( n13293, n12266, n13205 );
nor U13161 ( n13205, n13294, n15208 );
nand U13162 ( n13292, n13295, n7820 );
nor U13163 ( n13282, n15327, n12207 );
nand U13164 ( n1270, n13296, n13297 );
nor U13165 ( n13297, n13298, n13299 );
nor U13166 ( n13299, n12220, n10010 );
nand U13167 ( n10010, n13278, n13300 );
nand U13168 ( n13300, n13301, n13302 );
or U13169 ( n13278, n13302, n13301 );
xnor U13170 ( n13301, n13303, n12254 );
nand U13171 ( n13303, n13304, n13305 );
nand U13172 ( n13305, n12196, n7898 );
nand U13173 ( n13304, n10822, n7820 );
nor U13174 ( n13298, n12176, n13306 );
nand U13175 ( n13306, n11973, n11972 );
nand U13176 ( n11972, n13307, n13308 );
nor U13177 ( n13308, n13275, n13309 );
nor U13178 ( n13307, n13310, n13311 );
nor U13179 ( n13311, n13312, n13313 );
and U13180 ( n13310, n7820, n13314 );
nand U13181 ( n11973, n13274, n13315 );
nand U13182 ( n13315, n13272, n13316 );
not U13183 ( n13316, n13275 );
nor U13184 ( n13275, n7820, n13314 );
nand U13185 ( n13272, n7820, n13314 );
nand U13186 ( n13314, n13317, n13318 );
nand U13187 ( n13318, n13319, n9393 );
xnor U13188 ( n13319, n13226, n13225 );
nor U13189 ( n13225, n13320, n13321 );
nand U13190 ( n13317, n11979, n12742 );
xor U13191 ( n11979, n13268, n13322 );
nor U13192 ( n13322, n13323, n13324 );
nand U13193 ( n13324, n13325, n12765 );
nand U13194 ( n13325, n13326, n7919 );
nor U13195 ( n13323, n13226, n13327 );
nor U13196 ( n13274, n13312, n13328 );
nor U13197 ( n13328, n13309, n13329 );
nor U13198 ( n13296, n13330, n13331 );
nand U13199 ( n13331, n13332, n13333 );
nand U13200 ( n13333, n15208, n13334 );
nand U13201 ( n13334, n13335, n13336 );
or U13202 ( n13336, n12271, n13294 );
not U13203 ( n13335, n13295 );
nand U13204 ( n13295, n13337, n13338 );
nand U13205 ( n13338, n13339, n12342 );
nand U13206 ( n13337, n12333, n13213 );
not U13207 ( n13213, n13340 );
nand U13208 ( n13332, n13341, n7820 );
nand U13209 ( n13341, n13288, n13342 );
nand U13210 ( n13342, n12266, n13294 );
nand U13211 ( n13294, n13343, n13344 );
and U13212 ( n13288, n13345, n13346 );
nand U13213 ( n13346, n12333, n13340 );
nand U13214 ( n13340, n13347, n13343 );
nor U13215 ( n13343, n15206, n15207 );
nor U13216 ( n13345, n12345, n13348 );
nor U13217 ( n13348, n13339, n12336 );
nor U13218 ( n13339, n15207, n13216 );
not U13219 ( n13216, n13349 );
nor U13220 ( n13330, n15326, n12207 );
nand U13221 ( n1265, n13350, n13351 );
nor U13222 ( n13351, n13352, n13353 );
nor U13223 ( n13353, n12176, n12007 );
xor U13224 ( n12007, n13329, n13354 );
nor U13225 ( n13354, n13309, n13312 );
and U13226 ( n13312, n7844, n13355 );
nor U13227 ( n13309, n7844, n13355 );
nand U13228 ( n13355, n13356, n13357 );
nand U13229 ( n13357, n13358, n12742 );
nor U13230 ( n13358, n12699, n12004 );
and U13231 ( n12004, n13359, n13360 );
nand U13232 ( n13360, n13361, n13362 );
not U13233 ( n12699, n13268 );
nand U13234 ( n13268, n13363, n13361 );
nor U13235 ( n13363, n13364, n13359 );
and U13236 ( n13359, n13365, n13366 );
nand U13237 ( n13366, n13367, n13368 );
nand U13238 ( n13365, n13326, n7858 );
not U13239 ( n13364, n13362 );
nand U13240 ( n13356, n13369, n9393 );
xor U13241 ( n13369, n13320, n13321 );
not U13242 ( n13321, n13367 );
nand U13243 ( n13367, n13370, n13371 );
nor U13244 ( n13371, n13372, n13373 );
nand U13245 ( n13373, n13374, n13375 );
nor U13246 ( n13375, n13376, n13377 );
nor U13247 ( n13377, n15145, n13378 );
nor U13248 ( n13376, n15153, n13379 );
nor U13249 ( n13374, n13380, n13381 );
nor U13250 ( n13381, n15137, n13382 );
nor U13251 ( n13380, n15129, n13383 );
nand U13252 ( n13372, n13384, n13385 );
nor U13253 ( n13385, n13386, n13387 );
nor U13254 ( n13387, n15177, n13388 );
nor U13255 ( n13386, n15185, n13389 );
nor U13256 ( n13384, n13390, n13391 );
nor U13257 ( n13391, n15169, n13392 );
nor U13258 ( n13390, n15161, n13393 );
nor U13259 ( n13370, n13394, n13395 );
nand U13260 ( n13395, n13396, n13397 );
nor U13261 ( n13397, n13398, n13399 );
nor U13262 ( n13399, n15113, n13400 );
nor U13263 ( n13398, n15121, n13401 );
nor U13264 ( n13396, n13402, n13403 );
nor U13265 ( n13403, n15105, n13404 );
nor U13266 ( n13402, n15097, n13405 );
nand U13267 ( n13394, n13406, n13407 );
nor U13268 ( n13407, n13408, n13409 );
nor U13269 ( n13409, n15081, n13410 );
nor U13270 ( n13408, n15089, n13411 );
nor U13271 ( n13406, n13412, n13413 );
nor U13272 ( n13413, n15073, n13414 );
nor U13273 ( n13412, n15065, n13415 );
nand U13274 ( n13320, n13416, n13417 );
not U13275 ( n13329, n13313 );
nand U13276 ( n13313, n13418, n13419 );
nand U13277 ( n13419, n13420, n13421 );
nor U13278 ( n13352, n12220, n10031 );
nand U13279 ( n10031, n13302, n13422 );
nand U13280 ( n13422, n13423, n13424 );
or U13281 ( n13302, n13424, n13423 );
xnor U13282 ( n13423, n13425, n12254 );
nand U13283 ( n13425, n13426, n13427 );
nand U13284 ( n13427, n12196, n7899 );
nand U13285 ( n13426, n10822, n7844 );
nor U13286 ( n13350, n13428, n13429 );
nand U13287 ( n13429, n13430, n13431 );
nand U13288 ( n13431, n13432, n7844 );
nand U13289 ( n13432, n13433, n13434 );
nor U13290 ( n13433, n13435, n13436 );
nor U13291 ( n13436, n12440, n7827 );
nor U13292 ( n13435, n13349, n12336 );
nand U13293 ( n13430, n15207, n13437 );
nand U13294 ( n13437, n13438, n13439 );
nand U13295 ( n13439, n12342, n13349 );
nor U13296 ( n13349, n13440, n15206 );
nand U13297 ( n13438, n13441, n7827 );
nor U13298 ( n13428, n15325, n12207 );
nand U13299 ( n1260, n13442, n13443 );
nor U13300 ( n13443, n13444, n13445 );
nor U13301 ( n13445, n12176, n12030 );
xnor U13302 ( n12030, n13420, n13446 );
and U13303 ( n13446, n13421, n13418 );
nand U13304 ( n13418, n7827, n13447 );
or U13305 ( n13421, n7827, n13447 );
nand U13306 ( n13447, n13448, n13449 );
nand U13307 ( n13449, n13450, n9393 );
xor U13308 ( n13450, n13417, n13416 );
nor U13309 ( n13416, n13451, n13452 );
nand U13310 ( n13448, n12021, n12742 );
xor U13311 ( n12021, n13361, n13362 );
nand U13312 ( n13362, n13453, n13454 );
nand U13313 ( n13454, n13368, n13417 );
nand U13314 ( n13417, n13455, n13456 );
nor U13315 ( n13456, n13457, n13458 );
nand U13316 ( n13458, n13459, n13460 );
nor U13317 ( n13460, n13461, n13462 );
nor U13318 ( n13462, n15146, n13378 );
nor U13319 ( n13461, n15154, n13379 );
nor U13320 ( n13459, n13463, n13464 );
nor U13321 ( n13464, n15138, n13382 );
nor U13322 ( n13463, n15130, n13383 );
nand U13323 ( n13457, n13465, n13466 );
nor U13324 ( n13466, n13467, n13468 );
nor U13325 ( n13468, n15178, n13388 );
nor U13326 ( n13467, n15186, n13389 );
nor U13327 ( n13465, n13469, n13470 );
nor U13328 ( n13470, n15170, n13392 );
nor U13329 ( n13469, n15162, n13393 );
nor U13330 ( n13455, n13471, n13472 );
nand U13331 ( n13472, n13473, n13474 );
nor U13332 ( n13474, n13475, n13476 );
nor U13333 ( n13476, n15114, n13400 );
nor U13334 ( n13475, n15122, n13401 );
nor U13335 ( n13473, n13477, n13478 );
nor U13336 ( n13478, n15106, n13404 );
nor U13337 ( n13477, n15098, n13405 );
nand U13338 ( n13471, n13479, n13480 );
nor U13339 ( n13480, n13481, n13482 );
nor U13340 ( n13482, n15082, n13410 );
nor U13341 ( n13481, n15090, n13411 );
nor U13342 ( n13479, n13483, n13484 );
nor U13343 ( n13484, n15074, n13414 );
nor U13344 ( n13483, n15066, n13415 );
nand U13345 ( n13453, n13326, n7857 );
nor U13346 ( n13361, n13485, n13486 );
nand U13347 ( n13420, n13487, n13488 );
nand U13348 ( n13488, n13489, n7832 );
nor U13349 ( n13444, n12220, n10052 );
nand U13350 ( n10052, n13424, n13490 );
nand U13351 ( n13490, n13491, n13492 );
or U13352 ( n13424, n13492, n13491 );
xnor U13353 ( n13491, n13493, n12254 );
nand U13354 ( n13493, n13494, n13495 );
nand U13355 ( n13495, n12196, n7900 );
nand U13356 ( n13494, n10822, n7827 );
nor U13357 ( n13442, n13496, n13497 );
nand U13358 ( n13497, n13498, n13499 );
nand U13359 ( n13499, n15206, n13500 );
nand U13360 ( n13500, n13501, n13502 );
or U13361 ( n13502, n12336, n13440 );
not U13362 ( n13501, n13441 );
nand U13363 ( n13441, n13503, n13504 );
nand U13364 ( n13504, n13347, n12333 );
nand U13365 ( n13503, n12266, n13344 );
nand U13366 ( n13498, n13505, n7827 );
nand U13367 ( n13505, n13434, n13506 );
nand U13368 ( n13506, n12342, n13440 );
nand U13369 ( n13440, n13507, n13508 );
not U13370 ( n13507, n13509 );
and U13371 ( n13434, n13510, n13511 );
or U13372 ( n13511, n12271, n13344 );
nor U13373 ( n13344, n13509, n13512 );
nor U13374 ( n13510, n12345, n13513 );
nor U13375 ( n13513, n13347, n12347 );
nor U13376 ( n13347, n13514, n13509 );
nand U13377 ( n13509, n7808, n7832 );
nor U13378 ( n13496, n15324, n12207 );
nand U13379 ( n1255, n13515, n13516 );
nor U13380 ( n13516, n13517, n13518 );
nor U13381 ( n13518, n12176, n12062 );
nand U13382 ( n12062, n13519, n13520 );
nand U13383 ( n13520, n13521, n13522 );
nor U13384 ( n13519, n13523, n13524 );
nor U13385 ( n13524, n13525, n7832 );
nor U13386 ( n13525, n13526, n13521 );
not U13387 ( n13521, n13487 );
nand U13388 ( n13487, n13527, n13528 );
nand U13389 ( n13527, n15023, n13522 );
nor U13390 ( n13526, n13489, n13528 );
nor U13391 ( n13523, n15023, n13529 );
or U13392 ( n13529, n13528, n13522 );
not U13393 ( n13522, n13489 );
nand U13394 ( n13489, n13530, n13531 );
nand U13395 ( n13531, n13532, n9393 );
xor U13396 ( n13532, n13451, n13452 );
not U13397 ( n13452, n13533 );
nand U13398 ( n13530, n12041, n12742 );
xor U13399 ( n12041, n13485, n13486 );
and U13400 ( n13486, n13534, n13535 );
nand U13401 ( n13535, n13533, n13368 );
nand U13402 ( n13368, n13536, n13327 );
nor U13403 ( n13536, n12698, n13537 );
nand U13404 ( n13533, n13538, n13539 );
nor U13405 ( n13539, n13540, n13541 );
nand U13406 ( n13541, n13542, n13543 );
nor U13407 ( n13543, n13544, n13545 );
nor U13408 ( n13545, n15147, n13378 );
nor U13409 ( n13544, n15155, n13379 );
nor U13410 ( n13542, n13546, n13547 );
nor U13411 ( n13547, n15139, n13382 );
nor U13412 ( n13546, n15131, n13383 );
nand U13413 ( n13540, n13548, n13549 );
nor U13414 ( n13549, n13550, n13551 );
nor U13415 ( n13551, n15179, n13388 );
nor U13416 ( n13550, n15187, n13389 );
nor U13417 ( n13548, n13552, n13553 );
nor U13418 ( n13553, n15171, n13392 );
nor U13419 ( n13552, n15163, n13393 );
nor U13420 ( n13538, n13554, n13555 );
nand U13421 ( n13555, n13556, n13557 );
nor U13422 ( n13557, n13558, n13559 );
nor U13423 ( n13559, n15115, n13400 );
nor U13424 ( n13558, n15123, n13401 );
nor U13425 ( n13556, n13560, n13561 );
nor U13426 ( n13561, n15107, n13404 );
nor U13427 ( n13560, n15099, n13405 );
nand U13428 ( n13554, n13562, n13563 );
nor U13429 ( n13563, n13564, n13565 );
nor U13430 ( n13565, n15083, n13410 );
nor U13431 ( n13564, n15091, n13411 );
nor U13432 ( n13562, n13566, n13567 );
nor U13433 ( n13567, n15075, n13414 );
nor U13434 ( n13566, n15067, n13415 );
nand U13435 ( n13534, n13326, n7856 );
nand U13436 ( n13485, n13568, n13569 );
nor U13437 ( n13568, n13570, n13571 );
nand U13438 ( n13528, n13572, n13573 );
nand U13439 ( n13573, n13574, n7808 );
nand U13440 ( n13574, n13575, n13576 );
or U13441 ( n13572, n13576, n13575 );
not U13442 ( n13575, n13577 );
nor U13443 ( n13517, n12220, n10075 );
nand U13444 ( n10075, n13492, n13578 );
nand U13445 ( n13578, n13579, n13580 );
or U13446 ( n13492, n13580, n13579 );
xnor U13447 ( n13579, n13581, n12254 );
nand U13448 ( n13581, n13582, n13583 );
nand U13449 ( n13583, n12196, n7901 );
nand U13450 ( n13582, n10822, n7832 );
nor U13451 ( n13515, n13584, n13585 );
nand U13452 ( n13585, n13586, n13587 );
nand U13453 ( n13587, n13588, n7832 );
nand U13454 ( n13588, n13589, n13590 );
nand U13455 ( n13590, n15205, n12204 );
nand U13456 ( n12204, n12275, n12271 );
not U13457 ( n12275, n13591 );
not U13458 ( n13589, n13592 );
nand U13459 ( n13586, n13593, n15023 );
and U13460 ( n13593, n7808, n13594 );
nor U13461 ( n13584, n15323, n12207 );
nand U13462 ( n1250, n13595, n13596 );
nor U13463 ( n13596, n13597, n13598 );
nor U13464 ( n13598, n12220, n10099 );
nand U13465 ( n10099, n13580, n13599 );
nand U13466 ( n13599, n13600, n13601 );
or U13467 ( n13580, n13601, n13600 );
xnor U13468 ( n13600, n13602, n12254 );
nand U13469 ( n13602, n13603, n13604 );
nand U13470 ( n13604, n12196, n7902 );
nand U13471 ( n13603, n10822, n7808 );
or U13472 ( n13601, n13605, n13606 );
nor U13473 ( n13597, n12176, n12083 );
xor U13474 ( n12083, n13576, n13607 );
xor U13475 ( n13607, n7808, n13577 );
nand U13476 ( n13577, n13608, n13609 );
nand U13477 ( n13609, n13610, n9393 );
nor U13478 ( n13610, n13611, n13612 );
nor U13479 ( n13612, n13613, n13614 );
not U13480 ( n13611, n13451 );
nand U13481 ( n13451, n13614, n13613 );
nand U13482 ( n13608, n12075, n12742 );
nand U13483 ( n13576, n13615, n13616 );
nand U13484 ( n13616, n15204, n13617 );
nand U13485 ( n13617, n13618, n13619 );
or U13486 ( n13615, n13618, n13619 );
nor U13487 ( n13595, n13620, n13621 );
nand U13488 ( n13621, n13622, n13623 );
nand U13489 ( n13623, n15205, n13594 );
nand U13490 ( n13594, n13624, n13625 );
nand U13491 ( n13625, n12342, n13508 );
nor U13492 ( n13624, n13626, n13627 );
nor U13493 ( n13627, n13514, n12347 );
nor U13494 ( n13626, n13512, n12271 );
nand U13495 ( n13622, n13592, n7808 );
nand U13496 ( n13592, n13628, n13629 );
nor U13497 ( n13629, n12345, n13630 );
nor U13498 ( n13630, n13631, n12271 );
nor U13499 ( n13628, n13632, n13633 );
nor U13500 ( n13633, n12336, n13508 );
and U13501 ( n13632, n13514, n12333 );
nor U13502 ( n13620, n15322, n12207 );
nand U13503 ( n1245, n13634, n13635 );
nor U13504 ( n13635, n13636, n13637 );
nand U13505 ( n13637, n13638, n13639 );
nand U13506 ( n13639, n12342, n13640 );
nand U13507 ( n13640, n13508, n13514 );
nand U13508 ( n13514, n13631, n7817 );
not U13509 ( n13631, n13512 );
nand U13510 ( n13512, n7806, n7853 );
nand U13511 ( n13508, n15204, n13641 );
nand U13512 ( n13641, n7806, n7817 );
not U13513 ( n12342, n12336 );
nand U13514 ( n13638, n10119, n12188 );
xor U13515 ( n10119, n13605, n13606 );
xnor U13516 ( n13606, n13642, n12254 );
nand U13517 ( n13642, n13643, n13644 );
nand U13518 ( n13644, n12196, n7903 );
nand U13519 ( n13643, n10822, n7853 );
nor U13520 ( n13636, n12176, n12107 );
xor U13521 ( n12107, n13645, n13619 );
nand U13522 ( n13619, n13646, n13647 );
nor U13523 ( n13646, n13648, n13649 );
nor U13524 ( n13649, n9077, n12700 );
nor U13525 ( n13648, n13650, n13227 );
nor U13526 ( n13650, n13651, n13652 );
not U13527 ( n13652, n13614 );
nand U13528 ( n13614, n13653, n13654 );
nor U13529 ( n13651, n13653, n13654 );
nand U13530 ( n13654, n13655, n13656 );
xor U13531 ( n13645, n13618, n15204 );
nand U13532 ( n13618, n13657, n13658 );
nand U13533 ( n13658, n13659, n7806 );
or U13534 ( n13659, n13660, n13661 );
nand U13535 ( n13657, n13661, n13660 );
nor U13536 ( n13634, n13662, n13663 );
nand U13537 ( n13663, n13664, n13665 );
nand U13538 ( n13665, n13666, n7853 );
nand U13539 ( n13666, n13667, n13668 );
nand U13540 ( n13668, n12333, n15202 );
nor U13541 ( n13667, n12345, n13669 );
nor U13542 ( n13669, n12440, n7806 );
nor U13543 ( n12440, n12333, n12266 );
not U13544 ( n12333, n12347 );
nand U13545 ( n13664, n13670, n15204 );
nor U13546 ( n13670, n15203, n13671 );
nor U13547 ( n13671, n13672, n12266 );
not U13548 ( n12266, n12271 );
nor U13549 ( n13672, n15202, n12347 );
nor U13550 ( n13662, n15321, n12207 );
nand U13551 ( n1240, n13673, n13674 );
nor U13552 ( n13674, n13675, n13676 );
nor U13553 ( n13676, n12176, n12114 );
xor U13554 ( n12114, n13660, n13677 );
xor U13555 ( n13677, n15203, n13661 );
nor U13556 ( n13661, n13678, n15202 );
nand U13557 ( n13660, n13679, n13680 );
nor U13558 ( n13680, n9427, n13681 );
nor U13559 ( n13681, n12700, n13682 );
nor U13560 ( n13679, n12155, n13683 );
nand U13561 ( n13683, n13684, n13685 );
nand U13562 ( n13685, n13686, n13656 );
nand U13563 ( n13684, n13687, n13688 );
nor U13564 ( n13687, n13689, n13227 );
nor U13565 ( n13675, n12220, n10138 );
nand U13566 ( n10138, n13605, n13690 );
nand U13567 ( n13690, n13691, n13692 );
or U13568 ( n13605, n13692, n13691 );
and U13569 ( n13691, n10825, n13693 );
xnor U13570 ( n13692, n13694, n12254 );
nand U13571 ( n13694, n13695, n13696 );
nand U13572 ( n13696, n12196, n7904 );
nand U13573 ( n13695, n10822, n7806 );
nor U13574 ( n13673, n13697, n13698 );
nand U13575 ( n13698, n13699, n13700 );
nand U13576 ( n13700, n15203, n13701 );
nand U13577 ( n13701, n12271, n13702 );
nand U13578 ( n13702, n13591, n7817 );
nand U13579 ( n13699, n13703, n7806 );
nand U13580 ( n13703, n12409, n13704 );
nor U13581 ( n13697, n15320, n12207 );
nand U13582 ( n1235, n13705, n13706 );
nor U13583 ( n13706, n13707, n13708 );
nor U13584 ( n13708, n12220, n10166 );
xor U13585 ( n10166, n12196, n13693 );
xnor U13586 ( n13693, n13709, n12254 );
nand U13587 ( n13709, n13710, n13711 );
nand U13588 ( n13711, n12196, n7905 );
nand U13589 ( n13710, n10822, n7817 );
nand U13590 ( n13712, n13713, n9424 );
nand U13591 ( n12188, n13714, n13715 );
nand U13592 ( n13715, n13716, n9422 );
nand U13593 ( n13714, n13717, n10711 );
not U13594 ( n10711, n9173 );
nand U13595 ( n9173, n9440, n9393 );
nor U13596 ( n13707, n12176, n12139 );
xor U13597 ( n12139, n7817, n13678 );
and U13598 ( n13678, n13718, n13647 );
nand U13599 ( n13647, n9139, n10569 );
nor U13600 ( n13718, n13686, n13719 );
nor U13601 ( n13719, n12162, n12700 );
nor U13602 ( n13686, n13655, n13227 );
nand U13603 ( n13721, n13716, n10568 );
and U13604 ( n13716, n13722, n12168 );
not U13605 ( n12168, n12049 );
nand U13606 ( n12049, n13723, n7797 );
nor U13607 ( n13722, n12345, n13724 );
nand U13608 ( n13720, n13717, n13725 );
nand U13609 ( n13725, n13726, n13727 );
nor U13610 ( n13727, n9411, n13728 );
nor U13611 ( n13726, n13729, n10559 );
nor U13612 ( n10559, n10198, n10177 );
nor U13613 ( n13729, n13730, n9140 );
nor U13614 ( n13730, n13731, n13732 );
nor U13615 ( n13732, n12155, n13227 );
nor U13616 ( n13731, n9363, n13733 );
nand U13617 ( n13733, n13734, n9424 );
nor U13618 ( n13705, n13735, n13736 );
nand U13619 ( n13736, n13737, n13704 );
nand U13620 ( n13704, n15202, n13591 );
nand U13621 ( n13591, n12336, n12347 );
nand U13622 ( n12347, n13717, n13738 );
nand U13623 ( n13738, n13739, n13740 );
not U13624 ( n13740, n13741 );
nor U13625 ( n13739, n13742, n13743 );
nor U13626 ( n13743, n13744, n13724 );
not U13627 ( n13742, n13745 );
nand U13628 ( n12336, n13717, n11726 );
nand U13629 ( n13737, n13746, n7817 );
nand U13630 ( n13746, n12409, n12271 );
nand U13631 ( n12271, n13717, n10199 );
not U13632 ( n10199, n9418 );
nor U13633 ( n13717, n12345, n15061 );
not U13634 ( n12345, n12409 );
nor U13635 ( n13735, n15319, n12207 );
nand U13636 ( n12409, n13747, n13748 );
nor U13637 ( n13748, n13749, n13750 );
nor U13638 ( n13750, n13751, n10708 );
nand U13639 ( n10708, n9098, n9415 );
not U13640 ( n9098, n9109 );
nor U13641 ( n13751, n13752, n13753 );
nor U13642 ( n13753, READY_N, n13754 );
nor U13643 ( n13754, n13755, n13756 );
nor U13644 ( n13756, n13734, n10710 );
nor U13645 ( n13755, n13757, n10198 );
nor U13646 ( n13757, n9395, n10825 );
nor U13647 ( n13752, n13758, n10570 );
nor U13648 ( n13758, n13723, n9139 );
nor U13649 ( n13749, n9350, n13759 );
nand U13650 ( n13759, n13326, n10555 );
nor U13651 ( n13747, n13760, n10190 );
nor U13652 ( n10190, n7797, n12148 );
nor U13653 ( n13760, n13761, n9109 );
nor U13654 ( n13761, n13762, n13763 );
nand U13655 ( n13763, n13764, n13765 );
nand U13656 ( n13765, n13766, n10825 );
nor U13657 ( n13766, n10573, n9415 );
nand U13658 ( n13764, n13767, n10822 );
nor U13659 ( n13767, n9349, n13768 );
nand U13660 ( n13768, n10570, n9106 );
not U13661 ( n9106, READY_N );
nand U13662 ( n1230, n13769, n13770 );
nand U13663 ( n13770, n13771, n7803 );
nand U13664 ( n13769, n13772, n13773 );
nand U13665 ( n13772, n13774, n13775 );
nand U13666 ( n13775, n9383, n13776 );
nor U13667 ( n13774, n13777, n13778 );
nor U13668 ( n13778, n9386, n9087 );
nor U13669 ( n13777, n13779, n13780 );
nand U13670 ( n1225, n13781, n13782 );
nand U13671 ( n13782, n13771, n7825 );
nand U13672 ( n13781, n13783, n13773 );
nand U13673 ( n13783, n13784, n13785 );
nand U13674 ( n13785, n8231, n12119 );
nor U13675 ( n13784, n13786, n13787 );
nor U13676 ( n13787, n13779, n8490 );
nor U13677 ( n13786, n13788, n13789 );
nor U13678 ( n13788, n8242, n8324 );
nand U13679 ( n1220, n13790, n13791 );
nand U13680 ( n13791, n13771, n7826 );
nand U13681 ( n13790, n13792, n13773 );
nand U13682 ( n13792, n13793, n13794 );
nand U13683 ( n13794, n8231, n13795 );
nor U13684 ( n13793, n13796, n13797 );
nor U13685 ( n13797, n13779, n9070 );
nor U13686 ( n13796, n13798, n13789 );
xor U13687 ( n13798, n13799, n8747 );
nand U13688 ( n1215, n13800, n13801 );
nand U13689 ( n13801, n13771, n7804 );
not U13690 ( n13771, n13773 );
nand U13691 ( n13800, n13802, n13773 );
nand U13692 ( n13802, n13803, n13804 );
nand U13693 ( n13804, n8231, n12075 );
nor U13694 ( n13803, n13805, n13806 );
nor U13695 ( n13806, n13779, n8737 );
nor U13696 ( n13779, n7815, n15062 );
nor U13697 ( n13805, n13807, n13789 );
nor U13698 ( n13807, n13808, n13809 );
not U13699 ( n13809, n8333 );
nand U13700 ( n8333, n9078, n8748 );
nor U13701 ( n13808, n8748, n9078 );
nor U13702 ( n9078, n13799, n8990 );
not U13703 ( n8748, n9079 );
nor U13704 ( n1210, n15197, n13773 );
nand U13705 ( n13773, n13810, n13811 );
nand U13706 ( n13811, n13812, n9087 );
nand U13707 ( n9087, n13813, n13814 );
nand U13708 ( n13814, n13815, n9168 );
nand U13709 ( n9168, n13816, n13817 );
nand U13710 ( n13817, n13818, n7816 );
nand U13711 ( n13816, n15062, n9152 );
nand U13712 ( n9152, n13819, n13820 );
nand U13713 ( n13820, n13821, n7816 );
nand U13714 ( n13819, n13822, n9167 );
and U13715 ( n13815, n11773, n9169 );
nand U13716 ( n9169, n13823, n13824 );
nand U13717 ( n13824, n13818, n7800 );
nand U13718 ( n13823, n15062, n9157 );
nand U13719 ( n9157, n13825, n13826 );
nand U13720 ( n13826, n13821, n7800 );
nand U13721 ( n13825, n13827, n9167 );
not U13722 ( n13813, n9143 );
nand U13723 ( n9143, n13828, n13829 );
nand U13724 ( n13829, n15062, n13830 );
nand U13725 ( n13830, n13831, n13832 );
nand U13726 ( n13832, n10092, n9411 );
nand U13727 ( n13831, n13821, n7831 );
nand U13728 ( n13828, n13818, n7831 );
nor U13729 ( n13818, n7813, n15062 );
not U13730 ( n13812, n9086 );
nor U13731 ( n13810, n13833, n13834 );
nand U13732 ( n1205, n13835, n13836 );
nand U13733 ( n13836, n13837, n7798 );
nand U13734 ( n13835, n13838, n13839 );
nand U13735 ( n13838, n13840, n13841 );
nand U13736 ( n13841, n15202, n7799 );
nor U13737 ( n13840, n13842, n13843 );
and U13738 ( n13843, n15196, n9096 );
and U13739 ( n13842, n9161, n9105 );
nand U13740 ( n9161, n13844, n13845 );
nand U13741 ( n13845, n10178, n13846 );
not U13742 ( n10178, n13780 );
nor U13743 ( n13844, n13847, n13848 );
nor U13744 ( n13848, n7798, n10573 );
nor U13745 ( n13847, n15196, n9418 );
nand U13746 ( n1200, n13849, n13850 );
nand U13747 ( n13850, n13837, n7821 );
nand U13748 ( n13849, n13851, n13839 );
nand U13749 ( n13851, n13852, n13853 );
nand U13750 ( n13853, n9096, n13854 );
nor U13751 ( n13852, n13855, n13856 );
and U13752 ( n13856, n9166, n9105 );
nand U13753 ( n9166, n13857, n13858 );
nand U13754 ( n13858, n11727, n13854 );
nor U13755 ( n13857, n13859, n13860 );
nor U13756 ( n13860, n7821, n9418 );
nor U13757 ( n13859, n13861, n8490 );
nor U13758 ( n13855, n13862, n13863 );
nand U13759 ( n1195, n13864, n13865 );
nand U13760 ( n13865, n13837, n7800 );
nand U13761 ( n13864, n13866, n13839 );
nand U13762 ( n13866, n13867, n13868 );
nand U13763 ( n13868, n9096, n13869 );
nor U13764 ( n13867, n13870, n13871 );
and U13765 ( n13871, n13827, n9105 );
nand U13766 ( n13827, n13872, n13873 );
nor U13767 ( n13873, n13874, n13875 );
nor U13768 ( n13875, n13745, n13876 );
nor U13769 ( n13874, n13877, n13869 );
nor U13770 ( n13872, n13878, n13879 );
nor U13771 ( n13879, n13861, n9070 );
nor U13772 ( n13878, n13240, n9418 );
not U13773 ( n13240, n13250 );
xnor U13774 ( n13250, n7821, n15194 );
nor U13775 ( n13870, n13880, n13863 );
nand U13776 ( n13863, n7817, n7799 );
not U13777 ( n13880, n13862 );
xnor U13778 ( n13862, n7834, n15203 );
nand U13779 ( n1190, n13881, n13882 );
nand U13780 ( n13882, n13837, n7816 );
nand U13781 ( n13881, n13883, n13839 );
nand U13782 ( n13883, n13884, n13885 );
nand U13783 ( n13885, n9105, n13822 );
nand U13784 ( n13822, n13886, n13887 );
nor U13785 ( n13887, n13888, n13889 );
nor U13786 ( n13889, n13890, n13745 );
nand U13787 ( n13745, n13891, n13892 );
nor U13788 ( n13888, n13893, n13894 );
or U13789 ( n13894, n13877, n13895 );
nor U13790 ( n13877, n13728, n11726 );
nand U13791 ( n13893, n13896, n13897 );
nand U13792 ( n13897, n11345, n7816 );
nand U13793 ( n13896, n13898, n13899 );
nor U13794 ( n13886, n13900, n13901 );
nor U13795 ( n13901, n13241, n9418 );
not U13796 ( n13241, n13260 );
nand U13797 ( n13260, n13902, n11377 );
nor U13798 ( n13902, n13903, n13904 );
nor U13799 ( n13904, n15195, n11376 );
nor U13800 ( n13903, n15193, n7821 );
nor U13801 ( n13900, n13861, n8737 );
not U13802 ( n8737, n10107 );
not U13803 ( n13861, n13846 );
nand U13804 ( n13846, n13905, n13906 );
nor U13805 ( n13906, n9411, n9440 );
not U13806 ( n9411, n13907 );
nor U13807 ( n13905, n13908, n13741 );
nand U13808 ( n13741, n13909, n13910 );
and U13809 ( n13910, n13911, n13912 );
nor U13810 ( n13909, n13913, n13914 );
nand U13811 ( n13914, n13915, n13916 );
nand U13812 ( n13915, n12155, n9424 );
nor U13813 ( n13913, n13917, n9363 );
nand U13814 ( n13884, n9096, n13918 );
nand U13815 ( n1185, n13919, n13920 );
nand U13816 ( n13920, n13837, n7831 );
not U13817 ( n13837, n13839 );
nand U13818 ( n13919, n13921, n13839 );
nand U13819 ( n13839, n13922, n13923 );
nand U13820 ( n13923, n15063, n7815 );
nor U13821 ( n13922, n13833, n13924 );
nor U13822 ( n13924, n13821, n9109 );
nand U13823 ( n9109, n9120, n7814 );
not U13824 ( n13821, n9167 );
nand U13825 ( n9167, n13925, n13926 );
nor U13826 ( n13926, n13927, n13928 );
nand U13827 ( n13928, n13929, n13911 );
nand U13828 ( n13911, n13930, n10555 );
nor U13829 ( n13930, n9422, n9139 );
nand U13830 ( n13929, n10179, n13734 );
nor U13831 ( n13927, READY_N, n13931 );
nor U13832 ( n13931, n13932, n13933 );
nor U13833 ( n13933, n13907, n9349 );
nand U13834 ( n9349, n13934, n13935 );
nand U13835 ( n13935, n13936, n13937 );
nor U13836 ( n13937, n13938, n13939 );
nor U13837 ( n13936, n13940, n13941 );
not U13838 ( n13940, n13942 );
nor U13839 ( n13932, n9428, n13943 );
nor U13840 ( n13943, n13944, n13945 );
nor U13841 ( n13945, n9418, n10710 );
not U13842 ( n10710, n9395 );
nand U13843 ( n9418, n10179, n9348 );
nor U13844 ( n10179, n10822, n9424 );
nor U13845 ( n13944, n9434, n10198 );
nor U13846 ( n9434, n10160, n9395 );
nor U13847 ( n9395, n7805, n13946 );
nor U13848 ( n13925, n13762, n13947 );
nand U13849 ( n13947, n10363, n13948 );
nand U13850 ( n13948, n13728, n9415 );
not U13851 ( n13728, n9419 );
nand U13852 ( n9419, n13949, n11727 );
nor U13853 ( n13949, n13713, n9435 );
nand U13854 ( n10363, n9428, n11726 );
not U13855 ( n11726, n9429 );
nand U13856 ( n9429, n13950, n11727 );
not U13857 ( n11727, n10573 );
nand U13858 ( n10573, n13891, n13734 );
nor U13859 ( n13950, n9139, n9363 );
nand U13860 ( n13762, n13951, n13912 );
nand U13861 ( n13912, n9393, n13952 );
nand U13862 ( n13952, n13953, n10555 );
nor U13863 ( n13951, n13954, n13955 );
nor U13864 ( n13955, n13956, n10570 );
nor U13865 ( n13956, n13957, n13958 );
nor U13866 ( n13957, n13891, n9424 );
nor U13867 ( n13954, n13734, n13959 );
nor U13868 ( n13959, n9424, n13960 );
nor U13869 ( n13833, n9086, n15024 );
nand U13870 ( n9086, n9125, n7814 );
not U13871 ( n9125, n9386 );
nand U13872 ( n9386, n7797, n7799 );
nor U13873 ( n13921, n13907, n13961 );
nand U13874 ( n13961, n10092, n9105 );
xor U13875 ( n10092, n13962, n15192 );
nand U13876 ( n13962, n13963, n13964 );
nand U13877 ( n1180, n13965, n13966 );
nor U13878 ( n13966, n13967, n13968 );
nand U13879 ( n13968, n13969, n13970 );
nand U13880 ( n13970, n8131, n13971 );
nand U13881 ( n13969, n13972, n7916 );
nor U13882 ( n13967, n8135, n13973 );
nor U13883 ( n13965, n13974, n13975 );
nor U13884 ( n13975, n8139, n13976 );
nor U13885 ( n13974, n8141, n13977 );
nand U13886 ( n1175, n13978, n13979 );
nor U13887 ( n13979, n13980, n13981 );
nand U13888 ( n13981, n13982, n13983 );
nand U13889 ( n13983, n8148, n13971 );
nand U13890 ( n13982, n13972, n7917 );
nor U13891 ( n13980, n8149, n13973 );
nor U13892 ( n13978, n13984, n13985 );
nor U13893 ( n13985, n8152, n13976 );
nor U13894 ( n13984, n8153, n13977 );
nand U13895 ( n1170, n13986, n13987 );
nor U13896 ( n13987, n13988, n13989 );
nand U13897 ( n13989, n13990, n13991 );
nand U13898 ( n13991, n8160, n13971 );
nand U13899 ( n13990, n13972, n7859 );
nor U13900 ( n13988, n8161, n13973 );
nor U13901 ( n13986, n13992, n13993 );
nor U13902 ( n13993, n8164, n13976 );
nor U13903 ( n13992, n8165, n13977 );
nand U13904 ( n1165, n13994, n13995 );
nor U13905 ( n13995, n13996, n13997 );
nand U13906 ( n13997, n13998, n13999 );
nand U13907 ( n13999, n8172, n13971 );
nand U13908 ( n13998, n13972, n7918 );
nor U13909 ( n13996, n8173, n13973 );
nor U13910 ( n13994, n14000, n14001 );
nor U13911 ( n14001, n8176, n13976 );
nor U13912 ( n14000, n8177, n13977 );
nand U13913 ( n1160, n14002, n14003 );
nor U13914 ( n14003, n14004, n14005 );
nand U13915 ( n14005, n14006, n14007 );
nand U13916 ( n14007, n8184, n13971 );
nand U13917 ( n14006, n13972, n7856 );
nor U13918 ( n14004, n8185, n13973 );
nor U13919 ( n14002, n14008, n14009 );
nor U13920 ( n14009, n8188, n13976 );
nor U13921 ( n14008, n8189, n13977 );
nand U13922 ( n1155, n14010, n14011 );
nor U13923 ( n14011, n14012, n14013 );
nand U13924 ( n14013, n14014, n14015 );
nand U13925 ( n14015, n8089, n13971 );
nand U13926 ( n14014, n13972, n7857 );
nor U13927 ( n14012, n8196, n13973 );
nor U13928 ( n14010, n14016, n14017 );
nor U13929 ( n14017, n8093, n13976 );
nor U13930 ( n14016, n8098, n13977 );
nand U13931 ( n1150, n14018, n14019 );
nor U13932 ( n14019, n14020, n14021 );
nand U13933 ( n14021, n14022, n14023 );
nand U13934 ( n14023, n8106, n13971 );
nand U13935 ( n14022, n13972, n7858 );
nor U13936 ( n14020, n8205, n13973 );
nor U13937 ( n14018, n14024, n14025 );
nor U13938 ( n14025, n8108, n13976 );
nor U13939 ( n14024, n8111, n13977 );
nand U13940 ( n1145, n14026, n14027 );
nor U13941 ( n14027, n14028, n14029 );
nand U13942 ( n14029, n14030, n14031 );
nand U13943 ( n14031, n8118, n13971 );
nand U13944 ( n13971, n14032, n14033 );
nand U13945 ( n14033, n14034, n8218 );
nand U13946 ( n14032, n14035, n8482 );
nand U13947 ( n14030, n13972, n7919 );
nand U13948 ( n13972, n14036, n14037 );
nor U13949 ( n14037, n14038, n14039 );
and U13950 ( n14039, n7815, n13973 );
nor U13951 ( n14038, n14040, n14034 );
nand U13952 ( n14034, n13973, n14041 );
nand U13953 ( n14041, n14042, n8490 );
nor U13954 ( n14040, n14043, n8231 );
and U13955 ( n14043, n13976, n13977 );
nor U13956 ( n14036, n14044, n8235 );
nor U13957 ( n14044, n15061, n14035 );
nor U13958 ( n14028, n8119, n13973 );
nand U13959 ( n13973, n14045, n8494 );
nor U13960 ( n14026, n14046, n14047 );
nor U13961 ( n14047, n8124, n13976 );
nand U13962 ( n13976, n14048, n8498 );
nor U13963 ( n14046, n8121, n13977 );
nand U13964 ( n13977, n14049, n8500 );
nand U13965 ( n1140, n14050, n14051 );
nor U13966 ( n14051, n14052, n14053 );
nand U13967 ( n14053, n14054, n14055 );
nand U13968 ( n14055, n8131, n14056 );
nand U13969 ( n14054, n14057, n7995 );
nor U13970 ( n14052, n8135, n14058 );
nor U13971 ( n14050, n14059, n14060 );
nor U13972 ( n14060, n8139, n14061 );
nor U13973 ( n14059, n8141, n14062 );
nand U13974 ( n1135, n14063, n14064 );
nor U13975 ( n14064, n14065, n14066 );
nand U13976 ( n14066, n14067, n14068 );
nand U13977 ( n14068, n8148, n14056 );
nand U13978 ( n14067, n14057, n7996 );
nor U13979 ( n14065, n8149, n14058 );
nor U13980 ( n14063, n14069, n14070 );
nor U13981 ( n14070, n8152, n14061 );
nor U13982 ( n14069, n8153, n14062 );
nand U13983 ( n1130, n14071, n14072 );
nor U13984 ( n14072, n14073, n14074 );
nand U13985 ( n14074, n14075, n14076 );
nand U13986 ( n14076, n8160, n14056 );
nand U13987 ( n14075, n14057, n7997 );
nor U13988 ( n14073, n8161, n14058 );
nor U13989 ( n14071, n14077, n14078 );
nor U13990 ( n14078, n8164, n14061 );
nor U13991 ( n14077, n8165, n14062 );
nand U13992 ( n1125, n14079, n14080 );
nor U13993 ( n14080, n14081, n14082 );
nand U13994 ( n14082, n14083, n14084 );
nand U13995 ( n14084, n8172, n14056 );
nand U13996 ( n14083, n14057, n7998 );
nor U13997 ( n14081, n8173, n14058 );
nor U13998 ( n14079, n14085, n14086 );
nor U13999 ( n14086, n8176, n14061 );
nor U14000 ( n14085, n8177, n14062 );
nand U14001 ( n1120, n14087, n14088 );
nor U14002 ( n14088, n14089, n14090 );
nand U14003 ( n14090, n14091, n14092 );
nand U14004 ( n14092, n8184, n14056 );
nand U14005 ( n14091, n14057, n7999 );
nor U14006 ( n14089, n8185, n14058 );
nor U14007 ( n14087, n14093, n14094 );
nor U14008 ( n14094, n8188, n14061 );
nor U14009 ( n14093, n8189, n14062 );
nand U14010 ( n1115, n14095, n14096 );
nor U14011 ( n14096, n14097, n14098 );
nand U14012 ( n14098, n14099, n14100 );
nand U14013 ( n14100, n8089, n14056 );
nand U14014 ( n14099, n14057, n8000 );
nor U14015 ( n14097, n8196, n14058 );
nor U14016 ( n14095, n14101, n14102 );
nor U14017 ( n14102, n8093, n14061 );
nor U14018 ( n14101, n8098, n14062 );
nand U14019 ( n1110, n14103, n14104 );
nor U14020 ( n14104, n14105, n14106 );
nand U14021 ( n14106, n14107, n14108 );
nand U14022 ( n14108, n8106, n14056 );
nand U14023 ( n14107, n14057, n8001 );
nor U14024 ( n14105, n8205, n14058 );
nor U14025 ( n14103, n14109, n14110 );
nor U14026 ( n14110, n8108, n14061 );
nor U14027 ( n14109, n8111, n14062 );
nand U14028 ( n1105, n14111, n14112 );
nor U14029 ( n14112, n14113, n14114 );
nand U14030 ( n14114, n14115, n14116 );
nand U14031 ( n14116, n8118, n14056 );
nand U14032 ( n14056, n14117, n14118 );
nand U14033 ( n14118, n14119, n7797 );
nand U14034 ( n14117, n14120, n8218 );
nand U14035 ( n14115, n14057, n8068 );
nand U14036 ( n14057, n14121, n14122 );
nor U14037 ( n14122, n14123, n14124 );
nor U14038 ( n14124, n15061, n14119 );
nand U14039 ( n14119, n14058, n14125 );
nand U14040 ( n14125, n14035, n8224 );
nor U14041 ( n8224, n14126, n7803 );
nor U14042 ( n14123, n14127, n14120 );
nand U14043 ( n14120, n14058, n14128 );
nand U14044 ( n14128, n14042, n8228 );
nor U14045 ( n8228, n13780, n14129 );
nor U14046 ( n14127, n14130, n8231 );
nor U14047 ( n14130, n8232, n14131 );
nand U14048 ( n14131, n14062, n14061 );
nor U14049 ( n14121, n14132, n8235 );
and U14050 ( n14132, n7815, n14058 );
nor U14051 ( n14113, n8119, n14058 );
nand U14052 ( n14058, n14045, n8236 );
nor U14053 ( n14111, n14133, n14134 );
nor U14054 ( n14134, n8124, n14061 );
nand U14055 ( n14061, n14048, n8240 );
nor U14056 ( n14133, n8121, n14062 );
nand U14057 ( n14062, n14049, n8242 );
nor U14058 ( n8242, n14135, n13776 );
nand U14059 ( n1100, n14136, n14137 );
nor U14060 ( n14137, n14138, n14139 );
nand U14061 ( n14139, n14140, n14141 );
nand U14062 ( n14141, n8131, n14142 );
nand U14063 ( n14140, n14143, n8002 );
nor U14064 ( n14138, n8135, n14144 );
nor U14065 ( n14136, n14145, n14146 );
nor U14066 ( n14146, n8139, n14147 );
nor U14067 ( n14145, n8141, n14148 );
nand U14068 ( n1095, n14149, n14150 );
nor U14069 ( n14150, n14151, n14152 );
nand U14070 ( n14152, n14153, n14154 );
nand U14071 ( n14154, n8148, n14142 );
nand U14072 ( n14153, n14143, n8003 );
nor U14073 ( n14151, n8149, n14144 );
nor U14074 ( n14149, n14155, n14156 );
nor U14075 ( n14156, n8152, n14147 );
nor U14076 ( n14155, n8153, n14148 );
nand U14077 ( n1090, n14157, n14158 );
nor U14078 ( n14158, n14159, n14160 );
nand U14079 ( n14160, n14161, n14162 );
nand U14080 ( n14162, n8160, n14142 );
nand U14081 ( n14161, n14143, n8004 );
nor U14082 ( n14159, n8161, n14144 );
nor U14083 ( n14157, n14163, n14164 );
nor U14084 ( n14164, n8164, n14147 );
nor U14085 ( n14163, n8165, n14148 );
nand U14086 ( n1085, n14165, n14166 );
nor U14087 ( n14166, n14167, n14168 );
nand U14088 ( n14168, n14169, n14170 );
nand U14089 ( n14170, n8172, n14142 );
nand U14090 ( n14169, n14143, n8005 );
nor U14091 ( n14167, n8173, n14144 );
nor U14092 ( n14165, n14171, n14172 );
nor U14093 ( n14172, n8176, n14147 );
nor U14094 ( n14171, n8177, n14148 );
nand U14095 ( n1080, n14173, n14174 );
nor U14096 ( n14174, n14175, n14176 );
nand U14097 ( n14176, n14177, n14178 );
nand U14098 ( n14178, n8184, n14142 );
nand U14099 ( n14177, n14143, n8006 );
nor U14100 ( n14175, n8185, n14144 );
nor U14101 ( n14173, n14179, n14180 );
nor U14102 ( n14180, n8188, n14147 );
nor U14103 ( n14179, n8189, n14148 );
nand U14104 ( n1075, n14181, n14182 );
nor U14105 ( n14182, n14183, n14184 );
nand U14106 ( n14184, n14185, n14186 );
nand U14107 ( n14186, n8089, n14142 );
nand U14108 ( n14185, n14143, n8007 );
nor U14109 ( n14183, n8196, n14144 );
nor U14110 ( n14181, n14187, n14188 );
nor U14111 ( n14188, n8093, n14147 );
nor U14112 ( n14187, n8098, n14148 );
nand U14113 ( n1070, n14189, n14190 );
nor U14114 ( n14190, n14191, n14192 );
nand U14115 ( n14192, n14193, n14194 );
nand U14116 ( n14194, n8106, n14142 );
nand U14117 ( n14193, n14143, n8008 );
nor U14118 ( n14191, n8205, n14144 );
nor U14119 ( n14189, n14195, n14196 );
nor U14120 ( n14196, n8108, n14147 );
nor U14121 ( n14195, n8111, n14148 );
nand U14122 ( n1065, n14197, n14198 );
nor U14123 ( n14198, n14199, n14200 );
nand U14124 ( n14200, n14201, n14202 );
nand U14125 ( n14202, n8118, n14142 );
nand U14126 ( n14142, n14203, n14204 );
nand U14127 ( n14204, n14042, n8313 );
and U14128 ( n8313, n14129, n8218 );
nand U14129 ( n14203, n14035, n8314 );
nor U14130 ( n8314, n14205, n15061 );
nand U14131 ( n14201, n14143, n8069 );
nand U14132 ( n14143, n14206, n14035 );
nor U14133 ( n14206, n14207, n8317 );
nand U14134 ( n8317, n14208, n13834 );
not U14135 ( n13834, n8235 );
nor U14136 ( n14208, n8482, n14209 );
nor U14137 ( n14209, n14129, n14210 );
and U14138 ( n14207, n7815, n14144 );
nor U14139 ( n14199, n8119, n14144 );
nand U14140 ( n14144, n14045, n8320 );
nor U14141 ( n14197, n14211, n14212 );
nor U14142 ( n14212, n8124, n14147 );
nand U14143 ( n14147, n14048, n8323 );
nor U14144 ( n14211, n8121, n14148 );
nand U14145 ( n14148, n14049, n8324 );
nor U14146 ( n8324, n12162, n14213 );
nand U14147 ( n1060, n14214, n14215 );
nor U14148 ( n14215, n14216, n14217 );
nand U14149 ( n14217, n14218, n14219 );
nand U14150 ( n14219, n8131, n14220 );
nand U14151 ( n14218, n14221, n8009 );
nor U14152 ( n14216, n8135, n14222 );
nor U14153 ( n14214, n14223, n14224 );
nor U14154 ( n14224, n8139, n14225 );
nor U14155 ( n14223, n8141, n14226 );
nand U14156 ( n1055, n14227, n14228 );
nor U14157 ( n14228, n14229, n14230 );
nand U14158 ( n14230, n14231, n14232 );
nand U14159 ( n14232, n8148, n14220 );
nand U14160 ( n14231, n14221, n8010 );
nor U14161 ( n14229, n8149, n14222 );
nor U14162 ( n14227, n14233, n14234 );
nor U14163 ( n14234, n8152, n14225 );
nor U14164 ( n14233, n8153, n14226 );
nand U14165 ( n1050, n14235, n14236 );
nor U14166 ( n14236, n14237, n14238 );
nand U14167 ( n14238, n14239, n14240 );
nand U14168 ( n14240, n8160, n14220 );
nand U14169 ( n14239, n14221, n8011 );
nor U14170 ( n14237, n8161, n14222 );
nor U14171 ( n14235, n14241, n14242 );
nor U14172 ( n14242, n8164, n14225 );
nor U14173 ( n14241, n8165, n14226 );
nand U14174 ( n1045, n14243, n14244 );
nor U14175 ( n14244, n14245, n14246 );
nand U14176 ( n14246, n14247, n14248 );
nand U14177 ( n14248, n8172, n14220 );
nand U14178 ( n14247, n14221, n8012 );
nor U14179 ( n14245, n8173, n14222 );
nor U14180 ( n14243, n14249, n14250 );
nor U14181 ( n14250, n8176, n14225 );
nor U14182 ( n14249, n8177, n14226 );
nand U14183 ( n1040, n14251, n14252 );
nor U14184 ( n14252, n14253, n14254 );
nand U14185 ( n14254, n14255, n14256 );
nand U14186 ( n14256, n8184, n14220 );
nand U14187 ( n14255, n14221, n8013 );
nor U14188 ( n14253, n8185, n14222 );
nor U14189 ( n14251, n14257, n14258 );
nor U14190 ( n14258, n8188, n14225 );
nor U14191 ( n14257, n8189, n14226 );
nand U14192 ( n1035, n14259, n14260 );
nor U14193 ( n14260, n14261, n14262 );
nand U14194 ( n14262, n14263, n14264 );
nand U14195 ( n14264, n8089, n14220 );
not U14196 ( n10445, DATAI_5_ );
nand U14197 ( n14263, n14265, n8092 );
not U14198 ( n8092, n8196 );
nand U14199 ( n8196, n14266, n10483 );
nor U14200 ( n14261, n8093, n14225 );
nand U14201 ( n8093, DATAI_21_, n14267 );
nor U14202 ( n14259, n14268, n14269 );
nor U14203 ( n14269, n15162, n14270 );
nor U14204 ( n14268, n8098, n14226 );
nand U14205 ( n8098, DATAI_29_, n14267 );
nand U14206 ( n1030, n14271, n14272 );
nor U14207 ( n14272, n14273, n14274 );
nand U14208 ( n14274, n14275, n14276 );
nand U14209 ( n14276, n8106, n14220 );
not U14210 ( n10438, DATAI_6_ );
nand U14211 ( n14275, n14265, n8107 );
not U14212 ( n8107, n8205 );
nand U14213 ( n8205, n14266, n13744 );
nor U14214 ( n14273, n8108, n14225 );
nand U14215 ( n8108, DATAI_22_, n14267 );
nor U14216 ( n14271, n14277, n14278 );
nor U14217 ( n14278, n15161, n14270 );
nor U14218 ( n14277, n8111, n14226 );
nand U14219 ( n8111, DATAI_30_, n14267 );
nand U14220 ( n1025, n14279, n14280 );
nor U14221 ( n14280, n14281, n14282 );
nand U14222 ( n14282, n14283, n14284 );
nand U14223 ( n14284, n8118, n14220 );
nand U14224 ( n14220, n14285, n14286 );
nand U14225 ( n14286, n14287, n7797 );
nand U14226 ( n14285, n14288, n8218 );
not U14227 ( n10431, DATAI_7_ );
or U14228 ( n14283, n14270, n15160 );
not U14229 ( n14270, n14221 );
nand U14230 ( n14221, n14289, n14290 );
nor U14231 ( n14290, n14291, n14292 );
nor U14232 ( n14292, n15061, n14287 );
nand U14233 ( n14287, n14222, n14293 );
nand U14234 ( n14293, n14035, n8401 );
nor U14235 ( n8401, n7803, n14205 );
nor U14236 ( n14035, n14294, n8733 );
nor U14237 ( n14291, n14295, n14288 );
nand U14238 ( n14288, n14222, n14296 );
nand U14239 ( n14296, n14042, n8404 );
nor U14240 ( n8404, n8490, n13780 );
nor U14241 ( n14042, n8738, n10107 );
nor U14242 ( n14295, n14297, n8231 );
nor U14243 ( n14297, n8232, n14298 );
nand U14244 ( n14298, n14226, n14225 );
not U14245 ( n8232, n14267 );
nor U14246 ( n14289, n14299, n8235 );
nor U14247 ( n14299, n15060, n14265 );
not U14248 ( n14265, n14222 );
nor U14249 ( n14281, n8119, n14222 );
nand U14250 ( n14222, n14045, n8742 );
nor U14251 ( n14045, n7804, n7826 );
nand U14252 ( n8119, n14266, n9407 );
nor U14253 ( n14279, n14300, n14301 );
nor U14254 ( n14301, n8124, n14225 );
nand U14255 ( n14225, n14048, n8745 );
nor U14256 ( n14048, n13795, n12075 );
nand U14257 ( n8124, DATAI_23_, n14267 );
nor U14258 ( n14300, n8121, n14226 );
nand U14259 ( n14226, n14049, n8746 );
not U14260 ( n8746, n13799 );
nand U14261 ( n13799, n12162, n14135 );
nor U14262 ( n14049, n8747, n9079 );
nand U14263 ( n8121, DATAI_31_, n14267 );
nand U14264 ( n1020, n14302, n14303 );
nor U14265 ( n14303, n14304, n14305 );
nand U14266 ( n14305, n14306, n14307 );
nand U14267 ( n14307, n8131, n8090 );
not U14268 ( n10481, DATAI_0_ );
or U14269 ( n14306, n8135, n8120 );
nand U14270 ( n8135, n14266, n9424 );
nor U14271 ( n14304, n8094, n8139 );
nand U14272 ( n8139, DATAI_16_, n14267 );
nor U14273 ( n14302, n14308, n14309 );
nor U14274 ( n14309, n15159, n8097 );
nor U14275 ( n14308, n8099, n8141 );
nand U14276 ( n8141, DATAI_24_, n14267 );
nand U14277 ( n1015, n14310, n14311 );
nor U14278 ( n14311, n14312, n14313 );
nand U14279 ( n14313, n14314, n14315 );
nand U14280 ( n14315, n8148, n8090 );
not U14281 ( n10473, DATAI_1_ );
or U14282 ( n14314, n8149, n8120 );
nand U14283 ( n8149, n14266, n10825 );
nor U14284 ( n14312, n8094, n8152 );
nand U14285 ( n8152, DATAI_17_, n14267 );
nor U14286 ( n14310, n14316, n14317 );
nor U14287 ( n14317, n15158, n8097 );
nor U14288 ( n14316, n8099, n8153 );
nand U14289 ( n8153, DATAI_25_, n14267 );
nand U14290 ( n1010, n14318, n14319 );
nor U14291 ( n14319, n14320, n14321 );
nand U14292 ( n14321, n14322, n14323 );
nand U14293 ( n14323, n8160, n8090 );
not U14294 ( n10466, DATAI_2_ );
or U14295 ( n14322, n8161, n8120 );
nand U14296 ( n8161, n14266, n10570 );
nor U14297 ( n14320, n8094, n8164 );
nand U14298 ( n8164, DATAI_18_, n14267 );
nor U14299 ( n14318, n14324, n14325 );
nor U14300 ( n14325, n15157, n8097 );
nor U14301 ( n14324, n8099, n8165 );
nand U14302 ( n8165, DATAI_26_, n14267 );
nand U14303 ( n1005, n14326, n14327 );
nor U14304 ( n14327, n14328, n14329 );
nand U14305 ( n14329, n14330, n14331 );
nand U14306 ( n14331, n8172, n8090 );
not U14307 ( n10459, DATAI_3_ );
or U14308 ( n14330, n8173, n8120 );
nand U14309 ( n8173, n14266, n10569 );
nor U14310 ( n14328, n8094, n8176 );
nand U14311 ( n8176, DATAI_19_, n14267 );
nor U14312 ( n14326, n14332, n14333 );
nor U14313 ( n14333, n15156, n8097 );
nor U14314 ( n14332, n8099, n8177 );
nand U14315 ( n8177, DATAI_27_, n14267 );
nand U14316 ( n1000, n14334, n14335 );
nor U14317 ( n14335, n14336, n14337 );
nand U14318 ( n14337, n14338, n14339 );
nand U14319 ( n14339, n8184, n8090 );
nand U14320 ( n8090, n14340, n14341 );
nand U14321 ( n14341, n8218, n14342 );
nand U14322 ( n8218, n13789, n14210 );
nand U14323 ( n14340, n8482, n8225 );
nor U14324 ( n8482, n14126, n15061 );
not U14325 ( n10452, DATAI_4_ );
or U14326 ( n14338, n8097, n15155 );
and U14327 ( n8097, n14343, n14344 );
nor U14328 ( n14344, n14345, n14346 );
nor U14329 ( n14346, n15061, n8225 );
not U14330 ( n8225, n8319 );
nand U14331 ( n8319, n8734, n8733 );
nor U14332 ( n14345, n14347, n14342 );
nand U14333 ( n14342, n8120, n14348 );
nand U14334 ( n14348, n8229, n8490 );
not U14335 ( n8490, n14129 );
nor U14336 ( n8229, n9070, n10107 );
not U14337 ( n9070, n8738 );
nor U14338 ( n14347, n14349, n8231 );
not U14339 ( n8231, n14210 );
nand U14340 ( n14210, n15351, n9383 );
and U14341 ( n14349, n8094, n8099 );
nor U14342 ( n14343, n14350, n8235 );
nor U14343 ( n14350, n15060, n8091 );
not U14344 ( n8091, n8120 );
nor U14345 ( n14336, n8120, n8185 );
nand U14346 ( n8185, n14266, n10568 );
nor U14347 ( n14266, n8235, n15060 );
nand U14348 ( n8120, n8494, n8237 );
not U14349 ( n8494, n9165 );
nand U14350 ( n9165, n15200, n15201 );
nor U14351 ( n14334, n14351, n14352 );
nor U14352 ( n14352, n8094, n8188 );
nand U14353 ( n8188, DATAI_20_, n14267 );
nand U14354 ( n8094, n8241, n8498 );
nor U14355 ( n8498, n13776, n12119 );
nor U14356 ( n14351, n8099, n8189 );
nand U14357 ( n8189, DATAI_28_, n14267 );
nand U14358 ( n14353, n14354, n9119 );
nand U14359 ( n9119, n15061, n7799 );
nor U14360 ( n14354, n9096, n9120 );
nor U14361 ( n9096, n9428, n15060 );
not U14362 ( n9428, n9415 );
nand U14363 ( n9415, n14355, n14356 );
nand U14364 ( n14356, n14357, n13326 );
nor U14365 ( n14357, n13934, n14358 );
not U14366 ( n13934, n14359 );
nand U14367 ( n14355, n14360, n14361 );
nor U14368 ( n14361, n14362, n14363 );
nor U14369 ( n14363, n14364, n14365 );
nand U14370 ( n14365, n14359, n13271 );
nand U14371 ( n14359, n14366, n14367 );
nand U14372 ( n14367, n14368, n7831 );
or U14373 ( n14368, n15197, n14369 );
nand U14374 ( n14366, n15197, n14369 );
not U14375 ( n14364, n14358 );
nor U14376 ( n14362, n14370, n14358 );
nor U14377 ( n14370, n14371, n14372 );
and U14378 ( n14371, n13941, n13326 );
nor U14379 ( n14360, n14373, n14374 );
nor U14380 ( n14374, n13938, n14375 );
not U14381 ( n14375, n14372 );
nand U14382 ( n14372, n14376, n14377 );
nand U14383 ( n14377, n14378, n14379 );
nand U14384 ( n14379, n13941, n13271 );
xnor U14385 ( n13941, n14380, n14381 );
xor U14386 ( n14381, n15193, n15198 );
nor U14387 ( n14373, n14376, n14382 );
not U14388 ( n14382, n14378 );
nand U14389 ( n14378, n14383, n14384 );
nand U14390 ( n14384, n14385, n14386 );
nor U14391 ( n14385, n14387, n14388 );
not U14392 ( n14387, n14389 );
nand U14393 ( n14383, n14390, n14391 );
or U14394 ( n14391, n14392, n14393 );
nor U14395 ( n14390, n14394, n14395 );
nor U14396 ( n14395, n14396, n14389 );
nand U14397 ( n14389, n14397, n14398 );
or U14398 ( n14398, n10825, n14399 );
nand U14399 ( n14397, n13326, n13939 );
nor U14400 ( n14396, n13939, n14400 );
nand U14401 ( n14400, n14401, n7814 );
nand U14402 ( n14401, n9424, n10568 );
not U14403 ( n13939, n14386 );
xor U14404 ( n14386, n14402, n14403 );
xor U14405 ( n14403, n15194, n15199 );
nor U14406 ( n14394, n13942, n14404 );
nand U14407 ( n14404, n14405, n14358 );
nand U14408 ( n14358, n14406, n14407 );
nand U14409 ( n14407, n14408, n7814 );
nand U14410 ( n14408, n14409, n14410 );
nor U14411 ( n14409, n9393, n9427 );
nor U14412 ( n14406, n14411, n10562 );
nand U14413 ( n14405, n14392, n14393 );
nand U14414 ( n14393, n14412, n14413 );
nand U14415 ( n14413, n14414, n12742 );
not U14416 ( n12742, n12700 );
nand U14417 ( n12700, n10825, n10483 );
nor U14418 ( n14414, n14415, n13271 );
nand U14419 ( n14412, n14416, n14415 );
and U14420 ( n14415, n14417, n14418 );
nand U14421 ( n14418, n15196, n7803 );
nor U14422 ( n14416, n14419, n14388 );
and U14423 ( n14388, n13327, n14420 );
nand U14424 ( n14420, n9422, n7814 );
nor U14425 ( n14419, n14421, n14422 );
nor U14426 ( n14422, n14399, n10825 );
nor U14427 ( n14399, n10483, n10562 );
nor U14428 ( n14421, n9139, n14410 );
nand U14429 ( n14392, n14423, n14424 );
nor U14430 ( n14424, n14411, n9427 );
not U14431 ( n14411, n9397 );
nor U14432 ( n14423, n14425, n14426 );
nor U14433 ( n14426, n10822, n10568 );
nor U14434 ( n14425, n13942, n13271 );
xor U14435 ( n13942, n14417, n14427 );
xor U14436 ( n14427, n15195, n15200 );
and U14437 ( n14376, n14428, n14429 );
nand U14438 ( n14429, n13938, n13326 );
and U14439 ( n13938, n14430, n15192 );
nor U14440 ( n14430, n15197, n14369 );
and U14441 ( n14369, n14431, n14432 );
nand U14442 ( n14432, n15193, n14433 );
or U14443 ( n14433, n7804, n14380 );
nand U14444 ( n14431, n14380, n7804 );
nand U14445 ( n14380, n14434, n14435 );
nand U14446 ( n14435, n15194, n14436 );
or U14447 ( n14436, n7826, n14402 );
nand U14448 ( n14434, n14402, n7826 );
nand U14449 ( n14402, n14437, n14438 );
nand U14450 ( n14438, n15195, n14439 );
nand U14451 ( n14439, n15200, n14440 );
not U14452 ( n14440, n14417 );
nand U14453 ( n14437, n14417, n7825 );
nand U14454 ( n14417, n15201, n7798 );
nand U14455 ( n14428, n15063, n7831 );
nand U14456 ( n13789, n9383, n7830 );
nor U14457 ( n9383, n7815, n7797 );
nand U14458 ( n8099, n8500, n8243 );
nor U14459 ( n8243, n9079, n8990 );
not U14460 ( n8990, n8747 );
xnor U14461 ( n8747, n14441, n13795 );
nand U14462 ( n9079, n14442, n14443 );
nand U14463 ( n14443, n12075, n14441 );
nor U14464 ( n14442, n8497, n14444 );
not U14465 ( n14444, n8336 );
nand U14466 ( n8336, n8745, n8241 );
nor U14467 ( n8241, n9077, n12075 );
not U14468 ( n8745, n14441 );
nand U14469 ( n14441, n12119, n13776 );
nor U14470 ( n8497, n9076, n13795 );
not U14471 ( n13795, n9077 );
xor U14472 ( n9077, n14445, n14446 );
nand U14473 ( n14445, n14447, n14448 );
nand U14474 ( n14448, n14449, n14450 );
not U14475 ( n9076, n12075 );
xor U14476 ( n12075, n14451, n13571 );
and U14477 ( n13571, n14452, n14453 );
xor U14478 ( n14453, n12765, n14454 );
nand U14479 ( n14454, n14455, n14456 );
nand U14480 ( n14456, n10107, n15063 );
xor U14481 ( n10107, n13963, n13964 );
nand U14482 ( n13964, n14457, n14458 );
nand U14483 ( n14458, n9350, n7804 );
nor U14484 ( n14457, n14459, n14460 );
nor U14485 ( n14460, n15193, n14461 );
nor U14486 ( n14459, n8734, n12148 );
not U14487 ( n8734, n14294 );
nand U14488 ( n14294, n14462, n14463 );
nand U14489 ( n14463, n9164, n7804 );
nor U14490 ( n14462, n8493, n8408 );
not U14491 ( n8408, n8337 );
nand U14492 ( n8337, n8742, n8237 );
nor U14493 ( n8237, n7804, n15199 );
not U14494 ( n8742, n9164 );
nor U14495 ( n8493, n7826, n15198 );
and U14496 ( n13963, n14464, n14465 );
nor U14497 ( n14455, n14466, n14467 );
nor U14498 ( n14467, n12765, n13613 );
nor U14499 ( n14466, n14468, n14469 );
nor U14500 ( n14452, n14470, n14471 );
nor U14501 ( n14471, n15188, n13271 );
nor U14502 ( n14470, n14468, n13327 );
not U14503 ( n14468, n13613 );
nand U14504 ( n13613, n14472, n14473 );
nor U14505 ( n14473, n14474, n14475 );
nand U14506 ( n14475, n14476, n14477 );
nor U14507 ( n14477, n14478, n14479 );
nor U14508 ( n14479, n15084, n13410 );
nor U14509 ( n14478, n15092, n13411 );
nor U14510 ( n14476, n14480, n14481 );
nor U14511 ( n14481, n15076, n13414 );
nor U14512 ( n14480, n15068, n13415 );
nand U14513 ( n14474, n14482, n14483 );
nor U14514 ( n14483, n14484, n14485 );
nor U14515 ( n14485, n15116, n13400 );
nor U14516 ( n14484, n15124, n13401 );
nor U14517 ( n14482, n14486, n14487 );
nor U14518 ( n14487, n15108, n13404 );
nor U14519 ( n14486, n15100, n13405 );
nor U14520 ( n14472, n14488, n14489 );
nand U14521 ( n14489, n14490, n14491 );
nor U14522 ( n14491, n14492, n14493 );
nor U14523 ( n14493, n15180, n13388 );
nor U14524 ( n14492, n15188, n13389 );
nor U14525 ( n14490, n14494, n14495 );
nor U14526 ( n14495, n15172, n13392 );
nor U14527 ( n14494, n15164, n13393 );
nand U14528 ( n14488, n14496, n14497 );
nor U14529 ( n14497, n14498, n14499 );
nor U14530 ( n14499, n15148, n13378 );
nor U14531 ( n14498, n15156, n13379 );
nor U14532 ( n14496, n14500, n14501 );
nor U14533 ( n14501, n15140, n13382 );
nor U14534 ( n14500, n15132, n13383 );
nand U14535 ( n14451, n14446, n14447 );
not U14536 ( n14447, n13570 );
nor U14537 ( n13570, n14450, n14449 );
xnor U14538 ( n14449, n14502, n12765 );
nand U14539 ( n14502, n14503, n14504 );
nand U14540 ( n14504, n8738, n15063 );
xor U14541 ( n8738, n14464, n14465 );
nand U14542 ( n14465, n14505, n14506 );
nand U14543 ( n14506, n14507, n14508 );
or U14544 ( n14507, n14509, n14510 );
and U14545 ( n14464, n14511, n14512 );
nand U14546 ( n14512, n14513, n15194 );
nand U14547 ( n14511, n14461, n14513 );
and U14548 ( n14513, n14514, n14515 );
nand U14549 ( n14515, n8733, n9384 );
not U14550 ( n8733, n9067 );
xnor U14551 ( n9067, n9164, n15199 );
nand U14552 ( n9164, n7803, n7825 );
nand U14553 ( n14514, n9350, n7826 );
nor U14554 ( n14503, n14516, n14517 );
nor U14555 ( n14517, n12765, n14518 );
nor U14556 ( n14516, n13653, n14469 );
not U14557 ( n13653, n14518 );
nand U14558 ( n14450, n14519, n14520 );
nand U14559 ( n14520, n9347, n14518 );
nand U14560 ( n14518, n14521, n14522 );
nor U14561 ( n14522, n14523, n14524 );
nand U14562 ( n14524, n14525, n14526 );
nor U14563 ( n14526, n14527, n14528 );
nor U14564 ( n14528, n15149, n13378 );
nor U14565 ( n14527, n15157, n13379 );
nor U14566 ( n14525, n14529, n14530 );
nor U14567 ( n14530, n15141, n13382 );
nor U14568 ( n14529, n15133, n13383 );
nand U14569 ( n14523, n14531, n14532 );
nor U14570 ( n14532, n14533, n14534 );
nor U14571 ( n14534, n15181, n13388 );
nor U14572 ( n14533, n15189, n13389 );
nor U14573 ( n14531, n14535, n14536 );
nor U14574 ( n14536, n15173, n13392 );
nor U14575 ( n14535, n15165, n13393 );
nor U14576 ( n14521, n14537, n14538 );
nand U14577 ( n14538, n14539, n14540 );
nor U14578 ( n14540, n14541, n14542 );
nor U14579 ( n14542, n15117, n13400 );
nor U14580 ( n14541, n15125, n13401 );
nor U14581 ( n14539, n14543, n14544 );
nor U14582 ( n14544, n15109, n13404 );
nor U14583 ( n14543, n15101, n13405 );
nand U14584 ( n14537, n14545, n14546 );
nor U14585 ( n14546, n14547, n14548 );
nor U14586 ( n14548, n15085, n13410 );
nor U14587 ( n14547, n15093, n13411 );
nor U14588 ( n14545, n14549, n14550 );
nor U14589 ( n14550, n15077, n13414 );
nor U14590 ( n14549, n15069, n13415 );
nand U14591 ( n14519, n13326, n7859 );
not U14592 ( n13326, n13271 );
and U14593 ( n14446, n13569, n14551 );
nand U14594 ( n14551, n14552, n14553 );
nor U14595 ( n8500, n14135, n12162 );
not U14596 ( n14135, n14213 );
nor U14597 ( n14213, n8323, n8240 );
nor U14598 ( n8240, n12162, n12119 );
nor U14599 ( n8323, n13682, n13776 );
not U14600 ( n13776, n12162 );
xor U14601 ( n12162, n14554, n12698 );
nand U14602 ( n14554, n14555, n14556 );
nand U14603 ( n14556, n14557, n14558 );
not U14604 ( n13682, n12119 );
xnor U14605 ( n12119, n14559, n13569 );
xnor U14606 ( n13569, n14560, n12765 );
nand U14607 ( n14560, n14561, n14562 );
nand U14608 ( n14562, n14129, n15063 );
xnor U14609 ( n14129, n14563, n14508 );
nand U14610 ( n14508, n14564, n14565 );
nand U14611 ( n14565, n14566, n13908 );
not U14612 ( n13908, n13724 );
nand U14613 ( n13724, n14567, n13892 );
nor U14614 ( n14567, n10825, n10483 );
nor U14615 ( n14566, n15063, n10480 );
nand U14616 ( n14563, n14505, n14568 );
nand U14617 ( n14568, n14569, n14570 );
nand U14618 ( n14569, n14509, n14571 );
nand U14619 ( n14505, n14572, n14510 );
and U14620 ( n14572, n14509, n14571 );
nand U14621 ( n14571, n14573, n14461 );
not U14622 ( n14461, n14574 );
nand U14623 ( n14509, n14573, n15195 );
and U14624 ( n14573, n14575, n14576 );
nand U14625 ( n14576, n9350, n7825 );
nand U14626 ( n14575, n9384, n14126 );
not U14627 ( n14126, n14205 );
nor U14628 ( n14205, n8320, n8236 );
nor U14629 ( n8236, n7825, n15201 );
nor U14630 ( n8320, n7803, n15200 );
not U14631 ( n9384, n12148 );
nor U14632 ( n14561, n14577, n14578 );
nor U14633 ( n14578, n12765, n13656 );
nor U14634 ( n14577, n13688, n14469 );
not U14635 ( n13688, n13656 );
xnor U14636 ( n14559, n14553, n14552 );
and U14637 ( n14552, n14579, n14580 );
nand U14638 ( n14580, n9347, n13656 );
nand U14639 ( n13656, n14581, n14582 );
nor U14640 ( n14582, n14583, n14584 );
nand U14641 ( n14584, n14585, n14586 );
nor U14642 ( n14586, n14587, n14588 );
nor U14643 ( n14588, n15150, n13378 );
nor U14644 ( n14587, n15158, n13379 );
nor U14645 ( n14585, n14589, n14590 );
nor U14646 ( n14590, n15142, n13382 );
nor U14647 ( n14589, n15134, n13383 );
nand U14648 ( n14583, n14591, n14592 );
nor U14649 ( n14592, n14593, n14594 );
nor U14650 ( n14594, n15182, n13388 );
nor U14651 ( n14593, n15190, n13389 );
nor U14652 ( n14591, n14595, n14596 );
nor U14653 ( n14596, n15174, n13392 );
nor U14654 ( n14595, n15166, n13393 );
nor U14655 ( n14581, n14597, n14598 );
nand U14656 ( n14598, n14599, n14600 );
nor U14657 ( n14600, n14601, n14602 );
nor U14658 ( n14602, n15118, n13400 );
nor U14659 ( n14601, n15126, n13401 );
nor U14660 ( n14599, n14603, n14604 );
nor U14661 ( n14604, n15110, n13404 );
nor U14662 ( n14603, n15102, n13405 );
nand U14663 ( n14597, n14605, n14606 );
nor U14664 ( n14606, n14607, n14608 );
nor U14665 ( n14608, n15086, n13410 );
nor U14666 ( n14607, n15094, n13411 );
nor U14667 ( n14605, n14609, n14610 );
nor U14668 ( n14610, n15078, n13414 );
nor U14669 ( n14609, n15070, n13415 );
nor U14670 ( n14579, n13537, n14611 );
nor U14671 ( n14611, n15190, n13271 );
and U14672 ( n14553, n12765, n14555 );
or U14673 ( n14555, n14558, n14557 );
and U14674 ( n14557, n14612, n14613 );
nor U14675 ( n14613, n15063, n14614 );
nor U14676 ( n14614, n13689, n13327 );
nor U14677 ( n14612, n14615, n14616 );
nor U14678 ( n14616, n13226, n10568 );
nor U14679 ( n14615, n15191, n13271 );
xnor U14680 ( n14558, n12765, n14617 );
nor U14681 ( n14617, n14618, n14619 );
nand U14682 ( n14619, n14620, n14621 );
nand U14683 ( n14621, n13537, n13655 );
not U14684 ( n13537, n14469 );
nand U14685 ( n14469, n14622, n13226 );
nor U14686 ( n14622, n15063, n10568 );
nand U14687 ( n14620, n13689, n12698 );
not U14688 ( n12698, n12765 );
not U14689 ( n13689, n13655 );
nand U14690 ( n13655, n14623, n14624 );
nor U14691 ( n14624, n14625, n14626 );
nand U14692 ( n14626, n14627, n14628 );
nor U14693 ( n14628, n14629, n14630 );
nor U14694 ( n14630, n15151, n13378 );
nor U14695 ( n14629, n15159, n13379 );
nor U14696 ( n14627, n14631, n14632 );
nor U14697 ( n14632, n15143, n13382 );
nor U14698 ( n14631, n15135, n13383 );
nand U14699 ( n14625, n14633, n14634 );
nor U14700 ( n14634, n14635, n14636 );
nor U14701 ( n14636, n15183, n13388 );
nor U14702 ( n14635, n15191, n13389 );
nor U14703 ( n14633, n14637, n14638 );
nor U14704 ( n14638, n15175, n13392 );
nor U14705 ( n14637, n15167, n13393 );
nor U14706 ( n14623, n14639, n14640 );
nand U14707 ( n14640, n14641, n14642 );
nor U14708 ( n14642, n14643, n14644 );
nor U14709 ( n14644, n15119, n13400 );
nor U14710 ( n14643, n15127, n13401 );
nor U14711 ( n14641, n14645, n14646 );
nor U14712 ( n14646, n15111, n13404 );
nor U14713 ( n14645, n15103, n13405 );
nand U14714 ( n14639, n14647, n14648 );
nor U14715 ( n14648, n14649, n14650 );
nor U14716 ( n14650, n15087, n13410 );
nor U14717 ( n14649, n15095, n13411 );
nor U14718 ( n14647, n14651, n14652 );
nor U14719 ( n14652, n15079, n13414 );
nor U14720 ( n14651, n15071, n13415 );
nor U14721 ( n14618, n7814, n13780 );
nand U14722 ( n13780, n14570, n14653 );
nand U14723 ( n14653, n14654, n14655 );
not U14724 ( n14570, n14510 );
nor U14725 ( n14510, n14654, n14655 );
and U14726 ( n14655, n14656, n14657 );
nand U14727 ( n14657, n14574, n7798 );
nand U14728 ( n14574, n14658, n14659 );
nor U14729 ( n14659, n14660, n14661 );
nand U14730 ( n14661, n14662, n9397 );
nand U14731 ( n9397, n9347, n10825 );
not U14732 ( n9347, n13327 );
nand U14733 ( n14662, n10562, n14663 );
nor U14734 ( n10562, n10825, n13327 );
nand U14735 ( n13327, n9139, n7814 );
nor U14736 ( n14660, n15063, n14664 );
nor U14737 ( n14664, n14665, n14666 );
nand U14738 ( n14666, n14667, n14668 );
nand U14739 ( n14668, n12254, n14669 );
nand U14740 ( n9363, n10825, n10569 );
nor U14741 ( n14658, n14670, n14671 );
not U14742 ( n14671, n14564 );
nor U14743 ( n14564, n14672, n10195 );
nor U14744 ( n10195, n13907, n15063 );
nand U14745 ( n13907, n9348, n9364 );
not U14746 ( n9364, n9435 );
nand U14747 ( n9435, n10822, n9139 );
nor U14748 ( n9348, n13960, n13734 );
nand U14749 ( n13960, n13713, n14669 );
not U14750 ( n14669, n9140 );
nand U14751 ( n9140, n13723, n12153 );
not U14752 ( n12153, n14410 );
not U14753 ( n13723, n10480 );
nand U14754 ( n10480, n9407, n13744 );
and U14755 ( n14672, n14673, n9440 );
not U14756 ( n9440, n10198 );
nand U14757 ( n10198, n14674, n14675 );
nor U14758 ( n14675, n10483, n14676 );
nand U14759 ( n14676, n9422, n9407 );
nor U14760 ( n14674, n12155, n13744 );
nand U14761 ( n12155, n13734, n10569 );
nor U14762 ( n14673, n15063, n14677 );
nor U14763 ( n14677, n10160, n14678 );
nor U14764 ( n14678, n13946, n13227 );
nand U14765 ( n13946, n9179, n14679 );
nand U14766 ( n14679, n7802, n7819 );
nand U14767 ( n9179, n15025, n15026 );
not U14768 ( n10160, n10177 );
nand U14769 ( n10177, n9424, n10825 );
nor U14770 ( n14670, n10553, n13271 );
nand U14771 ( n13271, n14680, n9424 );
nor U14772 ( n14680, n15063, n9422 );
nor U14773 ( n14656, n14681, n14682 );
nor U14774 ( n14682, n15201, n9120 );
not U14775 ( n9120, n9350 );
nand U14776 ( n9350, n15062, n7797 );
nor U14777 ( n14681, n7803, n12148 );
nand U14778 ( n12148, n9105, n15063 );
and U14779 ( n14654, n14683, n14684 );
nor U14780 ( n14684, n14685, n14686 );
nand U14781 ( n14686, n13916, n14687 );
nand U14782 ( n14687, n14688, n10825 );
nand U14783 ( n14688, n14667, n14689 );
nand U14784 ( n14689, n10555, n10568 );
not U14785 ( n14667, n13958 );
nand U14786 ( n13958, n13917, n10569 );
and U14787 ( n13917, n13953, n14690 );
nand U14788 ( n14690, n10553, n9422 );
nand U14789 ( n13916, n9139, n14691 );
nand U14790 ( n14691, n14692, n14693 );
nand U14791 ( n14693, n14410, n10825 );
not U14792 ( n14692, n14663 );
nand U14793 ( n14663, n14694, n14695 );
nor U14794 ( n14695, n10361, n14696 );
nor U14795 ( n14696, n13713, n13891 );
and U14796 ( n13891, n14697, n10553 );
not U14797 ( n10553, n10555 );
nor U14798 ( n14697, n9422, n10361 );
not U14799 ( n13713, n10569 );
nor U14800 ( n14694, n14698, n14699 );
nand U14801 ( n14699, n14700, n14701 );
nand U14802 ( n14701, n14702, n13734 );
nor U14803 ( n14702, n9426, n9427 );
not U14804 ( n9427, n10483 );
nand U14805 ( n14700, n14410, n10570 );
nand U14806 ( n14410, n9422, n10483 );
nor U14807 ( n14698, n10568, n13744 );
not U14808 ( n9139, n9424 );
nand U14809 ( n14685, n14703, n7814 );
nand U14810 ( n14703, n9393, n14704 );
nand U14811 ( n14704, n10569, n10555 );
nand U14812 ( n10555, n9426, n10483 );
nor U14813 ( n14683, n14665, n14705 );
nand U14814 ( n14705, n9105, n14706 );
nand U14815 ( n14706, n13892, n9426 );
and U14816 ( n13892, n14707, n13734 );
not U14817 ( n13734, n10570 );
nor U14818 ( n14707, n9424, n10569 );
nand U14819 ( n10569, n14708, n14709 );
nor U14820 ( n14709, n14710, n14711 );
nand U14821 ( n14711, n14712, n14713 );
nor U14822 ( n14713, n14714, n14715 );
nor U14823 ( n14715, n15108, n14716 );
nor U14824 ( n14714, n15100, n14717 );
nor U14825 ( n14712, n14718, n14719 );
nor U14826 ( n14719, n15116, n14720 );
nor U14827 ( n14718, n15124, n14721 );
nand U14828 ( n14710, n14722, n14723 );
nor U14829 ( n14723, n14724, n14725 );
nor U14830 ( n14725, n15076, n14726 );
nor U14831 ( n14724, n15068, n14727 );
nor U14832 ( n14722, n14728, n14729 );
nor U14833 ( n14729, n15084, n14730 );
nor U14834 ( n14728, n15092, n14731 );
nor U14835 ( n14708, n14732, n14733 );
nand U14836 ( n14733, n14734, n14735 );
nor U14837 ( n14735, n14736, n14737 );
nor U14838 ( n14737, n15164, n14738 );
nor U14839 ( n14736, n15148, n14739 );
nor U14840 ( n14734, n14740, n14741 );
nor U14841 ( n14741, n15132, n14742 );
nor U14842 ( n14740, n15156, n14743 );
nand U14843 ( n14732, n14744, n14745 );
nor U14844 ( n14745, n14746, n14747 );
nor U14845 ( n14747, n15180, n14748 );
nor U14846 ( n14746, n15172, n14749 );
nor U14847 ( n14744, n14750, n14751 );
nor U14848 ( n14751, n15140, n14752 );
nor U14849 ( n14750, n15188, n14753 );
nor U14850 ( n9105, n7815, n7799 );
nand U14851 ( n14665, n14754, n14755 );
nand U14852 ( n14755, n9393, n14756 );
nand U14853 ( n14756, n13953, n9422 );
nor U14854 ( n13953, n10361, n10367 );
nor U14855 ( n10367, n10483, n9426 );
not U14856 ( n9426, n13744 );
nand U14857 ( n13744, n14757, n14758 );
nor U14858 ( n14758, n14759, n14760 );
nand U14859 ( n14760, n14761, n14762 );
nor U14860 ( n14762, n14763, n14764 );
nor U14861 ( n14764, n15105, n14716 );
nor U14862 ( n14763, n15097, n14717 );
nor U14863 ( n14761, n14765, n14766 );
nor U14864 ( n14766, n15113, n14720 );
nor U14865 ( n14765, n15121, n14721 );
nand U14866 ( n14759, n14767, n14768 );
nor U14867 ( n14768, n14769, n14770 );
nor U14868 ( n14770, n15073, n14726 );
nor U14869 ( n14769, n15065, n14727 );
nor U14870 ( n14767, n14771, n14772 );
nor U14871 ( n14772, n15081, n14730 );
nor U14872 ( n14771, n15089, n14731 );
nor U14873 ( n14757, n14773, n14774 );
nand U14874 ( n14774, n14775, n14776 );
nor U14875 ( n14776, n14777, n14778 );
nor U14876 ( n14778, n15161, n14738 );
nor U14877 ( n14777, n15145, n14739 );
nor U14878 ( n14775, n14779, n14780 );
nor U14879 ( n14780, n15129, n14742 );
nor U14880 ( n14779, n15153, n14743 );
nand U14881 ( n14773, n14781, n14782 );
nor U14882 ( n14782, n14783, n14784 );
nor U14883 ( n14784, n15177, n14748 );
nor U14884 ( n14783, n15169, n14749 );
nor U14885 ( n14781, n14785, n14786 );
nor U14886 ( n14786, n15137, n14752 );
nor U14887 ( n14785, n15185, n14753 );
nand U14888 ( n10483, n14787, n14788 );
nor U14889 ( n14788, n14789, n14790 );
nand U14890 ( n14790, n14791, n14792 );
nor U14891 ( n14792, n14793, n14794 );
nor U14892 ( n14794, n15106, n14716 );
nor U14893 ( n14793, n15098, n14717 );
nor U14894 ( n14791, n14795, n14796 );
nor U14895 ( n14796, n15114, n14720 );
nor U14896 ( n14795, n15122, n14721 );
nand U14897 ( n14789, n14797, n14798 );
nor U14898 ( n14798, n14799, n14800 );
nor U14899 ( n14800, n15074, n14726 );
nor U14900 ( n14799, n15066, n14727 );
nor U14901 ( n14797, n14801, n14802 );
nor U14902 ( n14802, n15082, n14730 );
nor U14903 ( n14801, n15090, n14731 );
nor U14904 ( n14787, n14803, n14804 );
nand U14905 ( n14804, n14805, n14806 );
nor U14906 ( n14806, n14807, n14808 );
nor U14907 ( n14808, n15162, n14738 );
nor U14908 ( n14807, n15146, n14739 );
nor U14909 ( n14805, n14809, n14810 );
nor U14910 ( n14810, n15130, n14742 );
nor U14911 ( n14809, n15154, n14743 );
nand U14912 ( n14803, n14811, n14812 );
nor U14913 ( n14812, n14813, n14814 );
nor U14914 ( n14814, n15178, n14748 );
nor U14915 ( n14813, n15170, n14749 );
nor U14916 ( n14811, n14815, n14816 );
nor U14917 ( n14816, n15138, n14752 );
nor U14918 ( n14815, n15186, n14753 );
not U14919 ( n10361, n9407 );
nand U14920 ( n9407, n14817, n14818 );
nor U14921 ( n14818, n14819, n14820 );
nand U14922 ( n14820, n14821, n14822 );
nor U14923 ( n14822, n14823, n14824 );
nor U14924 ( n14824, n15104, n14716 );
nor U14925 ( n14823, n15096, n14717 );
nor U14926 ( n14821, n14825, n14826 );
nor U14927 ( n14826, n15112, n14720 );
nor U14928 ( n14825, n15120, n14721 );
nand U14929 ( n14819, n14827, n14828 );
nor U14930 ( n14828, n14829, n14830 );
nor U14931 ( n14830, n15072, n14726 );
nor U14932 ( n14829, n15064, n14727 );
nor U14933 ( n14827, n14831, n14832 );
nor U14934 ( n14832, n15080, n14730 );
nor U14935 ( n14831, n15088, n14731 );
nor U14936 ( n14817, n14833, n14834 );
nand U14937 ( n14834, n14835, n14836 );
nor U14938 ( n14836, n14837, n14838 );
nor U14939 ( n14838, n15160, n14738 );
nor U14940 ( n14837, n15144, n14739 );
nor U14941 ( n14835, n14839, n14840 );
nor U14942 ( n14840, n15128, n14742 );
nor U14943 ( n14839, n15152, n14743 );
nand U14944 ( n14833, n14841, n14842 );
nor U14945 ( n14842, n14843, n14844 );
nor U14946 ( n14844, n15176, n14748 );
nor U14947 ( n14843, n15168, n14749 );
nor U14948 ( n14841, n14845, n14846 );
nor U14949 ( n14846, n15136, n14752 );
nor U14950 ( n14845, n15184, n14753 );
not U14951 ( n9393, n13227 );
nand U14952 ( n13227, n10822, n9424 );
nand U14953 ( n10825, n14847, n14848 );
nor U14954 ( n14848, n14849, n14850 );
nand U14955 ( n14850, n14851, n14852 );
nor U14956 ( n14852, n14853, n14854 );
nor U14957 ( n14854, n15110, n14716 );
nor U14958 ( n14853, n15102, n14717 );
nor U14959 ( n14851, n14855, n14856 );
nor U14960 ( n14856, n15118, n14720 );
nor U14961 ( n14855, n15126, n14721 );
nand U14962 ( n14849, n14857, n14858 );
nor U14963 ( n14858, n14859, n14860 );
nor U14964 ( n14860, n15078, n14726 );
nor U14965 ( n14859, n15070, n14727 );
nor U14966 ( n14857, n14861, n14862 );
nor U14967 ( n14862, n15086, n14730 );
nor U14968 ( n14861, n15094, n14731 );
nor U14969 ( n14847, n14863, n14864 );
nand U14970 ( n14864, n14865, n14866 );
nor U14971 ( n14866, n14867, n14868 );
nor U14972 ( n14868, n15166, n14738 );
nor U14973 ( n14867, n15150, n14739 );
nor U14974 ( n14865, n14869, n14870 );
nor U14975 ( n14870, n15134, n14742 );
nor U14976 ( n14869, n15158, n14743 );
nand U14977 ( n14863, n14871, n14872 );
nor U14978 ( n14872, n14873, n14874 );
nor U14979 ( n14874, n15182, n14748 );
nor U14980 ( n14873, n15174, n14749 );
nor U14981 ( n14871, n14875, n14876 );
nor U14982 ( n14876, n15142, n14752 );
nor U14983 ( n14875, n15190, n14753 );
nand U14984 ( n14754, n10570, n9424 );
nand U14985 ( n9424, n14877, n14878 );
nor U14986 ( n14878, n14879, n14880 );
nand U14987 ( n14880, n14881, n14882 );
nor U14988 ( n14882, n14883, n14884 );
nor U14989 ( n14884, n15111, n14716 );
nor U14990 ( n14883, n15103, n14717 );
nor U14991 ( n14881, n14885, n14886 );
nor U14992 ( n14886, n15119, n14720 );
nor U14993 ( n14885, n15127, n14721 );
nand U14994 ( n14879, n14887, n14888 );
nor U14995 ( n14888, n14889, n14890 );
nor U14996 ( n14890, n15079, n14726 );
nor U14997 ( n14889, n15071, n14727 );
nor U14998 ( n14887, n14891, n14892 );
nor U14999 ( n14892, n15087, n14730 );
nor U15000 ( n14891, n15095, n14731 );
nor U15001 ( n14877, n14893, n14894 );
nand U15002 ( n14894, n14895, n14896 );
nor U15003 ( n14896, n14897, n14898 );
nor U15004 ( n14898, n15167, n14738 );
nor U15005 ( n14897, n15151, n14739 );
nor U15006 ( n14895, n14899, n14900 );
nor U15007 ( n14900, n15135, n14742 );
nor U15008 ( n14899, n15159, n14743 );
nand U15009 ( n14893, n14901, n14902 );
nor U15010 ( n14902, n14903, n14904 );
nor U15011 ( n14904, n15183, n14748 );
nor U15012 ( n14903, n15175, n14749 );
nor U15013 ( n14901, n14905, n14906 );
nor U15014 ( n14906, n15143, n14752 );
nor U15015 ( n14905, n15191, n14753 );
nand U15016 ( n10570, n14907, n14908 );
nor U15017 ( n14908, n14909, n14910 );
nand U15018 ( n14910, n14911, n14912 );
nor U15019 ( n14912, n14913, n14914 );
nor U15020 ( n14914, n15109, n14716 );
nor U15021 ( n14913, n15101, n14717 );
nor U15022 ( n14911, n14915, n14916 );
nor U15023 ( n14916, n15117, n14720 );
nor U15024 ( n14915, n15125, n14721 );
nand U15025 ( n14909, n14917, n14918 );
nor U15026 ( n14918, n14919, n14920 );
nor U15027 ( n14920, n15077, n14726 );
nor U15028 ( n14919, n15069, n14727 );
nor U15029 ( n14917, n14921, n14922 );
nor U15030 ( n14922, n15085, n14730 );
nor U15031 ( n14921, n15093, n14731 );
nor U15032 ( n14907, n14923, n14924 );
nand U15033 ( n14924, n14925, n14926 );
nor U15034 ( n14926, n14927, n14928 );
nor U15035 ( n14928, n15165, n14738 );
nor U15036 ( n14927, n15149, n14739 );
nor U15037 ( n14925, n14929, n14930 );
nor U15038 ( n14930, n15133, n14742 );
nor U15039 ( n14929, n15157, n14743 );
nand U15040 ( n14923, n14931, n14932 );
nor U15041 ( n14932, n14933, n14934 );
nor U15042 ( n14934, n15181, n14748 );
nor U15043 ( n14933, n15173, n14749 );
nor U15044 ( n14931, n14935, n14936 );
nor U15045 ( n14936, n15141, n14752 );
nor U15046 ( n14935, n15189, n14753 );
nand U15047 ( n12765, n14937, n9422 );
not U15048 ( n9422, n10568 );
nand U15049 ( n10568, n14938, n14939 );
nor U15050 ( n14939, n14940, n14941 );
nand U15051 ( n14941, n14942, n14943 );
nor U15052 ( n14943, n14944, n14945 );
nor U15053 ( n14945, n15107, n14716 );
nand U15054 ( n14716, n14946, n11344 );
nor U15055 ( n14944, n15099, n14717 );
nand U15056 ( n14717, n14946, n11345 );
nor U15057 ( n14942, n14947, n14948 );
nor U15058 ( n14948, n15115, n14720 );
nand U15059 ( n14720, n14946, n11348 );
not U15060 ( n14946, n11377 );
nor U15061 ( n14947, n15123, n14721 );
nand U15062 ( n14721, n11358, n7816 );
nand U15063 ( n14940, n14949, n14950 );
nor U15064 ( n14950, n14951, n14952 );
nor U15065 ( n14952, n15075, n14726 );
nand U15066 ( n14726, n11344, n13895 );
nor U15067 ( n14951, n15067, n14727 );
nand U15068 ( n14727, n11345, n13895 );
nor U15069 ( n14949, n14953, n14954 );
nor U15070 ( n14954, n15083, n14730 );
nand U15071 ( n14730, n11348, n13895 );
nor U15072 ( n14953, n15091, n14731 );
nand U15073 ( n14731, n11349, n13895 );
nor U15074 ( n13895, n15193, n15194 );
nor U15075 ( n14938, n14955, n14956 );
nand U15076 ( n14956, n14957, n14958 );
nor U15077 ( n14958, n14959, n14960 );
nor U15078 ( n14960, n15163, n14738 );
nand U15079 ( n14738, n13898, n11345 );
nor U15080 ( n14959, n15147, n14739 );
nand U15081 ( n14739, n14961, n11348 );
nor U15082 ( n14957, n14962, n14963 );
nor U15083 ( n14963, n15131, n14742 );
nor U15084 ( n14962, n15155, n14743 );
nand U15085 ( n14743, n14961, n11349 );
not U15086 ( n11349, n11773 );
nand U15087 ( n14955, n14964, n14965 );
nor U15088 ( n14965, n14966, n14967 );
nor U15089 ( n14967, n15179, n14748 );
nand U15090 ( n14748, n13898, n11348 );
nor U15091 ( n11348, n7821, n15196 );
nor U15092 ( n14966, n15171, n14749 );
nand U15093 ( n14749, n13898, n11344 );
nor U15094 ( n13898, n7816, n7800 );
nor U15095 ( n14964, n14968, n14969 );
nor U15096 ( n14969, n15139, n14752 );
nand U15097 ( n14752, n14961, n11344 );
nor U15098 ( n11344, n7798, n15195 );
nor U15099 ( n14968, n15187, n14753 );
nand U15100 ( n14753, n15193, n11358 );
nor U15101 ( n11358, n7800, n11773 );
nor U15102 ( n14937, n15063, n13226 );
and U15103 ( n13226, n14970, n14971 );
nor U15104 ( n14971, n14972, n14973 );
nand U15105 ( n14973, n14974, n14975 );
nor U15106 ( n14975, n14976, n14977 );
nor U15107 ( n14977, n15080, n13410 );
nand U15108 ( n13410, n14978, n11742 );
nor U15109 ( n14976, n15088, n13411 );
nand U15110 ( n13411, n14978, n11741 );
nor U15111 ( n14974, n14979, n14980 );
nor U15112 ( n14980, n15072, n13414 );
nand U15113 ( n13414, n14978, n11738 );
nor U15114 ( n14979, n15064, n13415 );
nand U15115 ( n13415, n14978, n11737 );
nor U15116 ( n14978, n13876, n13890 );
nand U15117 ( n14972, n14981, n14982 );
nor U15118 ( n14982, n14983, n14984 );
nor U15119 ( n14984, n15112, n13400 );
nand U15120 ( n13400, n11742, n14985 );
nor U15121 ( n14983, n15120, n13401 );
nand U15122 ( n13401, n11741, n14985 );
nor U15123 ( n14981, n14986, n14987 );
nor U15124 ( n14987, n15104, n13404 );
nand U15125 ( n13404, n11738, n14985 );
nor U15126 ( n14986, n15096, n13405 );
nand U15127 ( n13405, n11737, n14985 );
nor U15128 ( n14985, n13869, n13890 );
not U15129 ( n13890, n13918 );
nor U15130 ( n14970, n14988, n14989 );
nand U15131 ( n14989, n14990, n14991 );
nor U15132 ( n14991, n14992, n14993 );
nor U15133 ( n14993, n15176, n13388 );
nand U15134 ( n13388, n14994, n11742 );
nor U15135 ( n14992, n15184, n13389 );
nand U15136 ( n13389, n14994, n11741 );
nor U15137 ( n14990, n14995, n14996 );
nor U15138 ( n14996, n15168, n13392 );
nand U15139 ( n13392, n14994, n11738 );
nor U15140 ( n14995, n15160, n13393 );
nand U15141 ( n13393, n14994, n11737 );
nor U15142 ( n14994, n13918, n13869 );
not U15143 ( n13869, n13876 );
nand U15144 ( n14988, n14997, n14998 );
nor U15145 ( n14998, n14999, n15000 );
nor U15146 ( n15000, n15144, n13378 );
nand U15147 ( n13378, n15001, n11742 );
nor U15148 ( n11742, n7798, n13854 );
nor U15149 ( n14999, n15152, n13379 );
nand U15150 ( n13379, n15001, n11741 );
nor U15151 ( n11741, n13854, n15196 );
not U15152 ( n13854, n15002 );
nor U15153 ( n14997, n15003, n15004 );
nor U15154 ( n15004, n15136, n13382 );
nand U15155 ( n13382, n15001, n11738 );
nor U15156 ( n11738, n15002, n15196 );
nor U15157 ( n15003, n15128, n13383 );
nand U15158 ( n13383, n15001, n11737 );
nor U15159 ( n11737, n15002, n7798 );
nand U15160 ( n15002, n13899, n11773 );
nand U15161 ( n11773, n15195, n15196 );
nor U15162 ( n15001, n13918, n13876 );
xnor U15163 ( n13876, n13899, n15194 );
nand U15164 ( n13918, n15005, n15006 );
nand U15165 ( n15006, n13899, n7816 );
and U15166 ( n15005, n11377, n14742 );
nand U15167 ( n14742, n14961, n11345 );
not U15168 ( n11345, n13899 );
nand U15169 ( n13899, n7821, n7798 );
not U15170 ( n14961, n11376 );
nand U15171 ( n11376, n15193, n7800 );
nand U15172 ( n11377, n15194, n7816 );
endmodule

