
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule
module b14_ori ( clk, reset, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
DATAI_1_, DATAI_0_, ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_,
ADDR_REG_16_, ADDR_REG_15_, ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_,
ADDR_REG_11_, ADDR_REG_10_, ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_,
ADDR_REG_6_, ADDR_REG_5_, ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_,
ADDR_REG_1_, ADDR_REG_0_, DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_,
DATAO_REG_28_, DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_,
DATAO_REG_24_, DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_,
DATAO_REG_20_, DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_,
DATAO_REG_16_, DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_,
DATAO_REG_12_, DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_,
DATAO_REG_8_, DATAO_REG_7_, DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_,
DATAO_REG_3_, DATAO_REG_2_, DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG
);
input clk, reset, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
DATAI_0_;
output ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_,
ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_,
ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_,
ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_,
DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_,
DATAO_REG_7_, DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_,
DATAO_REG_2_, DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG;
wire STATE_REG, n1337, n1327, n1322, n1317, n1312, n1307, n1302, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, n1297,
n1292, n1287, n1282, n1277, n1272, n1267, n1262, n1257, n1252, n1247,
n1242, n1237, n1232, n1227, n1222, n1217, n1212, n1207, n1202, n1197,
n1192, n1187, n1182, n1050, n1046, n1042, n1038, n1034, n1030, n1026,
n1022, n1018, n1014, n1010, n1006, n1002, n998, n994, n990, n986,
n982, n978, n974, n969, n964, n954, n949, n944, n939, n934, n929,
n924, n919, n914, n909, n904, n899, n894, n889, n884, n879, n874,
n869, n864, n859, n854, n849, n844, n839, n834, n829, n824, n819,
n814, D_REG_31_, n489, D_REG_30_, n484, D_REG_29_, n479, D_REG_28_,
n474, D_REG_27_, n469, D_REG_26_, n464, D_REG_25_, n459, D_REG_24_,
n454, D_REG_23_, n449, n444, D_REG_21_, n439, D_REG_20_, n434,
D_REG_19_, n429, D_REG_18_, n424, D_REG_17_, n419, D_REG_16_, n414,
D_REG_15_, n409, D_REG_14_, n404, D_REG_13_, n399, D_REG_12_, n394,
D_REG_11_, n389, D_REG_10_, n384, D_REG_9_, n379, D_REG_8_, n374,
n369, D_REG_6_, n364, D_REG_5_, n359, D_REG_4_, n354, D_REG_3_, n349,
D_REG_2_, n344, n329, n324, n319, n314, n309, n304, n299, n294, n289,
n284, n279, n274, n269, n264, n259, n254, n249, n244, n239, n234,
n229, n224, n219, n214, n209, n204, n199, n194, n189, n184, n179,
n174, n959, B_REG, REG2_REG_0_, n334, n339, n494, n499, n504, n509,
n514, n519, n524, n529, n534, n539, n544, n549, n554, n559, n564,
n569, n574, n579, n584, n589, n594, n599, n604, n609, n614, n619,
n624, n629, n634, n639, n644, n649, n654, n659, n664, n669, n674,
n679, n684, n689, n694, n699, n704, n709, n714, n719, n724, n729,
n734, n739, n744, n749, n754, n759, n764, n769, n774, n779, n784,
n789, n794, n799, n804, n809, n1054, n1058, n1062, n1066, n1070,
n1074, n1078, n1082, n1086, n1090, n1094, n1098, n1102, n1106, n1110,
n1114, n1118, n1122, n1126, n1130, n1134, n1138, n1142, n1146, n1150,
n1154, n1158, n1162, n1166, n1170, n1174, n1178, IR_REG_31_,
IR_REG_0_, IR_REG_1_, IR_REG_2_, IR_REG_3_, IR_REG_4_, IR_REG_5_,
IR_REG_6_, IR_REG_7_, IR_REG_8_, IR_REG_9_, IR_REG_10_, IR_REG_11_,
IR_REG_12_, IR_REG_13_, IR_REG_14_, IR_REG_15_, IR_REG_16_,
IR_REG_17_, IR_REG_18_, IR_REG_19_, IR_REG_20_, IR_REG_21_,
IR_REG_22_, IR_REG_23_, IR_REG_24_, IR_REG_25_, IR_REG_26_,
IR_REG_27_, IR_REG_28_, IR_REG_29_, IR_REG_30_, REG2_REG_1_,
REG1_REG_1_, REG0_REG_1_, REG3_REG_1_, REG2_REG_2_, REG1_REG_2_,
REG0_REG_2_, REG3_REG_2_, REG0_REG_0_, REG1_REG_0_, REG2_REG_3_,
REG1_REG_3_, REG0_REG_3_, REG2_REG_4_, REG1_REG_4_, REG0_REG_4_,
REG2_REG_5_, REG1_REG_5_, REG0_REG_5_, REG2_REG_6_, REG1_REG_6_,
REG0_REG_6_, REG2_REG_7_, REG1_REG_7_, REG0_REG_7_, REG2_REG_8_,
REG1_REG_8_, REG0_REG_8_, REG2_REG_9_, REG1_REG_9_, REG0_REG_9_,
REG2_REG_10_, REG1_REG_10_, REG0_REG_10_, REG2_REG_11_, REG1_REG_11_,
REG0_REG_11_, REG2_REG_12_, REG1_REG_12_, REG0_REG_12_, REG2_REG_13_,
REG1_REG_13_, REG0_REG_13_, REG2_REG_14_, REG1_REG_14_, REG0_REG_14_,
REG2_REG_15_, REG1_REG_15_, REG0_REG_15_, REG2_REG_16_, REG1_REG_16_,
REG0_REG_16_, REG2_REG_17_, REG1_REG_17_, REG0_REG_17_, REG2_REG_18_,
REG1_REG_18_, REG0_REG_18_, REG2_REG_19_, REG1_REG_19_, REG0_REG_19_,
REG1_REG_20_, REG0_REG_20_, REG1_REG_21_, REG0_REG_21_, REG1_REG_22_,
REG0_REG_22_, REG1_REG_23_, REG0_REG_23_, REG1_REG_24_, REG0_REG_24_,
REG1_REG_25_, REG0_REG_25_, REG1_REG_26_, REG0_REG_26_, REG1_REG_27_,
REG0_REG_27_, REG1_REG_28_, REG0_REG_28_, REG1_REG_29_, REG0_REG_29_,
REG1_REG_30_, REG0_REG_30_, REG1_REG_31_, REG0_REG_31_, REG3_REG_19_,
REG3_REG_18_, REG3_REG_17_, REG3_REG_16_, REG3_REG_15_, REG3_REG_14_,
REG3_REG_13_, REG3_REG_12_, REG3_REG_11_, REG3_REG_10_, REG3_REG_9_,
REG3_REG_8_, REG3_REG_7_, REG3_REG_6_, REG3_REG_5_, REG3_REG_4_,
REG3_REG_3_, REG3_REG_26_, REG3_REG_22_, REG3_REG_20_, REG3_REG_24_,
REG3_REG_25_, REG3_REG_21_, REG3_REG_28_, REG3_REG_23_, REG3_REG_27_,
D_REG_0_, D_REG_1_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
n13, n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
n42, n43, n44, n45, n46, n47, n49, n50, n51, n52, n53, n54, n55, n56,
n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70, n71,
n72, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n87, n88, n89,
n90, n92, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n106,
n107, n108, n109, n110, n111, n112, n113, n114, n116, n118, n119,
n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
n131, n132, n133, n135, n136, n137, n139, n140, n141, n142, n143,
n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
n166, n167, n168, n169, n170, n171, n172, n173, n175, n176, n177,
n178, n180, n181, n182, n183, n185, n186, n187, n188, n190, n191,
n192, n193, n195, n196, n197, n198, n200, n201, n202, n203, n205,
n206, n207, n208, n210, n211, n212, n213, n215, n216, n217, n218,
n220, n221, n222, n225, n226, n227, n228, n230, n231, n232, n233,
n235, n236, n237, n238, n240, n241, n242, n245, n247, n248, n250,
n251, n252, n253, n255, n256, n257, n258, n260, n261, n262, n263,
n265, n266, n267, n268, n270, n271, n272, n273, n275, n276, n278,
n280, n281, n282, n283, n285, n286, n287, n288, n290, n291, n292,
n293, n295, n296, n297, n298, n300, n301, n302, n303, n305, n306,
n307, n308, n310, n311, n312, n313, n315, n316, n317, n318, n320,
n321, n322, n323, n325, n326, n327, n328, n331, n332, n333, n335,
n336, n337, n338, n340, n341, n342, n343, n345, n346, n347, n388,
n473, n475, n476, n477, n478, n480, n481, n482, n483, n485, n486,
n487, n488, n491, n492, n493, n495, n496, n497, n498, n500, n501,
n502, n512, n513, n536, n537, n538, n540, n541, n542, n543, n545,
n546, n547, n548, n550, n551, n552, n553, n555, n556, n557, n558,
n560, n561, n562, n563, n565, n566, n567, n568, n570, n571, n572,
n573, n575, n576, n577, n578, n580, n581, n582, n583, n585, n586,
n587, n588, n590, n591, n592, n593, n595, n596, n597, n598, n600,
n601, n602, n603, n605, n606, n607, n608, n610, n611, n612, n613,
n615, n616, n617, n618, n620, n621, n622, n623, n625, n626, n627,
n628, n630, n631, n632, n633, n635, n636, n637, n638, n640, n641,
n642, n643, n645, n646, n647, n648, n650, n651, n652, n653, n655,
n656, n657, n658, n660, n661, n662, n663, n665, n666, n667, n668,
n670, n671, n672, n673, n675, n676, n677, n678, n680, n681, n682,
n683, n685, n686, n687, n688, n690, n691, n692, n693, n695, n696,
n697, n698, n700, n701, n702, n703, n705, n706, n707, n708, n710,
n711, n712, n713, n715, n716, n717, n718, n720, n721, n722, n723,
n725, n726, n727, n728, n730, n731, n732, n733, n735, n736, n737,
n738, n740, n741, n742, n743, n745, n746, n747, n748, n750, n751,
n752, n753, n755, n756, n757, n758, n760, n761, n762, n763, n765,
n766, n767, n768, n770, n771, n772, n773, n775, n776, n777, n778,
n780, n781, n782, n783, n785, n786, n788, n790, n791, n792, n793,
n795, n796, n797, n798, n800, n801, n802, n803, n805, n806, n807,
n808, n810, n811, n812, n813, n815, n816, n817, n818, n820, n821,
n822, n823, n825, n826, n827, n828, n830, n831, n832, n833, n835,
n836, n837, n838, n840, n841, n842, n843, n845, n846, n847, n848,
n850, n851, n852, n853, n855, n856, n857, n858, n860, n861, n862,
n863, n865, n866, n867, n868, n870, n871, n872, n873, n875, n876,
n877, n878, n880, n881, n882, n883, n885, n886, n887, n888, n890,
n891, n892, n893, n895, n896, n897, n898, n900, n901, n902, n903,
n905, n906, n907, n908, n910, n911, n912, n913, n915, n916, n917,
n918, n920, n921, n922, n923, n925, n926, n927, n928, n930, n931,
n932, n933, n935, n936, n937, n938, n940, n941, n942, n943, n945,
n946, n947, n948, n950, n951, n952, n953, n955, n956, n957, n958,
n960, n961, n962, n963, n965, n966, n967, n968, n970, n971, n972,
n973, n975, n976, n977, n979, n980, n981, n983, n984, n985, n987,
n988, n989, n991, n992, n993, n995, n996, n997, n999, n1000, n1001,
n1003, n1004, n1005, n1007, n1008, n1009, n1011, n1012, n1013, n1015,
n1016, n1017, n1019, n1020, n1021, n1023, n1024, n1025, n1027, n1028,
n1029, n1031, n1032, n1033, n1035, n1036, n1037, n1039, n1040, n1041,
n1043, n1044, n1045, n1047, n1048, n1049, n1051, n1052, n1053, n1055,
n1056, n1057, n1059, n1060, n1061, n1063, n1064, n1065, n1067, n1068,
n1069, n1071, n1072, n1073, n1075, n1076, n1077, n1079, n1080, n1081,
n1083, n1084, n1085, n1087, n1088, n1089, n1091, n1092, n1093, n1095,
n1096, n1097, n1099, n1100, n1101, n1103, n1104, n1105, n1107, n1108,
n1109, n1111, n1112, n1113, n1115, n1116, n1117, n1119, n1120, n1121,
n1123, n1124, n1125, n1127, n1128, n1129, n1131, n1132, n1133, n1135,
n1136, n1137, n1139, n1140, n1141, n1143, n1144, n1145, n1147, n1148,
n1149, n1151, n1152, n1153, n1155, n1156, n1157, n1159, n1160, n1161,
n1163, n1164, n1165, n1167, n1168, n1169, n1171, n1172, n1173, n1175,
n1176, n1177, n1179, n1180, n1181, n1183, n1184, n1185, n1186, n1188,
n1189, n1190, n1191, n1193, n1194, n1195, n1196, n1198, n1199, n1200,
n1201, n1203, n1204, n1205, n1206, n1208, n1209, n1210, n1211, n1213,
n1214, n1215, n1216, n1218, n1219, n1220, n1221, n1223, n1224, n1225,
n1226, n1228, n1229, n1230, n1231, n1233, n1234, n1235, n1236, n1238,
n1239, n1240, n1241, n1243, n1244, n1245, n1246, n1248, n1249, n1250,
n1251, n1253, n1254, n1255, n1256, n1258, n1259, n1260, n1261, n1263,
n1264, n1265, n1266, n1268, n1269, n1270, n1271, n1273, n1274, n1275,
n1276, n1278, n1279, n1280, n1281, n1283, n1284, n1285, n1286, n1288,
n1289, n1290, n1291, n1293, n1294, n1295, n1296, n1298, n1299, n1300,
n1301, n1303, n1304, n1305, n1306, n1308, n1309, n1310, n1311, n1313,
n1314, n1315, n1316, n1318, n1319, n1320, n1321, n1323, n1324, n1325,
n1326, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1498, n1499,
n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1538, n1539, n1540,
n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1590, n1591,
n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
n1722, n1723, n1724, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1764,
n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2027,
n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2036, n2037, n2038,
n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
n2129, n2130, n2131, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
n2251, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
n2824, n2825, n2826, n2827, n2828, n2830, n2831, n2832, n2833, n2834,
n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
n2845, n2846, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3175, n3176,
n3177, n3178, n3179, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3358,
n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
n3939, n3940, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
n4940, n4941, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
n5242, n5243, n5244, n5245, n5246, n5247, n5248;

dff STATE_REG_reg ( clk, reset, STATE_REG, n5246 );
not U_inv0 ( n4978, STATE_REG );
dff IR_REG_0__reg ( clk, reset, IR_REG_0_, n174 );
not U_inv1 ( n4979, IR_REG_0_ );
dff IR_REG_1__reg ( clk, reset, IR_REG_1_, n179 );
not U_inv2 ( n4989, IR_REG_1_ );
dff IR_REG_2__reg ( clk, reset, IR_REG_2_, n184 );
not U_inv3 ( n5088, IR_REG_2_ );
dff IR_REG_3__reg ( clk, reset, IR_REG_3_, n189 );
not U_inv4 ( n4990, IR_REG_3_ );
dff IR_REG_4__reg ( clk, reset, IR_REG_4_, n194 );
not U_inv5 ( n4980, IR_REG_4_ );
dff IR_REG_6__reg ( clk, reset, IR_REG_6_, n204 );
not U_inv6 ( n5000, IR_REG_6_ );
dff IR_REG_5__reg ( clk, reset, IR_REG_5_, n199 );
not U_inv7 ( n5001, IR_REG_5_ );
dff IR_REG_7__reg ( clk, reset, IR_REG_7_, n209 );
not U_inv8 ( n5086, IR_REG_7_ );
dff IR_REG_8__reg ( clk, reset, IR_REG_8_, n214 );
not U_inv9 ( n5014, IR_REG_8_ );
dff IR_REG_9__reg ( clk, reset, IR_REG_9_, n219 );
not U_inv10 ( n5085, IR_REG_9_ );
dff IR_REG_10__reg ( clk, reset, IR_REG_10_, n224 );
not U_inv11 ( n5021, IR_REG_10_ );
dff IR_REG_11__reg ( clk, reset, IR_REG_11_, n229 );
not U_inv12 ( n5084, IR_REG_11_ );
dff IR_REG_12__reg ( clk, reset, IR_REG_12_, n234 );
not U_inv13 ( n5017, IR_REG_12_ );
dff IR_REG_13__reg ( clk, reset, IR_REG_13_, n239 );
not U_inv14 ( n5083, IR_REG_13_ );
dff IR_REG_14__reg ( clk, reset, IR_REG_14_, n244 );
not U_inv15 ( n4982, IR_REG_14_ );
dff IR_REG_15__reg ( clk, reset, IR_REG_15_, n249 );
not U_inv16 ( n4984, IR_REG_15_ );
dff IR_REG_16__reg ( clk, reset, IR_REG_16_, n254 );
not U_inv17 ( n5034, IR_REG_16_ );
dff IR_REG_17__reg ( clk, reset, IR_REG_17_, n259 );
not U_inv18 ( n5080, IR_REG_17_ );
dff IR_REG_18__reg ( clk, reset, IR_REG_18_, n264 );
not U_inv19 ( n4981, IR_REG_18_ );
dff IR_REG_19__reg ( clk, reset, IR_REG_19_, n269 );
not U_inv20 ( n5078, IR_REG_19_ );
dff IR_REG_20__reg ( clk, reset, IR_REG_20_, n274 );
not U_inv21 ( n4985, IR_REG_20_ );
dff IR_REG_21__reg ( clk, reset, IR_REG_21_, n279 );
not U_inv22 ( n4983, IR_REG_21_ );
dff IR_REG_22__reg ( clk, reset, IR_REG_22_, n284 );
not U_inv23 ( n5077, IR_REG_22_ );
dff IR_REG_23__reg ( clk, reset, IR_REG_23_, n289 );
not U_inv24 ( n5063, IR_REG_23_ );
dff IR_REG_24__reg ( clk, reset, IR_REG_24_, n294 );
not U_inv25 ( n4986, IR_REG_24_ );
dff IR_REG_25__reg ( clk, reset, IR_REG_25_, n299 );
not U_inv26 ( n5082, IR_REG_25_ );
dff IR_REG_26__reg ( clk, reset, IR_REG_26_, n304 );
not U_inv27 ( n5079, IR_REG_26_ );
dff IR_REG_27__reg ( clk, reset, IR_REG_27_, n309 );
not U_inv28 ( n4987, IR_REG_27_ );
dff IR_REG_28__reg ( clk, reset, IR_REG_28_, n314 );
not U_inv29 ( n5081, IR_REG_28_ );
dff IR_REG_29__reg ( clk, reset, IR_REG_29_, n319 );
not U_inv30 ( n5087, IR_REG_29_ );
dff IR_REG_30__reg ( clk, reset, IR_REG_30_, n324 );
not U_inv31 ( n4988, IR_REG_30_ );
dff REG3_REG_12__reg ( clk, reset, REG3_REG_12_, n1272 );
not U_inv32 ( n5022, REG3_REG_12_ );
dff B_REG_reg ( clk, reset, B_REG, n1182 );
not U_inv33 ( n5058, B_REG );
dff D_REG_22__reg ( clk, reset, ex_wire0, n444 );
not U_inv34 ( n5064, ex_wire0 );
dff D_REG_7__reg ( clk, reset, ex_wire1, n369 );
not U_inv35 ( n5065, ex_wire1 );
dff D_REG_31__reg ( clk, reset, D_REG_31_, n489 );
dff D_REG_30__reg ( clk, reset, D_REG_30_, n484 );
dff D_REG_29__reg ( clk, reset, D_REG_29_, n479 );
dff D_REG_28__reg ( clk, reset, D_REG_28_, n474 );
dff D_REG_27__reg ( clk, reset, D_REG_27_, n469 );
dff D_REG_26__reg ( clk, reset, D_REG_26_, n464 );
dff D_REG_25__reg ( clk, reset, D_REG_25_, n459 );
dff D_REG_24__reg ( clk, reset, D_REG_24_, n454 );
dff D_REG_23__reg ( clk, reset, D_REG_23_, n449 );
dff D_REG_21__reg ( clk, reset, D_REG_21_, n439 );
dff D_REG_20__reg ( clk, reset, D_REG_20_, n434 );
dff D_REG_19__reg ( clk, reset, D_REG_19_, n429 );
dff D_REG_18__reg ( clk, reset, D_REG_18_, n424 );
dff D_REG_17__reg ( clk, reset, D_REG_17_, n419 );
dff D_REG_16__reg ( clk, reset, D_REG_16_, n414 );
dff D_REG_15__reg ( clk, reset, D_REG_15_, n409 );
dff D_REG_14__reg ( clk, reset, D_REG_14_, n404 );
dff D_REG_13__reg ( clk, reset, D_REG_13_, n399 );
dff D_REG_12__reg ( clk, reset, D_REG_12_, n394 );
dff D_REG_11__reg ( clk, reset, D_REG_11_, n389 );
dff D_REG_10__reg ( clk, reset, D_REG_10_, n384 );
dff D_REG_9__reg ( clk, reset, D_REG_9_, n379 );
dff D_REG_8__reg ( clk, reset, D_REG_8_, n374 );
dff D_REG_6__reg ( clk, reset, D_REG_6_, n364 );
dff D_REG_5__reg ( clk, reset, D_REG_5_, n359 );
dff D_REG_4__reg ( clk, reset, D_REG_4_, n354 );
dff D_REG_3__reg ( clk, reset, D_REG_3_, n349 );
dff D_REG_2__reg ( clk, reset, D_REG_2_, n344 );
dff D_REG_1__reg ( clk, reset, D_REG_1_, n339 );
dff D_REG_0__reg ( clk, reset, D_REG_0_, n334 );
dff REG2_REG_31__reg ( clk, reset, ex_wire2, n969 );
not U_inv36 ( n5073, ex_wire2 );
dff REG1_REG_31__reg ( clk, reset, REG1_REG_31_, n809 );
not U_inv37 ( n5072, REG1_REG_31_ );
dff REG0_REG_31__reg ( clk, reset, REG0_REG_31_, n649 );
dff REG1_REG_30__reg ( clk, reset, REG1_REG_30_, n804 );
not U_inv38 ( n5074, REG1_REG_30_ );
dff REG0_REG_30__reg ( clk, reset, REG0_REG_30_, n644 );
dff DATAO_REG_31__reg ( clk, reset, DATAO_REG_31_, n1178 );
dff REG2_REG_30__reg ( clk, reset, ex_wire3, n964 );
not U_inv39 ( n5075, ex_wire3 );
dff DATAO_REG_30__reg ( clk, reset, DATAO_REG_30_, n1174 );
dff REG3_REG_2__reg ( clk, reset, REG3_REG_2_, n1207 );
not U_inv40 ( n4995, REG3_REG_2_ );
dff REG2_REG_2__reg ( clk, reset, REG2_REG_2_, n824 );
not U_inv41 ( n4996, REG2_REG_2_ );
dff REG2_REG_1__reg ( clk, reset, REG2_REG_1_, n819 );
not U_inv42 ( n4991, REG2_REG_1_ );
dff REG2_REG_0__reg ( clk, reset, REG2_REG_0_, n814 );
not U_inv43 ( n4993, REG2_REG_0_ );
dff REG1_REG_0__reg ( clk, reset, REG1_REG_0_, n654 );
not U_inv44 ( n4994, REG1_REG_0_ );
dff REG3_REG_0__reg ( clk, reset, ex_wire4, n1232 );
not U_inv45 ( n4967, ex_wire4 );
dff REG0_REG_0__reg ( clk, reset, REG0_REG_0_, n494 );
dff DATAO_REG_0__reg ( clk, reset, DATAO_REG_0_, n1054 );
dff REG3_REG_1__reg ( clk, reset, REG3_REG_1_, n1282 );
not U_inv46 ( n4966, REG3_REG_1_ );
dff REG1_REG_1__reg ( clk, reset, REG1_REG_1_, n659 );
not U_inv47 ( n4992, REG1_REG_1_ );
dff REG0_REG_1__reg ( clk, reset, REG0_REG_1_, n499 );
dff DATAO_REG_1__reg ( clk, reset, DATAO_REG_1_, n1058 );
dff REG1_REG_3__reg ( clk, reset, REG1_REG_3_, n669 );
not U_inv48 ( n4999, REG1_REG_3_ );
dff REG0_REG_3__reg ( clk, reset, REG0_REG_3_, n509 );
dff REG1_REG_2__reg ( clk, reset, REG1_REG_2_, n664 );
not U_inv49 ( n4997, REG1_REG_2_ );
dff REG0_REG_2__reg ( clk, reset, REG0_REG_2_, n504 );
dff REG1_REG_4__reg ( clk, reset, REG1_REG_4_, n674 );
not U_inv50 ( n5006, REG1_REG_4_ );
dff REG0_REG_4__reg ( clk, reset, REG0_REG_4_, n514 );
dff REG3_REG_3__reg ( clk, reset, REG3_REG_3_, n1302 );
not U_inv51 ( n5076, REG3_REG_3_ );
dff REG1_REG_5__reg ( clk, reset, REG1_REG_5_, n679 );
not U_inv52 ( n5008, REG1_REG_5_ );
dff REG0_REG_5__reg ( clk, reset, REG0_REG_5_, n519 );
dff REG3_REG_4__reg ( clk, reset, REG3_REG_4_, n1242 );
not U_inv53 ( n5003, REG3_REG_4_ );
dff REG2_REG_4__reg ( clk, reset, REG2_REG_4_, n834 );
not U_inv54 ( n5005, REG2_REG_4_ );
dff REG1_REG_6__reg ( clk, reset, REG1_REG_6_, n684 );
not U_inv55 ( n5010, REG1_REG_6_ );
dff REG0_REG_6__reg ( clk, reset, REG0_REG_6_, n524 );
dff REG3_REG_5__reg ( clk, reset, REG3_REG_5_, n1257 );
not U_inv56 ( n5002, REG3_REG_5_ );
dff REG2_REG_5__reg ( clk, reset, REG2_REG_5_, n839 );
not U_inv57 ( n5007, REG2_REG_5_ );
dff REG3_REG_11__reg ( clk, reset, REG3_REG_11_, n1212 );
not U_inv58 ( n5018, REG3_REG_11_ );
dff REG2_REG_10__reg ( clk, reset, REG2_REG_10_, n864 );
not U_inv59 ( n5028, REG2_REG_10_ );
dff REG2_REG_9__reg ( clk, reset, REG2_REG_9_, n859 );
not U_inv60 ( n5023, REG2_REG_9_ );
dff REG2_REG_8__reg ( clk, reset, REG2_REG_8_, n854 );
not U_inv61 ( n5019, REG2_REG_8_ );
dff REG2_REG_7__reg ( clk, reset, REG2_REG_7_, n849 );
not U_inv62 ( n5011, REG2_REG_7_ );
dff REG3_REG_6__reg ( clk, reset, REG3_REG_6_, n1197 );
not U_inv63 ( n5004, REG3_REG_6_ );
dff REG2_REG_6__reg ( clk, reset, REG2_REG_6_, n844 );
not U_inv64 ( n5009, REG2_REG_6_ );
dff REG3_REG_7__reg ( clk, reset, REG3_REG_7_, n1327 );
not U_inv65 ( n5013, REG3_REG_7_ );
dff REG1_REG_7__reg ( clk, reset, REG1_REG_7_, n689 );
not U_inv66 ( n5012, REG1_REG_7_ );
dff REG0_REG_7__reg ( clk, reset, REG0_REG_7_, n529 );
dff REG1_REG_8__reg ( clk, reset, REG1_REG_8_, n694 );
not U_inv67 ( n5020, REG1_REG_8_ );
dff REG0_REG_8__reg ( clk, reset, REG0_REG_8_, n534 );
dff DATAO_REG_7__reg ( clk, reset, DATAO_REG_7_, n1082 );
dff REG3_REG_8__reg ( clk, reset, REG3_REG_8_, n1287 );
not U_inv68 ( n5016, REG3_REG_8_ );
dff DATAO_REG_8__reg ( clk, reset, DATAO_REG_8_, n1086 );
dff REG3_REG_9__reg ( clk, reset, REG3_REG_9_, n1237 );
not U_inv69 ( n5015, REG3_REG_9_ );
dff REG1_REG_9__reg ( clk, reset, REG1_REG_9_, n699 );
not U_inv70 ( n5024, REG1_REG_9_ );
dff REG0_REG_9__reg ( clk, reset, REG0_REG_9_, n539 );
dff DATAO_REG_9__reg ( clk, reset, DATAO_REG_9_, n1090 );
dff REG3_REG_10__reg ( clk, reset, REG3_REG_10_, n1307 );
not U_inv71 ( n5025, REG3_REG_10_ );
dff REG1_REG_10__reg ( clk, reset, REG1_REG_10_, n704 );
not U_inv72 ( n5029, REG1_REG_10_ );
dff REG0_REG_10__reg ( clk, reset, REG0_REG_10_, n544 );
dff DATAO_REG_10__reg ( clk, reset, DATAO_REG_10_, n1094 );
dff REG1_REG_12__reg ( clk, reset, REG1_REG_12_, n714 );
not U_inv73 ( n5027, REG1_REG_12_ );
dff REG0_REG_12__reg ( clk, reset, REG0_REG_12_, n554 );
dff REG1_REG_11__reg ( clk, reset, REG1_REG_11_, n709 );
not U_inv74 ( n5033, REG1_REG_11_ );
dff REG0_REG_11__reg ( clk, reset, REG0_REG_11_, n549 );
dff REG2_REG_11__reg ( clk, reset, REG2_REG_11_, n869 );
not U_inv75 ( n5031, REG2_REG_11_ );
dff REG2_REG_12__reg ( clk, reset, REG2_REG_12_, n874 );
not U_inv76 ( n5026, REG2_REG_12_ );
dff DATAO_REG_12__reg ( clk, reset, DATAO_REG_12_, n1102 );
dff DATAO_REG_11__reg ( clk, reset, DATAO_REG_11_, n1098 );
dff REG3_REG_15__reg ( clk, reset, REG3_REG_15_, n1187 );
not U_inv77 ( n4969, REG3_REG_15_ );
dff REG2_REG_14__reg ( clk, reset, REG2_REG_14_, n884 );
not U_inv78 ( n5035, REG2_REG_14_ );
dff REG1_REG_13__reg ( clk, reset, REG1_REG_13_, n719 );
not U_inv79 ( n5032, REG1_REG_13_ );
dff REG0_REG_13__reg ( clk, reset, REG0_REG_13_, n559 );
dff REG3_REG_13__reg ( clk, reset, REG3_REG_13_, n1222 );
not U_inv80 ( n4968, REG3_REG_13_ );
dff REG2_REG_13__reg ( clk, reset, REG2_REG_13_, n879 );
not U_inv81 ( n5030, REG2_REG_13_ );
dff REG3_REG_14__reg ( clk, reset, REG3_REG_14_, n1317 );
not U_inv82 ( n4970, REG3_REG_14_ );
dff REG1_REG_14__reg ( clk, reset, REG1_REG_14_, n724 );
not U_inv83 ( n5036, REG1_REG_14_ );
dff REG0_REG_14__reg ( clk, reset, REG0_REG_14_, n564 );
dff DATAO_REG_14__reg ( clk, reset, DATAO_REG_14_, n1110 );
dff REG1_REG_16__reg ( clk, reset, REG1_REG_16_, n734 );
not U_inv84 ( n5039, REG1_REG_16_ );
dff REG0_REG_16__reg ( clk, reset, REG0_REG_16_, n574 );
dff REG3_REG_26__reg ( clk, reset, REG3_REG_26_, n1192 );
dff REG2_REG_25__reg ( clk, reset, ex_wire5, n939 );
not U_inv85 ( n5061, ex_wire5 );
dff REG2_REG_24__reg ( clk, reset, ex_wire6, n934 );
not U_inv86 ( n5056, ex_wire6 );
dff REG2_REG_23__reg ( clk, reset, ex_wire7, n929 );
not U_inv87 ( n5054, ex_wire7 );
dff REG2_REG_22__reg ( clk, reset, ex_wire8, n924 );
not U_inv88 ( n5052, ex_wire8 );
dff REG2_REG_21__reg ( clk, reset, ex_wire9, n919 );
not U_inv89 ( n5049, ex_wire9 );
dff REG2_REG_20__reg ( clk, reset, ex_wire10, n914 );
not U_inv90 ( n5044, ex_wire10 );
dff REG2_REG_19__reg ( clk, reset, REG2_REG_19_, n909 );
not U_inv91 ( n5045, REG2_REG_19_ );
dff REG2_REG_18__reg ( clk, reset, REG2_REG_18_, n904 );
not U_inv92 ( n5048, REG2_REG_18_ );
dff REG2_REG_17__reg ( clk, reset, REG2_REG_17_, n899 );
not U_inv93 ( n5042, REG2_REG_17_ );
dff REG3_REG_16__reg ( clk, reset, REG3_REG_16_, n1262 );
not U_inv94 ( n4971, REG3_REG_16_ );
dff REG2_REG_16__reg ( clk, reset, REG2_REG_16_, n894 );
not U_inv95 ( n5038, REG2_REG_16_ );
dff REG3_REG_17__reg ( clk, reset, REG3_REG_17_, n1252 );
not U_inv96 ( n4972, REG3_REG_17_ );
dff REG1_REG_17__reg ( clk, reset, REG1_REG_17_, n739 );
not U_inv97 ( n5043, REG1_REG_17_ );
dff REG0_REG_17__reg ( clk, reset, REG0_REG_17_, n579 );
dff DATAO_REG_17__reg ( clk, reset, DATAO_REG_17_, n1122 );
dff REG3_REG_18__reg ( clk, reset, REG3_REG_18_, n1202 );
not U_inv98 ( n4974, REG3_REG_18_ );
dff REG1_REG_18__reg ( clk, reset, REG1_REG_18_, n744 );
not U_inv99 ( n5051, REG1_REG_18_ );
dff REG0_REG_18__reg ( clk, reset, REG0_REG_18_, n584 );
dff DATAO_REG_18__reg ( clk, reset, DATAO_REG_18_, n1126 );
dff REG3_REG_19__reg ( clk, reset, REG3_REG_19_, n1297 );
not U_inv100 ( n4973, REG3_REG_19_ );
dff REG1_REG_19__reg ( clk, reset, REG1_REG_19_, n749 );
not U_inv101 ( n5046, REG1_REG_19_ );
dff REG0_REG_19__reg ( clk, reset, REG0_REG_19_, n589 );
dff DATAO_REG_19__reg ( clk, reset, DATAO_REG_19_, n1130 );
dff REG3_REG_20__reg ( clk, reset, REG3_REG_20_, n1227 );
dff REG1_REG_20__reg ( clk, reset, REG1_REG_20_, n754 );
not U_inv102 ( n5047, REG1_REG_20_ );
dff REG0_REG_20__reg ( clk, reset, REG0_REG_20_, n594 );
dff DATAO_REG_20__reg ( clk, reset, DATAO_REG_20_, n1134 );
dff REG3_REG_21__reg ( clk, reset, REG3_REG_21_, n1277 );
not U_inv103 ( n5041, REG3_REG_21_ );
dff REG1_REG_21__reg ( clk, reset, REG1_REG_21_, n759 );
not U_inv104 ( n5050, REG1_REG_21_ );
dff REG0_REG_21__reg ( clk, reset, REG0_REG_21_, n599 );
dff DATAO_REG_21__reg ( clk, reset, DATAO_REG_21_, n1138 );
dff REG3_REG_22__reg ( clk, reset, REG3_REG_22_, n1217 );
dff REG1_REG_22__reg ( clk, reset, REG1_REG_22_, n764 );
not U_inv105 ( n5053, REG1_REG_22_ );
dff REG0_REG_22__reg ( clk, reset, REG0_REG_22_, n604 );
dff DATAO_REG_22__reg ( clk, reset, DATAO_REG_22_, n1142 );
dff REG3_REG_23__reg ( clk, reset, REG3_REG_23_, n1312 );
not U_inv106 ( n4975, REG3_REG_23_ );
dff REG1_REG_23__reg ( clk, reset, REG1_REG_23_, n769 );
not U_inv107 ( n5055, REG1_REG_23_ );
dff REG0_REG_23__reg ( clk, reset, REG0_REG_23_, n609 );
dff DATAO_REG_23__reg ( clk, reset, DATAO_REG_23_, n1146 );
dff REG3_REG_24__reg ( clk, reset, REG3_REG_24_, n1247 );
dff REG1_REG_24__reg ( clk, reset, REG1_REG_24_, n774 );
not U_inv108 ( n5057, REG1_REG_24_ );
dff REG0_REG_24__reg ( clk, reset, REG0_REG_24_, n614 );
dff DATAO_REG_24__reg ( clk, reset, DATAO_REG_24_, n1150 );
dff REG3_REG_25__reg ( clk, reset, REG3_REG_25_, n1267 );
not U_inv109 ( n4976, REG3_REG_25_ );
dff REG1_REG_25__reg ( clk, reset, REG1_REG_25_, n779 );
not U_inv110 ( n5062, REG1_REG_25_ );
dff REG0_REG_25__reg ( clk, reset, REG0_REG_25_, n619 );
dff DATAO_REG_25__reg ( clk, reset, DATAO_REG_25_, n1154 );
dff REG1_REG_27__reg ( clk, reset, REG1_REG_27_, n789 );
not U_inv111 ( n5069, REG1_REG_27_ );
dff REG0_REG_27__reg ( clk, reset, REG0_REG_27_, n629 );
dff REG1_REG_28__reg ( clk, reset, REG1_REG_28_, n794 );
not U_inv112 ( n5070, REG1_REG_28_ );
dff REG0_REG_28__reg ( clk, reset, REG0_REG_28_, n634 );
dff REG3_REG_27__reg ( clk, reset, REG3_REG_27_, n1322 );
not U_inv113 ( n4977, REG3_REG_27_ );
dff REG1_REG_29__reg ( clk, reset, REG1_REG_29_, n799 );
not U_inv114 ( n5071, REG1_REG_29_ );
dff REG0_REG_29__reg ( clk, reset, REG0_REG_29_, n639 );
dff REG3_REG_28__reg ( clk, reset, REG3_REG_28_, n1292 );
dff REG2_REG_29__reg ( clk, reset, ex_wire11, n959 );
not U_inv115 ( n5067, ex_wire11 );
dff DATAO_REG_29__reg ( clk, reset, DATAO_REG_29_, n1170 );
dff REG2_REG_28__reg ( clk, reset, ex_wire12, n954 );
not U_inv116 ( n5068, ex_wire12 );
dff DATAO_REG_28__reg ( clk, reset, DATAO_REG_28_, n1166 );
dff REG2_REG_27__reg ( clk, reset, ex_wire13, n949 );
not U_inv117 ( n5066, ex_wire13 );
dff DATAO_REG_27__reg ( clk, reset, DATAO_REG_27_, n1162 );
dff REG2_REG_26__reg ( clk, reset, ex_wire14, n944 );
not U_inv118 ( n5059, ex_wire14 );
dff REG1_REG_26__reg ( clk, reset, REG1_REG_26_, n784 );
not U_inv119 ( n5060, REG1_REG_26_ );
dff REG0_REG_26__reg ( clk, reset, REG0_REG_26_, n624 );
dff DATAO_REG_26__reg ( clk, reset, DATAO_REG_26_, n1158 );
dff DATAO_REG_16__reg ( clk, reset, DATAO_REG_16_, n1118 );
dff REG2_REG_15__reg ( clk, reset, REG2_REG_15_, n889 );
not U_inv120 ( n5037, REG2_REG_15_ );
dff REG1_REG_15__reg ( clk, reset, REG1_REG_15_, n729 );
not U_inv121 ( n5040, REG1_REG_15_ );
dff REG0_REG_15__reg ( clk, reset, REG0_REG_15_, n569 );
dff DATAO_REG_15__reg ( clk, reset, DATAO_REG_15_, n1114 );
dff DATAO_REG_6__reg ( clk, reset, DATAO_REG_6_, n1078 );
dff DATAO_REG_5__reg ( clk, reset, DATAO_REG_5_, n1074 );
dff DATAO_REG_4__reg ( clk, reset, DATAO_REG_4_, n1070 );
dff REG2_REG_3__reg ( clk, reset, REG2_REG_3_, n829 );
not U_inv122 ( n4998, REG2_REG_3_ );
dff DATAO_REG_3__reg ( clk, reset, DATAO_REG_3_, n1066 );
dff DATAO_REG_2__reg ( clk, reset, DATAO_REG_2_, n1062 );
dff DATAO_REG_13__reg ( clk, reset, DATAO_REG_13_, n1106 );
dff ADDR_REG_13__reg ( clk, reset, ADDR_REG_13_, n998 );
dff ADDR_REG_14__reg ( clk, reset, ADDR_REG_14_, n994 );
dff ADDR_REG_16__reg ( clk, reset, ADDR_REG_16_, n986 );
dff ADDR_REG_17__reg ( clk, reset, ADDR_REG_17_, n982 );
dff ADDR_REG_1__reg ( clk, reset, ADDR_REG_1_, n1046 );
dff ADDR_REG_2__reg ( clk, reset, ADDR_REG_2_, n1042 );
dff ADDR_REG_3__reg ( clk, reset, ADDR_REG_3_, n1038 );
dff ADDR_REG_4__reg ( clk, reset, ADDR_REG_4_, n1034 );
dff ADDR_REG_5__reg ( clk, reset, ADDR_REG_5_, n1030 );
dff ADDR_REG_6__reg ( clk, reset, ADDR_REG_6_, n1026 );
dff ADDR_REG_9__reg ( clk, reset, ADDR_REG_9_, n1014 );
dff ADDR_REG_15__reg ( clk, reset, ADDR_REG_15_, n990 );
dff ADDR_REG_18__reg ( clk, reset, ADDR_REG_18_, n978 );
dff ADDR_REG_19__reg ( clk, reset, ADDR_REG_19_, n974 );
dff ADDR_REG_0__reg ( clk, reset, ADDR_REG_0_, n1050 );
dff ADDR_REG_7__reg ( clk, reset, ADDR_REG_7_, n1022 );
dff ADDR_REG_8__reg ( clk, reset, ADDR_REG_8_, n1018 );
dff ADDR_REG_10__reg ( clk, reset, ADDR_REG_10_, n1010 );
dff ADDR_REG_11__reg ( clk, reset, ADDR_REG_11_, n1006 );
dff ADDR_REG_12__reg ( clk, reset, ADDR_REG_12_, n1002 );
dff RD_REG_reg ( clk, reset, RD_REG, n1337 );
dff WR_REG_reg ( clk, reset, WR_REG, n5142 );
dff IR_REG_31__reg ( clk, reset, IR_REG_31_, n329 );
xnor U4968 ( n1523, n1507, n328 );
buf U4969 ( n5233, n67 );
buf U4970 ( n5174, n5096 );
buf U4971 ( n5158, n5159 );
buf U4972 ( n5204, n5105 );
nor U4973 ( n1944, n105, n2402 );
buf U4974 ( n5206, n785 );
buf U4975 ( n5141, n5143 );
buf U4976 ( n5193, n5107 );
buf U4977 ( n5192, n5107 );
buf U4978 ( n5184, n5106 );
buf U4979 ( n5200, n5198 );
buf U4980 ( n5176, n2845 );
buf U4981 ( n5188, n5109 );
nor U4982 ( n1565, n3818, n122 );
nor U4983 ( n1554, n3817, n143 );
buf U4984 ( n5171, n3035 );
buf U4985 ( n5165, n5164 );
buf U4986 ( n5166, n5164 );
buf U4987 ( n5198, n1376 );
buf U4988 ( n5197, n5111 );
buf U4989 ( n5196, n5111 );
and U4990 ( n5089, n4667, n4668 );
buf U4991 ( n5147, n4313 );
or U4992 ( n4314, n4676, n332 );
buf U4993 ( n5136, n4328 );
buf U4994 ( n5151, n4310 );
buf U4995 ( n5210, n5212 );
nor U4996 ( n2615, n1266, n300 );
nor U4997 ( n3928, n312, n1047 );
buf U4998 ( n5164, n3050 );
buf U4999 ( n5247, n5248 );
buf U5000 ( n5235, n66 );
buf U5001 ( n5236, n66 );
buf U5002 ( n5237, n66 );
buf U5003 ( n5241, n64 );
buf U5004 ( n5242, n64 );
buf U5005 ( n5243, n64 );
and U5006 ( n4047, n4094, n2450 );
not U5007 ( n125, n1901 );
not U5008 ( n41, n2494 );
buf U5009 ( n5230, n5233 );
not U5010 ( n66, n741 );
not U5011 ( n64, n770 );
nand U5012 ( n1151, n5242, n1152 );
buf U5013 ( n5231, n5233 );
buf U5014 ( n5228, n5234 );
buf U5015 ( n5232, n5233 );
buf U5016 ( n5229, n5234 );
not U5017 ( n95, n2142 );
not U5018 ( n5173, n5174 );
not U5019 ( n5172, n5174 );
not U5020 ( n103, n2441 );
not U5021 ( n5155, n5097 );
not U5022 ( n3, n3260 );
not U5023 ( n5157, n5159 );
not U5024 ( n5, n3282 );
not U5025 ( n69, n3452 );
buf U5026 ( n5116, n5158 );
buf U5027 ( n5115, n5158 );
not U5028 ( n82, n3253 );
and U5029 ( n1791, n1840, n125 );
nor U5030 ( n1840, n255, n47 );
not U5031 ( n43, n1586 );
not U5032 ( n49, n2014 );
nor U5033 ( n1690, n1645, n1691 );
nor U5034 ( n2000, n273, n2003 );
not U5035 ( n45, n1579 );
not U5036 ( n46, n1572 );
nor U5037 ( n2450, n201, n193 );
nand U5038 ( n1752, n1753, n1754 );
nand U5039 ( n1753, n1755, n108 );
nand U5040 ( n1754, n1755, n105 );
nor U5041 ( n1755, n1756, n1757 );
nand U5042 ( n1616, n98, n1579 );
nor U5043 ( n1539, n1550, n1551 );
nor U5044 ( n1550, n1552, n1555 );
nor U5045 ( n1551, n1552, n1553 );
nand U5046 ( n1555, n108, n230 );
not U5047 ( n79, n3188 );
nor U5048 ( n1697, n1698, n1699 );
and U5049 ( n1698, n1702, n108 );
nand U5050 ( n1699, n1700, n1701 );
nand U5051 ( n1700, n105, n1702 );
not U5052 ( n42, n1799 );
nand U5053 ( n938, n2061, n2062 );
nor U5054 ( n2062, n2063, n2064 );
nor U5055 ( n2061, n2080, n2081 );
nor U5056 ( n2063, n2076, n2077 );
nor U5057 ( n2059, n140, n2079 );
nand U5058 ( n2078, n2059, n272 );
nand U5059 ( n1832, n24, n105 );
nor U5060 ( n1772, n1774, n1775 );
nor U5061 ( n1774, n1776, n1639 );
nor U5062 ( n1775, n111, n1648 );
nand U5063 ( n1831, n24, n108 );
and U5064 ( n1544, n1545, n26 );
nand U5065 ( n1694, n98, n1696 );
xor U5066 ( n792, n233, n25 );
nor U5067 ( n2064, n272, n2065 );
nor U5068 ( n2065, n2066, n2067 );
nand U5069 ( n2067, n2068, n2069 );
nand U5070 ( n2066, n2071, n2003 );
and U5071 ( n2073, n2179, n2180 );
nand U5072 ( n2179, n20, n108 );
nand U5073 ( n2180, n20, n105 );
nor U5074 ( n1972, n273, n1976 );
nor U5075 ( n1879, n47, n95 );
nor U5076 ( n1876, n1877, n1878 );
nor U5077 ( n1877, n97, n1794 );
and U5078 ( n1878, n125, n1879 );
nor U5079 ( n1898, n1899, n1900 );
nor U5080 ( n1899, n125, n97 );
nand U5081 ( n2094, n135, n2095 );
not U5082 ( n195, n2477 );
nor U5083 ( n1908, n47, n1901 );
or U5084 ( n2076, n2079, n140 );
nor U5085 ( n2164, n2073, n124 );
not U5086 ( n208, n2364 );
nand U5087 ( n4037, n4003, n4083 );
not U5088 ( n129, n4074 );
nor U5089 ( n2280, n51, n95 );
buf U5090 ( n5114, n5158 );
nor U5091 ( n4094, n4037, n4056 );
nor U5092 ( n1915, n1919, n261 );
nand U5093 ( n1901, n1921, n1915 );
nor U5094 ( n2321, n103, n19 );
nand U5095 ( n2319, n51, n2142 );
xor U5096 ( n1085, n218, n18 );
nand U5097 ( n2494, n2501, n2142 );
and U5098 ( n2548, n2441, n1196 );
and U5099 ( n2466, n2321, n2461 );
not U5100 ( n148, n2030 );
xor U5101 ( n1152, n19, n2461 );
not U5102 ( n266, n1919 );
nor U5103 ( n2617, n103, n2600 );
buf U5104 ( n5239, n65 );
buf U5105 ( n5238, n65 );
nand U5106 ( n2408, n40, n2142 );
nand U5107 ( n741, n5185, n5230 );
and U5108 ( n2587, n2441, n1219 );
buf U5109 ( n5240, n65 );
nand U5110 ( n770, n101, n5230 );
nand U5111 ( n1195, n1196, n5241 );
nand U5112 ( n1060, n5242, n1061 );
not U5113 ( n14, n2600 );
nor U5114 ( n2531, n2522, n2494 );
not U5115 ( n132, n1787 );
nor U5116 ( n2520, n2501, n2521 );
nand U5117 ( n2521, n2522, n2142 );
not U5118 ( n131, n1794 );
nor U5119 ( n2553, n2549, n2392 );
nor U5120 ( n2686, n103, n2675 );
not U5121 ( n38, n2653 );
not U5122 ( n39, n2586 );
nand U5123 ( n3930, n2522, n2461 );
not U5124 ( n13, n2675 );
nand U5125 ( n3919, n2775, n160 );
nand U5126 ( n3927, n218, n156 );
not U5127 ( n5202, n5204 );
not U5128 ( n5203, n5204 );
nor U5129 ( n3898, n3899, n3900 );
nand U5130 ( n3899, n256, n250 );
nand U5131 ( n3900, n268, n262 );
nand U5132 ( n3929, n213, n207 );
nor U5133 ( n2680, n2681, n2653 );
nor U5134 ( n2605, n2606, n2586 );
and U5135 ( n2712, n2441, n1298 );
nor U5136 ( n2779, n110, n2764 );
nand U5137 ( n1348, n2766, n2767 );
nor U5138 ( n2767, n2768, n2769 );
nor U5139 ( n2766, n2779, n2780 );
nor U5140 ( n2768, n2775, n2776 );
nor U5141 ( n2772, n104, n12 );
nand U5142 ( n2607, n2606, n2142 );
nand U5143 ( n2682, n2681, n2142 );
not U5144 ( n11, n2764 );
nand U5145 ( n2152, n133, n2142 );
buf U5146 ( n5234, n67 );
not U5147 ( n5140, n5141 );
buf U5148 ( n5226, n90 );
buf U5149 ( n5225, n90 );
buf U5150 ( n5227, n90 );
buf U5151 ( n5207, n5206 );
buf U5152 ( n5208, n5206 );
not U5153 ( n5191, n5192 );
not U5154 ( n5190, n5192 );
buf U5155 ( n5209, n5206 );
nand U5156 ( n2142, n96, n111 );
buf U5157 ( n5179, n5176 );
not U5158 ( n5183, n5184 );
not U5159 ( n5182, n5184 );
not U5160 ( n5180, n5108 );
buf U5161 ( n5119, n5193 );
buf U5162 ( n5220, n107 );
buf U5163 ( n5221, n107 );
buf U5164 ( n5118, n5193 );
buf U5165 ( n5117, n5193 );
buf U5166 ( n5222, n107 );
nand U5167 ( n2441, n104, n110 );
not U5168 ( n104, n2075 );
nor U5169 ( n2811, n5223, n5185 );
buf U5170 ( n5175, n5096 );
buf U5171 ( n5178, n5176 );
buf U5172 ( n5177, n5176 );
not U5173 ( n97, n1820 );
not U5174 ( n2, n3578 );
nand U5175 ( n3214, n3701, n3040 );
nor U5176 ( n3701, n3702, n3703 );
nor U5177 ( n3703, n3704, n3042 );
nor U5178 ( n3702, n3705, n3038 );
nand U5179 ( n3478, n3589, n3590 );
nand U5180 ( n3589, n3623, n3624 );
nand U5181 ( n3590, n3591, n82 );
nand U5182 ( n3623, n3625, n3255 );
nand U5183 ( n3387, n3731, n3732 );
nand U5184 ( n3732, n78, n3138 );
nor U5185 ( n3731, n3733, n3734 );
nor U5186 ( n3734, n88, n3735 );
nand U5187 ( n3136, n3510, n3132 );
nand U5188 ( n3358, n3322, n3324 );
nor U5189 ( n3192, n2, n3193 );
nor U5190 ( n3193, n80, n3190 );
nor U5191 ( n3591, n3153, n3436 );
nand U5192 ( n3084, n3680, n3681 );
nand U5193 ( n3680, n3767, n3768 );
nand U5194 ( n3681, n3682, n69 );
nand U5195 ( n3767, n3769, n3454 );
and U5196 ( n3067, n3181, n3182 );
nand U5197 ( n3182, n3183, n3184 );
nand U5198 ( n3181, n3192, n79 );
nand U5199 ( n3183, n3185, n3186 );
and U5200 ( n3682, n3463, n3462 );
nor U5201 ( n3560, n3188, n3561 );
nand U5202 ( n3561, n3186, n3562 );
nand U5203 ( n3562, n1, n3191 );
not U5204 ( n1, n3302 );
xor U5205 ( n3065, n3066, n3067 );
nand U5206 ( n3296, n3301, n3302 );
nand U5207 ( n3301, n3191, n3303 );
nor U5208 ( n3735, n78, n3138 );
not U5209 ( n78, n3133 );
xor U5210 ( n3372, n2, n3190 );
xnor U5211 ( n3097, n3098, n3099 );
nand U5212 ( n3260, n3434, n3435 );
or U5213 ( n3435, n3436, n3153 );
nor U5214 ( n3252, n3253, n3254 );
nand U5215 ( n3254, n3255, n3256 );
nand U5216 ( n3256, n3, n81 );
xnor U5217 ( n3477, n3478, n3479 );
nand U5218 ( n3428, n3433, n3260 );
nand U5219 ( n3433, n81, n3261 );
nand U5220 ( n3038, n72, n3046 );
not U5221 ( n72, n3704 );
nor U5222 ( n3353, n3354, n3355 );
nand U5223 ( n3355, n3356, n3324 );
nand U5224 ( n3356, n4, n3323 );
not U5225 ( n4, n3322 );
and U5226 ( n3352, n3354, n5090 );
and U5227 ( n5090, n3358, n3323 );
buf U5228 ( n5156, n5097 );
not U5229 ( n121, n2823 );
nand U5230 ( n3316, n3321, n3322 );
nand U5231 ( n3321, n3323, n3324 );
not U5232 ( n5186, n5188 );
nand U5233 ( n3452, n3768, n3283 );
nor U5234 ( n3769, n3459, n3771 );
nor U5235 ( n3771, n3452, n3460 );
nor U5236 ( n4657, n292, n5157 );
not U5237 ( n5187, n5188 );
nand U5238 ( n3282, n3460, n3461 );
nand U5239 ( n3461, n3462, n3463 );
nor U5240 ( n3451, n3452, n3453 );
nand U5241 ( n3453, n3454, n3455 );
nand U5242 ( n3455, n5, n75 );
nand U5243 ( n3276, n3281, n3282 );
nand U5244 ( n3281, n75, n3283 );
not U5245 ( n83, n3323 );
nand U5246 ( n4236, n4231, n2649 );
nand U5247 ( n3253, n3261, n3624 );
nor U5248 ( n3625, n3437, n3626 );
nor U5249 ( n3626, n3253, n3434 );
nor U5250 ( n3037, n3038, n3039 );
nand U5251 ( n3039, n3040, n3041 );
nand U5252 ( n3041, n6, n3042 );
not U5253 ( n6, n3047 );
nand U5254 ( n3538, n3543, n3047 );
nand U5255 ( n3543, n3042, n3046 );
and U5256 ( n4182, n2366, n2414 );
not U5257 ( n47, n2098 );
nor U5258 ( n1645, n1717, n242 );
nor U5259 ( n1691, n1692, n1715 );
and U5260 ( n1715, n1716, n1673 );
or U5261 ( n1716, n248, n1645 );
nor U5262 ( n1822, n1791, n260 );
not U5263 ( n50, n2327 );
nand U5264 ( n818, n1684, n1685 );
nor U5265 ( n1685, n1686, n1687 );
nor U5266 ( n1684, n1703, n1704 );
nor U5267 ( n1686, n1697, n1673 );
nand U5268 ( n1704, n1705, n1706 );
nand U5269 ( n1705, n1730, n1692 );
nand U5270 ( n1706, n1707, n1673 );
nor U5271 ( n1730, n1731, n111 );
nand U5272 ( n1799, n1822, n1837 );
nand U5273 ( n1837, n1838, n1797 );
nand U5274 ( n1707, n1708, n1709 );
nor U5275 ( n1708, n1723, n1724 );
nor U5276 ( n1709, n1710, n1711 );
nor U5277 ( n1723, n1620, n1702 );
nand U5278 ( n1586, n1636, n1644 );
nand U5279 ( n1644, n1645, n1646 );
nor U5280 ( n1611, n233, n1612 );
nor U5281 ( n1612, n1613, n1614 );
nand U5282 ( n1614, n1615, n1616 );
nand U5283 ( n1613, n1621, n1622 );
nor U5284 ( n1628, n1630, n1631 );
nand U5285 ( n1631, n1632, n1633 );
nand U5286 ( n1630, n1640, n1641 );
nand U5287 ( n1633, n98, n45 );
nor U5288 ( n1581, n1584, n1585 );
nor U5289 ( n1585, n1571, n1586 );
nor U5290 ( n1584, n43, n1573 );
nand U5291 ( n1561, n1574, n1575 );
nand U5292 ( n1575, n98, n1538 );
nand U5293 ( n1574, n112, n1580 );
nand U5294 ( n1580, n1581, n1568 );
not U5295 ( n183, n2649 );
nor U5296 ( n1976, n1916, n49 );
nand U5297 ( n2014, n1921, n2098 );
nor U5298 ( n2004, n1952, n111 );
nand U5299 ( n898, n1932, n1933 );
nor U5300 ( n1932, n1966, n1967 );
nor U5301 ( n1933, n1934, n1935 );
nor U5302 ( n1966, n320, n5127 );
nand U5303 ( n1935, n1936, n1937 );
nand U5304 ( n1936, n1949, n1950 );
nand U5305 ( n1937, n1938, n1930 );
nor U5306 ( n1949, n111, n1930 );
nand U5307 ( n1687, n1688, n1689 );
nand U5308 ( n1688, n1692, n1693 );
nand U5309 ( n1689, n1690, n112 );
nand U5310 ( n1693, n1694, n1695 );
not U5311 ( n168, n2683 );
nand U5312 ( n2003, n1820, n2070 );
nand U5313 ( n1639, n1790, n1783 );
nand U5314 ( n1790, n1784, n1793 );
nand U5315 ( n1793, n1786, n1794 );
nand U5316 ( n1783, n1791, n1792 );
nand U5317 ( n1579, n1636, n1637 );
nand U5318 ( n1637, n1638, n1639 );
not U5319 ( n167, n3985 );
nand U5320 ( n3188, n3303, n3184 );
nor U5321 ( n3185, n84, n3187 );
not U5322 ( n84, n3191 );
nor U5323 ( n3187, n3188, n3189 );
nand U5324 ( n3189, n80, n3190 );
nand U5325 ( n1648, n1782, n1783 );
nand U5326 ( n1782, n1784, n1785 );
nand U5327 ( n1785, n1786, n1787 );
nand U5328 ( n1572, n1636, n1647 );
nand U5329 ( n1647, n1638, n1648 );
nand U5330 ( n1538, n1576, n1568 );
nor U5331 ( n1576, n1577, n1578 );
nor U5332 ( n1578, n1579, n1571 );
nor U5333 ( n1577, n45, n1573 );
nand U5334 ( n2284, n205, n2302 );
nand U5335 ( n2302, n2303, n2304 );
or U5336 ( n1724, n5091, n5092 );
nor U5337 ( n5091, n1702, n1549 );
nor U5338 ( n5092, n1702, n110 );
nand U5339 ( n1702, n1663, n1727 );
nand U5340 ( n1727, n1659, n1728 );
nand U5341 ( n2664, n2665, n2666 );
not U5342 ( n193, n2495 );
nor U5343 ( n3129, n71, n3130 );
not U5344 ( n71, n3134 );
nand U5345 ( n3130, n3131, n3132 );
nand U5346 ( n3131, n7, n3133 );
not U5347 ( n7, n3510 );
nor U5348 ( n1567, n1569, n1570 );
nor U5349 ( n1570, n1571, n1572 );
nor U5350 ( n1569, n46, n1573 );
not U5351 ( n172, n2582 );
not U5352 ( n201, n4066 );
nor U5353 ( n1965, n1906, n2013 );
nor U5354 ( n2013, n2014, n273 );
not U5355 ( n24, n1728 );
nor U5356 ( n1756, n1760, n1761 );
nor U5357 ( n1760, n253, n24 );
nand U5358 ( n838, n1749, n1750 );
nor U5359 ( n1749, n1767, n1768 );
nor U5360 ( n1750, n1751, n1752 );
nor U5361 ( n1767, n323, n5128 );
not U5362 ( n26, n1546 );
nor U5363 ( n1640, n1652, n1653 );
nor U5364 ( n1652, n26, n110 );
nor U5365 ( n1653, n26, n1549 );
nand U5366 ( n1696, n1639, n1649 );
nor U5367 ( n3128, n3134, n3135 );
nand U5368 ( n3135, n3136, n3133 );
not U5369 ( n197, n2533 );
nand U5370 ( n1714, n1780, n1781 );
nand U5371 ( n1781, n1565, n1648 );
nand U5372 ( n1780, n99, n1639 );
nor U5373 ( n2410, n191, n2535 );
nor U5374 ( n1995, n268, n1996 );
nor U5375 ( n1996, n1997, n1947 );
nor U5376 ( n1997, n1944, n1958 );
nand U5377 ( n1552, n1558, n1559 );
nand U5378 ( n1559, n1547, n1546 );
nand U5379 ( n1558, n26, n1545 );
nand U5380 ( n1701, n1554, n1702 );
nand U5381 ( n858, n1813, n1814 );
nor U5382 ( n1813, n1841, n1842 );
nor U5383 ( n1814, n1815, n1816 );
nor U5384 ( n1842, n322, n5129 );
nor U5385 ( n1815, n250, n1828 );
nor U5386 ( n1828, n1829, n1830 );
nand U5387 ( n1830, n1831, n1832 );
nand U5388 ( n1829, n1833, n1834 );
nand U5389 ( n1768, n1769, n1770 );
nand U5390 ( n1770, n245, n1771 );
nand U5391 ( n1769, n1778, n1777 );
nand U5392 ( n1771, n1772, n1773 );
nand U5393 ( n1778, n1779, n44 );
not U5394 ( n44, n1714 );
nor U5395 ( n1779, n1788, n1789 );
and U5396 ( n1789, n1639, n98 );
not U5397 ( n20, n2058 );
nor U5398 ( n2079, n20, n2029 );
nor U5399 ( n2080, n2082, n2054 );
nor U5400 ( n2082, n2083, n2084 );
nand U5401 ( n2083, n2093, n2094 );
nand U5402 ( n2084, n2085, n2086 );
nor U5403 ( n2085, n2087, n2088 );
nor U5404 ( n2087, n104, n2057 );
and U5405 ( n2088, n2078, n1554 );
nor U5406 ( n1621, n1626, n1627 );
nor U5407 ( n1626, n1546, n110 );
nor U5408 ( n1627, n1546, n1549 );
and U5409 ( n1827, n1822, n1839 );
nand U5410 ( n1839, n132, n1797 );
nand U5411 ( n1773, n1717, n112 );
nor U5412 ( n1950, n271, n1951 );
nor U5413 ( n1951, n267, n1952 );
nand U5414 ( n1834, n24, n1554 );
nor U5415 ( n1757, n1758, n1759 );
nor U5416 ( n1758, n251, n1728 );
nor U5417 ( n1841, n1810, n1843 );
nor U5418 ( n1843, n1844, n1845 );
nand U5419 ( n1845, n1846, n1847 );
nor U5420 ( n1844, n24, n1620 );
nand U5421 ( n1540, n1541, n1542 );
nor U5422 ( n1541, n1548, n1549 );
nor U5423 ( n1542, n1543, n1544 );
and U5424 ( n1543, n1546, n1547 );
not U5425 ( n25, n1526 );
nor U5426 ( n1751, n110, n1762 );
nand U5427 ( n1762, n1746, n1747 );
or U5428 ( n1746, n1759, n5093 );
and U5429 ( n5093, n24, n1681 );
nor U5430 ( n2006, n2007, n2008 );
nand U5431 ( n2007, n2016, n2017 );
nand U5432 ( n2008, n2009, n2010 );
nor U5433 ( n2016, n2019, n2020 );
nand U5434 ( n2010, n1952, n1565 );
nand U5435 ( n1695, n99, n1696 );
and U5436 ( n1731, n1648, n1649 );
nand U5437 ( n1816, n1817, n1818 );
nand U5438 ( n1818, n1819, n1820 );
nand U5439 ( n1817, n250, n1824 );
xor U5440 ( n1819, n1821, n250 );
nand U5441 ( n1824, n1825, n1826 );
nand U5442 ( n1826, n1827, n1565 );
nand U5443 ( n1825, n42, n112 );
nand U5444 ( n3507, n3513, n3510 );
nand U5445 ( n3513, n3133, n3132 );
nand U5446 ( n1847, n1554, n1728 );
nand U5447 ( n1846, n105, n1728 );
nor U5448 ( n1867, n256, n1868 );
nor U5449 ( n1868, n1869, n1870 );
nand U5450 ( n1869, n1875, n1876 );
nand U5451 ( n1870, n1871, n1872 );
nand U5452 ( n878, n1864, n1865 );
nor U5453 ( n1864, n1893, n1894 );
nor U5454 ( n1865, n1866, n1867 );
nor U5455 ( n1894, n321, n5128 );
and U5456 ( n827, n1746, n1747 );
nor U5457 ( n2093, n2018, n2096 );
nor U5458 ( n2096, n1916, n2097 );
nand U5459 ( n2097, n112, n2014 );
and U5460 ( n2018, n1976, n1820 );
nand U5461 ( n1934, n1953, n1954 );
nand U5462 ( n1954, n1955, n262 );
nand U5463 ( n1953, n1961, n1904 );
nor U5464 ( n1955, n22, n1944 );
nor U5465 ( n1961, n261, n1962 );
nor U5466 ( n1962, n1963, n1964 );
nor U5467 ( n1963, n96, n1907 );
and U5468 ( n1964, n112, n1965 );
nor U5469 ( n761, n768, n770 );
nand U5470 ( n2071, n2072, n2057 );
nand U5471 ( n2072, n2073, n2074 );
nand U5472 ( n2074, n2075, n2029 );
nand U5473 ( n847, n1808, n1809 );
nand U5474 ( n1808, n24, n1811 );
or U5475 ( n1809, n1810, n24 );
not U5476 ( n75, n3459 );
nand U5477 ( n1821, n1822, n1823 );
nand U5478 ( n1823, n131, n1797 );
not U5479 ( n81, n3437 );
nand U5480 ( n2068, n1565, n2070 );
nand U5481 ( n1967, n1968, n1969 );
nand U5482 ( n1968, n1973, n1971 );
nand U5483 ( n1969, n1970, n1971 );
and U5484 ( n1971, n1974, n1904 );
nor U5485 ( n1973, n1972, n1975 );
nand U5486 ( n1872, n23, n108 );
nand U5487 ( n2077, n1554, n2078 );
nand U5488 ( n2009, n1965, n112 );
nand U5489 ( n2086, n1976, n1565 );
nor U5490 ( n2124, n2128, n2129 );
nor U5491 ( n2128, n136, n20 );
not U5492 ( n136, n2130 );
nand U5493 ( n2120, n2121, n2122 );
nand U5494 ( n2121, n2123, n108 );
nand U5495 ( n2122, n2123, n105 );
nor U5496 ( n2123, n2124, n2125 );
nand U5497 ( n958, n2117, n2118 );
nor U5498 ( n2117, n2135, n2136 );
nor U5499 ( n2118, n2119, n2120 );
nor U5500 ( n2135, n316, n5135 );
nor U5501 ( n1885, n23, n1620 );
xor U5502 ( n810, n1673, n1606 );
nand U5503 ( n2069, n112, n2070 );
or U5504 ( n2070, n1916, n49 );
nor U5505 ( n2242, n155, n153 );
nor U5506 ( n930, n2052, n2053 );
and U5507 ( n2053, n2054, n2055 );
and U5508 ( n2052, n2059, n272 );
nand U5509 ( n2055, n2056, n2057 );
nor U5510 ( n1900, n2098, n97 );
nor U5511 ( n1893, n1895, n1862 );
nor U5512 ( n1895, n1896, n1897 );
nor U5513 ( n1896, n1908, n1909 );
nor U5514 ( n1897, n131, n1898 );
nand U5515 ( n2364, n2359, n2398 );
nand U5516 ( n2136, n2137, n2138 );
nand U5517 ( n2137, n2149, n2150 );
nand U5518 ( n2138, n280, n2139 );
nand U5519 ( n2149, n2151, n2152 );
nand U5520 ( n2139, n2140, n2141 );
nand U5521 ( n2141, n126, n2142 );
nor U5522 ( n2140, n2144, n2145 );
nor U5523 ( n2144, n2098, n2147 );
and U5524 ( n2145, n2146, n1900 );
nand U5525 ( n2095, n2183, n2184 );
nand U5526 ( n2183, n108, n2058 );
nand U5527 ( n2184, n105, n2058 );
nand U5528 ( n2477, n2472, n2526 );
not U5529 ( n173, n2491 );
nor U5530 ( n2119, n110, n2131 );
nand U5531 ( n2131, n2114, n2115 );
nand U5532 ( n967, n2168, n2169 );
nand U5533 ( n2169, n2170, n2058 );
nand U5534 ( n2168, n20, n2171 );
nand U5535 ( n980, n2162, n2163 );
nor U5536 ( n2162, n2181, n2182 );
nor U5537 ( n2163, n2164, n2165 );
nor U5538 ( n2182, n315, n5135 );
nand U5539 ( n2165, n2166, n2167 );
nand U5540 ( n2166, n2172, n2173 );
nand U5541 ( n2167, n1554, n967 );
nand U5542 ( n2173, n1776, n2174 );
nand U5543 ( n1428, n2155, n2156 );
nor U5544 ( n2156, n2157, n2158 );
nor U5545 ( n2155, n2161, n980 );
nor U5546 ( n2157, n317, n5199 );
nand U5547 ( n975, n976, n977 );
nand U5548 ( n977, n5239, n979 );
nand U5549 ( n976, n5231, n980 );
nor U5550 ( n2020, n21, n1944 );
not U5551 ( n21, n1958 );
or U5552 ( n2115, n2129, n5094 );
and U5553 ( n5094, n2058, n2130 );
nand U5554 ( n2107, n2108, n2109 );
nand U5555 ( n2109, n951, n5223 );
nand U5556 ( n2108, n5218, n947 );
and U5557 ( n947, n2114, n2115 );
nor U5558 ( n737, n742, n743 );
nor U5559 ( n4045, n4053, n4054 );
nor U5560 ( n4054, n248, n1792 );
nor U5561 ( n4053, n4055, n4056 );
nor U5562 ( n4055, n4057, n4058 );
not U5563 ( n9, n3879 );
not U5564 ( n188, n4051 );
nand U5565 ( n4058, n4059, n1915 );
nor U5566 ( n4059, n4060, n4061 );
nor U5567 ( n4061, n276, n2101 );
nor U5568 ( n4060, n4062, n4037 );
nand U5569 ( n4024, n4025, n4026 );
nand U5570 ( n4026, n4027, n4028 );
nand U5571 ( n4025, n4040, n226 );
nor U5572 ( n4028, n4029, n4030 );
nand U5573 ( n2056, n135, n2058 );
nor U5574 ( n4040, n237, n4042 );
nor U5575 ( n4042, n4043, n4044 );
nand U5576 ( n4043, n4084, n4085 );
nand U5577 ( n4044, n4045, n4046 );
nand U5578 ( n2158, n2159, n2160 );
nand U5579 ( n2160, n5224, n979 );
nand U5580 ( n2159, n5218, n967 );
and U5581 ( n2181, n2095, n2170 );
xor U5582 ( n2172, n2098, n124 );
not U5583 ( n19, n2304 );
not U5584 ( n17, n2401 );
nand U5585 ( n1116, n2385, n2386 );
nor U5586 ( n2385, n2403, n2404 );
nor U5587 ( n2386, n2387, n2388 );
nor U5588 ( n2404, n307, n5131 );
nor U5589 ( n2387, n1944, n2394 );
nand U5590 ( n2394, n2382, n2383 );
nand U5591 ( n2383, n2395, n207 );
nor U5592 ( n2395, n2362, n2396 );
nor U5593 ( n2396, n215, n17 );
nand U5594 ( n1446, n2376, n2377 );
nor U5595 ( n2377, n2378, n2379 );
nor U5596 ( n2376, n2384, n1116 );
nor U5597 ( n2378, n310, n5200 );
nand U5598 ( n1111, n1112, n1113 );
nand U5599 ( n1113, n5239, n1115 );
nand U5600 ( n1112, n5231, n1116 );
nand U5601 ( n1003, n2203, n2204 );
nor U5602 ( n2204, n2205, n2206 );
nor U5603 ( n2203, n2209, n2210 );
nor U5604 ( n2206, n2178, n2207 );
nor U5605 ( n2209, n2201, n2211 );
nor U5606 ( n2211, n2212, n2213 );
and U5607 ( n2213, n2142, n2178 );
nor U5608 ( n2212, n1944, n2186 );
nand U5609 ( n1431, n2189, n2190 );
nor U5610 ( n2190, n2191, n2192 );
nor U5611 ( n2189, n2202, n1003 );
nor U5612 ( n2191, n316, n5199 );
nand U5613 ( n3932, n3933, n3934 );
nand U5614 ( n3934, n99, n3889 );
nand U5615 ( n3933, n9, n101 );
nand U5616 ( n4074, n2175, n2146 );
nor U5617 ( n4083, n4112, n4080 );
nand U5618 ( n4112, n2247, n2325 );
nand U5619 ( n4057, n4067, n4068 );
nor U5620 ( n4067, n4077, n4078 );
nor U5621 ( n4068, n255, n4069 );
nor U5622 ( n4078, n4079, n4080 );
nand U5623 ( n4073, n4075, n153 );
and U5624 ( n4075, n2214, n129 );
not U5625 ( n130, n4014 );
nor U5626 ( n2346, n2352, n2353 );
nor U5627 ( n2352, n2354, n2355 );
nor U5628 ( n2354, n95, n2327 );
nor U5629 ( n2355, n103, n18 );
not U5630 ( n18, n2351 );
nand U5631 ( n1443, n2333, n2334 );
nor U5632 ( n2334, n2335, n2336 );
nor U5633 ( n2333, n2343, n1093 );
nor U5634 ( n2335, n311, n5200 );
nor U5635 ( n2278, n2279, n2280 );
nor U5636 ( n2279, n95, n2247 );
not U5637 ( n51, n2291 );
nand U5638 ( n1437, n2257, n2258 );
nor U5639 ( n2258, n2259, n2260 );
nor U5640 ( n2257, n2270, n1048 );
nor U5641 ( n2259, n313, n5200 );
nand U5642 ( n1048, n2271, n2272 );
nor U5643 ( n2271, n2286, n2287 );
nor U5644 ( n2272, n2273, n2274 );
nor U5645 ( n2287, n311, n5132 );
nand U5646 ( n2379, n2380, n2381 );
nand U5647 ( n2381, n5224, n1115 );
nand U5648 ( n2380, n5218, n1103 );
and U5649 ( n1103, n2382, n2383 );
nor U5650 ( n2205, n1944, n2200 );
not U5651 ( n178, n4033 );
nor U5652 ( n3983, n186, n3986 );
nor U5653 ( n3986, n3987, n178 );
nor U5654 ( n3987, n181, n2683 );
nor U5655 ( n3967, n3968, n3969 );
nand U5656 ( n3968, n3990, n3991 );
nand U5657 ( n3969, n3970, n1904 );
nor U5658 ( n3990, n4009, n4010 );
nand U5659 ( n3976, n3977, n3978 );
nor U5660 ( n3977, n193, n3988 );
nand U5661 ( n3978, n3979, n3980 );
and U5662 ( n3988, n188, n2410 );
or U5663 ( n3885, n3889, n1975 );
not U5664 ( n140, n2057 );
nor U5665 ( n2348, n2349, n2350 );
nor U5666 ( n2349, n95, n50 );
nor U5667 ( n2350, n103, n2351 );
nor U5668 ( n4084, n242, n4091 );
nor U5669 ( n4091, n4092, n4093 );
nand U5670 ( n4092, n4051, n2582 );
nand U5671 ( n4093, n4047, n181 );
nand U5672 ( n1434, n2224, n2225 );
nor U5673 ( n2225, n2226, n2227 );
nor U5674 ( n2224, n2232, n1025 );
nor U5675 ( n2226, n315, n5200 );
nor U5676 ( n2235, n1944, n2248 );
nand U5677 ( n2248, n2230, n2231 );
not U5678 ( n255, n1797 );
nand U5679 ( n4056, n4036, n4108 );
nand U5680 ( n4108, n4109, n271 );
nor U5681 ( n4109, n261, n255 );
nand U5682 ( n1020, n1021, n1023 );
nand U5683 ( n1023, n5239, n1024 );
nand U5684 ( n1021, n5231, n1025 );
nand U5685 ( n989, n2199, n2200 );
or U5686 ( n2199, n2186, n2201 );
not U5687 ( n133, n2146 );
xor U5688 ( n912, n1958, n1990 );
nor U5689 ( n2442, n213, n2444 );
nor U5690 ( n2444, n2445, n2446 );
nor U5691 ( n2445, n95, n2439 );
nor U5692 ( n2446, n103, n2401 );
nand U5693 ( n1139, n2434, n2435 );
nor U5694 ( n2435, n2436, n2437 );
nor U5695 ( n2434, n2442, n2443 );
nor U5696 ( n2437, n2432, n2438 );
nand U5697 ( n1449, n2419, n2420 );
nor U5698 ( n2420, n2421, n2422 );
nor U5699 ( n2419, n2433, n1139 );
nor U5700 ( n2421, n308, n5200 );
not U5701 ( n206, n2366 );
nor U5702 ( n4003, n206, n212 );
not U5703 ( n212, n2414 );
nand U5704 ( n1919, n2012, n1907 );
nand U5705 ( n4000, n4012, n4013 );
nor U5706 ( n4013, n278, n4014 );
nor U5707 ( n4012, n1919, n4015 );
nor U5708 ( n3991, n260, n3992 );
nor U5709 ( n3992, n3993, n3994 );
nand U5710 ( n3993, n4004, n167 );
nand U5711 ( n3994, n123, n3979 );
not U5712 ( n123, n3974 );
xor U5713 ( n2237, n2217, n2238 );
not U5714 ( n157, n2247 );
not U5715 ( n261, n1903 );
nand U5716 ( n1440, n2295, n2296 );
nor U5717 ( n2296, n2297, n2298 );
nor U5718 ( n2295, n2305, n1071 );
nor U5719 ( n2297, n312, n5200 );
nor U5720 ( n2308, n2316, n2301 );
nor U5721 ( n2316, n2317, n2318 );
nor U5722 ( n2317, n103, n205 );
nand U5723 ( n2318, n2319, n2320 );
nand U5724 ( n2320, n2321, n2303 );
nand U5725 ( n1065, n1067, n1068 );
nand U5726 ( n1068, n5239, n1069 );
nand U5727 ( n1067, n5231, n1071 );
nor U5728 ( n2273, n103, n2268 );
nand U5729 ( n2227, n2228, n2229 );
nand U5730 ( n2229, n5224, n1024 );
nand U5731 ( n2228, n5218, n1012 );
and U5732 ( n1012, n2230, n2231 );
nor U5733 ( n2315, n2304, n103 );
nand U5734 ( n2030, n2251, n2036 );
not U5735 ( n278, n2101 );
nor U5736 ( n1921, n126, n278 );
nand U5737 ( n1125, n2429, n2430 );
nand U5738 ( n2429, n17, n2432 );
or U5739 ( n2430, n2431, n17 );
nand U5740 ( n4001, n2242, n4002 );
nand U5741 ( n4002, n4003, n203 );
nand U5742 ( n985, n987, n988 );
nand U5743 ( n988, n5203, n476 );
nand U5744 ( n987, n5242, n989 );
nand U5745 ( n4046, n4047, n4048 );
nand U5746 ( n4048, n4049, n4050 );
nand U5747 ( n4050, n176, n4051 );
nor U5748 ( n4049, n2535, n4052 );
and U5749 ( n2519, n2514, n5095 );
and U5750 ( n5095, n2515, n2441 );
nand U5751 ( n1455, n2504, n2505 );
nor U5752 ( n2505, n2506, n2507 );
nor U5753 ( n2504, n2516, n1184 );
nor U5754 ( n2506, n306, n5200 );
nand U5755 ( n2515, n2524, n2522 );
nor U5756 ( n2524, n2475, n2525 );
and U5757 ( n2525, n2526, n2527 );
nand U5758 ( n1184, n2517, n2518 );
nor U5759 ( n2517, n2531, n2532 );
nor U5760 ( n2518, n2519, n2520 );
nor U5761 ( n2532, n303, n5126 );
and U5762 ( n4086, n4094, n4104 );
nor U5763 ( n4104, n178, n4039 );
nand U5764 ( n1794, n1902, n1903 );
nand U5765 ( n1902, n1904, n1905 );
nand U5766 ( n1905, n1906, n1907 );
nor U5767 ( n2436, n2431, n2440 );
nand U5768 ( n2440, n2401, n2441 );
nand U5769 ( n1838, n1912, n1913 );
nand U5770 ( n1913, n1914, n1903 );
nand U5771 ( n1912, n1915, n1916 );
nor U5772 ( n2465, n2461, n2467 );
nor U5773 ( n2467, n2468, n2315 );
nor U5774 ( n2468, n191, n2492 );
nor U5775 ( n2492, n2493, n41 );
nand U5776 ( n1452, n2455, n2456 );
nor U5777 ( n2456, n2457, n2458 );
nor U5778 ( n2455, n2462, n1161 );
nor U5779 ( n2457, n307, n5200 );
nand U5780 ( n1161, n2463, n2464 );
nor U5781 ( n2463, n2496, n2497 );
nor U5782 ( n2464, n2465, n2466 );
nor U5783 ( n2497, n305, n5127 );
nand U5784 ( n2501, n2533, n2534 );
or U5785 ( n2534, n2373, n2535 );
nand U5786 ( n950, n951, n5238 );
not U5787 ( n37, n2750 );
and U5788 ( n3979, n3995, n2410 );
nor U5789 ( n3995, n190, n176 );
nand U5790 ( n1156, n1157, n1159 );
nand U5791 ( n1159, n5239, n1160 );
nand U5792 ( n1157, n5231, n1161 );
nand U5793 ( n1121, n1123, n1124 );
nand U5794 ( n1124, n5202, n498 );
nand U5795 ( n1123, n5242, n1125 );
and U5796 ( n1171, n2514, n2515 );
nand U5797 ( n1914, n1904, n1920 );
nand U5798 ( n1920, n276, n1907 );
xor U5799 ( n1196, n2549, n2527 );
nand U5800 ( n1205, n2545, n2546 );
nor U5801 ( n2545, n2553, n2554 );
nor U5802 ( n2546, n2547, n2548 );
nor U5803 ( n2554, n302, n5134 );
nand U5804 ( n1458, n2538, n2539 );
nor U5805 ( n2539, n2540, n2541 );
nor U5806 ( n2538, n2544, n1205 );
nor U5807 ( n2540, n305, n5200 );
nand U5808 ( n1031, n1032, n1033 );
nand U5809 ( n1033, n5203, n473 );
nand U5810 ( n1032, n5242, n1035 );
nand U5811 ( n1200, n1201, n1203 );
nand U5812 ( n1203, n5239, n1204 );
nand U5813 ( n1201, n5231, n1205 );
nor U5814 ( n4009, n4011, n4000 );
nor U5815 ( n4011, n4016, n4017 );
nand U5816 ( n4016, n4019, n2214 );
nand U5817 ( n4017, n129, n2246 );
nand U5818 ( n1787, n1917, n1903 );
nand U5819 ( n1917, n265, n1918 );
not U5820 ( n265, n1914 );
nand U5821 ( n1918, n266, n1916 );
xor U5822 ( n1061, n2284, n2301 );
nand U5823 ( n2298, n2299, n2300 );
nand U5824 ( n2299, n5223, n1069 );
nand U5825 ( n2300, n5218, n1061 );
not U5826 ( n40, n2373 );
nand U5827 ( n1167, n1168, n1169 );
nand U5828 ( n1169, n5202, n496 );
nand U5829 ( n1168, n1171, n5241 );
nand U5830 ( n2458, n2459, n2460 );
nand U5831 ( n2459, n5223, n1160 );
nand U5832 ( n2460, n5217, n1152 );
nand U5833 ( n3975, n3989, n2414 );
nor U5834 ( n3989, n201, n206 );
not U5835 ( n165, n2747 );
nand U5836 ( n2541, n2542, n2543 );
nand U5837 ( n2542, n5224, n1204 );
nand U5838 ( n2543, n5217, n1196 );
nor U5839 ( n4027, n4034, n4035 );
nand U5840 ( n4035, n4036, n127 );
nand U5841 ( n4034, n171, n4038 );
not U5842 ( n127, n4037 );
not U5843 ( n171, n4039 );
nand U5844 ( n1246, n2602, n2603 );
nor U5845 ( n2603, n2604, n2605 );
nor U5846 ( n2602, n2617, n2618 );
nor U5847 ( n2604, n2580, n2607 );
nand U5848 ( n2600, n2619, n2620 );
nand U5849 ( n2619, n2624, n2483 );
nand U5850 ( n2620, n2621, n2606 );
nor U5851 ( n2624, n2625, n2626 );
nand U5852 ( n1464, n2594, n2595 );
nor U5853 ( n2595, n2596, n2597 );
nor U5854 ( n2594, n2601, n1246 );
nor U5855 ( n2596, n302, n5200 );
nand U5856 ( n1241, n1243, n1244 );
nand U5857 ( n1244, n5240, n1245 );
nand U5858 ( n1243, n5231, n1246 );
not U5859 ( n65, n742 );
not U5860 ( n67, n756 );
buf U5861 ( n5224, n102 );
nand U5862 ( n2438, n2142, n2439 );
nand U5863 ( n1283, n1284, n1285 );
nand U5864 ( n1284, n5231, n1288 );
nand U5865 ( n1285, n5239, n1286 );
nor U5866 ( n2403, n207, n2405 );
nor U5867 ( n2405, n2406, n2407 );
nor U5868 ( n2406, n95, n2370 );
nor U5869 ( n2407, n2372, n2408 );
xnor U5870 ( n1219, n2579, n2551 );
nand U5871 ( n1226, n2573, n2574 );
nor U5872 ( n2574, n2575, n2576 );
nor U5873 ( n2573, n2587, n2588 );
nor U5874 ( n2576, n2577, n2578 );
nand U5875 ( n1461, n2562, n2563 );
nor U5876 ( n2563, n2564, n2565 );
nor U5877 ( n2562, n2572, n1226 );
nor U5878 ( n2564, n303, n5200 );
nand U5879 ( n1326, n1328, n1329 );
nand U5880 ( n1328, n5232, n1331 );
nand U5881 ( n1329, n5240, n1330 );
nand U5882 ( n1361, n1362, n1363 );
nand U5883 ( n1362, n5230, n1365 );
nand U5884 ( n1363, n5240, n1364 );
nand U5885 ( n2597, n2598, n2599 );
nand U5886 ( n2599, n5224, n1245 );
nand U5887 ( n2598, n5217, n14 );
nand U5888 ( n1379, n1380, n1381 );
nand U5889 ( n1380, n1383, n5230 );
nand U5890 ( n1381, n5242, n1382 );
nand U5891 ( n1251, n1253, n1254 );
nand U5892 ( n1254, n5202, n502 );
nand U5893 ( n1253, n5242, n1255 );
nand U5894 ( n4090, n164, n2719 );
nand U5895 ( n2392, n2142, n2373 );
nor U5896 ( n2388, n2389, n2390 );
nand U5897 ( n2390, n2391, n2370 );
nand U5898 ( n2391, n2392, n2393 );
nand U5899 ( n2393, n2142, n2372 );
not U5900 ( n273, n2012 );
nor U5901 ( n4122, n4102, n4124 );
nor U5902 ( n4124, n4125, n232 );
nor U5903 ( n4125, n237, n1646 );
nand U5904 ( n1268, n2640, n2641 );
nor U5905 ( n2641, n2642, n2643 );
nor U5906 ( n2640, n2654, n2655 );
nor U5907 ( n2643, n2644, n2645 );
nand U5908 ( n1467, n2629, n2630 );
nor U5909 ( n2630, n2631, n2632 );
nor U5910 ( n2629, n2639, n1268 );
nor U5911 ( n2631, n301, n5200 );
and U5912 ( n2654, n2441, n1255 );
and U5913 ( n4038, n4096, n4097 );
nor U5914 ( n4097, n168, n4098 );
nor U5915 ( n4096, n237, n4041 );
nand U5916 ( n4098, n2747, n2719 );
nor U5917 ( n2547, n2552, n2408 );
nor U5918 ( n2552, n197, n2535 );
not U5919 ( n267, n1907 );
not U5920 ( n232, n1588 );
nand U5921 ( n1662, n1663, n1664 );
not U5922 ( n242, n1649 );
nand U5923 ( n1664, n1659, n257 );
not U5924 ( n257, n1682 );
nor U5925 ( n1875, n1880, n1881 );
and U5926 ( n1881, n1838, n112 );
nor U5927 ( n1880, n111, n1787 );
nor U5928 ( n2606, n172, n176 );
nand U5929 ( n3888, n3893, n3894 );
nor U5930 ( n3894, n3895, n3896 );
nor U5931 ( n3893, n3913, n3914 );
nand U5932 ( n3896, n3897, n3898 );
nand U5933 ( n3917, n2606, n2579 );
nand U5934 ( n3914, n3915, n3916 );
nor U5935 ( n3915, n3919, n3920 );
nor U5936 ( n3916, n3917, n3918 );
nand U5937 ( n3920, n10, n2805 );
nand U5938 ( n1288, n2677, n2678 );
nor U5939 ( n2678, n2679, n2680 );
nor U5940 ( n2677, n2686, n2687 );
nor U5941 ( n2679, n2648, n2682 );
nand U5942 ( n2675, n2688, n2689 );
nand U5943 ( n2688, n2692, n2693 );
nand U5944 ( n2689, n2690, n2681 );
and U5945 ( n2693, n2662, n2665 );
nand U5946 ( n1470, n2669, n2670 );
nor U5947 ( n2670, n2671, n2672 );
nor U5948 ( n2669, n2676, n1288 );
nor U5949 ( n2671, n300, n5201 );
nor U5950 ( n2690, n170, n2691 );
and U5951 ( n2691, n2666, n2665 );
nand U5952 ( n2653, n2648, n2142 );
nand U5953 ( n2586, n2580, n2142 );
nor U5954 ( n2575, n2583, n2584 );
or U5955 ( n2584, n2579, n176 );
nor U5956 ( n2583, n2585, n39 );
nor U5957 ( n2585, n95, n2582 );
nor U5958 ( n2681, n186, n183 );
nand U5959 ( n3918, n2681, n2646 );
nor U5960 ( n2549, n2475, n198 );
not U5961 ( n198, n2526 );
or U5962 ( n3907, n2713, n2549 );
nor U5963 ( n2461, n203, n201 );
nand U5964 ( n3913, n3924, n3925 );
nor U5965 ( n3925, n3926, n3927 );
nor U5966 ( n3924, n3929, n3930 );
nand U5967 ( n3926, n2269, n147 );
nor U5968 ( n2522, n193, n191 );
nand U5969 ( n2578, n2579, n2558 );
nand U5970 ( n2672, n2673, n2674 );
nand U5971 ( n2674, n5224, n1286 );
nand U5972 ( n2673, n5217, n13 );
and U5973 ( n1638, n1649, n1646 );
nor U5974 ( n2775, n165, n164 );
not U5975 ( n156, n2301 );
not U5976 ( n160, n2746 );
not U5977 ( n272, n2054 );
nor U5978 ( n3897, n3903, n3904 );
nand U5979 ( n3904, n2201, n124 );
nand U5980 ( n3903, n280, n272 );
nor U5981 ( n1692, n1673, n248 );
not U5982 ( n147, n2238 );
not U5983 ( n268, n1990 );
nand U5984 ( n1077, n5203, n501 );
not U5985 ( n207, n2389 );
not U5986 ( n226, n4041 );
not U5987 ( n124, n2171 );
not U5988 ( n250, n1811 );
or U5989 ( n3911, n1777, n1673 );
not U5990 ( n213, n2432 );
not U5991 ( n262, n1930 );
not U5992 ( n256, n1862 );
not U5993 ( n218, n2353 );
xor U5994 ( n1298, n2666, n2713 );
nand U5995 ( n1473, n2698, n2699 );
nor U5996 ( n2699, n2700, n2701 );
nor U5997 ( n2698, n2708, n1310 );
nor U5998 ( n2700, n298, n5201 );
and U5999 ( n1679, n1664, n1681 );
not U6000 ( n10, n1382 );
not U6001 ( n280, n2150 );
not U6002 ( n233, n1629 );
xor U6003 ( n2718, n2616, n2713 );
not U6004 ( n135, n2029 );
nand U6005 ( n2127, n135, n2091 );
nor U6006 ( n2734, n95, n2743 );
nor U6007 ( n2743, n2744, n2745 );
nor U6008 ( n2744, n2751, n2752 );
nor U6009 ( n2745, n2746, n2721 );
nand U6010 ( n1476, n2725, n2726 );
nor U6011 ( n2726, n2727, n2728 );
nor U6012 ( n2725, n2731, n1331 );
nor U6013 ( n2727, n297, n5201 );
not U6014 ( n116, n2820 );
nand U6015 ( n1761, n245, n1681 );
not U6016 ( n245, n1777 );
nor U6017 ( n1545, n231, n235 );
not U6018 ( n235, n1522 );
nand U6019 ( n1553, n1554, n230 );
not U6020 ( n230, n1548 );
nand U6021 ( n1573, n231, n1588 );
nor U6022 ( n2493, n95, n2495 );
not U6023 ( n12, n2741 );
nand U6024 ( n2764, n2781, n2782 );
nand U6025 ( n2782, n2775, n12 );
or U6026 ( n2781, n2773, n12 );
nand U6027 ( n1479, n2755, n2756 );
nor U6028 ( n2756, n2757, n2758 );
nor U6029 ( n2755, n2765, n1348 );
nor U6030 ( n2757, n296, n5201 );
not U6031 ( n215, n2398 );
nand U6032 ( n2769, n2770, n2771 );
nand U6033 ( n2770, n2774, n2775 );
nand U6034 ( n2771, n2772, n2773 );
nor U6035 ( n2774, n95, n2750 );
nor U6036 ( n2776, n2777, n2778 );
nor U6037 ( n2777, n104, n2741 );
nor U6038 ( n2778, n95, n37 );
nor U6039 ( n2751, n165, n2750 );
not U6040 ( n251, n1681 );
and U6041 ( n3962, n1792, n1649 );
nor U6042 ( n2019, n97, n2012 );
nand U6043 ( n2728, n2729, n2730 );
nand U6044 ( n2730, n5224, n1330 );
nand U6045 ( n2729, n5217, n1319 );
not U6046 ( n180, n2646 );
nor U6047 ( n1974, n261, n276 );
nand U6048 ( n1759, n1659, n1680 );
nand U6049 ( n1482, n2789, n2790 );
nor U6050 ( n2790, n2791, n2792 );
nor U6051 ( n2789, n2795, n1365 );
nor U6052 ( n2791, n295, n5201 );
nand U6053 ( n2207, n2201, n2142 );
nor U6054 ( n2431, n2362, n215 );
nand U6055 ( n2644, n2142, n2649 );
nand U6056 ( n2577, n2582, n2142 );
nor U6057 ( n1810, n251, n253 );
buf U6058 ( n5205, n5105 );
not U6059 ( n57, n588 );
not U6060 ( n58, n4589 );
nand U6061 ( n2792, n2793, n2794 );
nand U6062 ( n2794, n5224, n1364 );
nand U6063 ( n2793, n5218, n1355 );
not U6064 ( n90, n3243 );
buf U6065 ( n5185, n5106 );
nor U6066 ( n785, n5199, n756 );
not U6067 ( n5195, n5196 );
not U6068 ( n5194, n5196 );
and U6069 ( n1383, n2812, n1382 );
nand U6070 ( n2812, n95, n103 );
not U6071 ( n96, n1941 );
nand U6072 ( n2845, n5244, n5215 );
and U6073 ( n5096, n5179, n5244 );
not U6074 ( n111, n1565 );
buf U6075 ( n5122, n5197 );
not U6076 ( n283, n3794 );
not U6077 ( n107, n3240 );
buf U6078 ( n5121, n5197 );
buf U6079 ( n5120, n5197 );
buf U6080 ( n5168, n5171 );
buf U6081 ( n5199, n5198 );
nor U6082 ( n3412, n293, n5165 );
buf U6083 ( n5169, n5171 );
nor U6084 ( n3395, n305, n5165 );
nor U6085 ( n3291, n325, n5166 );
nor U6086 ( n3246, n320, n5166 );
nor U6087 ( n3145, n317, n5166 );
nor U6088 ( n3380, n298, n5165 );
nor U6089 ( n3206, n303, n5166 );
nor U6090 ( n3347, n315, n5166 );
nor U6091 ( n3487, n307, n5165 );
nor U6092 ( n3331, n300, n5166 );
nor U6093 ( n3533, n301, n5165 );
nor U6094 ( n3123, n297, n5166 );
nor U6095 ( n3667, n312, n5165 );
nor U6096 ( n3311, n313, n5166 );
nor U6097 ( n3366, n323, n5166 );
nor U6098 ( n3471, n321, n5165 );
nor U6099 ( n3518, n316, n5165 );
nor U6100 ( n3160, n328, n5166 );
nor U6101 ( n3445, n310, n5165 );
nor U6102 ( n3271, n308, n5166 );
nor U6103 ( n3423, n318, n5165 );
nor U6104 ( n3554, n326, n5165 );
buf U6105 ( n5170, n5171 );
nor U6106 ( n3091, n322, n5167 );
nor U6107 ( n3030, n302, n5167 );
nor U6108 ( n3107, n306, n5167 );
nor U6109 ( n3059, n327, n5167 );
nor U6110 ( n3076, n311, n5167 );
not U6111 ( n110, n1554 );
nand U6112 ( n2075, n1620, n1549 );
nor U6113 ( n3812, n101, n1820 );
nand U6114 ( n3417, n3821, n5185 );
nor U6115 ( n3821, n3794, n2820 );
or U6116 ( n3239, n3055, n5123 );
nor U6117 ( n2655, n298, n5132 );
nor U6118 ( n2618, n300, n5133 );
nor U6119 ( n2443, n306, n5130 );
nor U6120 ( n2081, n317, n5126 );
nor U6121 ( n2687, n297, n5131 );
nor U6122 ( n1703, n325, n5129 );
nor U6123 ( n2210, n313, n5133 );
nor U6124 ( n2780, n293, n5130 );
not U6125 ( n101, n4020 );
nand U6126 ( n3529, n476, n3055 );
nand U6127 ( n3327, n473, n3055 );
nand U6128 ( n3087, n501, n3055 );
nand U6129 ( n3119, n496, n3055 );
nand U6130 ( n3218, n493, n3055 );
nand U6131 ( n3550, n502, n3055 );
nand U6132 ( n3287, n498, n3055 );
nand U6133 ( n3072, n3416, n3660 );
nand U6134 ( n3660, n3661, n5244 );
nand U6135 ( n3661, n63, n3662 );
nand U6136 ( n3662, n5185, n283 );
nor U6137 ( n3413, n3414, n3415 );
nand U6138 ( n3414, n3417, n5244 );
nand U6139 ( n3415, n63, n3416 );
nor U6140 ( n2813, n293, n5201 );
nand U6141 ( n2402, n1620, n110 );
not U6142 ( n105, n1549 );
nand U6143 ( n3416, n3797, n283 );
buf U6144 ( n5181, n5108 );
nor U6145 ( n3502, n293, n3240 );
buf U6146 ( n5223, n102 );
not U6147 ( n108, n1620 );
nor U6148 ( n3222, n292, n3240 );
buf U6149 ( n5142, n5143 );
buf U6150 ( n5217, n113 );
buf U6151 ( n5218, n113 );
buf U6152 ( n5219, n113 );
buf U6153 ( n5201, n5198 );
nor U6154 ( n1776, n98, n99 );
nor U6155 ( n2174, n1565, n112 );
not U6156 ( n98, n1975 );
or U6157 ( n5097, n5162, n4658 );
xnor U6158 ( n3238, n5160, n3751 );
nor U6159 ( n3751, n3752, n3753 );
nor U6160 ( n3753, n293, n5157 );
nor U6161 ( n3752, n163, n5155 );
nand U6162 ( n1820, n1975, n1619 );
nor U6163 ( n3746, n3237, n3238 );
nand U6164 ( n3525, n3597, n3598 );
nand U6165 ( n3598, n83, n3359 );
nor U6166 ( n3597, n3599, n3600 );
nor U6167 ( n3600, n89, n3601 );
nand U6168 ( n3510, n3742, n3743 );
nand U6169 ( n3743, n3238, n3237 );
nor U6170 ( n3742, n3744, n3745 );
nor U6171 ( n3745, n3746, n3747 );
nand U6172 ( n3322, n3609, n3610 );
nand U6173 ( n3609, n3614, n3613 );
nand U6174 ( n3610, n3611, n3612 );
or U6175 ( n3611, n3613, n3614 );
nor U6176 ( n4671, n106, n143 );
nor U6177 ( n3733, n3736, n3136 );
nor U6178 ( n3736, n3138, n3137 );
nor U6179 ( n3599, n3603, n3358 );
nor U6180 ( n3603, n3359, n3602 );
nor U6181 ( n3705, n3716, n3717 );
and U6182 ( n3717, n3339, n3336 );
nor U6183 ( n3716, n3338, n3546 );
nand U6184 ( n3578, n3579, n3580 );
nand U6185 ( n3579, n3096, n3098 );
nand U6186 ( n3580, n3581, n3099 );
or U6187 ( n3581, n3098, n3096 );
and U6188 ( n3153, n3592, n3593 );
nand U6189 ( n3592, n3523, n3525 );
nand U6190 ( n3593, n3594, n3526 );
or U6191 ( n3594, n3525, n3523 );
and U6192 ( n3338, n3723, n3724 );
nand U6193 ( n3723, n3387, n3388 );
nand U6194 ( n3724, n3385, n3725 );
or U6195 ( n3725, n3388, n3387 );
nand U6196 ( n4669, n4670, n97 );
nor U6197 ( n4670, n92, n3814 );
not U6198 ( n144, n2928 );
xor U6199 ( n3166, n3167, n3168 );
nand U6200 ( n3167, n3194, n3195 );
nand U6201 ( n3168, n3169, n3170 );
nand U6202 ( n3194, n5114, n811 );
not U6203 ( n5162, n5089 );
nand U6204 ( n3169, n3067, n3171 );
nand U6205 ( n3171, n3064, n3066 );
nand U6206 ( n3161, n3162, n3163 );
nand U6207 ( n3162, n5220, n832 );
nand U6208 ( n3163, n3164, n5168 );
xor U6209 ( n3164, n3165, n3166 );
nand U6210 ( n3402, n3693, n3694 );
nand U6211 ( n3693, n3214, n3213 );
nand U6212 ( n3694, n3211, n3695 );
or U6213 ( n3695, n3213, n3214 );
nand U6214 ( n3114, n3688, n3689 );
nand U6215 ( n3688, n3400, n3402 );
nand U6216 ( n3689, n3690, n3403 );
or U6217 ( n3690, n3402, n3400 );
nand U6218 ( n3463, n3683, n3684 );
nand U6219 ( n3683, n3112, n3114 );
nand U6220 ( n3684, n3685, n3115 );
or U6221 ( n3685, n3114, n3112 );
nand U6222 ( n3612, n3675, n3676 );
nand U6223 ( n3675, n3081, n3084 );
nand U6224 ( n3676, n3677, n3083 );
or U6225 ( n3677, n3084, n3081 );
nand U6226 ( n3098, n3584, n3585 );
nand U6227 ( n3584, n3476, n3478 );
nand U6228 ( n3585, n3586, n3479 );
or U6229 ( n3586, n3478, n3476 );
nand U6230 ( n3302, n3573, n3574 );
nand U6231 ( n3573, n80, n3578 );
nand U6232 ( n3574, n3575, n3190 );
nand U6233 ( n3575, n2, n3371 );
nand U6234 ( n3555, n3556, n3557 );
nand U6235 ( n3556, n5222, n867 );
nand U6236 ( n3557, n3558, n5168 );
nor U6237 ( n3558, n3559, n3560 );
nand U6238 ( n1975, n4671, n122 );
nor U6239 ( n3559, n3565, n3566 );
xor U6240 ( n3565, n3564, n3563 );
nand U6241 ( n3566, n3567, n3191 );
nand U6242 ( n3567, n3302, n3303 );
nand U6243 ( n3060, n3061, n3062 );
nand U6244 ( n3061, n5220, n851 );
nand U6245 ( n3062, n5168, n3063 );
xnor U6246 ( n3063, n3064, n3065 );
nor U6247 ( n4656, n36, n5155 );
nand U6248 ( n3292, n3293, n3294 );
nand U6249 ( n3293, n5220, n891 );
nand U6250 ( n3294, n5169, n3295 );
nand U6251 ( n3295, n3296, n3297 );
nand U6252 ( n3297, n3298, n1 );
xor U6253 ( n3298, n3299, n3300 );
not U6254 ( n92, n2824 );
xnor U6255 ( n3512, n5160, n3737 );
nor U6256 ( n3737, n3738, n3739 );
nor U6257 ( n3739, n295, n5157 );
nor U6258 ( n3738, n166, n5155 );
nand U6259 ( n3133, n3512, n3511 );
nand U6260 ( n3367, n3368, n3369 );
nand U6261 ( n3368, n5221, n907 );
nand U6262 ( n3369, n5169, n3370 );
xor U6263 ( n3370, n3371, n3372 );
not U6264 ( n282, n4305 );
not U6265 ( n291, n4933 );
or U6266 ( n3132, n3511, n3512 );
xor U6267 ( n3138, n5161, n3758 );
nor U6268 ( n3758, n3759, n3760 );
nor U6269 ( n3760, n296, n5157 );
nor U6270 ( n3759, n161, n5155 );
nand U6271 ( n3092, n3093, n3094 );
nand U6272 ( n3093, n5220, n931 );
nand U6273 ( n3094, n5170, n3095 );
xnor U6274 ( n3095, n3096, n3097 );
buf U6275 ( n5213, n5210 );
buf U6276 ( n5214, n5210 );
nand U6277 ( n3247, n3248, n3249 );
nand U6278 ( n3248, n5220, n972 );
nand U6279 ( n3249, n3250, n5168 );
nor U6280 ( n3250, n3251, n3252 );
nor U6281 ( n3251, n3257, n3258 );
xor U6282 ( n3257, n3262, n3263 );
nand U6283 ( n3258, n3259, n81 );
nand U6284 ( n3259, n3260, n3261 );
nand U6285 ( n3472, n3473, n3474 );
nand U6286 ( n3473, n5221, n952 );
nand U6287 ( n3474, n5168, n3475 );
xnor U6288 ( n3475, n3476, n3477 );
xnor U6289 ( n3336, n5160, n3718 );
nor U6290 ( n3718, n3719, n3720 );
nor U6291 ( n3720, n298, n5157 );
nor U6292 ( n3719, n185, n5155 );
nor U6293 ( n3546, n3339, n3336 );
xnor U6294 ( n3385, n5160, n3726 );
nor U6295 ( n3726, n3727, n3728 );
nor U6296 ( n3728, n297, n5157 );
nor U6297 ( n3727, n169, n5155 );
nand U6298 ( n3424, n3425, n3426 );
nand U6299 ( n3425, n5221, n995 );
nand U6300 ( n3426, n5169, n3427 );
nand U6301 ( n3427, n3428, n3429 );
nand U6302 ( n3429, n3430, n3 );
xor U6303 ( n3430, n3431, n3432 );
xnor U6304 ( n3542, n5160, n3706 );
nor U6305 ( n3706, n3707, n3708 );
nor U6306 ( n3708, n300, n3179 );
nor U6307 ( n3707, n177, n5155 );
or U6308 ( n3046, n3541, n3542 );
xnor U6309 ( n3151, n3152, n3153 );
nand U6310 ( n3146, n3147, n3148 );
nand U6311 ( n3147, n5220, n1017 );
nand U6312 ( n3148, n5169, n3149 );
xor U6313 ( n3149, n3150, n3151 );
nand U6314 ( n1297, n3143, n3144 );
nor U6315 ( n3143, n733, n3154 );
nor U6316 ( n3144, n3145, n3146 );
nand U6317 ( n3154, n3155, n3156 );
nand U6318 ( n3042, n3542, n3541 );
xnor U6319 ( n3524, n3525, n3526 );
nand U6320 ( n3519, n3520, n3521 );
nand U6321 ( n3520, n5221, n1040 );
nand U6322 ( n3521, n5169, n3522 );
xnor U6323 ( n3522, n3523, n3524 );
nand U6324 ( n1202, n3516, n3517 );
nor U6325 ( n3516, n648, n3527 );
nor U6326 ( n3517, n3518, n3519 );
nand U6327 ( n3527, n3528, n3529 );
nand U6328 ( n3348, n3349, n3350 );
nand U6329 ( n3349, n5221, n1063 );
nand U6330 ( n3350, n3351, n5168 );
nor U6331 ( n3351, n3352, n3353 );
nand U6332 ( n1252, n3345, n3346 );
nor U6333 ( n3345, n630, n3360 );
nor U6334 ( n3346, n3347, n3348 );
nand U6335 ( n3360, n3361, n3362 );
xor U6336 ( n3211, n5161, n3696 );
nor U6337 ( n3696, n3697, n3698 );
nor U6338 ( n3698, n302, n3179 );
nor U6339 ( n3697, n187, n5155 );
nor U6340 ( n3704, n3049, n3048 );
nand U6341 ( n4020, n4664, n143 );
nor U6342 ( n4664, n106, n122 );
not U6343 ( n5159, n3179 );
nand U6344 ( n3179, n4663, n4305 );
nand U6345 ( n4663, n4020, n4304 );
nand U6346 ( n1262, n3309, n3310 );
nor U6347 ( n3309, n611, n3325 );
nor U6348 ( n3310, n3311, n3312 );
nand U6349 ( n3325, n3326, n3327 );
nand U6350 ( n3312, n3313, n3314 );
nand U6351 ( n3313, n5221, n1080 );
nand U6352 ( n3314, n5169, n3315 );
nand U6353 ( n3315, n3316, n3317 );
nand U6354 ( n3317, n3318, n4 );
xor U6355 ( n3318, n3319, n3320 );
xor U6356 ( n3672, n3612, n3613 );
nand U6357 ( n3668, n3669, n3670 );
nand U6358 ( n3669, n5222, n1108 );
nand U6359 ( n3670, n5169, n3671 );
xor U6360 ( n3671, n3614, n3672 );
nand U6361 ( n1187, n3665, n3666 );
nor U6362 ( n3665, n592, n3799 );
nor U6363 ( n3666, n3667, n3668 );
nand U6364 ( n3799, n3800, n3801 );
nand U6365 ( n2823, n143, n122 );
xnor U6366 ( n3400, n5160, n3761 );
nor U6367 ( n3761, n3762, n3763 );
nor U6368 ( n3763, n303, n5157 );
nor U6369 ( n3762, n200, n5155 );
nand U6370 ( n3283, n3279, n3280 );
xor U6371 ( n3280, n5160, n3784 );
nor U6372 ( n3784, n3785, n3786 );
nor U6373 ( n3786, n307, n5157 );
nor U6374 ( n3785, n216, n5155 );
nand U6375 ( n4684, n4658, n3817 );
not U6376 ( n5160, n5161 );
nor U6377 ( n4662, n36, n5157 );
xor U6378 ( n3082, n3083, n3084 );
nand U6379 ( n3077, n3078, n3079 );
nand U6380 ( n3078, n5220, n1131 );
nand U6381 ( n3079, n5170, n3080 );
xor U6382 ( n3080, n3081, n3082 );
nand U6383 ( n1317, n3074, n3075 );
nor U6384 ( n3074, n572, n3085 );
nor U6385 ( n3075, n3076, n3077 );
nand U6386 ( n3085, n3086, n3087 );
nand U6387 ( n3446, n3447, n3448 );
nand U6388 ( n3447, n5221, n1153 );
nand U6389 ( n3448, n3449, n5168 );
nor U6390 ( n3449, n3450, n3451 );
nand U6391 ( n1222, n3443, n3444 );
nor U6392 ( n3443, n553, n3465 );
nor U6393 ( n3444, n3445, n3446 );
nand U6394 ( n3465, n3466, n3467 );
nand U6395 ( n3460, n3492, n3494 );
xnor U6396 ( n3492, n5160, n3774 );
nor U6397 ( n3774, n3775, n3776 );
nor U6398 ( n3776, n306, n5157 );
nor U6399 ( n3775, n202, n5155 );
xnor U6400 ( n3112, n5160, n3764 );
nor U6401 ( n3764, n3765, n3766 );
nor U6402 ( n3766, n305, n5157 );
nor U6403 ( n3765, n196, n5155 );
nor U6404 ( n3459, n3280, n3279 );
nor U6405 ( n3450, n3456, n3457 );
xor U6406 ( n3456, n3464, n87 );
nand U6407 ( n3457, n3458, n75 );
nand U6408 ( n3458, n3282, n3283 );
nand U6409 ( n3040, n3048, n3049 );
or U6410 ( n3462, n3494, n3492 );
nand U6411 ( n1272, n3269, n3270 );
nor U6412 ( n3269, n3284, n3285 );
nor U6413 ( n3270, n3271, n3272 );
nand U6414 ( n3285, n3286, n3287 );
nand U6415 ( n3272, n3273, n3274 );
nand U6416 ( n3273, n5220, n1176 );
nand U6417 ( n3274, n5169, n3275 );
nand U6418 ( n3275, n3276, n3277 );
nand U6419 ( n3277, n3278, n5 );
xor U6420 ( n3278, n3279, n3280 );
xnor U6421 ( n3493, n3463, n3494 );
nand U6422 ( n3488, n3489, n3490 );
nand U6423 ( n3489, n5221, n1198 );
nand U6424 ( n3490, n5168, n3491 );
xnor U6425 ( n3491, n3492, n3493 );
nand U6426 ( n1212, n3485, n3486 );
nor U6427 ( n3485, n3495, n3496 );
nor U6428 ( n3486, n3487, n3488 );
nand U6429 ( n3496, n3497, n3498 );
not U6430 ( n88, n3137 );
not U6431 ( n293, n1375 );
buf U6432 ( n5150, n5147 );
buf U6433 ( n5189, n5109 );
buf U6434 ( n5137, n5136 );
nor U6435 ( n4255, n1342, n161 );
nand U6436 ( n4249, n2719, n4253 );
nand U6437 ( n4253, n4254, n166 );
nor U6438 ( n4254, n295, n4255 );
nand U6439 ( n4138, n1646, n4139 );
nand U6440 ( n4139, n4140, n1650 );
nor U6441 ( n4140, n4141, n4142 );
nor U6442 ( n4142, n247, n325 );
nand U6443 ( n4178, n4187, n2369 );
nor U6444 ( n4187, n4188, n4189 );
nor U6445 ( n4189, n1153, n4190 );
nor U6446 ( n4188, n4191, n4192 );
nand U6447 ( n4150, n1903, n4151 );
nand U6448 ( n4151, n4152, n3901 );
nor U6449 ( n4152, n4153, n4154 );
nor U6450 ( n4154, n270, n320 );
nor U6451 ( n4170, n4171, n3928 );
nor U6452 ( n4171, n4172, n4173 );
nor U6453 ( n4172, n152, n1063 );
nand U6454 ( n4173, n2292, n4174 );
nand U6455 ( n4235, n4247, n4248 );
nand U6456 ( n4248, n4249, n1324 );
nor U6457 ( n4247, n4250, n4251 );
nor U6458 ( n4250, n4256, n4257 );
nor U6459 ( n4210, n4213, n4214 );
nand U6460 ( n4214, n4215, n4209 );
nand U6461 ( n4213, n4228, n4229 );
nor U6462 ( n4215, n4223, n4224 );
nor U6463 ( n4129, n4120, n4130 );
nand U6464 ( n4130, n4131, n4132 );
nand U6465 ( n4131, n328, n228 );
nand U6466 ( n4132, n4133, n4134 );
nor U6467 ( n4165, n4167, n4168 );
nor U6468 ( n4167, n145, n1017 );
nand U6469 ( n4168, n2216, n4169 );
nand U6470 ( n4169, n4170, n2214 );
nand U6471 ( n3880, n3881, n3882 );
nor U6472 ( n3882, n3883, n3884 );
nor U6473 ( n3881, n3931, n3932 );
nand U6474 ( n3884, n3885, n3886 );
nor U6475 ( n3931, n1377, n4126 );
nand U6476 ( n4126, n3960, n4127 );
nand U6477 ( n4127, n4128, n3949 );
nor U6478 ( n4128, n4129, n4103 );
buf U6479 ( n5154, n5151 );
xnor U6480 ( n3113, n3114, n3115 );
nand U6481 ( n3921, n163, n1375 );
nand U6482 ( n3108, n3109, n3110 );
nand U6483 ( n3109, n5220, n1214 );
nand U6484 ( n3110, n5170, n3111 );
xnor U6485 ( n3111, n3112, n3113 );
nand U6486 ( n1307, n3105, n3106 );
nor U6487 ( n3105, n3116, n3117 );
nor U6488 ( n3106, n3107, n3108 );
nand U6489 ( n3117, n3118, n3119 );
not U6490 ( n292, n2798 );
xnor U6491 ( n3081, n5160, n3787 );
nor U6492 ( n3787, n3788, n3789 );
nor U6493 ( n3789, n310, n5157 );
nor U6494 ( n3788, n222, n5155 );
nand U6495 ( n3768, n87, n3464 );
xnor U6496 ( n3614, n3175, n3790 );
nor U6497 ( n3790, n3791, n3792 );
nor U6498 ( n3792, n311, n5157 );
nor U6499 ( n3791, n158, n5155 );
nand U6500 ( n2719, n161, n1342 );
nand U6501 ( n3323, n3320, n3319 );
xnor U6502 ( n3320, n3175, n3604 );
nor U6503 ( n3604, n3605, n3606 );
nor U6504 ( n3606, n312, n3179 );
nor U6505 ( n3605, n152, n5155 );
nor U6506 ( n3601, n83, n3359 );
buf U6507 ( n5146, n4314 );
not U6508 ( n295, n1359 );
or U6509 ( n3324, n3319, n3320 );
xnor U6510 ( n3401, n3402, n3403 );
nand U6511 ( n3396, n3397, n3398 );
nand U6512 ( n3397, n5221, n1239 );
nand U6513 ( n3398, n5169, n3399 );
xnor U6514 ( n3399, n3400, n3401 );
nand U6515 ( n1237, n3393, n3394 );
nor U6516 ( n3393, n3404, n3405 );
nor U6517 ( n3394, n3395, n3396 );
nand U6518 ( n3405, n3406, n3407 );
not U6519 ( n296, n1342 );
nand U6520 ( n3454, n70, n3770 );
not U6521 ( n70, n3464 );
nand U6522 ( n4257, n2749, n2685 );
nand U6523 ( n2582, n175, n1260 );
and U6524 ( n4231, n2582, n4240 );
nand U6525 ( n4240, n177, n1280 );
xor U6526 ( n3212, n3213, n3214 );
nand U6527 ( n3207, n3208, n3209 );
nand U6528 ( n3208, n5220, n1260 );
nand U6529 ( n3209, n5169, n3210 );
xor U6530 ( n3210, n3211, n3212 );
nand U6531 ( n1287, n3204, n3205 );
nor U6532 ( n3204, n3215, n3216 );
nor U6533 ( n3205, n3206, n3207 );
nand U6534 ( n3216, n3217, n3218 );
nand U6535 ( n2649, n185, n1303 );
nand U6536 ( n3261, n3431, n3432 );
nand U6537 ( n4229, n4230, n4231 );
nor U6538 ( n4230, n185, n1303 );
or U6539 ( n3624, n3262, n3263 );
nand U6540 ( n3047, n3544, n3545 );
nand U6541 ( n3544, n3336, n3339 );
or U6542 ( n3545, n3546, n3338 );
nand U6543 ( n3031, n3032, n3033 );
nand U6544 ( n3032, n5220, n1280 );
nand U6545 ( n3033, n3034, n5168 );
nor U6546 ( n3034, n3036, n3037 );
nand U6547 ( n1327, n3028, n3029 );
nor U6548 ( n3028, n3051, n3052 );
nor U6549 ( n3029, n3030, n3031 );
nand U6550 ( n3052, n3053, n3054 );
nor U6551 ( n4224, n175, n1260 );
nor U6552 ( n4223, n187, n1239 );
nand U6553 ( n3434, n3150, n3152 );
xnor U6554 ( n3150, n3175, n3629 );
nor U6555 ( n3629, n3630, n3631 );
nor U6556 ( n3631, n316, n3179 );
nor U6557 ( n3630, n137, n5155 );
xnor U6558 ( n3523, n3175, n3620 );
nor U6559 ( n3620, n3621, n3622 );
nor U6560 ( n3622, n315, n3179 );
nor U6561 ( n3621, n145, n5155 );
nor U6562 ( n3036, n3043, n3044 );
xor U6563 ( n3043, n3048, n3049 );
nand U6564 ( n3044, n3045, n3042 );
nand U6565 ( n3045, n3046, n3047 );
nor U6566 ( n3437, n3432, n3431 );
buf U6567 ( n5215, n5210 );
nand U6568 ( n3534, n3535, n3536 );
nand U6569 ( n3535, n5221, n1303 );
nand U6570 ( n3536, n5168, n3537 );
nand U6571 ( n3537, n3538, n3539 );
nand U6572 ( n3539, n3540, n6 );
xor U6573 ( n3540, n3541, n3542 );
nand U6574 ( n1197, n3531, n3532 );
nor U6575 ( n3531, n3547, n3548 );
nor U6576 ( n3532, n3533, n3534 );
nand U6577 ( n3548, n3549, n3550 );
nor U6578 ( n3436, n3152, n3150 );
not U6579 ( n298, n1303 );
not U6580 ( n297, n1324 );
nand U6581 ( n4212, n2452, n1214 );
nand U6582 ( n3255, n3263, n3262 );
nand U6583 ( n2366, n210, n1131 );
nand U6584 ( n2414, n216, n1153 );
xor U6585 ( n3337, n3338, n3339 );
nand U6586 ( n3332, n3333, n3334 );
nand U6587 ( n3333, n5221, n1324 );
nand U6588 ( n3334, n5169, n3335 );
xnor U6589 ( n3335, n3336, n3337 );
nand U6590 ( n1257, n3329, n3330 );
nor U6591 ( n3329, n3340, n3341 );
nor U6592 ( n3330, n3331, n3332 );
nand U6593 ( n3341, n3342, n3343 );
not U6594 ( n300, n1280 );
nor U6595 ( n4534, n3551, n5137 );
nand U6596 ( n2098, n2175, n2176 );
nand U6597 ( n2176, n2177, n2178 );
nand U6598 ( n2750, n3921, n4008 );
nand U6599 ( n4008, n3922, n2804 );
nand U6600 ( n2373, n2555, n2556 );
nand U6601 ( n2555, n2557, n2558 );
nor U6602 ( n2557, n172, n2559 );
nand U6603 ( n2178, n2214, n2215 );
nand U6604 ( n2215, n2216, n2217 );
nand U6605 ( n2327, n2366, n2367 );
nand U6606 ( n2367, n2368, n2369 );
nand U6607 ( n2368, n2370, n2371 );
or U6608 ( n2371, n2372, n2373 );
nand U6609 ( n2721, n2747, n2748 );
nand U6610 ( n2748, n2749, n2750 );
nand U6611 ( n2217, n2239, n2240 );
nand U6612 ( n2239, n2244, n2245 );
nand U6613 ( n2240, n2241, n2242 );
nand U6614 ( n2244, n2246, n2247 );
and U6615 ( n1717, n1796, n1798 );
nand U6616 ( n1798, n1799, n1792 );
nand U6617 ( n2558, n2580, n2581 );
nand U6618 ( n1404, n1667, n1668 );
nor U6619 ( n1668, n1669, n1670 );
nor U6620 ( n1667, n1683, n818 );
nor U6621 ( n1669, n327, n5199 );
nand U6622 ( n1711, n1712, n1713 );
nand U6623 ( n1713, n1714, n1649 );
or U6624 ( n1712, n1625, n1691 );
nor U6625 ( n2241, n50, n220 );
not U6626 ( n220, n2243 );
nand U6627 ( n2616, n2719, n2720 );
nand U6628 ( n2720, n2721, n2722 );
nand U6629 ( n2580, n2608, n2609 );
nand U6630 ( n2609, n2610, n2611 );
nand U6631 ( n2608, n167, n2616 );
nand U6632 ( n2611, n2612, n2613 );
buf U6633 ( n5153, n5151 );
nand U6634 ( n798, n1608, n1609 );
nand U6635 ( n1609, n60, n832 );
nor U6636 ( n1608, n1610, n1611 );
nor U6637 ( n1610, n1628, n1629 );
nand U6638 ( n1401, n1592, n1593 );
nor U6639 ( n1593, n1594, n1595 );
nor U6640 ( n1592, n1607, n798 );
nor U6641 ( n1594, n328, n5199 );
nor U6642 ( n1622, n1623, n1624 );
nor U6643 ( n1623, n46, n111 );
nor U6644 ( n1624, n43, n1625 );
nand U6645 ( n4179, n2243, n4180 );
nand U6646 ( n4180, n4181, n4182 );
nor U6647 ( n4181, n202, n1176 );
nand U6648 ( n813, n815, n816 );
nand U6649 ( n816, n817, n5239 );
nand U6650 ( n815, n5231, n818 );
nand U6651 ( n949, n800, n801 );
nor U6652 ( n801, n802, n803 );
nor U6653 ( n800, n812, n813 );
nand U6654 ( n803, n805, n806 );
nand U6655 ( n954, n777, n778 );
nor U6656 ( n778, n780, n781 );
nor U6657 ( n777, n793, n795 );
nand U6658 ( n781, n782, n783 );
nand U6659 ( n795, n796, n797 );
nand U6660 ( n797, n236, n5235 );
nand U6661 ( n796, n5230, n798 );
nor U6662 ( n1641, n1642, n1643 );
nor U6663 ( n1642, n1572, n111 );
nor U6664 ( n1643, n1586, n1625 );
nand U6665 ( n767, n1528, n1529 );
nor U6666 ( n1529, n1530, n1531 );
nor U6667 ( n1528, n1561, n1562 );
nand U6668 ( n1530, n1539, n1540 );
nand U6669 ( n1398, n1512, n1513 );
nor U6670 ( n1513, n1514, n1515 );
nor U6671 ( n1512, n1527, n767 );
nor U6672 ( n1514, n1493, n776 );
nor U6673 ( n2612, n183, n2615 );
xnor U6674 ( n3386, n3387, n3388 );
nand U6675 ( n1242, n3378, n3379 );
nor U6676 ( n3378, n3389, n3390 );
nor U6677 ( n3379, n3380, n3381 );
nand U6678 ( n3390, n3391, n3392 );
nand U6679 ( n3381, n3382, n3383 );
nand U6680 ( n3382, n5221, n1342 );
nand U6681 ( n3383, n5169, n3384 );
xnor U6682 ( n3384, n3385, n3386 );
nand U6683 ( n1947, n1998, n1999 );
nor U6684 ( n1999, n2000, n2001 );
nor U6685 ( n1998, n2004, n2005 );
nor U6686 ( n2001, n97, n2002 );
nor U6687 ( n1942, n267, n1945 );
nor U6688 ( n1945, n1946, n1947 );
nor U6689 ( n1946, n111, n1948 );
and U6690 ( n1952, n2002, n2011 );
nand U6691 ( n2011, n2070, n2012 );
nand U6692 ( n1416, n1924, n1925 );
nor U6693 ( n1925, n1926, n1927 );
nor U6694 ( n1924, n1931, n898 );
nor U6695 ( n1926, n322, n5199 );
nand U6696 ( n1938, n1939, n1940 );
nand U6697 ( n1940, n271, n1941 );
nor U6698 ( n1939, n1942, n1943 );
nor U6699 ( n1943, n1944, n1891 );
nand U6700 ( n893, n895, n896 );
nand U6701 ( n896, n897, n5239 );
nand U6702 ( n895, n5231, n898 );
nand U6703 ( n929, n880, n881 );
nor U6704 ( n881, n882, n883 );
nor U6705 ( n880, n892, n893 );
nand U6706 ( n883, n885, n886 );
nand U6707 ( n2747, n166, n1359 );
not U6708 ( n87, n3770 );
nand U6709 ( n2683, n169, n1324 );
nand U6710 ( n2613, n168, n2614 );
nor U6711 ( n1615, n1617, n1618 );
nor U6712 ( n1617, n1546, n1620 );
nor U6713 ( n1618, n45, n1619 );
not U6714 ( n305, n1198 );
buf U6715 ( n5149, n5147 );
nand U6716 ( n3985, n4005, n2610 );
and U6717 ( n4005, n2614, n2685 );
nor U6718 ( n4498, n3120, n5137 );
or U6719 ( n3303, n3299, n3300 );
or U6720 ( n3184, n3564, n3563 );
nor U6721 ( n1632, n1634, n1635 );
nor U6722 ( n1634, n26, n1620 );
nor U6723 ( n1635, n1579, n1619 );
not U6724 ( n303, n1214 );
not U6725 ( n80, n3371 );
nand U6726 ( n1728, n1682, n1848 );
nand U6727 ( n1848, n1660, n1657 );
nand U6728 ( n2666, n2714, n2715 );
nand U6729 ( n2715, n2716, n2717 );
nand U6730 ( n1958, n2021, n2022 );
and U6731 ( n2021, n2031, n2032 );
nand U6732 ( n2022, n2023, n2024 );
nand U6733 ( n2032, n2033, n2034 );
nand U6734 ( n2741, n2783, n2784 );
nand U6735 ( n2784, n2785, n2786 );
nand U6736 ( n2716, n2739, n2740 );
nand U6737 ( n2740, n2741, n2742 );
nor U6738 ( n2785, n292, n36 );
nor U6739 ( n2480, n2481, n2482 );
nand U6740 ( n2482, n2483, n195 );
nand U6741 ( n2481, n2484, n2485 );
nand U6742 ( n2304, n2469, n2470 );
nand U6743 ( n2470, n2471, n2472 );
nor U6744 ( n2469, n2479, n2480 );
nand U6745 ( n2471, n2473, n2474 );
nand U6746 ( n2495, n196, n1198 );
nand U6747 ( n2370, n2411, n2412 );
nand U6748 ( n2412, n2413, n2414 );
nand U6749 ( n2413, n2415, n2416 );
nand U6750 ( n2415, n2450, n2451 );
nand U6751 ( n2451, n197, n2452 );
nand U6752 ( n3124, n3125, n3126 );
nand U6753 ( n3125, n5220, n1359 );
nand U6754 ( n3126, n3127, n5168 );
nor U6755 ( n3127, n3128, n3129 );
nand U6756 ( n1302, n3121, n3122 );
nor U6757 ( n3121, n3139, n3140 );
nor U6758 ( n3122, n3123, n3124 );
nand U6759 ( n3140, n3141, n3142 );
nand U6760 ( n1562, n1563, n1564 );
nand U6761 ( n1563, n60, n811 );
nand U6762 ( n1564, n1565, n1566 );
nand U6763 ( n1566, n1567, n1568 );
nand U6764 ( n4066, n202, n1176 );
nor U6765 ( n2005, n1965, n1625 );
nand U6766 ( n1407, n1735, n1736 );
nor U6767 ( n1736, n1737, n1738 );
nor U6768 ( n1735, n1748, n838 );
nor U6769 ( n1737, n326, n5199 );
nand U6770 ( n2247, n158, n1080 );
nand U6771 ( n2786, n293, n163 );
nand U6772 ( n3191, n3300, n3299 );
nand U6773 ( n1546, n1654, n1655 );
and U6774 ( n1654, n1603, n1661 );
nand U6775 ( n1655, n1656, n1657 );
nand U6776 ( n1661, n1662, n1605 );
nand U6777 ( n1710, n1718, n1719 );
nand U6778 ( n1718, n248, n1722 );
nand U6779 ( n1719, n98, n1720 );
nand U6780 ( n1722, n1619, n111 );
nand U6781 ( n1720, n1721, n1696 );
nand U6782 ( n835, n836, n837 );
nand U6783 ( n837, n247, n5235 );
nand U6784 ( n836, n5231, n838 );
nand U6785 ( n944, n820, n821 );
nor U6786 ( n821, n822, n823 );
nor U6787 ( n820, n833, n835 );
nand U6788 ( n822, n828, n830 );
nor U6789 ( n4516, n3219, n5137 );
nand U6790 ( n2533, n200, n1214 );
nor U6791 ( n2535, n1214, n200 );
nand U6792 ( n2372, n2409, n2410 );
nor U6793 ( n2409, n217, n203 );
not U6794 ( n217, n2411 );
buf U6795 ( n5145, n4314 );
nand U6796 ( n1419, n1979, n1980 );
nor U6797 ( n1980, n1981, n1982 );
nor U6798 ( n1979, n1991, n918 );
nor U6799 ( n1981, n321, n5199 );
nand U6800 ( n918, n1992, n1993 );
nand U6801 ( n1993, n60, n952 );
nor U6802 ( n1992, n1994, n1995 );
nor U6803 ( n1994, n2006, n1990 );
nand U6804 ( n924, n900, n901 );
nor U6805 ( n901, n902, n903 );
nor U6806 ( n900, n913, n915 );
nand U6807 ( n903, n905, n906 );
nand U6808 ( n915, n916, n917 );
nand U6809 ( n917, n270, n5235 );
nand U6810 ( n916, n5231, n918 );
nor U6811 ( n1788, n1717, n1625 );
nor U6812 ( n1833, n1835, n1836 );
nor U6813 ( n1835, n1827, n111 );
nor U6814 ( n1836, n42, n1625 );
nand U6815 ( n1410, n1802, n1803 );
nor U6816 ( n1803, n1804, n1805 );
nor U6817 ( n1802, n1812, n858 );
nor U6818 ( n1804, n325, n5199 );
nand U6819 ( n853, n855, n856 );
nand U6820 ( n856, n857, n5239 );
nand U6821 ( n855, n5231, n858 );
nand U6822 ( n939, n840, n841 );
nor U6823 ( n841, n842, n843 );
nor U6824 ( n840, n852, n853 );
nand U6825 ( n842, n848, n850 );
nand U6826 ( n2186, n2218, n2219 );
and U6827 ( n2218, n2220, n2221 );
nand U6828 ( n2219, n148, n2024 );
nand U6829 ( n2221, n154, n2036 );
nand U6830 ( n1422, n2046, n2047 );
nor U6831 ( n2047, n2048, n2049 );
nor U6832 ( n2046, n2060, n938 );
nor U6833 ( n2048, n320, n5199 );
nand U6834 ( n2058, n2043, n2185 );
nand U6835 ( n2185, n2186, n2027 );
not U6836 ( n302, n1239 );
not U6837 ( n306, n1176 );
nand U6838 ( n933, n935, n936 );
nand U6839 ( n936, n937, n5238 );
nand U6840 ( n935, n5231, n938 );
nand U6841 ( n919, n920, n921 );
nor U6842 ( n921, n922, n923 );
nor U6843 ( n920, n932, n933 );
nand U6844 ( n923, n925, n926 );
not U6845 ( n191, n2452 );
nand U6846 ( n3508, n3509, n7 );
xor U6847 ( n3509, n3511, n3512 );
nor U6848 ( n1515, n768, n1516 );
nand U6849 ( n1606, n1674, n1675 );
nand U6850 ( n1674, n1677, n1678 );
nand U6851 ( n1675, n1676, n1659 );
nand U6852 ( n1677, n1679, n1680 );
nand U6853 ( n1526, n1603, n1604 );
nand U6854 ( n1604, n1605, n1606 );
and U6855 ( n768, n1517, n1518 );
nand U6856 ( n1517, n1523, n1524 );
nand U6857 ( n1518, n231, n1519 );
nand U6858 ( n1524, n1522, n1525 );
nand U6859 ( n1519, n1520, n1521 );
nand U6860 ( n1521, n25, n1522 );
and U6861 ( n1676, n1657, n1660 );
nand U6862 ( n2742, n295, n166 );
nand U6863 ( n3186, n3563, n3564 );
not U6864 ( n203, n2416 );
nand U6865 ( n1525, n1520, n1526 );
nand U6866 ( n1595, n1596, n1597 );
nand U6867 ( n1597, n791, n5223 );
nand U6868 ( n1596, n5217, n792 );
buf U6869 ( n5138, n5136 );
nor U6870 ( n4480, n3288, n5138 );
nor U6871 ( n1871, n1873, n1874 );
nor U6872 ( n1873, n110, n1657 );
nor U6873 ( n1874, n1549, n1657 );
nand U6874 ( n1413, n1851, n1852 );
nor U6875 ( n1852, n1853, n1854 );
nor U6876 ( n1851, n1863, n878 );
nor U6877 ( n1853, n323, n5199 );
not U6878 ( n307, n1153 );
nand U6879 ( n1738, n1739, n1740 );
nand U6880 ( n1740, n831, n5223 );
nand U6881 ( n1739, n5219, n827 );
nand U6882 ( n875, n876, n877 );
nand U6883 ( n877, n258, n5235 );
nand U6884 ( n876, n5231, n878 );
nand U6885 ( n934, n860, n861 );
nor U6886 ( n861, n862, n863 );
nor U6887 ( n860, n873, n875 );
nand U6888 ( n863, n865, n866 );
or U6889 ( n1747, n1761, n5098 );
and U6890 ( n5098, n1728, n1764 );
nand U6891 ( n2717, n296, n161 );
nand U6892 ( n1805, n1806, n1807 );
nand U6893 ( n1807, n857, n5223 );
nand U6894 ( n1806, n5218, n847 );
nand U6895 ( n2017, n2018, n2002 );
nand U6896 ( n2214, n149, n1040 );
nor U6897 ( n1970, n1972, n1619 );
xor U6898 ( n3134, n3137, n3138 );
not U6899 ( n23, n1657 );
nand U6900 ( n780, n788, n790 );
nand U6901 ( n790, n791, n5238 );
nand U6902 ( n788, n5241, n792 );
nand U6903 ( n1425, n2104, n2105 );
nor U6904 ( n2105, n2106, n2107 );
nor U6905 ( n2104, n2116, n958 );
nor U6906 ( n2106, n318, n5199 );
not U6907 ( n310, n1108 );
nand U6908 ( n955, n956, n957 );
nand U6909 ( n957, n281, n5235 );
nand U6910 ( n956, n5231, n958 );
nand U6911 ( n914, n940, n941 );
nor U6912 ( n941, n942, n943 );
nor U6913 ( n940, n953, n955 );
nand U6914 ( n942, n948, n950 );
nor U6915 ( n1866, n1882, n1883 );
and U6916 ( n1883, n1682, n1660 );
nor U6917 ( n1882, n1885, n1886 );
nand U6918 ( n1886, n1887, n1888 );
nand U6919 ( n3228, n77, n3229 );
not U6920 ( n77, n3233 );
nand U6921 ( n3229, n3230, n3231 );
nand U6922 ( n3231, n3232, n5160 );
or U6923 ( n3170, n3064, n3066 );
nand U6924 ( n823, n825, n826 );
nand U6925 ( n826, n5203, n486 );
nand U6926 ( n825, n827, n5241 );
nand U6927 ( n3227, n3233, n3234 );
nand U6928 ( n3234, n3232, n3235 );
nand U6929 ( n3235, n5161, n3230 );
nor U6930 ( n4462, n3088, n5138 );
nand U6931 ( n1888, n1554, n1657 );
nand U6932 ( n1670, n1671, n1672 );
nand U6933 ( n1671, n817, n5223 );
nand U6934 ( n1672, n5219, n810 );
nand U6935 ( n1887, n105, n1657 );
nand U6936 ( n2665, n297, n169 );
nand U6937 ( n843, n845, n846 );
nand U6938 ( n845, n252, n5235 );
nand U6939 ( n846, n5243, n847 );
not U6940 ( n308, n1131 );
not U6941 ( n155, n2292 );
nor U6942 ( n2246, n3928, n4018 );
and U6943 ( n4018, n221, n2242 );
not U6944 ( n221, n2325 );
nand U6945 ( n2049, n2050, n2051 );
nand U6946 ( n2050, n937, n5223 );
nand U6947 ( n2051, n930, n5217 );
not U6948 ( n153, n2245 );
nor U6949 ( n2363, n2364, n2365 );
nand U6950 ( n2359, n308, n210 );
not U6951 ( n205, n2312 );
nand U6952 ( n2398, n307, n216 );
xor U6953 ( n3233, n3237, n3238 );
nor U6954 ( n2125, n2126, n2127 );
nor U6955 ( n2126, n139, n2058 );
not U6956 ( n139, n2092 );
nand U6957 ( n2526, n303, n200 );
nor U6958 ( n2479, n2486, n2487 );
nand U6959 ( n2486, n2485, n2491 );
nand U6960 ( n2487, n195, n2488 );
nand U6961 ( n2488, n2489, n2490 );
nand U6962 ( n743, n1494, n1495 );
nand U6963 ( n1495, n225, n1496 );
or U6964 ( n1494, n1496, n225 );
nand U6965 ( n1496, n1504, n1505 );
nor U6966 ( n1504, n227, n228 );
and U6967 ( n1987, n2112, n137 );
nor U6968 ( n2112, n281, n2113 );
and U6969 ( n1600, n1745, n1743 );
nor U6970 ( n1745, n247, n252 );
and U6971 ( n1859, n1989, n1987 );
nor U6972 ( n1989, n270, n275 );
and U6973 ( n1743, n1861, n1859 );
nor U6974 ( n1861, n258, n263 );
and U6975 ( n1505, n1602, n1600 );
nor U6976 ( n1602, n236, n240 );
nand U6977 ( n1391, n1490, n1491 );
nand U6978 ( n1491, n5185, n225 );
nor U6979 ( n1490, n61, n1492 );
nor U6980 ( n1492, n1493, n743 );
nand U6981 ( n2325, n222, n1108 );
nor U6982 ( n2483, n173, n2623 );
nand U6983 ( n2491, n301, n175 );
nand U6984 ( n2662, n298, n185 );
or U6985 ( n2114, n2127, n5099 );
and U6986 ( n5099, n20, n2092 );
nor U6987 ( n2473, n2475, n2476 );
nor U6988 ( n2476, n2477, n2478 );
nand U6989 ( n2472, n305, n196 );
nor U6990 ( n2362, n307, n216 );
nand U6991 ( n909, n960, n961 );
nor U6992 ( n961, n962, n963 );
nor U6993 ( n960, n973, n975 );
nand U6994 ( n962, n970, n971 );
nand U6995 ( n802, n807, n808 );
nand U6996 ( n807, n5209, n811 );
nand U6997 ( n808, n5243, n810 );
nand U6998 ( n1395, n1500, n1501 );
nand U6999 ( n1501, n227, n5185 );
nor U7000 ( n1500, n61, n1502 );
nor U7001 ( n1502, n1493, n753 );
nand U7002 ( n2151, n1879, n2143 );
nand U7003 ( n922, n927, n928 );
nand U7004 ( n927, n5208, n931 );
nand U7005 ( n928, n930, n5241 );
and U7006 ( n3419, n3420, n5168 );
xor U7007 ( n776, n1505, n228 );
nor U7008 ( n2475, n303, n200 );
not U7009 ( n301, n1260 );
xor U7010 ( n872, n1657, n1862 );
nand U7011 ( n1854, n1855, n1856 );
nand U7012 ( n1856, n871, n5223 );
nand U7013 ( n1855, n5218, n872 );
nand U7014 ( n2146, n137, n995 );
nand U7015 ( n4039, n4105, n4106 );
nor U7016 ( n4106, n172, n4107 );
nor U7017 ( n4105, n2615, n188 );
nand U7018 ( n4107, n2495, n4066 );
nor U7019 ( n4051, n2559, n197 );
nand U7020 ( n3879, n4021, n4022 );
nor U7021 ( n4021, n4116, n4117 );
nor U7022 ( n4022, n4023, n4024 );
nor U7023 ( n4117, n225, n331 );
nor U7024 ( n4062, n4063, n4064 );
nand U7025 ( n4064, n4065, n2416 );
nor U7026 ( n4063, n4039, n2614 );
nand U7027 ( n4065, n191, n4066 );
not U7028 ( n22, n1891 );
nand U7029 ( n772, n773, n775 );
nand U7030 ( n775, n228, n5235 );
or U7031 ( n773, n776, n742 );
nor U7032 ( n750, n742, n753 );
nand U7033 ( n2485, n302, n187 );
not U7034 ( n89, n3602 );
not U7035 ( n311, n1080 );
nand U7036 ( n862, n868, n870 );
nand U7037 ( n870, n871, n5239 );
nand U7038 ( n868, n5243, n872 );
nand U7039 ( n943, n945, n946 );
nand U7040 ( n946, n5203, n478 );
nand U7041 ( n945, n947, n5241 );
and U7042 ( n2303, n2322, n208 );
nor U7043 ( n2322, n2323, n2324 );
nand U7044 ( n2401, n2365, n2447 );
or U7045 ( n2447, n19, n2324 );
nand U7046 ( n879, n1095, n1096 );
nor U7047 ( n1096, n1097, n1099 );
nor U7048 ( n1095, n1109, n1111 );
nand U7049 ( n1097, n1105, n1107 );
not U7050 ( n312, n1063 );
nor U7051 ( n4444, n3328, n5138 );
xor U7052 ( n890, n1891, n1930 );
nand U7053 ( n1927, n1928, n1929 );
nand U7054 ( n1928, n897, n5223 );
nand U7055 ( n1929, n5218, n890 );
nand U7056 ( n904, n981, n983 );
nor U7057 ( n983, n984, n985 );
nor U7058 ( n981, n996, n997 );
nand U7059 ( n984, n991, n992 );
nand U7060 ( n4080, n4113, n4114 );
nor U7061 ( n4114, n276, n4115 );
nor U7062 ( n4113, n3928, n4074 );
nand U7063 ( n4115, n2099, n2214 );
nor U7064 ( n4069, n4070, n4071 );
nand U7065 ( n4071, n2002, n2099 );
nor U7066 ( n4070, n4015, n4072 );
nand U7067 ( n4072, n4073, n130 );
nand U7068 ( n2175, n145, n1017 );
nand U7069 ( n830, n831, n5239 );
nor U7070 ( n4014, n2216, n4074 );
nand U7071 ( n1093, n2344, n2345 );
nand U7072 ( n2345, n60, n1131 );
nor U7073 ( n2344, n2346, n2347 );
nor U7074 ( n2347, n218, n2348 );
nand U7075 ( n2351, n2330, n2356 );
nand U7076 ( n2356, n2357, n208 );
nor U7077 ( n2357, n2324, n19 );
nand U7078 ( n2382, n2397, n208 );
nor U7079 ( n2397, n2399, n2400 );
nor U7080 ( n2400, n210, n308 );
nor U7081 ( n2399, n2362, n2401 );
nor U7082 ( n2274, n2269, n2275 );
nor U7083 ( n2275, n2276, n2277 );
nor U7084 ( n2277, n103, n2024 );
nor U7085 ( n2276, n155, n2278 );
nand U7086 ( n2291, n2325, n2326 );
nand U7087 ( n2326, n2243, n2327 );
nand U7088 ( n2029, n2089, n2130 );
nand U7089 ( n2130, n316, n137 );
nor U7090 ( n2042, n2029, n2043 );
nand U7091 ( n2031, n2039, n2028 );
nand U7092 ( n2039, n2040, n2041 );
nand U7093 ( n2041, n275, n952 );
nor U7094 ( n2040, n140, n2042 );
nand U7095 ( n884, n1072, n1073 );
nor U7096 ( n1073, n1075, n1076 );
nor U7097 ( n1072, n1087, n1088 );
nand U7098 ( n1076, n1077, n1079 );
nor U7099 ( n4077, n4082, n128 );
nor U7100 ( n4082, n3998, n211 );
not U7101 ( n128, n4083 );
not U7102 ( n211, n2369 );
nand U7103 ( n894, n1027, n1028 );
nor U7104 ( n1028, n1029, n1031 );
nor U7105 ( n1027, n1041, n1043 );
nand U7106 ( n1029, n1036, n1037 );
nand U7107 ( n2200, n2208, n2186 );
nand U7108 ( n2208, n2027, n2043 );
nor U7109 ( n3970, n3971, n3972 );
nor U7110 ( n3972, n267, n2002 );
nor U7111 ( n3971, n3973, n3974 );
nor U7112 ( n3973, n3975, n3976 );
nand U7113 ( n4033, n183, n2610 );
nor U7114 ( n3946, n3955, n3956 );
nand U7115 ( n3956, n3954, n3957 );
nand U7116 ( n3955, n3962, n3963 );
nand U7117 ( n3957, n327, n3953 );
nand U7118 ( n3963, n3964, n1796 );
nand U7119 ( n3964, n3965, n3966 );
nand U7120 ( n3966, n261, n3902 );
nor U7121 ( n3965, n255, n3967 );
nand U7122 ( n3889, n3935, n3936 );
nor U7123 ( n3936, n3937, n3938 );
nor U7124 ( n3935, n3946, n3947 );
nand U7125 ( n3938, n3939, n3940 );
nand U7126 ( n3980, n3981, n3982 );
nor U7127 ( n3982, n172, n2615 );
nor U7128 ( n3981, n3983, n3984 );
nor U7129 ( n3984, n3985, n2719 );
not U7130 ( n276, n2002 );
nand U7131 ( n2057, n2089, n2090 );
nand U7132 ( n2090, n2091, n2092 );
nand U7133 ( n2091, n281, n972 );
nand U7134 ( n3262, n3635, n3636 );
nand U7135 ( n3636, n5114, n275 );
nand U7136 ( n3635, n5162, n952 );
and U7137 ( n3431, n3637, n3638 );
nand U7138 ( n3638, n5115, n281 );
nand U7139 ( n3637, n5162, n972 );
nand U7140 ( n1982, n1983, n1984 );
nand U7141 ( n1983, n5218, n912 );
nand U7142 ( n1984, n911, n5223 );
nand U7143 ( n1025, n2233, n2234 );
nand U7144 ( n2234, n60, n1063 );
nor U7145 ( n2233, n2235, n2236 );
nor U7146 ( n2236, n95, n2237 );
or U7147 ( n2230, n5100, n5101 );
nand U7148 ( n5100, n148, n2220 );
nor U7149 ( n5101, n2024, n154 );
nand U7150 ( n2231, n2249, n2250 );
nor U7151 ( n2249, n2238, n154 );
nand U7152 ( n2250, n2251, n2024 );
nand U7153 ( n1797, n322, n258 );
and U7154 ( n4036, n4110, n1786 );
nor U7155 ( n4110, n248, n4111 );
nor U7156 ( n4111, n255, n3901 );
nand U7157 ( n882, n887, n888 );
nand U7158 ( n887, n5208, n891 );
nand U7159 ( n888, n5243, n890 );
nand U7160 ( n899, n1004, n1005 );
nor U7161 ( n1005, n1007, n1008 );
nor U7162 ( n1004, n1019, n1020 );
nand U7163 ( n1007, n1015, n1016 );
nand U7164 ( n2192, n2193, n2194 );
nand U7165 ( n2194, n993, n5223 );
nand U7166 ( n2193, n5218, n989 );
nand U7167 ( n4015, n4076, n2143 );
or U7168 ( n4076, n2177, n133 );
nand U7169 ( n1907, n270, n320 );
nand U7170 ( n874, n1117, n1119 );
nor U7171 ( n1119, n1120, n1121 );
nor U7172 ( n1117, n1132, n1133 );
nand U7173 ( n1120, n1127, n1128 );
nor U7174 ( n3998, n2411, n206 );
xor U7175 ( n3354, n3359, n89 );
nand U7176 ( n3974, n3996, n3997 );
nor U7177 ( n3997, n3998, n3999 );
nor U7178 ( n3996, n4000, n4001 );
nand U7179 ( n3999, n2243, n2369 );
not U7180 ( n313, n1040 );
nor U7181 ( n4079, n4081, n155 );
nor U7182 ( n4081, n157, n2243 );
nor U7183 ( n3877, n3818, n3879 );
nor U7184 ( n2033, n2037, n2029 );
nor U7185 ( n2037, n154, n2038 );
nor U7186 ( n2038, n149, n313 );
nand U7187 ( n2012, n275, n318 );
nor U7188 ( n2023, n5102, n5103 );
or U7189 ( n5102, n2029, n2030 );
nand U7190 ( n5103, n2027, n2028 );
nand U7191 ( n1903, n263, n321 );
nand U7192 ( n1071, n2306, n2307 );
nand U7193 ( n2307, n60, n1108 );
nor U7194 ( n2306, n2308, n2309 );
nor U7195 ( n2309, n156, n2310 );
nand U7196 ( n889, n1049, n1051 );
nor U7197 ( n1051, n1052, n1053 );
nor U7198 ( n1049, n1064, n1065 );
nand U7199 ( n1052, n1059, n1060 );
nand U7200 ( n2268, n2281, n2024 );
nand U7201 ( n2281, n2254, n2251 );
not U7202 ( n35, n2113 );
nor U7203 ( n951, n1987, n2110 );
and U7204 ( n2110, n281, n2111 );
nand U7205 ( n2111, n137, n35 );
nand U7206 ( n2336, n2337, n2338 );
nand U7207 ( n2338, n1084, n5223 );
nand U7208 ( n2337, n5218, n1085 );
nor U7209 ( n2310, n2311, n2280 );
nor U7210 ( n2311, n2312, n2313 );
nor U7211 ( n2313, n2314, n2315 );
nor U7212 ( n2314, n2303, n103 );
nand U7213 ( n2036, n313, n149 );
nand U7214 ( n902, n908, n910 );
nand U7215 ( n908, n5242, n912 );
nand U7216 ( n910, n911, n5239 );
nand U7217 ( n2027, n315, n145 );
and U7218 ( n2034, n2028, n5104 );
and U7219 ( n5104, n2036, n2027 );
nand U7220 ( n2251, n312, n152 );
nand U7221 ( n2101, n281, n317 );
nand U7222 ( n2422, n2423, n2424 );
nand U7223 ( n2424, n1129, n5223 );
nand U7224 ( n2423, n5217, n1125 );
not U7225 ( n154, n2254 );
nand U7226 ( n2527, n2478, n2550 );
nand U7227 ( n2550, n2551, n2485 );
nand U7228 ( n2551, n2589, n2489 );
nor U7229 ( n2589, n2590, n2591 );
nor U7230 ( n2591, n173, n2490 );
and U7231 ( n2590, n2484, n2483 );
nand U7232 ( n4085, n4086, n4087 );
nand U7233 ( n4087, n2685, n4088 );
nand U7234 ( n4088, n4089, n2683 );
nand U7235 ( n4089, n2722, n4090 );
nand U7236 ( n1916, n2099, n2100 );
nand U7237 ( n2100, n133, n2101 );
nand U7238 ( n1906, n2002, n2015 );
nand U7239 ( n2015, n2012, n1916 );
nand U7240 ( n2514, n2528, n195 );
nor U7241 ( n2528, n2529, n2530 );
nor U7242 ( n2530, n196, n305 );
nor U7243 ( n2529, n2475, n2527 );
nand U7244 ( n1035, n2267, n2268 );
or U7245 ( n2267, n2024, n2269 );
nand U7246 ( n2260, n2261, n2262 );
nand U7247 ( n2262, n1039, n5223 );
nand U7248 ( n2261, n5218, n1035 );
nand U7249 ( n864, n1163, n1164 );
nor U7250 ( n1164, n1165, n1167 );
nor U7251 ( n1163, n1177, n1179 );
nand U7252 ( n1165, n1172, n1173 );
not U7253 ( n181, n2610 );
not U7254 ( n315, n1017 );
xor U7255 ( n979, n35, n137 );
not U7256 ( n5163, n5089 );
nor U7257 ( n4426, n3530, n5138 );
nor U7258 ( n4004, n162, n4006 );
not U7259 ( n162, n2722 );
nor U7260 ( n4006, n4007, n165 );
nor U7261 ( n4007, n37, n164 );
nand U7262 ( n869, n1140, n1141 );
nor U7263 ( n1141, n1143, n1144 );
nor U7264 ( n1140, n1155, n1156 );
nand U7265 ( n1143, n1149, n1151 );
not U7266 ( n126, n2143 );
nand U7267 ( n1075, n1081, n1083 );
nand U7268 ( n1083, n1084, n5238 );
nand U7269 ( n1081, n5242, n1085 );
not U7270 ( n248, n1721 );
nor U7271 ( n2286, n2288, n2289 );
nand U7272 ( n2288, n2247, n2142 );
nand U7273 ( n2289, n2269, n2290 );
nand U7274 ( n2290, n2291, n2292 );
nand U7275 ( n2507, n2508, n2509 );
nand U7276 ( n2509, n1175, n5223 );
nand U7277 ( n2508, n5217, n1171 );
not U7278 ( n34, n2198 );
nand U7279 ( n859, n1185, n1186 );
nor U7280 ( n1186, n1188, n1189 );
nor U7281 ( n1185, n1199, n1200 );
nand U7282 ( n1188, n1194, n1195 );
and U7283 ( n1786, n3902, n1796 );
nand U7284 ( n3195, n236, n5156 );
not U7285 ( n186, n2614 );
xor U7286 ( n1024, n34, n149 );
not U7287 ( n271, n1948 );
nand U7288 ( n992, n993, n5238 );
not U7289 ( n316, n995 );
buf U7290 ( n5152, n5151 );
nand U7291 ( n2439, n2448, n2416 );
nand U7292 ( n2448, n192, n2449 );
not U7293 ( n192, n2415 );
nand U7294 ( n2449, n40, n2410 );
and U7295 ( n1904, n3901, n1948 );
not U7296 ( n317, n972 );
buf U7297 ( n5148, n5147 );
nor U7298 ( n4052, n197, n2556 );
not U7299 ( n33, n2266 );
nor U7300 ( n4023, n3922, n4095 );
nand U7301 ( n4095, n4086, n4038 );
not U7302 ( n15, n2484 );
nor U7303 ( n2621, n182, n2622 );
nor U7304 ( n2622, n2623, n15 );
not U7305 ( n190, n2556 );
not U7306 ( n322, n891 );
not U7307 ( n176, n2581 );
nand U7308 ( n849, n1228, n1229 );
nor U7309 ( n1229, n1230, n1231 );
nor U7310 ( n1228, n1240, n1241 );
nand U7311 ( n1230, n1236, n1238 );
not U7312 ( n164, n2749 );
nand U7313 ( n4019, n157, n2245 );
nand U7314 ( n742, n1374, n5230 );
nand U7315 ( n756, n116, n1384 );
nand U7316 ( n1384, n1385, n1377 );
nand U7317 ( n1385, n1386, n286 );
nor U7318 ( n1386, n1387, n1388 );
not U7319 ( n102, n1493 );
nand U7320 ( n1209, n1215, n1216 );
nand U7321 ( n1215, n5242, n1219 );
nand U7322 ( n1216, n1218, n5238 );
nand U7323 ( n1291, n1299, n1300 );
nand U7324 ( n1299, n5207, n1303 );
nand U7325 ( n1300, n1301, n5238 );
nand U7326 ( n1037, n1039, n5238 );
nand U7327 ( n1128, n1129, n5238 );
nand U7328 ( n1173, n1175, n5238 );
nand U7329 ( n1250, n1256, n1258 );
nand U7330 ( n1256, n5207, n1260 );
nand U7331 ( n1258, n1259, n5238 );
nand U7332 ( n1334, n1339, n1340 );
nand U7333 ( n1339, n5207, n1342 );
nand U7334 ( n1340, n1341, n5238 );
nand U7335 ( n839, n1269, n1270 );
nor U7336 ( n1270, n1271, n1273 );
nor U7337 ( n1269, n1281, n1283 );
nand U7338 ( n1271, n1278, n1279 );
nand U7339 ( n805, n240, n5235 );
nand U7340 ( n925, n275, n5235 );
nand U7341 ( n885, n263, n5235 );
not U7342 ( n320, n931 );
nand U7343 ( n829, n1311, n1313 );
nor U7344 ( n1313, n1314, n1315 );
nor U7345 ( n1311, n1325, n1326 );
nand U7346 ( n1314, n1321, n1323 );
not U7347 ( n318, n952 );
nor U7348 ( n2496, n2498, n2499 );
nand U7349 ( n2498, n2495, n2142 );
nand U7350 ( n2499, n2461, n2500 );
nand U7351 ( n2500, n2501, n2452 );
nor U7352 ( n2625, n182, n2484 );
not U7353 ( n321, n907 );
xor U7354 ( n1069, n33, n158 );
buf U7355 ( n5139, n5136 );
not U7356 ( n32, n2342 );
not U7357 ( n346, n4881 );
nand U7358 ( n2565, n2566, n2567 );
nand U7359 ( n2567, n1218, n5223 );
nand U7360 ( n2566, n5217, n1219 );
not U7361 ( n260, n3902 );
nand U7362 ( n1646, n240, n326 );
nor U7363 ( n4116, n4101, n4118 );
nor U7364 ( n4118, n4119, n4120 );
nor U7365 ( n4119, n4103, n4121 );
nor U7366 ( n4121, n4122, n4123 );
nor U7367 ( n1909, n1910, n1911 );
nor U7368 ( n1911, n1625, n1838 );
nor U7369 ( n1910, n132, n111 );
not U7370 ( n237, n1587 );
nand U7371 ( n1255, n2656, n2657 );
nand U7372 ( n2657, n2658, n2484 );
nand U7373 ( n2656, n15, n180 );
or U7374 ( n2658, n182, n2623 );
nor U7375 ( n4102, n328, n228 );
nand U7376 ( n4041, n4099, n4100 );
nor U7377 ( n4100, n241, n4101 );
nor U7378 ( n4099, n4102, n4103 );
not U7379 ( n241, n1650 );
nand U7380 ( n3479, n3587, n3588 );
nand U7381 ( n3588, n5114, n270 );
nand U7382 ( n3587, n5163, n931 );
nor U7383 ( n4010, n1919, n2099 );
buf U7384 ( n5144, n4314 );
nand U7385 ( n1588, n236, n327 );
nand U7386 ( n1792, n252, n323 );
xor U7387 ( n1115, n32, n210 );
nand U7388 ( n1784, n1795, n1796 );
nand U7389 ( n1795, n1797, n1792 );
nand U7390 ( n3564, n3654, n3655 );
nand U7391 ( n3655, n5115, n247 );
nand U7392 ( n3654, n5162, n851 );
nand U7393 ( n1681, n252, n867 );
nand U7394 ( n1663, n1678, n1729 );
nand U7395 ( n1729, n1680, n1681 );
nand U7396 ( n4029, n4032, n4033 );
and U7397 ( n4032, n3921, n1948 );
nand U7398 ( n1680, n247, n851 );
nand U7399 ( n1649, n247, n325 );
nand U7400 ( n1682, n258, n891 );
nand U7401 ( n3299, n3571, n3572 );
nand U7402 ( n3572, n5114, n252 );
nand U7403 ( n3571, n5163, n867 );
not U7404 ( n31, n2428 );
nand U7405 ( n2632, n2633, n2634 );
nand U7406 ( n2634, n1259, n5223 );
nand U7407 ( n2633, n5217, n1255 );
not U7408 ( n287, n2836 );
and U7409 ( n1659, n1678, n1764 );
nor U7410 ( n2692, n2694, n2695 );
nor U7411 ( n2695, n185, n298 );
nor U7412 ( n2694, n170, n2666 );
nand U7413 ( n2648, n2683, n2684 );
nand U7414 ( n2684, n2685, n2616 );
nor U7415 ( n2642, n2650, n2651 );
nand U7416 ( n2651, n180, n2614 );
nor U7417 ( n2650, n2652, n38 );
nor U7418 ( n2652, n95, n2649 );
nand U7419 ( n3190, n3576, n3577 );
nand U7420 ( n3577, n5114, n258 );
nand U7421 ( n3576, n5163, n891 );
nand U7422 ( n3895, n3905, n3906 );
nor U7423 ( n3905, n3910, n3911 );
nor U7424 ( n3906, n3907, n3908 );
nand U7425 ( n3910, n233, n3912 );
xor U7426 ( n1160, n31, n202 );
nand U7427 ( n3099, n3582, n3583 );
nand U7428 ( n3583, n5114, n263 );
nand U7429 ( n3582, n5163, n907 );
nand U7430 ( n2645, n2646, n2647 );
nand U7431 ( n2647, n2648, n2614 );
and U7432 ( n1636, n1650, n1651 );
nand U7433 ( n1651, n248, n1646 );
nand U7434 ( n2301, n2247, n2292 );
or U7435 ( n5105, n1377, n756 );
nand U7436 ( n2746, n2719, n2722 );
nand U7437 ( n2054, n2002, n2012 );
nand U7438 ( n1673, n1650, n1646 );
not U7439 ( n30, n2513 );
nand U7440 ( n926, n5203, n480 );
nand U7441 ( n886, n5203, n482 );
nand U7442 ( n2238, n2216, n2214 );
and U7443 ( n1656, n1658, n1659 );
and U7444 ( n1658, n1660, n1605 );
nand U7445 ( n1990, n1907, n1948 );
nand U7446 ( n1210, n1211, n1213 );
nand U7447 ( n1213, n5207, n1214 );
nand U7448 ( n1211, n5202, n493 );
nand U7449 ( n905, n5203, n481 );
nand U7450 ( n865, n5203, n483 );
nand U7451 ( n1015, n5203, n475 );
nand U7452 ( n970, n5203, n477 );
nand U7453 ( n848, n5203, n485 );
nand U7454 ( n1105, n5202, n500 );
nand U7455 ( n1236, n5202, n492 );
nand U7456 ( n1278, n5202, n512 );
nand U7457 ( n2389, n2369, n2366 );
nand U7458 ( n2171, n2143, n2146 );
nand U7459 ( n1811, n1796, n1792 );
nand U7460 ( n2432, n2411, n2414 );
nand U7461 ( n1930, n1903, n3901 );
nand U7462 ( n1862, n3902, n1797 );
nand U7463 ( n806, n5203, n487 );
nand U7464 ( n782, n5202, n488 );
nand U7465 ( n2353, n2243, n2325 );
nor U7466 ( n2646, n2615, n181 );
nand U7467 ( n1310, n2709, n2710 );
nand U7468 ( n2710, n60, n1342 );
nor U7469 ( n2709, n2711, n2712 );
nor U7470 ( n2711, n95, n2718 );
and U7471 ( n2713, n2663, n2665 );
and U7472 ( n3959, n3960, n3961 );
nand U7473 ( n3961, n227, n3942 );
and U7474 ( n3954, n1646, n3958 );
nand U7475 ( n3958, n3945, n3943 );
nor U7476 ( n2579, n2559, n190 );
nand U7477 ( n1382, n2804, n3923 );
nand U7478 ( n2150, n2101, n2099 );
nand U7479 ( n3945, n3959, n786 );
nand U7480 ( n3923, n36, n2798 );
nor U7481 ( n2269, n3928, n153 );
nand U7482 ( n1629, n1587, n1588 );
nand U7483 ( n4030, n3923, n4031 );
nand U7484 ( n4031, n106, n2804 );
nand U7485 ( n1777, n1721, n1649 );
and U7486 ( n2201, n2175, n2177 );
nand U7487 ( n1603, n240, n832 );
and U7488 ( n2805, n3921, n3922 );
xor U7489 ( n1204, n30, n200 );
nand U7490 ( n3947, n3948, n3949 );
nand U7491 ( n3948, n3950, n3951 );
nand U7492 ( n3950, n1650, n1721 );
nand U7493 ( n3951, n3952, n3953 );
nand U7494 ( n3952, n3954, n811 );
not U7495 ( n29, n2571 );
not U7496 ( n326, n832 );
nand U7497 ( n2701, n2702, n2703 );
nand U7498 ( n2703, n1301, n5223 );
nand U7499 ( n2702, n5217, n1298 );
nand U7500 ( n1331, n2732, n2733 );
nand U7501 ( n2733, n60, n1359 );
nor U7502 ( n2732, n2734, n2735 );
and U7503 ( n2735, n2441, n1319 );
nand U7504 ( n2820, n4910, n118 );
nor U7505 ( n4910, n5123, n282 );
not U7506 ( n231, n1523 );
nand U7507 ( n1319, n2736, n2737 );
or U7508 ( n2736, n2716, n160 );
nand U7509 ( n2737, n2738, n2716 );
nand U7510 ( n2738, n2717, n2714 );
not U7511 ( n327, n811 );
nand U7512 ( n1522, n236, n811 );
not U7513 ( n325, n851 );
nand U7514 ( n1548, n1556, n1557 );
nand U7515 ( n1557, n238, n1523 );
nand U7516 ( n1556, n235, n231 );
nand U7517 ( n2129, n280, n2092 );
not U7518 ( n323, n867 );
xor U7519 ( n1245, n29, n175 );
not U7520 ( n328, n786 );
nand U7521 ( n2752, n2746, n2749 );
nand U7522 ( n2147, n2148, n2146 );
nand U7523 ( n2148, n111, n1625 );
nor U7524 ( n1387, n121, n3806 );
nand U7525 ( n3066, n3172, n3173 );
nand U7526 ( n3173, n5114, n240 );
nand U7527 ( n3172, n5163, n832 );
not U7528 ( n28, n2638 );
not U7529 ( n238, n1520 );
nand U7530 ( n2758, n2759, n2760 );
nand U7531 ( n2760, n1341, n5223 );
nand U7532 ( n2759, n5217, n11 );
nand U7533 ( n1571, n1523, n1587 );
nor U7534 ( n3937, n3944, n1587 );
and U7535 ( n3944, n3943, n3945 );
nor U7536 ( n1547, n1523, n238 );
and U7537 ( n1568, n1582, n1583 );
nand U7538 ( n1582, n232, n1523 );
nand U7539 ( n1583, n237, n231 );
or U7540 ( n3939, n3943, n328 );
not U7541 ( n182, n2490 );
nor U7542 ( n2626, n175, n301 );
not U7543 ( n170, n2663 );
nand U7544 ( n2835, n288, n333 );
xor U7545 ( n1286, n28, n185 );
nand U7546 ( n2170, n2092, n2130 );
not U7547 ( n253, n1764 );
nor U7548 ( n2800, n95, n2803 );
xnor U7549 ( n2803, n2804, n2805 );
nand U7550 ( n1365, n2796, n2797 );
nand U7551 ( n2797, n60, n2798 );
nor U7552 ( n2796, n2800, n2801 );
and U7553 ( n2801, n2441, n1355 );
nand U7554 ( n2773, n2742, n2739 );
not U7555 ( n27, n2707 );
xnor U7556 ( n1355, n2802, n2785 );
nand U7557 ( n2802, n2783, n2786 );
not U7558 ( n59, n4593 );
nand U7559 ( n4835, n4907, n4908 );
nand U7560 ( n4907, n4911, n4909 );
nand U7561 ( n4908, n116, n4909 );
nor U7562 ( n4911, n5123, n118 );
not U7563 ( n5143, n4315 );
nand U7564 ( n4315, n4693, n118 );
nor U7565 ( n4693, n5123, n4305 );
nand U7566 ( n3949, n331, n225 );
xor U7567 ( n1330, n27, n161 );
nand U7568 ( n588, n290, n4835 );
nand U7569 ( n4589, n4303, n4835 );
nand U7570 ( n3243, n116, n3823 );
nand U7571 ( n3823, n1377, n3824 );
nand U7572 ( n3824, n3794, n5185 );
and U7573 ( n5106, n92, n114 );
nand U7574 ( n3200, n3201, n3202 );
nand U7575 ( n3202, n488, n3072 );
nand U7576 ( n3201, n5225, n236 );
nand U7577 ( n3374, n3375, n3376 );
nand U7578 ( n3376, n483, n3072 );
nand U7579 ( n3375, n5226, n258 );
nand U7580 ( n3481, n3482, n3483 );
nand U7581 ( n3483, n481, n3072 );
nand U7582 ( n3482, n5226, n270 );
nand U7583 ( n3439, n3440, n3441 );
nand U7584 ( n3441, n478, n3072 );
nand U7585 ( n3440, n5226, n281 );
nand U7586 ( n3305, n3306, n3307 );
nand U7587 ( n3307, n485, n3072 );
nand U7588 ( n3306, n5225, n252 );
nand U7589 ( n3265, n3266, n3267 );
nand U7590 ( n3267, n480, n3072 );
nand U7591 ( n3266, n5225, n275 );
nand U7592 ( n3069, n3070, n3071 );
nand U7593 ( n3071, n487, n3072 );
nand U7594 ( n3070, n5225, n240 );
nand U7595 ( n3101, n3102, n3103 );
nand U7596 ( n3103, n482, n3072 );
nand U7597 ( n3102, n5225, n263 );
nand U7598 ( n3657, n3658, n3659 );
nand U7599 ( n3659, n486, n3072 );
nand U7600 ( n3658, n5227, n247 );
nor U7601 ( n2814, n10, n1516 );
nand U7602 ( n1485, n2808, n2809 );
nor U7603 ( n2809, n1383, n2810 );
nor U7604 ( n2808, n2813, n2814 );
nor U7605 ( n2810, n36, n2811 );
xor U7606 ( n1364, n163, n36 );
nand U7607 ( n1279, n5207, n1280 );
nand U7608 ( n1323, n5207, n1324 );
nand U7609 ( n1107, n5208, n1108 );
nand U7610 ( n906, n5208, n907 );
nand U7611 ( n1079, n5208, n1080 );
nand U7612 ( n1016, n5208, n1017 );
nand U7613 ( n971, n5208, n972 );
nand U7614 ( n1358, n5207, n1359 );
nand U7615 ( n1238, n5207, n1239 );
nand U7616 ( n1172, n5207, n1176 );
nand U7617 ( n1127, n5208, n1131 );
nand U7618 ( n1059, n5208, n1063 );
and U7619 ( n5107, n1486, n286 );
nand U7620 ( n1036, n5208, n1040 );
nand U7621 ( n948, n5208, n952 );
nand U7622 ( n1149, n5207, n1153 );
nand U7623 ( n991, n5208, n995 );
nand U7624 ( n1194, n5207, n1198 );
nand U7625 ( n866, n5209, n867 );
nand U7626 ( n783, n5209, n786 );
nand U7627 ( n850, n5209, n851 );
nand U7628 ( n828, n5209, n832 );
nor U7629 ( n4794, n337, n588 );
nor U7630 ( n4781, n338, n588 );
nor U7631 ( n4769, n341, n588 );
nor U7632 ( n4744, n345, n588 );
nor U7633 ( n4731, n343, n588 );
nor U7634 ( n652, n122, n588 );
nor U7635 ( n633, n146, n588 );
nor U7636 ( n576, n159, n588 );
nand U7637 ( n1941, n97, n1625 );
nor U7638 ( n2544, n200, n5183 );
nor U7639 ( n2676, n185, n5183 );
not U7640 ( n5244, n4978 );
nor U7641 ( n2843, n2846, n5173 );
nor U7642 ( n2863, n2865, n5173 );
nor U7643 ( n2882, n2884, n5173 );
nor U7644 ( n2907, n2909, n5173 );
nor U7645 ( n2919, n2921, n5173 );
nor U7646 ( n2931, n2933, n5173 );
nor U7647 ( n2943, n2945, n5173 );
nor U7648 ( n2955, n2957, n5173 );
nor U7649 ( n2601, n175, n5183 );
nor U7650 ( n2462, n202, n5183 );
nor U7651 ( n2991, n2993, n5172 );
nor U7652 ( n3007, n3009, n5173 );
nor U7653 ( n2967, n2969, n5172 );
nor U7654 ( n2979, n2981, n5173 );
nor U7655 ( n3001, n5172, n3003 );
or U7656 ( n3003, n3004, n346 );
nor U7657 ( n2202, n145, n5182 );
nor U7658 ( n2516, n196, n5183 );
and U7659 ( n5108, n116, n2836 );
nor U7660 ( n2731, n161, n5182 );
nor U7661 ( n2232, n149, n5183 );
nor U7662 ( n2384, n210, n5183 );
nor U7663 ( n2795, n163, n5183 );
nor U7664 ( n2270, n152, n5183 );
nor U7665 ( n2765, n166, n5182 );
not U7666 ( n56, n4909 );
nor U7667 ( n2572, n187, n5183 );
nor U7668 ( n2305, n158, n5183 );
nor U7669 ( n2433, n216, n5183 );
nor U7670 ( n2639, n177, n5183 );
nor U7671 ( n2343, n222, n5183 );
nor U7672 ( n2161, n137, n5182 );
nor U7673 ( n2708, n169, n5183 );
nand U7674 ( n2822, n2823, n2824 );
buf U7675 ( n5123, n5245 );
nor U7676 ( n3794, n1388, n286 );
nand U7677 ( n3240, n3796, n3797 );
nor U7678 ( n3796, n290, n283 );
nor U7679 ( n3242, n163, n3243 );
nor U7680 ( n3515, n166, n3243 );
not U7681 ( n61, n757 );
nor U7682 ( n3418, n36, n3243 );
not U7683 ( n112, n1625 );
and U7684 ( n3035, n3793, n3794 );
nor U7685 ( n3793, n3795, n2820 );
not U7686 ( n62, n3806 );
nand U7687 ( n1376, n62, n290 );
buf U7688 ( n5167, n5164 );
nor U7689 ( n745, n756, n757 );
nand U7690 ( n1620, n109, n114 );
not U7691 ( n109, n4304 );
nand U7692 ( n1549, n3814, n106 );
nand U7693 ( n3055, n3802, n3803 );
nand U7694 ( n3803, n3663, n5244 );
and U7695 ( n3802, n3417, n3416 );
nor U7696 ( n2588, n301, n5134 );
nand U7697 ( n3156, n477, n3055 );
nand U7698 ( n3362, n475, n3055 );
nand U7699 ( n3467, n500, n3055 );
nand U7700 ( n3801, n491, n3055 );
nand U7701 ( n3407, n495, n3055 );
nand U7702 ( n3054, n492, n3055 );
nand U7703 ( n3498, n497, n3055 );
nand U7704 ( n3343, n512, n3055 );
not U7705 ( n63, n3663 );
and U7706 ( n3797, n3820, n109 );
nor U7707 ( n3820, n114, n2820 );
nand U7708 ( n1337, n3025, n3026 );
nand U7709 ( n3026, n3027, n5187 );
nor U7710 ( n3027, n282, n62 );
and U7711 ( n3019, n3021, n5175 );
and U7712 ( n2996, n2998, n5175 );
not U7713 ( n113, n1516 );
not U7714 ( n99, n1619 );
not U7715 ( n60, n1732 );
buf U7716 ( n5133, n1732 );
buf U7717 ( n5132, n1732 );
buf U7718 ( n5129, n5125 );
buf U7719 ( n5127, n5125 );
buf U7720 ( n5126, n5125 );
buf U7721 ( n5131, n5125 );
buf U7722 ( n5130, n5125 );
buf U7723 ( n5128, n5125 );
buf U7724 ( n5135, n1732 );
buf U7725 ( n5134, n1732 );
nand U7726 ( n4302, n109, n4303 );
not U7727 ( n476, n3530 );
not U7728 ( n473, n3328 );
buf U7729 ( n5124, n5245 );
not U7730 ( n501, n3088 );
not U7731 ( n498, n3288 );
not U7732 ( n496, n3120 );
not U7733 ( n493, n3219 );
not U7734 ( n502, n3551 );
nand U7735 ( n1619, n4671, n695 );
not U7736 ( n106, n2825 );
nand U7737 ( n2928, n4951, n151 );
nand U7738 ( n4668, n4658, n695 );
nand U7739 ( n4667, n4305, n4669 );
nand U7740 ( n4881, n4888, n4980 );
nor U7741 ( n3744, n3236, n3749 );
nand U7742 ( n3749, n3750, n76 );
nand U7743 ( n3750, n8, n5161 );
not U7744 ( n76, n3746 );
not U7745 ( n342, n2988 );
not U7746 ( n340, n2976 );
not U7747 ( n335, n2952 );
not U7748 ( n120, n2916 );
not U7749 ( n151, n2940 );
not U7750 ( n336, n2964 );
not U7751 ( n143, n2816 );
xor U7752 ( n2909, n2916, n4985 );
nand U7753 ( n1322, n3057, n3058 );
nor U7754 ( n3057, n3068, n3069 );
nor U7755 ( n3058, n3059, n3060 );
nor U7756 ( n3068, STATE_REG, n4977 );
nand U7757 ( n1267, n3289, n3290 );
nor U7758 ( n3289, n3304, n3305 );
nor U7759 ( n3290, n3291, n3292 );
nor U7760 ( n3304, STATE_REG, n4976 );
not U7761 ( n122, n695 );
nand U7762 ( n3818, n143, n2826 );
nor U7763 ( n3814, n3818, n695 );
nand U7764 ( n2824, n106, n2816 );
nand U7765 ( n4305, n4923, n3871 );
nor U7766 ( n4923, n333, n3829 );
nor U7767 ( n4658, n2825, n282 );
nand U7768 ( n4278, n335, n4982 );
nand U7769 ( n4933, n4944, n4945 );
nor U7770 ( n4945, n4946, n4947 );
nor U7771 ( n4944, n4950, n4278 );
nand U7772 ( n4947, n4948, n4981 );
nand U7773 ( n2879, n4940, n291 );
xor U7774 ( n2884, n4933, n4986 );
not U7775 ( n333, n3868 );
nand U7776 ( n1312, n3089, n3090 );
nor U7777 ( n3089, n3100, n3101 );
nor U7778 ( n3090, n3091, n3092 );
nor U7779 ( n3100, STATE_REG, n4975 );
nand U7780 ( n1277, n3244, n3245 );
nor U7781 ( n3244, n3264, n3265 );
nor U7782 ( n3245, n3246, n3247 );
nor U7783 ( n3264, STATE_REG, n5041 );
buf U7784 ( n5216, n5211 );
buf U7785 ( n5211, n5212 );
nand U7786 ( n4950, n4951, n4984 );
xnor U7787 ( n3048, n3711, n5161 );
nand U7788 ( n3711, n3712, n3713 );
nand U7789 ( n3712, n5115, n1260 );
nand U7790 ( n3713, n5156, n1235 );
nand U7791 ( n4304, n121, n2825 );
not U7792 ( n163, n1356 );
xor U7793 ( n2865, n2872, n4987 );
and U7794 ( n5109, n4650, n290 );
not U7795 ( n290, n2799 );
nand U7796 ( n3237, n3754, n3755 );
nand U7797 ( n3755, n5116, n1356 );
nand U7798 ( n3754, n5162, n1375 );
not U7799 ( n5161, n3175 );
nand U7800 ( n3175, n4684, n4685 );
nand U7801 ( n4685, n2816, n2825 );
not U7802 ( n36, n1373 );
not U7803 ( n8, n3748 );
nand U7804 ( n3817, n122, n2826 );
nand U7805 ( n3747, n3748, n5160 );
nand U7806 ( n3511, n3740, n3741 );
nand U7807 ( n3741, n5116, n1347 );
nand U7808 ( n3740, n5162, n1359 );
not U7809 ( n166, n1347 );
not U7810 ( n161, n1320 );
nand U7811 ( n3137, n3756, n3757 );
nand U7812 ( n3757, n5116, n1320 );
nand U7813 ( n3756, n5162, n1342 );
xor U7814 ( n2846, n4988, n2840 );
nand U7815 ( n4313, n332, n4676 );
nand U7816 ( n1375, n4573, n4574 );
nor U7817 ( n4574, n4575, n4576 );
nor U7818 ( n4573, n4577, n4578 );
nor U7819 ( n4575, n4991, n5146 );
nor U7820 ( n4577, n4992, n5150 );
not U7821 ( n332, n4677 );
nor U7822 ( n4576, n5137, n4966 );
nand U7823 ( n4328, n4676, n4677 );
nor U7824 ( n4251, n4252, n1309 );
nor U7825 ( n4252, n1324, n4249 );
nor U7826 ( n4141, n4143, n4144 );
nor U7827 ( n4143, n851, n1766 );
nand U7828 ( n4144, n1792, n4145 );
nand U7829 ( n4145, n4146, n1796 );
nor U7830 ( n4158, n4159, n4160 );
nor U7831 ( n4160, n281, n317 );
nor U7832 ( n4159, n4161, n4162 );
nor U7833 ( n4161, n972, n2134 );
nor U7834 ( n4153, n4155, n4156 );
nor U7835 ( n4155, n931, n1960 );
nand U7836 ( n4156, n2012, n4157 );
nand U7837 ( n4157, n4158, n2002 );
nor U7838 ( n4146, n4147, n4148 );
nor U7839 ( n4148, n258, n322 );
nor U7840 ( n4147, n4149, n4150 );
nor U7841 ( n4149, n1884, n891 );
nand U7842 ( n3874, n3875, n3876 );
nand U7843 ( n3876, n3877, n3878 );
nand U7844 ( n3875, n3880, n3808 );
nor U7845 ( n3878, n118, n122 );
nand U7846 ( n4191, n4207, n4208 );
nand U7847 ( n4208, n2559, n4209 );
nor U7848 ( n4207, n4210, n4211 );
nor U7849 ( n4211, n1193, n4212 );
nand U7850 ( n4174, n4175, n2247 );
nor U7851 ( n4175, n4176, n4177 );
nor U7852 ( n4177, n310, n1092 );
nor U7853 ( n4176, n4178, n4179 );
nand U7854 ( n4162, n2143, n4163 );
nand U7855 ( n4163, n4164, n2146 );
nor U7856 ( n4164, n4165, n4166 );
nor U7857 ( n4166, n315, n1001 );
nor U7858 ( n4228, n4232, n4233 );
nor U7859 ( n4233, n1280, n4234 );
nor U7860 ( n4232, n4235, n4236 );
nand U7861 ( n4234, n2582, n1266 );
nor U7862 ( n4133, n4135, n4136 );
nor U7863 ( n4136, n236, n327 );
nor U7864 ( n4135, n4137, n4138 );
nor U7865 ( n4137, n811, n1560 );
nor U7866 ( n4310, n4677, n4676 );
nand U7867 ( n4256, n4264, n3922 );
nor U7868 ( n4264, n4255, n4265 );
nor U7869 ( n4265, n2798, n4266 );
nand U7870 ( n4266, n3921, n1373 );
nand U7871 ( n2798, n4672, n4673 );
nor U7872 ( n4673, n4674, n4675 );
nor U7873 ( n4672, n4678, n4679 );
nor U7874 ( n4674, n4993, n5146 );
nor U7875 ( n4678, n4994, n5150 );
nor U7876 ( n4675, n5137, n4967 );
xor U7877 ( n3464, n3777, n5161 );
nand U7878 ( n3777, n3778, n3779 );
nand U7879 ( n3778, n5116, n1131 );
nand U7880 ( n3779, n5156, n1104 );
nand U7881 ( n3388, n3729, n3730 );
nand U7882 ( n3730, n5115, n1309 );
nand U7883 ( n3729, n5162, n1324 );
nor U7884 ( n4569, n4997, n5150 );
nand U7885 ( n1359, n4565, n4566 );
nor U7886 ( n4566, n4567, n4568 );
nor U7887 ( n4565, n4569, n4570 );
nor U7888 ( n4567, n4996, n5146 );
nor U7889 ( n4568, n5137, n4995 );
not U7890 ( n185, n1276 );
nand U7891 ( n3339, n3721, n3722 );
nand U7892 ( n3722, n5115, n1276 );
nand U7893 ( n3721, n5162, n1303 );
nand U7894 ( n1342, n4557, n4558 );
nor U7895 ( n4558, n4559, n4560 );
nor U7896 ( n4557, n4561, n4562 );
nor U7897 ( n4559, n4998, n5146 );
not U7898 ( n169, n1309 );
nand U7899 ( n2685, n297, n1309 );
nand U7900 ( n3049, n3714, n3715 );
nand U7901 ( n3715, n5115, n1235 );
nand U7902 ( n3714, n5162, n1260 );
not U7903 ( n175, n1235 );
nand U7904 ( n2749, n295, n1347 );
nand U7905 ( n3922, n293, n1356 );
nand U7906 ( n3541, n3709, n3710 );
nand U7907 ( n3710, n5115, n1266 );
nand U7908 ( n3709, n5162, n1280 );
not U7909 ( n177, n1266 );
xor U7910 ( n3432, n3175, n3639 );
nor U7911 ( n3639, n3640, n3641 );
nor U7912 ( n3641, n317, n3179 );
nor U7913 ( n3640, n5155, n2134 );
xnor U7914 ( n3263, n3175, n3632 );
nor U7915 ( n3632, n3633, n3634 );
nor U7916 ( n3634, n318, n3179 );
nor U7917 ( n3633, n5155, n1988 );
not U7918 ( n187, n1225 );
nand U7919 ( n2452, n305, n1183 );
and U7920 ( n4209, n2452, n4216 );
nand U7921 ( n4216, n303, n1193 );
nand U7922 ( n1303, n4541, n4542 );
nor U7923 ( n4542, n4543, n4544 );
nor U7924 ( n4541, n4545, n4546 );
nor U7925 ( n4544, n5007, n5146 );
nor U7926 ( n4553, n5006, n5150 );
nand U7927 ( n1324, n4549, n4550 );
nor U7928 ( n4550, n4551, n4552 );
nor U7929 ( n4549, n4553, n4554 );
nor U7930 ( n4552, n5005, n5146 );
not U7931 ( n210, n1104 );
nand U7932 ( n4192, n4193, n4182 );
nor U7933 ( n4193, n4202, n4203 );
nor U7934 ( n4203, n305, n1183 );
nor U7935 ( n4202, n306, n1148 );
not U7936 ( n216, n1137 );
nor U7937 ( n4543, n3344, n5137 );
nand U7938 ( n3213, n3699, n3700 );
nand U7939 ( n3700, n5115, n1225 );
nand U7940 ( n3699, n5162, n1239 );
nor U7941 ( n4551, n513, n5137 );
not U7942 ( n513, n1296 );
nand U7943 ( n1280, n4532, n4533 );
nor U7944 ( n4533, n4534, n4535 );
nor U7945 ( n4532, n4537, n4538 );
nor U7946 ( n4535, n5009, n5146 );
nor U7947 ( n4537, n5010, n5150 );
nand U7948 ( n4190, n2366, n1137 );
nor U7949 ( n2559, n302, n1225 );
xnor U7950 ( n3359, n3617, n5161 );
nand U7951 ( n3617, n3618, n3619 );
nand U7952 ( n3618, n5114, n1040 );
nand U7953 ( n3619, n5156, n1013 );
not U7954 ( n200, n1193 );
nand U7955 ( n1260, n4523, n4524 );
nor U7956 ( n4524, n4525, n4526 );
nor U7957 ( n4523, n4528, n4529 );
nor U7958 ( n4526, n5011, n5146 );
nor U7959 ( n4528, n5012, n5150 );
nand U7960 ( n2804, n292, n1373 );
not U7961 ( n202, n1148 );
nand U7962 ( n762, n763, n765 );
or U7963 ( n765, n5205, n766 );
nand U7964 ( n763, n5230, n767 );
nand U7965 ( n959, n758, n760 );
nor U7966 ( n758, n771, n772 );
nor U7967 ( n760, n761, n762 );
nor U7968 ( n771, n5228, n5067 );
xnor U7969 ( n3476, n3175, n3642 );
nor U7970 ( n3642, n3643, n3644 );
nor U7971 ( n3644, n320, n3179 );
nor U7972 ( n3643, n5155, n1960 );
nor U7973 ( n4525, n3056, n5137 );
nand U7974 ( n3770, n3780, n3781 );
nand U7975 ( n3781, n5116, n1104 );
nand U7976 ( n3780, n5162, n1131 );
and U7977 ( n3279, n3782, n3783 );
nand U7978 ( n3783, n5116, n1137 );
nand U7979 ( n3782, n5162, n1153 );
nand U7980 ( n3403, n3691, n3692 );
nand U7981 ( n3692, n5115, n1193 );
nand U7982 ( n3691, n5162, n1214 );
nand U7983 ( n1198, n4496, n4497 );
nor U7984 ( n4497, n4498, n4499 );
nor U7985 ( n4496, n4501, n4502 );
nor U7986 ( n4499, n5028, n5145 );
nand U7987 ( n2243, n310, n1092 );
nand U7988 ( n2614, n298, n1276 );
xnor U7989 ( n3300, n3175, n3568 );
nor U7990 ( n3568, n3569, n3570 );
nor U7991 ( n3570, n323, n3179 );
nor U7992 ( n3569, n5155, n1744 );
xnor U7993 ( n3563, n5160, n3651 );
nor U7994 ( n3651, n3652, n3653 );
nor U7995 ( n3653, n325, n3179 );
nor U7996 ( n3652, n5155, n1766 );
nand U7997 ( n1214, n4505, n4506 );
nor U7998 ( n4506, n4507, n4508 );
nor U7999 ( n4505, n4510, n4511 );
nor U8000 ( n4508, n5023, n5145 );
nand U8001 ( n2369, n308, n1104 );
nor U8002 ( n4507, n3408, n5137 );
nand U8003 ( n1531, n1532, n1533 );
nand U8004 ( n1533, n1508, n1534 );
nand U8005 ( n1532, n99, n1538 );
xor U8006 ( n3371, n3175, n3648 );
nor U8007 ( n3648, n3649, n3650 );
nor U8008 ( n3650, n322, n3179 );
nor U8009 ( n3649, n5155, n1884 );
nand U8010 ( n3494, n3772, n3773 );
nand U8011 ( n3773, n5116, n1148 );
nand U8012 ( n3772, n5162, n1176 );
xnor U8013 ( n3096, n3175, n3645 );
nor U8014 ( n3645, n3646, n3647 );
nor U8015 ( n3647, n321, n3179 );
nor U8016 ( n3646, n5155, n1860 );
not U8017 ( n196, n1183 );
nand U8018 ( n2024, n2282, n2283 );
nand U8019 ( n2282, n1080, n1057 );
nand U8020 ( n2283, n2284, n2285 );
nand U8021 ( n2285, n311, n158 );
nand U8022 ( n2484, n2659, n2660 );
nand U8023 ( n2659, n1303, n1276 );
nand U8024 ( n2660, n2661, n2662 );
nand U8025 ( n2661, n2663, n2664 );
nand U8026 ( n1657, n1889, n1890 );
nand U8027 ( n1889, n263, n907 );
nand U8028 ( n1890, n1891, n1892 );
nand U8029 ( n1892, n321, n1860 );
nand U8030 ( n1891, n1956, n1957 );
nand U8031 ( n1956, n270, n931 );
nand U8032 ( n1957, n1958, n1959 );
nand U8033 ( n1959, n320, n1960 );
nand U8034 ( n2610, n300, n1266 );
nand U8035 ( n2722, n296, n1320 );
not U8036 ( n158, n1057 );
nand U8037 ( n1239, n4514, n4515 );
nor U8038 ( n4515, n4516, n4517 );
nor U8039 ( n4514, n4519, n4520 );
nor U8040 ( n4517, n5019, n5145 );
nand U8041 ( n3115, n3686, n3687 );
nand U8042 ( n3687, n5115, n1183 );
nand U8043 ( n3686, n5162, n1198 );
nand U8044 ( n1176, n4487, n4488 );
nor U8045 ( n4488, n4489, n4490 );
nor U8046 ( n4487, n4492, n4493 );
nor U8047 ( n4490, n5031, n5145 );
nor U8048 ( n4492, n5033, n5149 );
nor U8049 ( n4489, n3499, n5137 );
nand U8050 ( n1207, n3500, n3501 );
nor U8051 ( n3500, n3514, n3515 );
nor U8052 ( n3501, n3502, n3503 );
nor U8053 ( n3514, n296, n5165 );
nand U8054 ( n2416, n306, n1148 );
not U8055 ( n152, n1047 );
nand U8056 ( n2783, n1375, n1356 );
nand U8057 ( n1131, n4469, n4470 );
nor U8058 ( n4470, n4471, n4472 );
nor U8059 ( n4469, n4474, n4475 );
nor U8060 ( n4472, n5030, n5145 );
nand U8061 ( n2292, n311, n1057 );
nand U8062 ( n1153, n4478, n4479 );
nor U8063 ( n4479, n4480, n4481 );
nor U8064 ( n4478, n4483, n4484 );
nor U8065 ( n4481, n5026, n5145 );
nand U8066 ( n2411, n307, n1137 );
nor U8067 ( n4471, n3468, n5138 );
nand U8068 ( n2581, n301, n1235 );
nand U8069 ( n2739, n1359, n1347 );
not U8070 ( n149, n1013 );
nand U8071 ( n2556, n302, n1225 );
xnor U8072 ( n3064, n5160, n3176 );
nor U8073 ( n3176, n3177, n3178 );
nor U8074 ( n3178, n326, n3179 );
nor U8075 ( n3177, n5155, n1601 );
xor U8076 ( n3420, n4652, n3236 );
xor U8077 ( n4652, n3175, n8 );
nor U8078 ( n4646, n3420, n4651 );
nand U8079 ( n4651, n4650, n2799 );
nand U8080 ( n4642, n4643, n4615 );
nand U8081 ( n4643, n59, n4694 );
xnor U8082 ( n4694, n4695, n4696 );
xor U8083 ( n4696, n5006, n4260 );
nand U8084 ( n4613, n4614, n4615 );
nand U8085 ( n4614, n59, n4616 );
xnor U8086 ( n4616, n4617, n4618 );
xor U8087 ( n4618, n4997, n4263 );
nand U8088 ( n1034, n4639, n4640 );
nor U8089 ( n4639, n3389, n4700 );
nor U8090 ( n4640, n4641, n4642 );
nand U8091 ( n4700, n4701, n4702 );
nand U8092 ( n1042, n4610, n4611 );
nor U8093 ( n4610, n4622, n4623 );
nor U8094 ( n4611, n4612, n4613 );
nor U8095 ( n4622, STATE_REG, n4995 );
nand U8096 ( n4615, n4644, n4645 );
nor U8097 ( n4644, n4692, n5140 );
nor U8098 ( n4645, n4646, n4647 );
and U8099 ( n4692, n4303, n4606 );
not U8100 ( n222, n1092 );
nand U8101 ( n1108, n4460, n4461 );
nor U8102 ( n4461, n4462, n4463 );
nor U8103 ( n4460, n4465, n4466 );
nor U8104 ( n4463, n5035, n5145 );
nor U8105 ( n4465, n5036, n5149 );
nand U8106 ( n3232, n3236, n8 );
nand U8107 ( n1282, n3220, n3221 );
nor U8108 ( n3220, n3241, n3242 );
nor U8109 ( n3221, n3222, n3223 );
nor U8110 ( n3241, n295, n5166 );
or U8111 ( n3230, n3236, n8 );
nand U8112 ( n2245, n312, n1047 );
nand U8113 ( n2714, n1342, n1320 );
nand U8114 ( n2330, n2358, n2359 );
nand U8115 ( n2358, n2360, n2361 );
nand U8116 ( n2361, n1131, n1104 );
nor U8117 ( n2360, n2362, n2363 );
nor U8118 ( n2312, n2323, n2328 );
and U8119 ( n2328, n2329, n2330 );
nand U8120 ( n2329, n1108, n1092 );
not U8121 ( n145, n1001 );
nand U8122 ( n3083, n3678, n3679 );
nand U8123 ( n3679, n5115, n1092 );
nand U8124 ( n3678, n5162, n1108 );
nand U8125 ( n3613, n3673, n3674 );
nand U8126 ( n3674, n5115, n1057 );
nand U8127 ( n3673, n5162, n1080 );
nand U8128 ( n2216, n313, n1013 );
nand U8129 ( n2513, n2570, n175 );
nor U8130 ( n2570, n2571, n1225 );
nand U8131 ( n2638, n2706, n161 );
nor U8132 ( n2706, n2707, n1309 );
nand U8133 ( n2428, n2512, n196 );
nor U8134 ( n2512, n2513, n1193 );
nand U8135 ( n2113, n2197, n145 );
nor U8136 ( n2197, n2198, n1013 );
nand U8137 ( n2198, n2265, n152 );
nor U8138 ( n2265, n2266, n1057 );
nand U8139 ( n2707, n2763, n36 );
nor U8140 ( n2763, n1356, n1347 );
nand U8141 ( n2571, n2637, n177 );
nor U8142 ( n2637, n2638, n1276 );
nand U8143 ( n2266, n2341, n222 );
nor U8144 ( n2341, n2342, n1104 );
nand U8145 ( n2342, n2427, n216 );
nor U8146 ( n2427, n2428, n1148 );
nand U8147 ( n3319, n3607, n3608 );
nand U8148 ( n3608, n5114, n1047 );
nand U8149 ( n3607, n5162, n1063 );
nand U8150 ( n753, n1503, n1496 );
nand U8151 ( n1503, n227, n1506 );
nand U8152 ( n1506, n1505, n1507 );
nand U8153 ( n2663, n1324, n1309 );
nand U8154 ( n2365, n1176, n1148 );
nand U8155 ( n1232, n3409, n3410 );
nor U8156 ( n3410, n3411, n3412 );
nor U8157 ( n3409, n3418, n3419 );
nor U8158 ( n3411, n3413, n4967 );
nor U8159 ( n2623, n1280, n1266 );
nor U8160 ( n791, n1505, n1598 );
and U8161 ( n1598, n236, n1599 );
nand U8162 ( n1599, n1600, n1601 );
not U8163 ( n137, n968 );
nand U8164 ( n969, n735, n736 );
nor U8165 ( n735, n745, n746 );
nor U8166 ( n736, n737, n738 );
nor U8167 ( n746, n5230, n5073 );
nor U8168 ( n3883, n3890, n695 );
nor U8169 ( n3890, n3891, n3892 );
nor U8170 ( n3892, n2824, n3888 );
nor U8171 ( n3891, n9, n2816 );
nand U8172 ( n3602, n3615, n3616 );
nand U8173 ( n3616, n5114, n1013 );
nand U8174 ( n3615, n5162, n1040 );
nand U8175 ( n964, n747, n748 );
nor U8176 ( n747, n745, n755 );
nor U8177 ( n748, n750, n751 );
nor U8178 ( n755, n5228, n5075 );
nand U8179 ( n2490, n1280, n1266 );
xor U8180 ( n817, n1601, n1600 );
nand U8181 ( n2478, n1239, n1225 );
nor U8182 ( n831, n1600, n1741 );
and U8183 ( n1741, n247, n1742 );
nand U8184 ( n1742, n1743, n1744 );
nand U8185 ( n1080, n4451, n4452 );
nor U8186 ( n4452, n4453, n4454 );
nor U8187 ( n4451, n4456, n4457 );
nor U8188 ( n4454, n5037, n5145 );
nor U8189 ( n4456, n5040, n5149 );
nor U8190 ( n4453, n3822, n5138 );
nand U8191 ( n2489, n1260, n1235 );
nand U8192 ( n1063, n4442, n4443 );
nor U8193 ( n4443, n4444, n4445 );
nor U8194 ( n4442, n4447, n4448 );
nor U8195 ( n4445, n5038, n5145 );
nor U8196 ( n4447, n5039, n5149 );
nand U8197 ( n963, n965, n966 );
nand U8198 ( n965, n5235, n968 );
nand U8199 ( n966, n5242, n967 );
xor U8200 ( n857, n1743, n1744 );
nand U8201 ( n997, n999, n1000 );
nand U8202 ( n1000, n5235, n1001 );
nand U8203 ( n999, n5231, n1003 );
nand U8204 ( n2143, n316, n968 );
nor U8205 ( n871, n1743, n1857 );
and U8206 ( n1857, n258, n1858 );
nand U8207 ( n1858, n1859, n1860 );
nor U8208 ( n2324, n1176, n1148 );
nand U8209 ( n1088, n1089, n1091 );
nand U8210 ( n1091, n5236, n1092 );
nand U8211 ( n1089, n5231, n1093 );
nor U8212 ( n2323, n1108, n1092 );
nand U8213 ( n1043, n1044, n1045 );
nand U8214 ( n1045, n5236, n1047 );
nand U8215 ( n1044, n5231, n1048 );
not U8216 ( n281, n2134 );
nand U8217 ( n2002, n952, n1988 );
nand U8218 ( n2474, n1198, n1183 );
xor U8219 ( n897, n1860, n1859 );
nor U8220 ( n911, n1859, n1985 );
and U8221 ( n1985, n270, n1986 );
nand U8222 ( n1986, n1987, n1988 );
not U8223 ( n258, n1884 );
nor U8224 ( n657, n658, n660 );
nor U8225 ( n660, n661, n662 );
nor U8226 ( n658, n142, n667 );
nand U8227 ( n662, n663, n665 );
nand U8228 ( n663, n150, n146 );
not U8229 ( n150, n645 );
nand U8230 ( n653, n655, n656 );
nand U8231 ( n655, n696, n59 );
nand U8232 ( n656, n657, n58 );
nor U8233 ( n696, n697, n698 );
nand U8234 ( n2092, n995, n968 );
not U8235 ( n270, n1960 );
nand U8236 ( n1133, n1135, n1136 );
nand U8237 ( n1136, n5236, n1137 );
nand U8238 ( n1135, n5231, n1139 );
nand U8239 ( n1040, n4433, n4434 );
nor U8240 ( n4434, n4435, n4436 );
nor U8241 ( n4433, n4438, n4439 );
nor U8242 ( n4436, n5042, n5145 );
nand U8243 ( n1099, n1100, n1101 );
nand U8244 ( n1100, n5236, n1104 );
nand U8245 ( n1101, n1103, n5241 );
not U8246 ( n275, n1988 );
nor U8247 ( n4435, n3363, n5138 );
nand U8248 ( n2099, n972, n2134 );
not U8249 ( n263, n1860 );
xor U8250 ( n937, n1987, n1988 );
nand U8251 ( n3152, n3627, n3628 );
nand U8252 ( n3628, n5114, n968 );
nand U8253 ( n3627, n5162, n995 );
nand U8254 ( n666, n642, n645 );
nand U8255 ( n665, n666, n5048 );
xor U8256 ( n3021, n4989, n4979 );
not U8257 ( n347, n4269 );
nand U8258 ( n702, n52, n146 );
not U8259 ( n52, n640 );
not U8260 ( n54, n4806 );
not U8261 ( n55, n4813 );
not U8262 ( n53, n731 );
nand U8263 ( n2089, n317, n2134 );
nand U8264 ( n2254, n1063, n1047 );
nand U8265 ( n2043, n1017, n1001 );
nand U8266 ( n1179, n1180, n1181 );
nand U8267 ( n1181, n5236, n1183 );
nand U8268 ( n1180, n5231, n1184 );
nor U8269 ( n698, n700, n701 );
nand U8270 ( n701, n702, n703 );
nand U8271 ( n703, n705, n5051 );
nand U8272 ( n705, n642, n640 );
nand U8273 ( n2177, n315, n1001 );
nand U8274 ( n1017, n4424, n4425 );
nor U8275 ( n4425, n4426, n4427 );
nor U8276 ( n4424, n4429, n4430 );
nor U8277 ( n4427, n5048, n5145 );
nor U8278 ( n4429, n5051, n5149 );
nand U8279 ( n3526, n3595, n3596 );
nand U8280 ( n3596, n5114, n1001 );
nand U8281 ( n3595, n5163, n1017 );
nor U8282 ( n993, n35, n2195 );
and U8283 ( n2195, n1001, n2196 );
nand U8284 ( n2196, n149, n34 );
nand U8285 ( n1008, n1009, n1011 );
nand U8286 ( n1009, n5236, n1013 );
nand U8287 ( n1011, n1012, n5241 );
nand U8288 ( n1721, n851, n1766 );
nand U8289 ( n3901, n907, n1860 );
nand U8290 ( n635, n636, n637 );
nand U8291 ( n637, n59, n638 );
nand U8292 ( n636, n58, n643 );
xor U8293 ( n638, n640, n641 );
nand U8294 ( n2028, n318, n1988 );
nand U8295 ( n1796, n867, n1744 );
nand U8296 ( n1948, n931, n1960 );
xor U8297 ( n3009, n3016, n4990 );
nand U8298 ( n995, n4415, n4416 );
nor U8299 ( n4416, n4417, n4418 );
nor U8300 ( n4415, n4420, n4421 );
nor U8301 ( n4418, n5045, n5145 );
nand U8302 ( n3902, n891, n1884 );
nor U8303 ( n4417, n3157, n5138 );
nor U8304 ( n1039, n34, n2263 );
and U8305 ( n2263, n1047, n2264 );
nand U8306 ( n2264, n158, n33 );
nand U8307 ( n972, n4406, n4407 );
nor U8308 ( n4407, n4408, n4409 );
nor U8309 ( n4406, n4411, n4412 );
nor U8310 ( n4409, n5144, n5044 );
nand U8311 ( n891, n4370, n4371 );
nor U8312 ( n4371, n4372, n4373 );
nor U8313 ( n4370, n4375, n4376 );
nor U8314 ( n4373, n5144, n5056 );
nand U8315 ( n1493, n4295, n106 );
nor U8316 ( n4295, n2816, n2826 );
nand U8317 ( n1377, n5224, n695 );
nand U8318 ( n824, n1332, n1333 );
nor U8319 ( n1332, n1343, n1344 );
nor U8320 ( n1333, n1334, n1335 );
nor U8321 ( n1343, n5228, n4996 );
nand U8322 ( n844, n1248, n1249 );
nor U8323 ( n1248, n1261, n1263 );
nor U8324 ( n1249, n1250, n1251 );
nor U8325 ( n1261, n5228, n5009 );
nand U8326 ( n854, n1206, n1208 );
nor U8327 ( n1206, n1220, n1221 );
nor U8328 ( n1208, n1209, n1210 );
nor U8329 ( n1220, n5229, n5019 );
nand U8330 ( n834, n1289, n1290 );
nor U8331 ( n1289, n1304, n1305 );
nor U8332 ( n1290, n1291, n1293 );
nor U8333 ( n1304, n5228, n5005 );
nand U8334 ( n1189, n1190, n1191 );
nand U8335 ( n1191, n5202, n495 );
nand U8336 ( n1190, n5236, n1193 );
nand U8337 ( n1053, n1055, n1056 );
nand U8338 ( n1056, n5203, n491 );
nand U8339 ( n1055, n5236, n1057 );
nand U8340 ( n1273, n1274, n1275 );
nand U8341 ( n1275, n13, n5241 );
nand U8342 ( n1274, n5236, n1276 );
nand U8343 ( n1263, n1264, n1265 );
nand U8344 ( n1264, n5231, n1268 );
nand U8345 ( n1265, n5236, n1266 );
nand U8346 ( n1231, n1233, n1234 );
nand U8347 ( n1234, n14, n5241 );
nand U8348 ( n1233, n5236, n1235 );
nand U8349 ( n1144, n1145, n1147 );
nand U8350 ( n1147, n5202, n497 );
nand U8351 ( n1145, n5236, n1148 );
nand U8352 ( n1221, n1223, n1224 );
nand U8353 ( n1223, n5231, n1226 );
nand U8354 ( n1224, n5236, n1225 );
nand U8355 ( n931, n4388, n4389 );
nor U8356 ( n4389, n4390, n4391 );
nor U8357 ( n4388, n4393, n4394 );
nor U8358 ( n4391, n5144, n5052 );
nor U8359 ( n4408, n3442, n5138 );
nand U8360 ( n819, n1349, n1350 );
nor U8361 ( n1350, n1351, n1352 );
nor U8362 ( n1349, n1360, n1361 );
nand U8363 ( n1351, n1357, n1358 );
nand U8364 ( n1344, n1345, n1346 );
nand U8365 ( n1345, n5232, n1348 );
nand U8366 ( n1346, n5237, n1347 );
nand U8367 ( n1352, n1353, n1354 );
nand U8368 ( n1354, n5242, n1355 );
nand U8369 ( n1353, n5237, n1356 );
nand U8370 ( n1315, n1316, n1318 );
nand U8371 ( n1318, n5242, n1319 );
nand U8372 ( n1316, n5237, n1320 );
nand U8373 ( n1305, n1306, n1308 );
nand U8374 ( n1306, n5232, n1310 );
nand U8375 ( n1308, n5237, n1309 );
nand U8376 ( n1293, n1294, n1295 );
nand U8377 ( n1295, n5202, n1296 );
nand U8378 ( n1294, n1298, n5241 );
nand U8379 ( n952, n4397, n4398 );
nor U8380 ( n4398, n4399, n4400 );
nor U8381 ( n4397, n4402, n4403 );
nor U8382 ( n4400, n5144, n5049 );
nand U8383 ( n814, n1366, n1367 );
nor U8384 ( n1367, n1368, n1369 );
nor U8385 ( n1366, n1378, n1379 );
nor U8386 ( n1368, n5205, n4967 );
nand U8387 ( n907, n4379, n4380 );
nor U8388 ( n4380, n4381, n4382 );
nor U8389 ( n4379, n4384, n4385 );
nor U8390 ( n4382, n5144, n5054 );
nor U8391 ( n4372, n3377, n5139 );
nand U8392 ( n616, n617, n618 );
nand U8393 ( n618, n59, n620 );
nand U8394 ( n617, n58, n625 );
xor U8395 ( n620, n621, n622 );
nor U8396 ( n4399, n3268, n5138 );
nor U8397 ( n1084, n33, n2339 );
and U8398 ( n2339, n1092, n2340 );
nand U8399 ( n2340, n210, n32 );
nor U8400 ( n4390, n3484, n5138 );
nor U8401 ( n2998, n4880, n4869 );
nor U8402 ( n4880, n5001, n346 );
nand U8403 ( n2220, n1040, n1013 );
nor U8404 ( n4381, n3104, n5138 );
not U8405 ( n240, n1601 );
nand U8406 ( n1587, n811, n1560 );
not U8407 ( n228, n1507 );
not U8408 ( n236, n1560 );
not U8409 ( n252, n1744 );
nor U8410 ( n1129, n32, n2425 );
and U8411 ( n2425, n1137, n2426 );
nand U8412 ( n2426, n202, n31 );
nand U8413 ( n1650, n832, n1601 );
not U8414 ( n247, n1766 );
xnor U8415 ( n2993, n5000, n4869 );
nor U8416 ( n3004, n4980, n4888 );
nor U8417 ( n4887, n4888, n3004 );
nand U8418 ( n851, n4352, n4353 );
nor U8419 ( n4353, n4354, n4355 );
nor U8420 ( n4352, n4357, n4358 );
nor U8421 ( n4355, n5144, n5059 );
nand U8422 ( n597, n598, n600 );
nand U8423 ( n600, n59, n601 );
nand U8424 ( n598, n58, n606 );
xnor U8425 ( n601, n602, n603 );
nor U8426 ( n4101, n1509, n740 );
nand U8427 ( n2836, n3866, n3867 );
nand U8428 ( n3867, n3868, n5058 );
nor U8429 ( n3866, n288, n3869 );
nor U8430 ( n3869, n5058, n3870 );
nand U8431 ( n1388, n285, n2828 );
not U8432 ( n285, n2827 );
nand U8433 ( n3833, n3834, n3835 );
nand U8434 ( n3834, n287, n3839 );
nand U8435 ( n3835, n287, n3836 );
nand U8436 ( n3839, n3840, n3841 );
nand U8437 ( n3870, n333, n3829 );
nand U8438 ( n2827, n3830, n3831 );
nor U8439 ( n3830, n3849, n3850 );
nor U8440 ( n3831, n3832, n3833 );
nand U8441 ( n3849, n3859, n3860 );
xor U8442 ( n2957, n2964, n5017 );
nand U8443 ( n3850, n3851, n3852 );
nand U8444 ( n3851, n287, n3856 );
nand U8445 ( n3852, n287, n3853 );
nand U8446 ( n3856, n3857, n3858 );
nand U8447 ( n1764, n323, n1744 );
not U8448 ( n288, n3871 );
nand U8449 ( n3832, n3842, n3843 );
nand U8450 ( n3842, n287, n3847 );
nand U8451 ( n3843, n287, n3844 );
nand U8452 ( n3847, n3848, n5065 );
xor U8453 ( n2969, n5021, n2976 );
nand U8454 ( n1678, n325, n1766 );
and U8455 ( n4103, n1534, n752 );
nor U8456 ( n4354, n3664, n5139 );
nand U8457 ( n867, n4361, n4362 );
nor U8458 ( n4362, n4363, n4364 );
nor U8459 ( n4361, n4366, n4367 );
nor U8460 ( n4364, n5144, n5061 );
xor U8461 ( n2981, n2988, n5014 );
nor U8462 ( n1175, n31, n2510 );
and U8463 ( n2510, n1183, n2511 );
nand U8464 ( n2511, n200, n30 );
nand U8465 ( n3886, n3887, n92 );
and U8466 ( n3887, n695, n3888 );
nand U8467 ( n1321, n5202, n5076 );
nor U8468 ( n4363, n3308, n5139 );
nand U8469 ( n1660, n322, n1884 );
nand U8470 ( n1605, n326, n1601 );
not U8471 ( n227, n752 );
nand U8472 ( n3943, n3959, n1507 );
nand U8473 ( n3953, n3954, n1560 );
xor U8474 ( n2945, n2952, n4982 );
xor U8475 ( n581, n582, n583 );
xor U8476 ( n583, n5037, n159 );
nand U8477 ( n577, n578, n580 );
nand U8478 ( n578, n59, n585 );
nand U8479 ( n580, n58, n581 );
xor U8480 ( n585, n586, n587 );
nor U8481 ( n4123, n1507, n786 );
nor U8482 ( n1218, n30, n2568 );
and U8483 ( n2568, n1225, n2569 );
nand U8484 ( n2569, n175, n29 );
xor U8485 ( n3120, n5025, n4491 );
nor U8486 ( n4527, n5002, n4536 );
nor U8487 ( n4509, n5013, n4518 );
nor U8488 ( n4491, n5015, n4500 );
nand U8489 ( n3960, n1509, n740 );
nand U8490 ( n832, n4343, n4344 );
nor U8491 ( n4344, n4345, n4346 );
nor U8492 ( n4343, n4348, n4349 );
nor U8493 ( n4346, n5144, n5066 );
nor U8494 ( n4473, n5018, n4482 );
not U8495 ( n286, n1487 );
not U8496 ( n118, n3808 );
nor U8497 ( n2891, n5063, n2892 );
nor U8498 ( n4921, n2892, n2891 );
nor U8499 ( n4606, n4993, n4979 );
nand U8500 ( n811, n4334, n4335 );
nor U8501 ( n4335, n4336, n4337 );
nor U8502 ( n4334, n4339, n4340 );
nor U8503 ( n4337, n5144, n5068 );
nand U8504 ( n3908, n3909, n1523 );
xor U8505 ( n3909, n740, n1509 );
xor U8506 ( n2933, n2940, n5034 );
xor U8507 ( n3551, n5004, n4527 );
nor U8508 ( n4345, n3073, n5139 );
nand U8509 ( n786, n4324, n4325 );
nor U8510 ( n4325, n4326, n4327 );
nor U8511 ( n4324, n4330, n4331 );
nor U8512 ( n4327, n5144, n5067 );
xor U8513 ( n3088, n4970, n4455 );
nor U8514 ( n4455, n4464, n4968 );
nand U8515 ( n1369, n1370, n1371 );
nand U8516 ( n1370, n5207, n1375 );
nand U8517 ( n1371, n1372, n1373 );
nand U8518 ( n1372, n742, n741 );
nor U8519 ( n1259, n29, n2635 );
and U8520 ( n2635, n1266, n2636 );
nand U8521 ( n2636, n185, n28 );
xor U8522 ( n3288, n5022, n4473 );
nor U8523 ( n4336, n3203, n5139 );
nor U8524 ( n4120, n752, n1534 );
nand U8525 ( n558, n560, n561 );
nand U8526 ( n560, n59, n567 );
nand U8527 ( n561, n58, n562 );
xnor U8528 ( n567, n568, n570 );
nand U8529 ( n1520, n327, n1560 );
nand U8530 ( n3806, n2825, n2826 );
xor U8531 ( n3912, n752, n1534 );
nand U8532 ( n2832, n288, n3829 );
nor U8533 ( n738, n740, n741 );
nor U8534 ( n751, n741, n752 );
nor U8535 ( n4326, n766, n5139 );
xor U8536 ( n2921, n2928, n4981 );
nor U8537 ( n4401, n4410, n4973 );
nor U8538 ( n4383, n5041, n4392 );
nor U8539 ( n4365, n4975, n4374 );
nor U8540 ( n4437, n4446, n4969 );
nor U8541 ( n4419, n4428, n4972 );
not U8542 ( n225, n740 );
nor U8543 ( n1301, n28, n2704 );
and U8544 ( n2704, n1309, n2705 );
nand U8545 ( n2705, n161, n27 );
nor U8546 ( n996, n5230, n5048 );
nor U8547 ( n1064, n5230, n5037 );
nor U8548 ( n1019, n5230, n5042 );
nor U8549 ( n973, n5230, n5045 );
nor U8550 ( n953, n5230, n5044 );
nor U8551 ( n913, n5230, n5052 );
nor U8552 ( n892, n5230, n5054 );
xor U8553 ( n3219, n5016, n4509 );
nand U8554 ( n4909, n4915, n3025 );
nor U8555 ( n4915, n4917, n4918 );
nor U8556 ( n4918, n4305, n3808 );
nor U8557 ( n4917, n62, n5189 );
nand U8558 ( n4593, n4650, n4835 );
nand U8559 ( n4588, n59, n4994 );
and U8560 ( n3025, n4916, n5244 );
nand U8561 ( n4916, n5187, n3808 );
nand U8562 ( n1050, n4581, n4582 );
nor U8563 ( n4581, n4594, n4595 );
nor U8564 ( n4582, n4583, n4584 );
nor U8565 ( n4595, n5244, n4967 );
nor U8566 ( n1378, n5228, n4993 );
nor U8567 ( n1132, n5229, n5026 );
nor U8568 ( n1155, n5229, n5031 );
nor U8569 ( n1240, n5228, n5011 );
nor U8570 ( n1177, n5229, n5028 );
nor U8571 ( n1360, n5228, n4991 );
nor U8572 ( n1325, n5228, n4998 );
nor U8573 ( n1041, n5229, n5038 );
nor U8574 ( n1109, n5229, n5030 );
nor U8575 ( n1087, n5229, n5035 );
nor U8576 ( n1199, n5229, n5023 );
nor U8577 ( n1281, n5228, n5007 );
nor U8578 ( n833, n5228, n5059 );
nor U8579 ( n812, n5229, n5066 );
nor U8580 ( n793, n5228, n5068 );
nor U8581 ( n932, n5229, n5049 );
nor U8582 ( n873, n5229, n5056 );
nor U8583 ( n852, n5229, n5061 );
or U8584 ( n3940, n5110, n3942 );
or U8585 ( n5110, n227, n740 );
nand U8586 ( n4134, n786, n1507 );
xor U8587 ( n3165, n3175, n3196 );
nor U8588 ( n3196, n3197, n3198 );
nor U8589 ( n3198, n327, n5089 );
nor U8590 ( n3197, n1560, n3179 );
nor U8591 ( n4347, n4976, n4356 );
xor U8592 ( n3328, n4971, n4437 );
nand U8593 ( n540, n541, n542 );
nand U8594 ( n541, n59, n548 );
nand U8595 ( n542, n58, n543 );
xor U8596 ( n548, n550, n551 );
nand U8597 ( n3942, n1534, n1509 );
nand U8598 ( n4599, n4600, n4601 );
nand U8599 ( n4601, n4602, n59 );
nand U8600 ( n4600, n57, n4269 );
xor U8601 ( n4602, n4269, n4603 );
nand U8602 ( n1046, n4596, n4597 );
nor U8603 ( n4596, n4608, n4609 );
nor U8604 ( n4597, n4598, n4599 );
nor U8605 ( n4609, STATE_REG, n4966 );
nand U8606 ( n4702, n57, n4260 );
nor U8607 ( n1341, n27, n2761 );
and U8608 ( n2761, n1347, n2762 );
nand U8609 ( n2762, n36, n163 );
nand U8610 ( n4770, n4771, n4772 );
nand U8611 ( n4771, n59, n4776 );
nand U8612 ( n4772, n58, n4773 );
xor U8613 ( n4776, n341, n4777 );
nand U8614 ( n4745, n4746, n4747 );
nand U8615 ( n4746, n59, n4751 );
nand U8616 ( n4747, n58, n4748 );
xor U8617 ( n4751, n345, n4752 );
nand U8618 ( n4706, n4707, n4708 );
nand U8619 ( n4707, n59, n4712 );
nand U8620 ( n4708, n58, n4709 );
xor U8621 ( n4712, n4239, n4713 );
nand U8622 ( n4629, n4630, n4631 );
nand U8623 ( n4630, n59, n4635 );
nand U8624 ( n4631, n58, n4632 );
xor U8625 ( n4635, n4272, n4636 );
nand U8626 ( n4795, n4796, n4797 );
nand U8627 ( n4797, n59, n4798 );
nand U8628 ( n4796, n58, n4836 );
xor U8629 ( n4798, n337, n4799 );
nand U8630 ( n4782, n4783, n4784 );
nand U8631 ( n4784, n59, n4785 );
nand U8632 ( n4783, n58, n4788 );
xor U8633 ( n4785, n4786, n4787 );
nand U8634 ( n4732, n4733, n4734 );
nand U8635 ( n4734, n59, n4735 );
nand U8636 ( n4733, n58, n4738 );
xor U8637 ( n4735, n4736, n4737 );
nand U8638 ( n4757, n4758, n4759 );
nand U8639 ( n4759, n59, n4760 );
nand U8640 ( n4758, n58, n4763 );
xor U8641 ( n4760, n4761, n4762 );
nand U8642 ( n4719, n4720, n4721 );
nand U8643 ( n4721, n59, n4722 );
nand U8644 ( n4720, n58, n4725 );
xnor U8645 ( n4722, n4723, n4724 );
and U8646 ( n4718, n4243, n57 );
and U8647 ( n615, n623, n57 );
and U8648 ( n596, n605, n57 );
and U8649 ( n557, n566, n57 );
and U8650 ( n538, n547, n57 );
and U8651 ( n4756, n4219, n57 );
and U8652 ( n4705, n4239, n57 );
and U8653 ( n4628, n4272, n57 );
nand U8654 ( n3361, n5226, n1013 );
nand U8655 ( n3466, n5226, n1104 );
nand U8656 ( n3528, n5226, n1001 );
nand U8657 ( n3326, n5226, n1047 );
nand U8658 ( n3118, n5225, n1183 );
nand U8659 ( n3406, n5226, n1193 );
nand U8660 ( n3342, n5226, n1276 );
nand U8661 ( n3053, n5225, n1235 );
nand U8662 ( n3286, n5225, n1137 );
nand U8663 ( n3155, n5225, n968 );
nand U8664 ( n3141, n5225, n1320 );
nand U8665 ( n3497, n5226, n1148 );
nand U8666 ( n3549, n5226, n1266 );
nand U8667 ( n3086, n5225, n1092 );
nand U8668 ( n3217, n5225, n1225 );
nand U8669 ( n3391, n5226, n1309 );
nand U8670 ( n3800, n5227, n1057 );
nor U8671 ( n4329, n4338, n4977 );
xor U8672 ( n3530, n4974, n4419 );
and U8673 ( n5111, n1486, n1487 );
and U8674 ( n1486, n2817, n2818 );
nor U8675 ( n2818, n2819, n2820 );
nor U8676 ( n2817, n2827, n2828 );
nor U8677 ( n2819, n2821, n2822 );
not U8678 ( n114, n2826 );
not U8679 ( n345, n4227 );
xnor U8680 ( n4836, n693, n4837 );
xor U8681 ( n4837, n5026, n692 );
nor U8682 ( n4598, n4589, n4605 );
xor U8683 ( n4605, n4606, n4607 );
xor U8684 ( n4607, n4991, n4269 );
nor U8685 ( n2895, n2897, n5173 );
and U8686 ( n1508, n62, n1535 );
nand U8687 ( n1535, n1536, n5186 );
nand U8688 ( n1536, n290, n5058 );
nor U8689 ( n2900, n5173, n2902 );
nand U8690 ( n2902, n2903, n2904 );
nor U8691 ( n2924, n5173, n2926 );
nand U8692 ( n2926, n2927, n2928 );
nor U8693 ( n2936, n5173, n2938 );
nand U8694 ( n2938, n2939, n2940 );
nor U8695 ( n2850, n5172, n2852 );
nand U8696 ( n2852, n2853, n2840 );
nor U8697 ( n2856, n5172, n2858 );
nand U8698 ( n2858, n2859, n2860 );
nor U8699 ( n2868, n5172, n2870 );
nand U8700 ( n2870, n2871, n2872 );
nor U8701 ( n2875, n5172, n2877 );
nand U8702 ( n2877, n2878, n2879 );
nor U8703 ( n2887, n5172, n2889 );
nand U8704 ( n2889, n2890, n119 );
nand U8705 ( n2890, n2892, n5063 );
not U8706 ( n119, n2891 );
nor U8707 ( n2912, n5172, n2914 );
nand U8708 ( n2914, n2915, n2916 );
nor U8709 ( n2948, n5172, n2950 );
nand U8710 ( n2950, n2951, n2952 );
nor U8711 ( n2960, n5172, n2962 );
nand U8712 ( n2962, n2963, n2964 );
nor U8713 ( n2972, n5172, n2974 );
nand U8714 ( n2974, n2975, n2976 );
nor U8715 ( n2984, n5172, n2986 );
nand U8716 ( n2986, n2987, n2988 );
nor U8717 ( n3012, n5172, n3014 );
nand U8718 ( n3014, n3015, n3016 );
not U8719 ( n331, n1509 );
nor U8720 ( n1607, n5182, n1560 );
nor U8721 ( n1812, n5182, n1744 );
nor U8722 ( n2060, n5182, n1988 );
nor U8723 ( n1683, n5182, n1601 );
nor U8724 ( n1931, n5182, n1860 );
nor U8725 ( n1527, n5182, n1507 );
nor U8726 ( n1748, n5182, n1766 );
nor U8727 ( n1991, n5182, n1960 );
nor U8728 ( n2116, n5182, n2134 );
nor U8729 ( n1863, n5182, n1884 );
nand U8730 ( n1625, n3819, n695 );
nor U8731 ( n3819, n114, n143 );
xor U8732 ( n2821, n2825, n2826 );
buf U8733 ( n5245, n5247 );
nand U8734 ( n757, n1508, n1509 );
xor U8735 ( n4788, n4789, n4790 );
xor U8736 ( n4790, n5031, n338 );
nor U8737 ( n3813, n3815, n2825 );
nor U8738 ( n3815, n112, n3816 );
nand U8739 ( n3816, n111, n110 );
and U8740 ( n3795, n3809, n3810 );
nor U8741 ( n3810, n1374, n3811 );
nor U8742 ( n3809, n3813, n2075 );
nor U8743 ( n3811, n3812, n2826 );
nand U8744 ( n3050, n3798, n3797 );
nor U8745 ( n3798, n2799, n283 );
not U8746 ( n341, n4222 );
nand U8747 ( n3663, n3804, n3805 );
nor U8748 ( n3805, n282, n1387 );
nor U8749 ( n3804, n3807, n3808 );
nor U8750 ( n3807, n3795, n3794 );
nand U8751 ( n3392, n1296, n3055 );
nand U8752 ( n3142, n3055, n5076 );
xnor U8753 ( n4773, n4774, n4775 );
xor U8754 ( n4775, n5028, n4222 );
nor U8755 ( n1374, n1493, n695 );
nor U8756 ( n369, n5181, n5065 );
nor U8757 ( n444, n5181, n5064 );
nand U8758 ( n1516, n2815, n114 );
nor U8759 ( n2815, n122, n2816 );
not U8760 ( n337, n692 );
xnor U8761 ( n4748, n4749, n4750 );
xor U8762 ( n4750, n5019, n4227 );
xor U8763 ( n4738, n4739, n4740 );
xor U8764 ( n4740, n5011, n343 );
nand U8765 ( n1732, n62, n2799 );
nand U8766 ( n5125, n62, n2799 );
xnor U8767 ( n4725, n4726, n4727 );
xor U8768 ( n4727, n5009, n4243 );
nor U8769 ( n4297, n5123, n4299 );
nor U8770 ( n4299, n4300, n3808 );
nor U8771 ( n4300, n4301, n4302 );
nand U8772 ( n4301, n2826, n4305 );
nor U8773 ( n4303, n290, n4650 );
not U8774 ( n488, n3203 );
not U8775 ( n487, n3073 );
not U8776 ( n486, n3664 );
not U8777 ( n142, n661 );
nand U8778 ( n4298, n2826, n3808 );
not U8779 ( n146, n642 );
not U8780 ( n485, n3308 );
not U8781 ( n483, n3377 );
not U8782 ( n482, n3104 );
not U8783 ( n159, n590 );
xor U8784 ( n587, n5040, n159 );
not U8785 ( n481, n3484 );
xor U8786 ( n603, n5039, n605 );
not U8787 ( n480, n3268 );
xor U8788 ( n570, n5036, n566 );
nor U8789 ( n3139, n5244, n5076 );
nor U8790 ( n733, n5244, n4973 );
nor U8791 ( n630, n5244, n4972 );
nor U8792 ( n553, n5244, n4968 );
nor U8793 ( n592, n5244, n4969 );
nor U8794 ( n3404, n5244, n5015 );
nor U8795 ( n3051, n5244, n5013 );
nor U8796 ( n3495, n5244, n5018 );
nor U8797 ( n3340, n5244, n5002 );
nor U8798 ( n648, n5244, n4974 );
nor U8799 ( n611, n5244, n4971 );
nor U8800 ( n572, n5244, n4970 );
nor U8801 ( n3116, n5244, n5025 );
nor U8802 ( n3215, n5244, n5016 );
nor U8803 ( n3547, n5244, n5004 );
nor U8804 ( n3284, n5244, n5022 );
not U8805 ( n478, n3442 );
nor U8806 ( n3389, n5244, n5003 );
xor U8807 ( n4787, n5033, n338 );
xor U8808 ( n4737, n5012, n343 );
not U8809 ( n338, n4206 );
not U8810 ( n343, n4246 );
xor U8811 ( n4724, n5010, n4243 );
not U8812 ( n477, n3157 );
not U8813 ( n475, n3363 );
not U8814 ( n491, n3822 );
buf U8815 ( n5246, n5247 );
not U8816 ( n500, n3468 );
not U8817 ( n497, n3499 );
not U8818 ( n495, n3408 );
not U8819 ( n492, n3056 );
xor U8820 ( n4603, n4992, n4604 );
not U8821 ( n512, n3344 );
nor U8822 ( n4869, n4881, IR_REG_5_ );
nand U8823 ( n3016, n4965, n4979 );
nor U8824 ( n4965, IR_REG_2_, IR_REG_1_ );
nor U8825 ( n4888, n3016, IR_REG_3_ );
nand U8826 ( n2976, n4963, n342 );
nor U8827 ( n4963, IR_REG_9_, IR_REG_8_ );
nand U8828 ( n2988, n4964, n4869 );
nor U8829 ( n4964, IR_REG_7_, IR_REG_6_ );
nand U8830 ( n2916, n4959, n144 );
nor U8831 ( n4959, IR_REG_19_, IR_REG_18_ );
nand U8832 ( n2964, n4962, n340 );
nor U8833 ( n4962, IR_REG_11_, IR_REG_10_ );
nand U8834 ( n2940, n4960, n335 );
nor U8835 ( n4960, IR_REG_15_, IR_REG_14_ );
nand U8836 ( n2952, n4961, n336 );
nor U8837 ( n4961, IR_REG_13_, IR_REG_12_ );
nand U8838 ( n2825, n4954, n4955 );
nand U8839 ( n4954, IR_REG_21_, n5214 );
nand U8840 ( n4955, n4956, IR_REG_31_ );
and U8841 ( n4956, n2904, n2903 );
nand U8842 ( n2903, IR_REG_21_, n4957 );
nand U8843 ( n4957, n120, n4985 );
nand U8844 ( n1292, n3158, n3159 );
nor U8845 ( n3158, n3199, n3200 );
nor U8846 ( n3159, n3160, n3161 );
and U8847 ( n3199, n5246, REG3_REG_28_ );
nand U8848 ( n2904, n4958, n120 );
nor U8849 ( n4958, IR_REG_21_, IR_REG_20_ );
nand U8850 ( n1192, n3552, n3553 );
nor U8851 ( n3552, n3656, n3657 );
nor U8852 ( n3553, n3554, n3555 );
and U8853 ( n3656, n5246, REG3_REG_26_ );
nand U8854 ( n2816, n4686, n4687 );
nand U8855 ( n4686, IR_REG_20_, n5214 );
or U8856 ( n4687, n2909, n5213 );
xor U8857 ( n3236, n4653, n5161 );
nand U8858 ( n4653, n4654, n4655 );
nand U8859 ( n4655, REG1_REG_0_, n282 );
nor U8860 ( n4654, n4656, n4657 );
nand U8861 ( n2915, IR_REG_19_, n4691 );
nand U8862 ( n4691, n144, n4981 );
nand U8863 ( n695, n4688, n4689 );
nand U8864 ( n4688, IR_REG_19_, n5214 );
nand U8865 ( n4689, n4690, IR_REG_31_ );
and U8866 ( n4690, n2916, n2915 );
xnor U8867 ( n2897, n2904, IR_REG_22_ );
nand U8868 ( n2826, n4952, n4953 );
nand U8869 ( n4952, IR_REG_22_, n5216 );
or U8870 ( n4953, n2897, n5213 );
nand U8871 ( n1247, n3364, n3365 );
nor U8872 ( n3364, n3373, n3374 );
nor U8873 ( n3365, n3366, n3367 );
and U8874 ( n3373, n5246, REG3_REG_24_ );
and U8875 ( n3829, n4927, n4928 );
nand U8876 ( n4927, IR_REG_25_, n5216 );
nand U8877 ( n4928, n4929, IR_REG_31_ );
and U8878 ( n4929, n2879, n2878 );
nand U8879 ( n2878, IR_REG_25_, n4930 );
nand U8880 ( n4930, n291, n4986 );
nand U8881 ( n3871, n4924, n4925 );
nand U8882 ( n4924, IR_REG_26_, n5216 );
nand U8883 ( n4925, n4926, IR_REG_31_ );
and U8884 ( n4926, n2872, n2871 );
or U8885 ( n2872, n2879, IR_REG_26_ );
nand U8886 ( n3868, n4931, n4932 );
nand U8887 ( n4931, IR_REG_24_, n5216 );
or U8888 ( n4932, n2884, n5213 );
nand U8889 ( n2871, IR_REG_26_, n2879 );
buf U8890 ( n5212, n388 );
not U8891 ( n388, IR_REG_31_ );
nand U8892 ( n1217, n3469, n3470 );
nor U8893 ( n3469, n3480, n3481 );
nor U8894 ( n3470, n3471, n3472 );
and U8895 ( n3480, n5246, REG3_REG_22_ );
nand U8896 ( n1227, n3421, n3422 );
nor U8897 ( n3421, n3438, n3439 );
nor U8898 ( n3422, n3423, n3424 );
and U8899 ( n3438, n5246, REG3_REG_20_ );
nor U8900 ( n4951, IR_REG_17_, IR_REG_16_ );
nand U8901 ( n4946, n4949, n4983 );
nor U8902 ( n4949, IR_REG_23_, IR_REG_22_ );
nor U8903 ( n4948, IR_REG_20_, IR_REG_19_ );
nor U8904 ( n4650, n5112, n5113 );
and U8905 ( n5112, IR_REG_27_, n5216 );
nor U8906 ( n5113, n2865, n5213 );
nand U8907 ( n1356, n4267, n4268 );
nand U8908 ( n4268, n5189, n4269 );
nand U8909 ( n4267, DATAI_1_, n5186 );
nand U8910 ( n2799, n4934, n4935 );
nand U8911 ( n4934, IR_REG_28_, n5216 );
nand U8912 ( n4935, n4936, IR_REG_31_ );
and U8913 ( n4936, n2860, n2859 );
nand U8914 ( n2860, n4939, n4938 );
nor U8915 ( n4939, IR_REG_28_, n4933 );
nand U8916 ( n2859, IR_REG_28_, n4937 );
nand U8917 ( n4937, n4938, n291 );
nand U8918 ( n3748, n4659, n4660 );
nand U8919 ( n4660, IR_REG_0_, n282 );
nor U8920 ( n4659, n4661, n4662 );
nor U8921 ( n4661, n292, n5089 );
nand U8922 ( n1373, n4665, n4666 );
nand U8923 ( n4666, n5189, IR_REG_0_ );
nand U8924 ( n4665, DATAI_0_, n5187 );
nor U8925 ( n4940, IR_REG_25_, IR_REG_24_ );
nand U8926 ( n1347, n4261, n4262 );
nand U8927 ( n4262, n5189, n4263 );
nand U8928 ( n4261, DATAI_2_, n5186 );
nand U8929 ( n1320, n4270, n4271 );
nand U8930 ( n4271, n5189, n4272 );
nand U8931 ( n4270, DATAI_3_, n5186 );
nand U8932 ( n4677, n4682, n4683 );
nand U8933 ( n4682, IR_REG_30_, n5214 );
or U8934 ( n4683, n2846, n5213 );
or U8935 ( n2840, n2860, IR_REG_29_ );
nand U8936 ( n1182, n3872, n3873 );
nand U8937 ( n3872, B_REG, n4296 );
nand U8938 ( n3873, n3874, n5244 );
nand U8939 ( n4296, n4297, n4298 );
and U8940 ( n4578, n5154, REG0_REG_1_ );
and U8941 ( n4679, n5154, REG0_REG_0_ );
nand U8942 ( n4676, n4680, n4681 );
nand U8943 ( n4680, IR_REG_29_, n5215 );
nand U8944 ( n4681, IR_REG_31_, n2853 );
nand U8945 ( n2853, IR_REG_29_, n2860 );
nand U8946 ( n1276, n4237, n4238 );
nand U8947 ( n4238, n5189, n4239 );
nand U8948 ( n4237, DATAI_5_, n5187 );
and U8949 ( n4570, n5154, REG0_REG_2_ );
nor U8950 ( n4561, n4999, n5150 );
nand U8951 ( n1309, n4258, n4259 );
nand U8952 ( n4259, n5189, n4260 );
nand U8953 ( n4258, DATAI_4_, n5186 );
nand U8954 ( n1235, n4244, n4245 );
nand U8955 ( n4245, n5189, n4246 );
nand U8956 ( n4244, DATAI_7_, n5187 );
nor U8957 ( n4560, REG3_REG_3_, n5137 );
and U8958 ( n4562, n5154, REG0_REG_3_ );
nand U8959 ( n1266, n4241, n4242 );
nand U8960 ( n4242, n5189, n4243 );
nand U8961 ( n4241, DATAI_6_, n5187 );
nand U8962 ( n1225, n4225, n4226 );
nand U8963 ( n4226, n5189, n4227 );
nand U8964 ( n4225, DATAI_8_, n5187 );
and U8965 ( n4938, n4940, n4941 );
nor U8966 ( n4941, IR_REG_27_, IR_REG_26_ );
nand U8967 ( n1183, n4220, n4221 );
nand U8968 ( n4221, n5189, n4222 );
nand U8969 ( n4220, DATAI_10_, n5187 );
nand U8970 ( n1193, n4217, n4218 );
nand U8971 ( n4218, n5189, n4219 );
nand U8972 ( n4217, DATAI_9_, n5187 );
nor U8973 ( n4545, n5008, n5150 );
nand U8974 ( n1104, n4196, n4197 );
nand U8975 ( n4197, n5189, n547 );
nand U8976 ( n4196, DATAI_13_, n5187 );
nand U8977 ( n1137, n4194, n4195 );
nand U8978 ( n4195, n5189, n692 );
nand U8979 ( n4194, DATAI_12_, n5187 );
and U8980 ( n4554, n5154, REG0_REG_4_ );
and U8981 ( n4546, n5154, REG0_REG_5_ );
nand U8982 ( n1148, n4204, n4205 );
nand U8983 ( n4205, n5189, n4206 );
nand U8984 ( n4204, DATAI_11_, n5187 );
nand U8985 ( n629, n1665, n1666 );
nand U8986 ( n1665, REG0_REG_27_, n5191 );
nand U8987 ( n1666, n5117, n1404 );
nand U8988 ( n789, n1402, n1403 );
nand U8989 ( n1402, REG1_REG_27_, n5195 );
nand U8990 ( n1403, n5120, n1404 );
and U8991 ( n4538, n5153, REG0_REG_6_ );
nand U8992 ( n634, n1590, n1591 );
nand U8993 ( n1590, REG0_REG_28_, n5190 );
nand U8994 ( n1591, n5117, n1401 );
nand U8995 ( n794, n1399, n1400 );
nand U8996 ( n1399, REG1_REG_28_, n5194 );
nand U8997 ( n1400, n5120, n1401 );
nand U8998 ( n639, n1510, n1511 );
nand U8999 ( n1510, REG0_REG_29_, n5191 );
nand U9000 ( n1511, n5117, n1398 );
nand U9001 ( n799, n1396, n1397 );
nand U9002 ( n1396, REG1_REG_29_, n5195 );
nand U9003 ( n1397, n5120, n1398 );
and U9004 ( n4529, n5153, REG0_REG_7_ );
nand U9005 ( n609, n1922, n1923 );
nand U9006 ( n1922, REG0_REG_23_, n5191 );
nand U9007 ( n1923, n5117, n1416 );
nand U9008 ( n769, n1414, n1415 );
nand U9009 ( n1414, REG1_REG_23_, n5195 );
nand U9010 ( n1415, n5120, n1416 );
and U9011 ( n4502, n5153, REG0_REG_10_ );
nor U9012 ( n4501, n5029, n5149 );
nand U9013 ( n1092, n4183, n4184 );
nand U9014 ( n4184, n5189, n566 );
nand U9015 ( n4183, DATAI_14_, n5187 );
and U9016 ( n4511, n5153, REG0_REG_9_ );
nor U9017 ( n4510, n5024, n5149 );
nand U9018 ( n624, n1733, n1734 );
nand U9019 ( n1733, REG0_REG_26_, n5190 );
nand U9020 ( n1734, n5117, n1407 );
nand U9021 ( n784, n1405, n1406 );
nand U9022 ( n1405, REG1_REG_26_, n5194 );
nand U9023 ( n1406, n5120, n1407 );
nand U9024 ( n1057, n4273, n4274 );
nand U9025 ( n4274, n5189, n590 );
nand U9026 ( n4273, DATAI_15_, n5186 );
and U9027 ( n4520, n5153, REG0_REG_8_ );
nor U9028 ( n4519, n5020, n5149 );
nand U9029 ( n604, n1977, n1978 );
nand U9030 ( n1977, REG0_REG_22_, n5191 );
nand U9031 ( n1978, n5117, n1419 );
nand U9032 ( n764, n1417, n1418 );
nand U9033 ( n1417, REG1_REG_22_, n5195 );
nand U9034 ( n1418, n5120, n1419 );
nand U9035 ( n619, n1800, n1801 );
nand U9036 ( n1800, REG0_REG_25_, n5191 );
nand U9037 ( n1801, n5117, n1410 );
nand U9038 ( n779, n1408, n1409 );
nand U9039 ( n1408, REG1_REG_25_, n5195 );
nand U9040 ( n1409, n5120, n1410 );
nand U9041 ( n599, n2044, n2045 );
nand U9042 ( n2044, REG0_REG_21_, n5191 );
nand U9043 ( n2045, n5117, n1422 );
nand U9044 ( n759, n1420, n1421 );
nand U9045 ( n1420, REG1_REG_21_, n5195 );
nand U9046 ( n1421, n5120, n1422 );
and U9047 ( n4493, n5153, REG0_REG_11_ );
nand U9048 ( n3503, n3504, n3505 );
nand U9049 ( n3504, REG3_REG_2_, n3239 );
nand U9050 ( n3505, n5168, n3506 );
nand U9051 ( n3506, n3507, n3508 );
nand U9052 ( n1047, n4279, n4280 );
nand U9053 ( n4280, n5189, n605 );
nand U9054 ( n4279, DATAI_16_, n5186 );
and U9055 ( n4475, n5153, REG0_REG_13_ );
nor U9056 ( n4474, n5032, n5149 );
and U9057 ( n4484, n5153, REG0_REG_12_ );
nor U9058 ( n4483, n5027, n5149 );
nand U9059 ( n4269, n4905, n4906 );
nand U9060 ( n4906, IR_REG_31_, n3021 );
nand U9061 ( n4905, IR_REG_1_, n5215 );
nand U9062 ( n614, n1849, n1850 );
nand U9063 ( n1849, REG0_REG_24_, n5190 );
nand U9064 ( n1850, n5117, n1413 );
nand U9065 ( n774, n1411, n1412 );
nand U9066 ( n1411, REG1_REG_24_, n5194 );
nand U9067 ( n1412, n5120, n1413 );
nand U9068 ( n1013, n4283, n4284 );
nand U9069 ( n4284, n5189, n623 );
nand U9070 ( n4283, DATAI_17_, n5186 );
nand U9071 ( n594, n2102, n2103 );
nand U9072 ( n2102, REG0_REG_20_, n5191 );
nand U9073 ( n2103, n5117, n1425 );
nand U9074 ( n754, n1423, n1424 );
nand U9075 ( n1423, REG1_REG_20_, n5195 );
nand U9076 ( n1424, n5120, n1425 );
and U9077 ( n4466, n5153, REG0_REG_14_ );
nand U9078 ( n3223, n3224, n3225 );
nand U9079 ( n3224, REG3_REG_1_, n3239 );
nand U9080 ( n3225, n5169, n3226 );
nand U9081 ( n3226, n3227, n3228 );
nand U9082 ( n1001, n4289, n4290 );
nand U9083 ( n4290, n5189, n642 );
nand U9084 ( n4289, DATAI_18_, n5186 );
nand U9085 ( n649, n1488, n1489 );
nand U9086 ( n1488, REG0_REG_31_, n5191 );
nand U9087 ( n1489, n5117, n1391 );
nand U9088 ( n809, n1389, n1390 );
nand U9089 ( n1389, REG1_REG_31_, n5195 );
nand U9090 ( n1390, n5120, n1391 );
nand U9091 ( n589, n2153, n2154 );
nand U9092 ( n2153, REG0_REG_19_, n5191 );
nand U9093 ( n2154, n5118, n1428 );
nand U9094 ( n749, n1426, n1427 );
nand U9095 ( n1426, REG1_REG_19_, n5195 );
nand U9096 ( n1427, n5121, n1428 );
nand U9097 ( n4263, n4898, n4899 );
nand U9098 ( n4899, n4900, IR_REG_31_ );
nand U9099 ( n4898, IR_REG_2_, n5215 );
and U9100 ( n4900, n3016, n3015 );
nand U9101 ( n4272, n4893, n4894 );
nand U9102 ( n4893, IR_REG_3_, n5215 );
or U9103 ( n4894, n3009, n5213 );
nand U9104 ( n644, n1498, n1499 );
nand U9105 ( n1498, REG0_REG_30_, n5190 );
nand U9106 ( n1499, n5117, n1395 );
nand U9107 ( n804, n1393, n1394 );
nand U9108 ( n1393, REG1_REG_30_, n5194 );
nand U9109 ( n1394, n5120, n1395 );
nand U9110 ( n968, n4293, n4294 );
nand U9111 ( n4294, n5189, n695 );
nand U9112 ( n4293, DATAI_19_, n5186 );
and U9113 ( n4457, n5153, REG0_REG_15_ );
nand U9114 ( n719, n1444, n1445 );
nand U9115 ( n1444, REG1_REG_13_, n5195 );
nand U9116 ( n1445, n5121, n1446 );
nand U9117 ( n559, n2374, n2375 );
nand U9118 ( n2374, REG0_REG_13_, n5191 );
nand U9119 ( n2375, n5118, n1446 );
and U9120 ( n4448, n5153, REG0_REG_16_ );
nand U9121 ( n744, n1429, n1430 );
nand U9122 ( n1429, REG1_REG_18_, n5195 );
nand U9123 ( n1430, n5121, n1431 );
nand U9124 ( n584, n2187, n2188 );
nand U9125 ( n2187, REG0_REG_18_, n5191 );
nand U9126 ( n2188, n5118, n1431 );
nand U9127 ( n564, n2331, n2332 );
nand U9128 ( n2331, REG0_REG_14_, n5191 );
nand U9129 ( n2332, n5118, n1443 );
nand U9130 ( n724, n1441, n1442 );
nand U9131 ( n1441, REG1_REG_14_, n5195 );
nand U9132 ( n1442, n5121, n1443 );
nand U9133 ( n574, n2255, n2256 );
nand U9134 ( n2255, REG0_REG_16_, n5191 );
nand U9135 ( n2256, n5118, n1437 );
nand U9136 ( n734, n1435, n1436 );
nand U9137 ( n1435, REG1_REG_16_, n5195 );
nand U9138 ( n1436, n5121, n1437 );
nand U9139 ( n2134, DATAI_20_, n5186 );
nand U9140 ( n1988, DATAI_21_, n5186 );
nand U9141 ( n739, n1432, n1433 );
nand U9142 ( n1432, REG1_REG_17_, n5195 );
nand U9143 ( n1433, n5121, n1434 );
nand U9144 ( n579, n2222, n2223 );
nand U9145 ( n2222, REG0_REG_17_, n5191 );
nand U9146 ( n2223, n5118, n1434 );
nand U9147 ( n1884, DATAI_24_, n5187 );
nand U9148 ( n4699, n4890, n4891 );
nand U9149 ( n4890, n4633, n4272 );
nand U9150 ( n4891, REG2_REG_3_, n4892 );
or U9151 ( n4892, n4272, n4633 );
nand U9152 ( n645, n670, n671 );
nand U9153 ( n670, n626, n623 );
nand U9154 ( n671, REG2_REG_17_, n672 );
or U9155 ( n672, n626, n623 );
nand U9156 ( n4633, n4895, n4896 );
nand U9157 ( n4895, n4621, n4263 );
nand U9158 ( n4896, REG2_REG_2_, n4897 );
or U9159 ( n4897, n4263, n4621 );
nand U9160 ( n4710, n4882, n4883 );
nand U9161 ( n4882, n4699, n4260 );
nand U9162 ( n4883, REG2_REG_4_, n4884 );
or U9163 ( n4884, n4260, n4699 );
nand U9164 ( n4739, n4870, n4871 );
nand U9165 ( n4870, n4726, n4243 );
nand U9166 ( n4871, REG2_REG_6_, n4872 );
or U9167 ( n4872, n4243, n4726 );
nand U9168 ( n4764, n4857, n4858 );
nand U9169 ( n4857, n4749, n4227 );
nand U9170 ( n4858, REG2_REG_8_, n4859 );
or U9171 ( n4859, n4227, n4749 );
nand U9172 ( n4789, n4845, n4846 );
nand U9173 ( n4845, n4774, n4222 );
nand U9174 ( n4846, REG2_REG_10_, n4847 );
or U9175 ( n4847, n4222, n4774 );
nand U9176 ( n545, n688, n690 );
nand U9177 ( n688, n693, n692 );
nand U9178 ( n690, REG2_REG_12_, n691 );
or U9179 ( n691, n692, n693 );
nand U9180 ( n4774, n4850, n4851 );
nand U9181 ( n4850, n4764, n4219 );
nand U9182 ( n4851, REG2_REG_9_, n4852 );
or U9183 ( n4852, n4219, n4764 );
nand U9184 ( n563, n685, n686 );
nand U9185 ( n685, n545, n547 );
nand U9186 ( n686, REG2_REG_13_, n687 );
or U9187 ( n687, n545, n547 );
nand U9188 ( n582, n681, n682 );
nand U9189 ( n681, n563, n566 );
nand U9190 ( n682, REG2_REG_14_, n683 );
or U9191 ( n683, n563, n566 );
nand U9192 ( n667, n666, n668 );
nand U9193 ( n668, REG2_REG_18_, n663 );
nand U9194 ( n4749, n4862, n4863 );
nand U9195 ( n4862, n4739, n4246 );
nand U9196 ( n4863, REG2_REG_7_, n4864 );
or U9197 ( n4864, n4246, n4739 );
nand U9198 ( n607, n677, n678 );
nand U9199 ( n677, n582, n590 );
nand U9200 ( n678, REG2_REG_15_, n680 );
or U9201 ( n680, n582, n590 );
nand U9202 ( n4726, n4875, n4876 );
nand U9203 ( n4875, n4710, n4239 );
nand U9204 ( n4876, REG2_REG_5_, n4877 );
or U9205 ( n4877, n4239, n4710 );
nand U9206 ( n4621, n4902, n4903 );
nand U9207 ( n4902, n4606, n4269 );
nand U9208 ( n4903, REG2_REG_1_, n4904 );
or U9209 ( n4904, n4269, n4606 );
nand U9210 ( n626, n673, n675 );
nand U9211 ( n673, n607, n605 );
nand U9212 ( n675, REG2_REG_16_, n676 );
or U9213 ( n676, n607, n605 );
nand U9214 ( n693, n4838, n4839 );
nand U9215 ( n4838, n4789, n4206 );
nand U9216 ( n4839, REG2_REG_11_, n4840 );
or U9217 ( n4840, n4206, n4789 );
nand U9218 ( n974, n650, n651 );
nor U9219 ( n650, n732, n733 );
nor U9220 ( n651, n652, n653 );
and U9221 ( n732, ADDR_REG_19_, n56 );
nand U9222 ( n714, n1447, n1448 );
nand U9223 ( n1447, REG1_REG_12_, n5195 );
nand U9224 ( n1448, n5121, n1449 );
nand U9225 ( n554, n2417, n2418 );
nand U9226 ( n2417, REG0_REG_12_, n5191 );
nand U9227 ( n2418, n5118, n1449 );
nand U9228 ( n1960, DATAI_22_, n5186 );
and U9229 ( n4439, n5153, REG0_REG_17_ );
nor U9230 ( n4438, n5043, n5149 );
nand U9231 ( n1860, DATAI_23_, n5187 );
nand U9232 ( n569, n2293, n2294 );
nand U9233 ( n2293, REG0_REG_15_, n5191 );
nand U9234 ( n2294, n5118, n1440 );
nand U9235 ( n729, n1438, n1439 );
nand U9236 ( n1438, REG1_REG_15_, n5195 );
nand U9237 ( n1439, n5121, n1440 );
nand U9238 ( n4714, n4823, n4824 );
nand U9239 ( n4823, n4695, n4260 );
nand U9240 ( n4824, REG1_REG_4_, n4825 );
or U9241 ( n4825, n4695, n4260 );
nand U9242 ( n4637, n4829, n4830 );
nand U9243 ( n4829, n4617, n4263 );
nand U9244 ( n4830, REG1_REG_2_, n4831 );
or U9245 ( n4831, n4617, n4263 );
nand U9246 ( n4786, n4803, n4804 );
nand U9247 ( n4803, n4222, n4806 );
nand U9248 ( n4804, REG1_REG_10_, n4805 );
nand U9249 ( n4805, n54, n341 );
nand U9250 ( n4761, n4810, n4811 );
nand U9251 ( n4810, n4227, n4813 );
nand U9252 ( n4811, REG1_REG_8_, n4812 );
nand U9253 ( n4812, n55, n345 );
nand U9254 ( n4723, n4820, n4821 );
nand U9255 ( n4820, n4239, n4714 );
nand U9256 ( n4821, REG1_REG_5_, n4822 );
or U9257 ( n4822, n4714, n4239 );
nand U9258 ( n568, n723, n725 );
nand U9259 ( n723, n550, n547 );
nand U9260 ( n725, REG1_REG_13_, n726 );
or U9261 ( n726, n550, n547 );
nand U9262 ( n4617, n4832, n4833 );
or U9263 ( n4832, n4604, n347 );
nand U9264 ( n4833, REG1_REG_1_, n4834 );
nand U9265 ( n4834, n347, n4604 );
nand U9266 ( n602, n716, n717 );
nand U9267 ( n716, n586, n590 );
nand U9268 ( n717, REG1_REG_15_, n718 );
or U9269 ( n718, n586, n590 );
nand U9270 ( n4813, n4814, n4815 );
nand U9271 ( n4814, n4736, n4246 );
nand U9272 ( n4815, REG1_REG_7_, n4816 );
or U9273 ( n4816, n4736, n4246 );
nand U9274 ( n731, n4800, n4801 );
nand U9275 ( n4800, n4786, n4206 );
nand U9276 ( n4801, REG1_REG_11_, n4802 );
or U9277 ( n4802, n4786, n4206 );
nand U9278 ( n4806, n4807, n4808 );
nand U9279 ( n4807, n4761, n4219 );
nand U9280 ( n4808, REG1_REG_9_, n4809 );
or U9281 ( n4809, n4761, n4219 );
nor U9282 ( n697, n141, n706 );
not U9283 ( n141, n700 );
nand U9284 ( n706, n705, n707 );
nand U9285 ( n707, REG1_REG_18_, n702 );
nand U9286 ( n640, n708, n710 );
nand U9287 ( n708, n621, n623 );
nand U9288 ( n710, REG1_REG_17_, n711 );
or U9289 ( n711, n621, n623 );
nand U9290 ( n550, n727, n728 );
nand U9291 ( n727, n692, n731 );
nand U9292 ( n728, REG1_REG_12_, n730 );
nand U9293 ( n730, n53, n337 );
nand U9294 ( n4736, n4817, n4818 );
nand U9295 ( n4817, n4723, n4243 );
nand U9296 ( n4818, REG1_REG_6_, n4819 );
or U9297 ( n4819, n4723, n4243 );
nand U9298 ( n586, n720, n721 );
nand U9299 ( n720, n568, n566 );
nand U9300 ( n721, REG1_REG_14_, n722 );
or U9301 ( n722, n568, n566 );
nand U9302 ( n621, n712, n713 );
nand U9303 ( n712, n602, n605 );
nand U9304 ( n713, REG1_REG_16_, n715 );
or U9305 ( n715, n602, n605 );
nand U9306 ( n4695, n4826, n4827 );
nand U9307 ( n4826, n4272, n4637 );
nand U9308 ( n4827, REG1_REG_3_, n4828 );
or U9309 ( n4828, n4637, n4272 );
nand U9310 ( n4239, n4878, n4879 );
nand U9311 ( n4879, n2998, IR_REG_31_ );
nand U9312 ( n4878, IR_REG_5_, n5215 );
nand U9313 ( n704, n1453, n1454 );
nand U9314 ( n1453, REG1_REG_10_, n5194 );
nand U9315 ( n1454, n5121, n1455 );
nand U9316 ( n544, n2502, n2503 );
nand U9317 ( n2502, REG0_REG_10_, n5190 );
nand U9318 ( n2503, n5118, n1455 );
and U9319 ( n4430, n5153, REG0_REG_18_ );
nand U9320 ( n549, n2453, n2454 );
nand U9321 ( n2453, REG0_REG_11_, n5190 );
nand U9322 ( n2454, n5118, n1452 );
nand U9323 ( n709, n1450, n1451 );
nand U9324 ( n1450, REG1_REG_11_, n5194 );
nand U9325 ( n1451, n5121, n1452 );
nand U9326 ( n1766, DATAI_26_, n5187 );
nand U9327 ( n4243, n4873, n4874 );
nand U9328 ( n4873, IR_REG_6_, n5215 );
or U9329 ( n4874, n2993, n5213 );
nand U9330 ( n699, n1456, n1457 );
nand U9331 ( n1456, REG1_REG_9_, n5194 );
nand U9332 ( n1457, n5121, n1458 );
nand U9333 ( n539, n2536, n2537 );
nand U9334 ( n2536, REG0_REG_9_, n5190 );
nand U9335 ( n2537, n5118, n1458 );
nand U9336 ( n4246, n4865, n4866 );
nand U9337 ( n4866, n4867, IR_REG_31_ );
nand U9338 ( n4865, IR_REG_7_, n5215 );
and U9339 ( n4867, n2988, n2987 );
xor U9340 ( n643, n645, n646 );
xor U9341 ( n646, n642, REG2_REG_18_ );
nand U9342 ( n978, n631, n632 );
nor U9343 ( n631, n647, n648 );
nor U9344 ( n632, n633, n635 );
and U9345 ( n647, ADDR_REG_18_, n56 );
nand U9346 ( n1744, DATAI_25_, n5187 );
nand U9347 ( n3015, IR_REG_2_, n4901 );
nand U9348 ( n4901, n4979, n4989 );
and U9349 ( n4421, n5152, REG0_REG_19_ );
nor U9350 ( n4420, n5046, n5149 );
nor U9351 ( n4411, n5148, n5047 );
nand U9352 ( n529, n2592, n2593 );
nand U9353 ( n2592, REG0_REG_7_, n5190 );
nand U9354 ( n2593, n5119, n1464 );
nand U9355 ( n689, n1462, n1463 );
nand U9356 ( n1462, REG1_REG_7_, n5194 );
nand U9357 ( n1463, n5122, n1464 );
nor U9358 ( n4375, n5148, n5057 );
and U9359 ( n4412, n5152, REG0_REG_20_ );
nand U9360 ( n694, n1459, n1460 );
nand U9361 ( n1459, REG1_REG_8_, n5194 );
nand U9362 ( n1460, n5121, n1461 );
nand U9363 ( n534, n2560, n2561 );
nand U9364 ( n2560, REG0_REG_8_, n5190 );
nand U9365 ( n2561, n5118, n1461 );
nor U9366 ( n4393, n5148, n5053 );
nor U9367 ( n4402, n5148, n5050 );
nand U9368 ( n1335, n1336, n1338 );
nand U9369 ( n1338, REG3_REG_2_, n5202 );
nand U9370 ( n1336, n11, n5241 );
nor U9371 ( n4384, n5148, n5055 );
nand U9372 ( n4227, n4860, n4861 );
nand U9373 ( n4860, IR_REG_8_, n5215 );
or U9374 ( n4861, n2981, n5214 );
and U9375 ( n4403, n5152, REG0_REG_21_ );
xor U9376 ( n625, n626, n627 );
xor U9377 ( n627, n623, REG2_REG_17_ );
nand U9378 ( n982, n612, n613 );
nor U9379 ( n612, n628, n630 );
nor U9380 ( n613, n615, n616 );
and U9381 ( n628, ADDR_REG_17_, n56 );
and U9382 ( n4376, n5152, REG0_REG_24_ );
nand U9383 ( n1601, DATAI_27_, n5187 );
and U9384 ( n4394, n5152, REG0_REG_22_ );
nand U9385 ( n4222, n4848, n4849 );
nand U9386 ( n4848, IR_REG_10_, n5215 );
or U9387 ( n4849, n2969, n5213 );
nand U9388 ( n1560, DATAI_28_, n5187 );
nand U9389 ( n524, n2627, n2628 );
nand U9390 ( n2627, REG0_REG_6_, n5190 );
nand U9391 ( n2628, n5119, n1467 );
nand U9392 ( n684, n1465, n1466 );
nand U9393 ( n1465, REG1_REG_6_, n5194 );
nand U9394 ( n1466, n5122, n1467 );
nand U9395 ( n1507, DATAI_29_, n5187 );
and U9396 ( n4385, n5152, REG0_REG_23_ );
nand U9397 ( n547, n4198, n4199 );
nand U9398 ( n4198, IR_REG_13_, n5214 );
nand U9399 ( n4199, n4200, IR_REG_31_ );
and U9400 ( n4200, n2952, n2951 );
nand U9401 ( n2951, IR_REG_13_, n4201 );
nand U9402 ( n4201, n336, n5017 );
nand U9403 ( n2987, IR_REG_7_, n4868 );
nand U9404 ( n4868, n4869, n5000 );
nand U9405 ( n4219, n4853, n4854 );
nand U9406 ( n4854, n4855, IR_REG_31_ );
nand U9407 ( n4853, IR_REG_9_, n5215 );
and U9408 ( n4855, n2976, n2975 );
nand U9409 ( n4260, n4885, n4886 );
nand U9410 ( n4885, IR_REG_4_, n4889 );
nand U9411 ( n4886, n4887, IR_REG_31_ );
nand U9412 ( n4889, n3004, IR_REG_31_ );
nor U9413 ( n4357, n5148, n5060 );
nand U9414 ( n692, n4912, n4913 );
nand U9415 ( n4912, IR_REG_12_, n5215 );
or U9416 ( n4913, n2957, n5213 );
xor U9417 ( n606, n607, n608 );
xor U9418 ( n608, n605, REG2_REG_16_ );
nand U9419 ( n986, n593, n595 );
nor U9420 ( n593, n610, n611 );
nor U9421 ( n595, n596, n597 );
and U9422 ( n610, ADDR_REG_16_, n56 );
nand U9423 ( n740, DATAI_31_, n5187 );
nand U9424 ( n679, n1468, n1469 );
nand U9425 ( n1468, REG1_REG_5_, n5194 );
nand U9426 ( n1469, n5122, n1470 );
nand U9427 ( n519, n2667, n2668 );
nand U9428 ( n2667, REG0_REG_5_, n5190 );
nand U9429 ( n2668, n5119, n1470 );
nand U9430 ( n752, DATAI_30_, n5187 );
nand U9431 ( n3860, n287, n3861 );
nand U9432 ( n3861, n3862, n5064 );
nor U9433 ( n3862, D_REG_24_, D_REG_23_ );
nand U9434 ( n3859, n287, n3863 );
nand U9435 ( n3863, n3864, n3865 );
nor U9436 ( n3864, D_REG_19_, D_REG_18_ );
nor U9437 ( n3865, D_REG_21_, D_REG_20_ );
and U9438 ( n4358, n5152, REG0_REG_26_ );
nor U9439 ( n4366, n5148, n5062 );
nand U9440 ( n4206, n4841, n4842 );
nand U9441 ( n4842, n4843, IR_REG_31_ );
nand U9442 ( n4841, IR_REG_11_, n5214 );
and U9443 ( n4843, n2964, n2963 );
nand U9444 ( n2975, IR_REG_9_, n4856 );
nand U9445 ( n4856, n342, n5014 );
nand U9446 ( n1357, REG3_REG_1_, n5202 );
nand U9447 ( n2828, n3827, n3828 );
nand U9448 ( n3828, n2832, n2836 );
nand U9449 ( n3827, D_REG_1_, n287 );
and U9450 ( n4367, n5152, REG0_REG_25_ );
nand U9451 ( n2963, IR_REG_11_, n4844 );
nand U9452 ( n4844, n340, n5021 );
nand U9453 ( n514, n2696, n2697 );
nand U9454 ( n2696, REG0_REG_4_, n5190 );
nand U9455 ( n2697, n5119, n1473 );
nand U9456 ( n674, n1471, n1472 );
nand U9457 ( n1471, REG1_REG_4_, n5194 );
nand U9458 ( n1472, n5122, n1473 );
nand U9459 ( n566, n4185, n4186 );
nand U9460 ( n4185, IR_REG_14_, n5214 );
or U9461 ( n4186, n2945, n5213 );
nand U9462 ( n990, n573, n575 );
nor U9463 ( n573, n591, n592 );
nor U9464 ( n575, n576, n577 );
and U9465 ( n591, ADDR_REG_15_, n56 );
nand U9466 ( n590, n4275, n4276 );
nand U9467 ( n4275, IR_REG_15_, n5214 );
nand U9468 ( n4276, n4277, IR_REG_31_ );
and U9469 ( n4277, n2940, n2939 );
nand U9470 ( n2939, IR_REG_15_, n4278 );
nand U9471 ( n4536, REG3_REG_4_, REG3_REG_3_ );
nand U9472 ( n4518, REG3_REG_6_, n4527 );
nand U9473 ( n4500, REG3_REG_8_, n4509 );
nor U9474 ( n4348, n5148, n5069 );
xor U9475 ( n3468, n4464, REG3_REG_13_ );
nand U9476 ( n4464, REG3_REG_12_, n4473 );
nand U9477 ( n4482, REG3_REG_10_, n4491 );
nand U9478 ( n1487, n3825, n3826 );
nand U9479 ( n3826, n2835, n2836 );
nand U9480 ( n3825, D_REG_0_, n287 );
nand U9481 ( n669, n1474, n1475 );
nand U9482 ( n1474, REG1_REG_3_, n5194 );
nand U9483 ( n1475, n5122, n1476 );
nand U9484 ( n509, n2723, n2724 );
nand U9485 ( n2723, REG0_REG_3_, n5190 );
nand U9486 ( n2724, n5119, n1476 );
nand U9487 ( n3808, n4919, n4920 );
nand U9488 ( n4919, IR_REG_23_, n4922 );
nand U9489 ( n4920, n4921, IR_REG_31_ );
nand U9490 ( n4922, n2891, IR_REG_31_ );
nor U9491 ( n2892, n2904, IR_REG_22_ );
nor U9492 ( n4339, n5148, n5070 );
nand U9493 ( n605, n4281, n4282 );
nand U9494 ( n4281, IR_REG_16_, n5214 );
or U9495 ( n4282, n2933, n5213 );
xor U9496 ( n3408, n4500, REG3_REG_9_ );
xor U9497 ( n3499, n4482, REG3_REG_11_ );
nand U9498 ( n504, n2753, n2754 );
nand U9499 ( n2753, REG0_REG_2_, n5190 );
nand U9500 ( n2754, n5119, n1479 );
nand U9501 ( n664, n1477, n1478 );
nand U9502 ( n1477, REG1_REG_2_, n5194 );
nand U9503 ( n1478, n5122, n1479 );
xor U9504 ( n3344, n4536, REG3_REG_5_ );
nor U9505 ( n4330, n5148, n5071 );
xnor U9506 ( n1296, n5003, REG3_REG_3_ );
nand U9507 ( n623, n4285, n4286 );
nand U9508 ( n4285, IR_REG_17_, n5214 );
nand U9509 ( n4286, n4287, IR_REG_31_ );
and U9510 ( n4287, n2928, n2927 );
nand U9511 ( n2927, IR_REG_17_, n4288 );
nand U9512 ( n4288, n151, n5034 );
xor U9513 ( n3056, n4518, REG3_REG_7_ );
and U9514 ( n4349, n5152, REG0_REG_27_ );
and U9515 ( n4340, n5152, REG0_REG_28_ );
xor U9516 ( n562, n563, n565 );
xor U9517 ( n565, n566, REG2_REG_14_ );
nand U9518 ( n994, n555, n556 );
nor U9519 ( n555, n571, n572 );
nor U9520 ( n556, n557, n558 );
and U9521 ( n571, ADDR_REG_14_, n56 );
nand U9522 ( n1509, n4308, n4309 );
nand U9523 ( n4309, REG0_REG_31_, n5152 );
nor U9524 ( n4308, n4311, n4312 );
nor U9525 ( n4311, n5144, n5073 );
nor U9526 ( n4312, n5148, n5072 );
and U9527 ( n4331, n5152, REG0_REG_29_ );
nand U9528 ( n1534, n4318, n4319 );
nand U9529 ( n4319, REG0_REG_30_, n5152 );
nor U9530 ( n4318, n4320, n4321 );
nor U9531 ( n4320, n5144, n5075 );
nor U9532 ( n4321, n5148, n5074 );
nand U9533 ( n642, n4291, n4292 );
nand U9534 ( n4291, IR_REG_18_, n5214 );
or U9535 ( n4292, n2921, n5213 );
xnor U9536 ( n3377, REG3_REG_24_, n4365 );
nand U9537 ( n4446, n4455, REG3_REG_14_ );
nand U9538 ( n4428, n4437, REG3_REG_16_ );
nand U9539 ( n4410, n4419, REG3_REG_18_ );
nand U9540 ( n4392, REG3_REG_20_, n4401 );
nand U9541 ( n4374, REG3_REG_22_, n4383 );
nand U9542 ( n499, n2787, n2788 );
nand U9543 ( n2787, REG0_REG_1_, n5190 );
nand U9544 ( n2788, n5119, n1482 );
nand U9545 ( n659, n1480, n1481 );
nand U9546 ( n1480, REG1_REG_1_, n5194 );
nand U9547 ( n1481, n5122, n1482 );
nand U9548 ( n4604, REG1_REG_0_, IR_REG_0_ );
nor U9549 ( n4584, n4585, n4979 );
nor U9550 ( n4585, n4586, n4587 );
nor U9551 ( n4586, REG2_REG_0_, n4589 );
nand U9552 ( n4587, n4588, n588 );
xor U9553 ( n3822, n4446, REG3_REG_15_ );
xnor U9554 ( n3664, REG3_REG_26_, n4347 );
nand U9555 ( n4356, REG3_REG_24_, n4365 );
xor U9556 ( n543, n545, n546 );
xor U9557 ( n546, n547, REG2_REG_13_ );
nand U9558 ( n998, n536, n537 );
nor U9559 ( n536, n552, n553 );
nor U9560 ( n537, n538, n540 );
and U9561 ( n552, ADDR_REG_13_, n56 );
nand U9562 ( n4623, n4624, n4625 );
nand U9563 ( n4624, ADDR_REG_2_, n56 );
nand U9564 ( n4625, n57, n4263 );
xor U9565 ( n3363, n4428, REG3_REG_17_ );
xor U9566 ( n3104, n4374, REG3_REG_23_ );
nand U9567 ( n1010, n4767, n4768 );
nor U9568 ( n4767, n4778, n3116 );
nor U9569 ( n4768, n4769, n4770 );
and U9570 ( n4778, ADDR_REG_10_, n56 );
nand U9571 ( n1018, n4742, n4743 );
nor U9572 ( n4742, n4753, n3215 );
nor U9573 ( n4743, n4744, n4745 );
and U9574 ( n4753, ADDR_REG_8_, n56 );
nand U9575 ( n1030, n4703, n4704 );
nor U9576 ( n4703, n4715, n3340 );
nor U9577 ( n4704, n4705, n4706 );
and U9578 ( n4715, ADDR_REG_5_, n56 );
nand U9579 ( n1038, n4626, n4627 );
nor U9580 ( n4626, n4638, n3139 );
nor U9581 ( n4627, n4628, n4629 );
and U9582 ( n4638, ADDR_REG_3_, n56 );
nor U9583 ( n4583, IR_REG_0_, n4590 );
nor U9584 ( n4590, n4591, n4592 );
nor U9585 ( n4591, n4994, n4593 );
nor U9586 ( n4592, n4993, n4589 );
nand U9587 ( n1002, n4792, n4793 );
nor U9588 ( n4792, n4914, n3284 );
nor U9589 ( n4793, n4794, n4795 );
and U9590 ( n4914, ADDR_REG_12_, n56 );
nand U9591 ( n1006, n4779, n4780 );
nor U9592 ( n4779, n4791, n3495 );
nor U9593 ( n4780, n4781, n4782 );
and U9594 ( n4791, ADDR_REG_11_, n56 );
nand U9595 ( n1022, n4729, n4730 );
nor U9596 ( n4729, n4741, n3051 );
nor U9597 ( n4730, n4731, n4732 );
and U9598 ( n4741, ADDR_REG_7_, n56 );
nand U9599 ( n1014, n4754, n4755 );
nor U9600 ( n4754, n4766, n3404 );
nor U9601 ( n4755, n4756, n4757 );
and U9602 ( n4766, ADDR_REG_9_, n56 );
nand U9603 ( n1026, n4716, n4717 );
nor U9604 ( n4716, n4728, n3547 );
nor U9605 ( n4717, n4718, n4719 );
and U9606 ( n4728, ADDR_REG_6_, n56 );
xnor U9607 ( n3484, REG3_REG_22_, n4383 );
xnor U9608 ( n3203, REG3_REG_28_, n4329 );
nand U9609 ( n4338, REG3_REG_26_, n4347 );
nand U9610 ( n494, n2806, n2807 );
nand U9611 ( n2806, REG0_REG_0_, n5190 );
nand U9612 ( n2807, n5119, n1485 );
nand U9613 ( n654, n1483, n1484 );
nand U9614 ( n1483, REG1_REG_0_, n5194 );
nand U9615 ( n1484, n5122, n1485 );
xor U9616 ( n4799, REG1_REG_12_, n53 );
xor U9617 ( n3308, n4356, REG3_REG_25_ );
xor U9618 ( n3268, n4392, REG3_REG_21_ );
xor U9619 ( n3073, n4338, REG3_REG_27_ );
xor U9620 ( n3157, n4410, REG3_REG_19_ );
nand U9621 ( n1078, n4530, n4531 );
nand U9622 ( n4531, n5142, n1280 );
nand U9623 ( n4530, DATAO_REG_6_, n5140 );
nand U9624 ( n1098, n4485, n4486 );
nand U9625 ( n4486, n5142, n1176 );
nand U9626 ( n4485, DATAO_REG_11_, n5140 );
nand U9627 ( n1066, n4555, n4556 );
nand U9628 ( n4556, n5142, n1342 );
nand U9629 ( n4555, DATAO_REG_3_, n5140 );
nand U9630 ( n1070, n4547, n4548 );
nand U9631 ( n4548, n5142, n1324 );
nand U9632 ( n4547, DATAO_REG_4_, n5140 );
nand U9633 ( n1110, n4458, n4459 );
nand U9634 ( n4459, n5142, n1108 );
nand U9635 ( n4458, DATAO_REG_14_, n5140 );
nand U9636 ( n1082, n4521, n4522 );
nand U9637 ( n4522, n5142, n1260 );
nand U9638 ( n4521, DATAO_REG_7_, n5140 );
nand U9639 ( n1106, n4467, n4468 );
nand U9640 ( n4468, n5142, n1131 );
nand U9641 ( n4467, DATAO_REG_13_, n5140 );
nand U9642 ( n1090, n4503, n4504 );
nand U9643 ( n4504, n5142, n1214 );
nand U9644 ( n4503, DATAO_REG_9_, n5140 );
nand U9645 ( n1074, n4539, n4540 );
nand U9646 ( n4540, n5142, n1303 );
nand U9647 ( n4539, DATAO_REG_5_, n5140 );
nand U9648 ( n1118, n4440, n4441 );
nand U9649 ( n4441, n5142, n1063 );
nand U9650 ( n4440, DATAO_REG_16_, n5140 );
nand U9651 ( n1126, n4422, n4423 );
nand U9652 ( n4423, n5141, n1017 );
nand U9653 ( n4422, DATAO_REG_18_, n5140 );
nand U9654 ( n1062, n4563, n4564 );
nand U9655 ( n4564, n5142, n1359 );
nand U9656 ( n4563, DATAO_REG_2_, n5140 );
nand U9657 ( n1122, n4431, n4432 );
nand U9658 ( n4432, n5141, n1040 );
nand U9659 ( n4431, DATAO_REG_17_, n5140 );
nand U9660 ( n1102, n4476, n4477 );
nand U9661 ( n4477, n5142, n1153 );
nand U9662 ( n4476, DATAO_REG_12_, n5140 );
nand U9663 ( n1086, n4512, n4513 );
nand U9664 ( n4513, n5142, n1239 );
nand U9665 ( n4512, DATAO_REG_8_, n5140 );
nand U9666 ( n1114, n4449, n4450 );
nand U9667 ( n4450, n5142, n1080 );
nand U9668 ( n4449, DATAO_REG_15_, n5140 );
nand U9669 ( n1094, n4494, n4495 );
nand U9670 ( n4495, n5142, n1198 );
nand U9671 ( n4494, DATAO_REG_10_, n5140 );
nand U9672 ( n1058, n4571, n4572 );
nand U9673 ( n4572, n5142, n1375 );
nand U9674 ( n4571, DATAO_REG_1_, n5140 );
nand U9675 ( n1054, n4579, n4580 );
nand U9676 ( n4580, n5142, n2798 );
nand U9677 ( n4579, DATAO_REG_0_, n5140 );
xnor U9678 ( n3442, REG3_REG_20_, n4401 );
nand U9679 ( n1166, n4332, n4333 );
nand U9680 ( n4333, n5141, n811 );
nand U9681 ( n4332, DATAO_REG_28_, n5140 );
nand U9682 ( n1158, n4350, n4351 );
nand U9683 ( n4351, n5141, n851 );
nand U9684 ( n4350, DATAO_REG_26_, n4315 );
nand U9685 ( n1142, n4386, n4387 );
nand U9686 ( n4387, n5141, n931 );
nand U9687 ( n4386, DATAO_REG_22_, n4315 );
nand U9688 ( n1134, n4404, n4405 );
nand U9689 ( n4405, n5141, n972 );
nand U9690 ( n4404, DATAO_REG_20_, n4315 );
nand U9691 ( n1150, n4368, n4369 );
nand U9692 ( n4369, n5141, n891 );
nand U9693 ( n4368, DATAO_REG_24_, n4315 );
nand U9694 ( n1162, n4341, n4342 );
nand U9695 ( n4342, n5141, n832 );
nand U9696 ( n4341, DATAO_REG_27_, n4315 );
nand U9697 ( n1138, n4395, n4396 );
nand U9698 ( n4396, n5141, n952 );
nand U9699 ( n4395, DATAO_REG_21_, n4315 );
nand U9700 ( n1178, n4306, n4307 );
nand U9701 ( n4307, n5142, n1509 );
nand U9702 ( n4306, DATAO_REG_31_, n4315 );
nand U9703 ( n1154, n4359, n4360 );
nand U9704 ( n4360, n5141, n867 );
nand U9705 ( n4359, DATAO_REG_25_, n4315 );
nand U9706 ( n1146, n4377, n4378 );
nand U9707 ( n4378, n5141, n907 );
nand U9708 ( n4377, DATAO_REG_23_, n4315 );
nand U9709 ( n1130, n4413, n4414 );
nand U9710 ( n4414, n5141, n995 );
nand U9711 ( n4413, DATAO_REG_19_, n4315 );
nand U9712 ( n1174, n4316, n4317 );
nand U9713 ( n4317, n5141, n1534 );
nand U9714 ( n4316, DATAO_REG_30_, n4315 );
nand U9715 ( n1170, n4322, n4323 );
nand U9716 ( n4323, n5141, n786 );
nand U9717 ( n4322, DATAO_REG_29_, n4315 );
nand U9718 ( n766, n4329, REG3_REG_28_ );
nor U9719 ( n4641, n4697, n4589 );
xnor U9720 ( n4697, n4698, n4699 );
xor U9721 ( n4698, n4260, REG2_REG_4_ );
nor U9722 ( n4612, n4619, n4589 );
xnor U9723 ( n4619, n4620, n4621 );
xor U9724 ( n4620, n4263, REG2_REG_2_ );
nand U9725 ( n284, n2893, n2894 );
nand U9726 ( n2894, DATAI_22_, n5123 );
nor U9727 ( n2893, n2895, n2896 );
nor U9728 ( n2896, n5077, n5177 );
not U9729 ( n5248, STATE_REG );
nand U9730 ( n309, n2861, n2862 );
nand U9731 ( n2862, DATAI_27_, n5123 );
nor U9732 ( n2861, n2863, n2864 );
nor U9733 ( n2864, n4987, n5177 );
nand U9734 ( n274, n2905, n2906 );
nand U9735 ( n2906, DATAI_20_, n5123 );
nor U9736 ( n2905, n2907, n2908 );
nor U9737 ( n2908, n4985, n5177 );
nand U9738 ( n264, n2917, n2918 );
nand U9739 ( n2918, DATAI_18_, n5123 );
nor U9740 ( n2917, n2919, n2920 );
nor U9741 ( n2920, n4981, n5178 );
nand U9742 ( n324, n2841, n2842 );
nand U9743 ( n2842, DATAI_30_, n5123 );
nor U9744 ( n2841, n2843, n2844 );
nor U9745 ( n2844, n4988, n5177 );
nand U9746 ( n294, n2880, n2881 );
nand U9747 ( n2881, DATAI_24_, n5123 );
nor U9748 ( n2880, n2882, n2883 );
nor U9749 ( n2883, n4986, n5177 );
nand U9750 ( n254, n2929, n2930 );
nand U9751 ( n2930, DATAI_16_, n5124 );
nor U9752 ( n2929, n2931, n2932 );
nor U9753 ( n2932, n5034, n5178 );
nand U9754 ( n244, n2941, n2942 );
nand U9755 ( n2942, DATAI_14_, n5124 );
nor U9756 ( n2941, n2943, n2944 );
nor U9757 ( n2944, n4982, n5178 );
nand U9758 ( n234, n2953, n2954 );
nand U9759 ( n2954, DATAI_12_, n5124 );
nor U9760 ( n2953, n2955, n2956 );
nor U9761 ( n2956, n5017, n5178 );
nand U9762 ( n189, n3005, n3006 );
nand U9763 ( n3006, DATAI_3_, n5246 );
nor U9764 ( n3005, n3007, n3008 );
nor U9765 ( n3008, n4990, n5179 );
nand U9766 ( n204, n2989, n2990 );
nand U9767 ( n2990, DATAI_6_, n5124 );
nor U9768 ( n2989, n2991, n2992 );
nor U9769 ( n2992, n5000, n5179 );
nand U9770 ( n224, n2965, n2966 );
nand U9771 ( n2966, DATAI_10_, n5124 );
nor U9772 ( n2965, n2967, n2968 );
nor U9773 ( n2968, n5021, n5178 );
nand U9774 ( n214, n2977, n2978 );
nand U9775 ( n2978, DATAI_8_, n5124 );
nor U9776 ( n2977, n2979, n2980 );
nor U9777 ( n2980, n5014, n5178 );
nand U9778 ( n279, n2898, n2899 );
nand U9779 ( n2899, DATAI_21_, n5123 );
nor U9780 ( n2898, n2900, n2901 );
nor U9781 ( n2901, n4983, n5177 );
nand U9782 ( n259, n2922, n2923 );
nand U9783 ( n2923, DATAI_17_, n5124 );
nor U9784 ( n2922, n2924, n2925 );
nor U9785 ( n2925, n5080, n5178 );
nand U9786 ( n249, n2934, n2935 );
nand U9787 ( n2935, DATAI_15_, n5124 );
nor U9788 ( n2934, n2936, n2937 );
nor U9789 ( n2937, n4984, n5178 );
nand U9790 ( n319, n2848, n2849 );
nand U9791 ( n2849, DATAI_29_, n5123 );
nor U9792 ( n2848, n2850, n2851 );
nor U9793 ( n2851, n5087, n5177 );
nand U9794 ( n304, n2866, n2867 );
nand U9795 ( n2867, DATAI_26_, n5123 );
nor U9796 ( n2866, n2868, n2869 );
nor U9797 ( n2869, n5079, n5177 );
nand U9798 ( n314, n2854, n2855 );
nand U9799 ( n2855, DATAI_28_, n5123 );
nor U9800 ( n2854, n2856, n2857 );
nor U9801 ( n2857, n5081, n5177 );
nand U9802 ( n299, n2873, n2874 );
nand U9803 ( n2874, DATAI_25_, n5123 );
nor U9804 ( n2873, n2875, n2876 );
nor U9805 ( n2876, n5082, n5177 );
nand U9806 ( n289, n2885, n2886 );
nand U9807 ( n2886, DATAI_23_, n5123 );
nor U9808 ( n2885, n2887, n2888 );
nor U9809 ( n2888, n5063, n5177 );
nand U9810 ( n269, n2910, n2911 );
nand U9811 ( n2911, DATAI_19_, n5123 );
nor U9812 ( n2910, n2912, n2913 );
nor U9813 ( n2913, n5078, n5177 );
nand U9814 ( n239, n2946, n2947 );
nand U9815 ( n2947, DATAI_13_, n5124 );
nor U9816 ( n2946, n2948, n2949 );
nor U9817 ( n2949, n5083, n5178 );
nand U9818 ( n229, n2958, n2959 );
nand U9819 ( n2959, DATAI_11_, n5124 );
nor U9820 ( n2958, n2960, n2961 );
nor U9821 ( n2961, n5084, n5178 );
nand U9822 ( n219, n2970, n2971 );
nand U9823 ( n2971, DATAI_9_, n5124 );
nor U9824 ( n2970, n2972, n2973 );
nor U9825 ( n2973, n5085, n5178 );
nand U9826 ( n209, n2982, n2983 );
nand U9827 ( n2983, DATAI_7_, n5124 );
nor U9828 ( n2982, n2984, n2985 );
nor U9829 ( n2985, n5086, n5178 );
nand U9830 ( n194, n2999, n3000 );
nand U9831 ( n3000, DATAI_4_, n5124 );
nor U9832 ( n2999, n3001, n3002 );
nor U9833 ( n3002, n4980, n5179 );
nand U9834 ( n184, n3010, n3011 );
nand U9835 ( n3011, DATAI_2_, n5246 );
nor U9836 ( n3010, n3012, n3013 );
nor U9837 ( n3013, n5088, n5179 );
nand U9838 ( n334, n2833, n2834 );
nand U9839 ( n2834, n5181, n2835 );
nand U9840 ( n2833, D_REG_0_, n5180 );
nand U9841 ( n339, n2830, n2831 );
nand U9842 ( n2831, n5181, n2832 );
nand U9843 ( n2830, D_REG_1_, n5180 );
nand U9844 ( n4701, ADDR_REG_4_, n56 );
and U9845 ( n344, n5180, D_REG_2_ );
and U9846 ( n354, n5180, D_REG_4_ );
and U9847 ( n364, n5180, D_REG_6_ );
and U9848 ( n379, n5180, D_REG_9_ );
and U9849 ( n389, n5180, D_REG_11_ );
and U9850 ( n399, n5180, D_REG_13_ );
and U9851 ( n409, n5180, D_REG_15_ );
and U9852 ( n419, n5180, D_REG_17_ );
and U9853 ( n429, n5180, D_REG_19_ );
and U9854 ( n439, n5180, D_REG_21_ );
and U9855 ( n454, n5180, D_REG_24_ );
and U9856 ( n464, n5180, D_REG_26_ );
and U9857 ( n349, n5180, D_REG_3_ );
and U9858 ( n359, n5180, D_REG_5_ );
and U9859 ( n374, n5180, D_REG_8_ );
and U9860 ( n384, n5180, D_REG_10_ );
and U9861 ( n394, n5180, D_REG_12_ );
and U9862 ( n404, n5180, D_REG_14_ );
and U9863 ( n414, n5180, D_REG_16_ );
and U9864 ( n424, n5180, D_REG_18_ );
and U9865 ( n434, n5180, D_REG_20_ );
and U9866 ( n449, n5180, D_REG_23_ );
and U9867 ( n459, n5180, D_REG_25_ );
and U9868 ( n469, n5180, D_REG_27_ );
and U9869 ( n4594, ADDR_REG_0_, n56 );
and U9870 ( n4608, ADDR_REG_1_, n56 );
and U9871 ( n474, n5180, D_REG_28_ );
and U9872 ( n489, n5180, D_REG_31_ );
and U9873 ( n479, n5180, D_REG_29_ );
and U9874 ( n484, n5180, D_REG_30_ );
nand U9875 ( n174, n3022, n3023 );
nand U9876 ( n3022, DATAI_0_, n5246 );
nand U9877 ( n3023, IR_REG_0_, n3024 );
nand U9878 ( n3024, n5179, n5172 );
xor U9879 ( n4777, REG1_REG_10_, n54 );
xor U9880 ( n4763, n4764, n4765 );
xor U9881 ( n4765, n4219, REG2_REG_9_ );
nand U9882 ( n199, n2994, n2995 );
nand U9883 ( n2995, DATAI_5_, n5124 );
nor U9884 ( n2994, n2996, n2997 );
nor U9885 ( n2997, n5001, n5179 );
nand U9886 ( n179, n3017, n3018 );
nand U9887 ( n3018, DATAI_1_, n5246 );
nor U9888 ( n3017, n3019, n3020 );
nor U9889 ( n3020, n4989, n5179 );
nand U9890 ( n329, n2837, n2838 );
nand U9891 ( n2837, DATAI_31_, n5124 );
nand U9892 ( n2838, n2839, n5175 );
nor U9893 ( n2839, IR_REG_30_, n2840 );
xor U9894 ( n4752, REG1_REG_8_, n55 );
nand U9895 ( n3836, n3837, n3838 );
nor U9896 ( n3837, D_REG_4_, D_REG_3_ );
nor U9897 ( n3838, D_REG_6_, D_REG_5_ );
nor U9898 ( n3841, D_REG_17_, D_REG_16_ );
nand U9899 ( n3853, n3854, n3855 );
nor U9900 ( n3854, D_REG_26_, D_REG_25_ );
nor U9901 ( n3855, D_REG_28_, D_REG_27_ );
nor U9902 ( n3858, D_REG_13_, D_REG_12_ );
nor U9903 ( n3840, D_REG_15_, D_REG_14_ );
nand U9904 ( n3844, n3845, n3846 );
nor U9905 ( n3845, D_REG_2_, D_REG_29_ );
nor U9906 ( n3846, D_REG_31_, D_REG_30_ );
nor U9907 ( n3857, D_REG_11_, D_REG_10_ );
nor U9908 ( n3848, D_REG_9_, D_REG_8_ );
xor U9909 ( n4713, n4714, REG1_REG_5_ );
nor U9910 ( n4647, IR_REG_0_, n4648 );
nor U9911 ( n4648, n4649, n290 );
nor U9912 ( n4649, REG2_REG_0_, n4650 );
xor U9913 ( n4709, n4710, n4711 );
xor U9914 ( n4711, n4239, REG2_REG_5_ );
xnor U9915 ( n661, n695, REG2_REG_19_ );
xnor U9916 ( n700, n695, REG1_REG_19_ );
xor U9917 ( n4636, n4637, REG1_REG_3_ );
xor U9918 ( n641, n642, REG1_REG_18_ );
xor U9919 ( n622, n623, REG1_REG_17_ );
xor U9920 ( n4632, n4633, n4634 );
xor U9921 ( n4634, n4272, REG2_REG_3_ );
xor U9922 ( n551, n547, REG1_REG_13_ );
xor U9923 ( n4762, n4219, REG1_REG_9_ );
endmodule

