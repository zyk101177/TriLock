
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule



module b12_ori ( clk, reset, START, K_3_, K_2_, K_1_, K_0_, NLOSS_REG, NL_REG_3_,
NL_REG_2_, NL_REG_1_, NL_REG_0_, SPEAKER_REG );
input clk, reset, START, K_3_, K_2_, K_1_, K_0_;
output NLOSS_REG, NL_REG_3_, NL_REG_2_, NL_REG_1_, NL_REG_0_, SPEAKER_REG;
wire ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, n558, n563, n568, n596, n601, n606, n611, n616, n591, n586, n553,
n549, n535, n520, n515, n510, n505, n500, n480, n475, n470, n460,
n455, n445, n440, n435, n430, n410, n405, n400, n395, n390, n385,
n380, n375, n370, n365, n361, n357, n353, n349, n344, n339, n334,
n329, n324, n319, n314, n309, n304, n299, n294, n289, n284, n279,
n274, n269, n264, n259, n254, n249, n244, n239, n234, n229, n224,
n219, n214, n209, n204, n199, n194, n189, n184, n179, n174, n169,
n164, n159, n154, n149, n144, n139, n134, n129, n124, n119, n114,
n109, n104, n99, n94, n89, n84, n79, n74, n69, n64, n59, n54, n49,
n44, n39, n34, n29, GAMMA_REG_4_, GAMMA_REG_3_, GAMMA_REG_1_,
GAMMA_REG_2_, n573, n415, n420, n425, n450, n465, n485, n490, n495,
n525, n530, n540, n545, NUM_REG_1_, NUM_REG_0_, n1, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
n2145, n2146, n2147, n2148, n2149, n2150, n2151;

dff COUNT_REG_0__reg ( clk, reset, ex_wire0, n1 );
not U_inv0 ( n1, ex_wire0 );
dff COUNT_REG_1__reg ( clk, reset, ex_wire1, n573 );
not U_inv1 ( n2106, ex_wire1 );
dff NUM_REG_1__reg ( clk, reset, NUM_REG_1_, n573 );
dff NUM_REG_0__reg ( clk, reset, NUM_REG_0_, n1 );
dff GAMMA_REG_0__reg ( clk, reset, ex_wire2, n616 );
not U_inv2 ( n2117, ex_wire2 );
dff COUNT_REG2_4__reg ( clk, reset, n1102, n460 );
not U_inv3 ( n2115, n1102 );
dff MAX_REG_0__reg ( clk, reset, ex_wire3, n410 );
not U_inv4 ( n2132, ex_wire3 );
dff MAX_REG_1__reg ( clk, reset, ex_wire4, n405 );
not U_inv5 ( n2131, ex_wire4 );
dff MAX_REG_2__reg ( clk, reset, n1093, n400 );
not U_inv6 ( n2130, n1093 );
dff MAX_REG_3__reg ( clk, reset, n1089, n395 );
not U_inv7 ( n2129, n1089 );
dff MAX_REG_4__reg ( clk, reset, n1100, n390 );
not U_inv8 ( n2128, n1100 );
dff SCAN_REG_3__reg ( clk, reset, n1098, n370 );
not U_inv9 ( n2124, n1098 );
dff SCAN_REG_4__reg ( clk, reset, n1173, n365 );
not U_inv10 ( n2123, n1173 );
dff ADDRESS_REG_4__reg ( clk, reset, ex_wire5, n500 );
not U_inv11 ( n2145, ex_wire5 );
dff MEMORY_REG_24__0__reg ( clk, reset, n1171, n104 );
dff DATA_OUT_REG_0__reg ( clk, reset, n1083, n591 );
not U_inv12 ( n2151, n1083 );
dff GAMMA_REG_2__reg ( clk, reset, GAMMA_REG_2_, n606 );
dff SCAN_REG_0__reg ( clk, reset, ex_wire6, n385 );
not U_inv13 ( n2127, ex_wire6 );
dff SCAN_REG_1__reg ( clk, reset, n1099, n380 );
not U_inv14 ( n2126, n1099 );
dff SCAN_REG_2__reg ( clk, reset, n1088, n375 );
not U_inv15 ( n2125, n1088 );
dff GAMMA_REG_3__reg ( clk, reset, GAMMA_REG_3_, n601 );
dff GAMMA_REG_1__reg ( clk, reset, GAMMA_REG_1_, n611 );
dff IND_REG_0__reg ( clk, reset, n1091, n420 );
not U_inv16 ( n2133, n1091 );
dff IND_REG_1__reg ( clk, reset, n1084, n415 );
dff GAMMA_REG_4__reg ( clk, reset, GAMMA_REG_4_, n596 );
dff DATA_IN_REG_0__reg ( clk, reset, ex_wire7, n530 );
not U_inv17 ( n2122, ex_wire7 );
dff DATA_IN_REG_1__reg ( clk, reset, ex_wire8, n525 );
not U_inv18 ( n2118, ex_wire8 );
dff WR_REG_reg ( clk, reset, ex_wire9, n553 );
not U_inv19 ( n2121, ex_wire9 );
dff MEMORY_REG_24__1__reg ( clk, reset, n1116, n99 );
dff ADDRESS_REG_0__reg ( clk, reset, n1096, n520 );
not U_inv20 ( n2147, n1096 );
dff ADDRESS_REG_1__reg ( clk, reset, n1085, n515 );
not U_inv21 ( n2119, n1085 );
dff ADDRESS_REG_2__reg ( clk, reset, n1087, n510 );
not U_inv22 ( n2120, n1087 );
dff MEMORY_REG_25__0__reg ( clk, reset, n1111, n94 );
dff MEMORY_REG_25__1__reg ( clk, reset, n1115, n89 );
dff MEMORY_REG_28__0__reg ( clk, reset, n1108, n64 );
dff MEMORY_REG_28__1__reg ( clk, reset, n1112, n59 );
dff MEMORY_REG_29__0__reg ( clk, reset, n1117, n54 );
dff MEMORY_REG_29__1__reg ( clk, reset, n1118, n49 );
dff ADDRESS_REG_3__reg ( clk, reset, n1092, n505 );
not U_inv23 ( n2146, n1092 );
dff MEMORY_REG_27__0__reg ( clk, reset, n1110, n74 );
dff MEMORY_REG_27__1__reg ( clk, reset, n1114, n69 );
dff MEMORY_REG_26__0__reg ( clk, reset, n1109, n84 );
dff MEMORY_REG_26__1__reg ( clk, reset, n1113, n79 );
dff MEMORY_REG_30__0__reg ( clk, reset, n1119, n44 );
dff MEMORY_REG_30__1__reg ( clk, reset, n1120, n39 );
dff MEMORY_REG_31__0__reg ( clk, reset, n1122, n34 );
dff MEMORY_REG_31__1__reg ( clk, reset, n1133, n29 );
dff MEMORY_REG_0__0__reg ( clk, reset, n1121, n344 );
dff MEMORY_REG_0__1__reg ( clk, reset, n1123, n339 );
dff MEMORY_REG_1__0__reg ( clk, reset, n1124, n334 );
dff MEMORY_REG_1__1__reg ( clk, reset, n1125, n329 );
dff MEMORY_REG_4__0__reg ( clk, reset, n1130, n304 );
dff MEMORY_REG_4__1__reg ( clk, reset, n1131, n299 );
dff MEMORY_REG_5__0__reg ( clk, reset, n1132, n294 );
dff MEMORY_REG_5__1__reg ( clk, reset, n1134, n289 );
dff MEMORY_REG_10__0__reg ( clk, reset, n1143, n244 );
dff MEMORY_REG_10__1__reg ( clk, reset, n1144, n239 );
dff MEMORY_REG_11__0__reg ( clk, reset, n1145, n234 );
dff MEMORY_REG_11__1__reg ( clk, reset, n1146, n229 );
dff MEMORY_REG_14__0__reg ( clk, reset, n1151, n204 );
dff MEMORY_REG_14__1__reg ( clk, reset, n1152, n199 );
dff MEMORY_REG_15__0__reg ( clk, reset, n1153, n194 );
dff MEMORY_REG_15__1__reg ( clk, reset, n1154, n189 );
dff MEMORY_REG_2__0__reg ( clk, reset, n1126, n324 );
dff MEMORY_REG_2__1__reg ( clk, reset, n1127, n319 );
dff MEMORY_REG_3__0__reg ( clk, reset, n1128, n314 );
dff MEMORY_REG_3__1__reg ( clk, reset, n1129, n309 );
dff MEMORY_REG_6__0__reg ( clk, reset, n1135, n284 );
dff MEMORY_REG_6__1__reg ( clk, reset, n1136, n279 );
dff MEMORY_REG_7__0__reg ( clk, reset, n1137, n274 );
dff MEMORY_REG_7__1__reg ( clk, reset, n1138, n269 );
dff MEMORY_REG_8__0__reg ( clk, reset, n1139, n264 );
dff MEMORY_REG_8__1__reg ( clk, reset, n1140, n259 );
dff MEMORY_REG_9__0__reg ( clk, reset, n1141, n254 );
dff MEMORY_REG_9__1__reg ( clk, reset, n1142, n249 );
dff MEMORY_REG_12__0__reg ( clk, reset, n1147, n224 );
dff MEMORY_REG_12__1__reg ( clk, reset, n1148, n219 );
dff MEMORY_REG_13__0__reg ( clk, reset, n1149, n214 );
dff MEMORY_REG_13__1__reg ( clk, reset, n1150, n209 );
dff MEMORY_REG_16__0__reg ( clk, reset, n1155, n184 );
dff MEMORY_REG_16__1__reg ( clk, reset, n1156, n179 );
dff MEMORY_REG_17__0__reg ( clk, reset, n1157, n174 );
dff MEMORY_REG_17__1__reg ( clk, reset, n1158, n169 );
dff MEMORY_REG_20__0__reg ( clk, reset, n1163, n144 );
dff MEMORY_REG_20__1__reg ( clk, reset, n1164, n139 );
dff MEMORY_REG_21__0__reg ( clk, reset, n1165, n134 );
dff MEMORY_REG_21__1__reg ( clk, reset, n1166, n129 );
dff MEMORY_REG_18__0__reg ( clk, reset, n1159, n164 );
dff MEMORY_REG_18__1__reg ( clk, reset, n1160, n159 );
dff MEMORY_REG_19__0__reg ( clk, reset, n1161, n154 );
dff MEMORY_REG_19__1__reg ( clk, reset, n1162, n149 );
dff MEMORY_REG_22__0__reg ( clk, reset, n1167, n124 );
dff MEMORY_REG_22__1__reg ( clk, reset, n1168, n119 );
dff MEMORY_REG_23__0__reg ( clk, reset, n1169, n114 );
dff MEMORY_REG_23__1__reg ( clk, reset, n1170, n109 );
dff DATA_OUT_REG_1__reg ( clk, reset, n1090, n586 );
not U_inv24 ( n2150, n1090 );
dff SOUND_REG_2__reg ( clk, reset, n1097, n485 );
not U_inv25 ( n2143, n1097 );
dff SOUND_REG_1__reg ( clk, reset, n1086, n490 );
not U_inv26 ( n2144, n1086 );
dff NLOSS_REG_reg ( clk, reset, NLOSS_REG, n545 );
dff SOUND_REG_0__reg ( clk, reset, n1094, n495 );
dff TIMEBASE_REG_0__reg ( clk, reset, n1106, n450 );
not U_inv27 ( n2139, n1106 );
dff COUNT_REG2_0__reg ( clk, reset, ex_wire10, n480 );
not U_inv28 ( n2116, ex_wire10 );
dff TIMEBASE_REG_1__reg ( clk, reset, n1107, n445 );
not U_inv29 ( n2138, n1107 );
dff COUNT_REG2_1__reg ( clk, reset, ex_wire11, n475 );
not U_inv30 ( n2142, ex_wire11 );
dff TIMEBASE_REG_2__reg ( clk, reset, n1105, n440 );
not U_inv31 ( n2137, n1105 );
dff COUNT_REG2_2__reg ( clk, reset, ex_wire12, n470 );
not U_inv32 ( n2141, ex_wire12 );
dff TIMEBASE_REG_3__reg ( clk, reset, n1104, n435 );
not U_inv33 ( n2136, n1104 );
dff COUNT_REG2_3__reg ( clk, reset, n1103, n465 );
not U_inv34 ( n2114, n1103 );
dff TIMEBASE_REG_4__reg ( clk, reset, ex_wire13, n430 );
not U_inv35 ( n2135, ex_wire13 );
dff TIMEBASE_REG_5__reg ( clk, reset, n1095, n425 );
not U_inv36 ( n2134, n1095 );
dff COUNT_REG2_5__reg ( clk, reset, n1174, n455 );
not U_inv37 ( n2140, n1174 );
dff PLAY_REG_reg ( clk, reset, ex_wire14, n540 );
not U_inv38 ( n2148, ex_wire14 );
dff COUNTER_REG_0__reg ( clk, reset, ex_wire15, n568 );
not U_inv39 ( n2149, ex_wire15 );
dff COUNTER_REG_1__reg ( clk, reset, n1101, n563 );
not U_inv40 ( n2109, n1101 );
dff COUNTER_REG_2__reg ( clk, reset, n1172, n558 );
dff SPEAKER_REG_reg ( clk, reset, SPEAKER_REG, n549 );
not U_inv41 ( n2107, SPEAKER_REG );
dff S_REG_reg ( clk, reset, ex_wire16, n535 );
not U_inv42 ( n2108, ex_wire16 );
dff NL_REG_0__reg ( clk, reset, NL_REG_0_, n361 );
not U_inv43 ( n2110, NL_REG_0_ );
dff NL_REG_1__reg ( clk, reset, NL_REG_1_, n357 );
not U_inv44 ( n2111, NL_REG_1_ );
dff NL_REG_2__reg ( clk, reset, NL_REG_2_, n353 );
not U_inv45 ( n2112, NL_REG_2_ );
dff NL_REG_3__reg ( clk, reset, NL_REG_3_, n349 );
not U_inv46 ( n2113, NL_REG_3_ );
not U1085 ( n1187, n2121 );
nor U1086 ( n1183, n2122, n2121 );
nor U1087 ( n1178, n2121, n2118 );
nand U1088 ( n99, n1175, n1176 );
nand U1089 ( n1176, n1177, n1116 );
nand U1090 ( n1175, n1178, n1179 );
nand U1091 ( n94, n1180, n1181 );
nand U1092 ( n1181, n1182, n1111 );
nand U1093 ( n1180, n1183, n1184 );
nand U1094 ( n89, n1185, n1186 );
nand U1095 ( n1186, n1182, n1115 );
nand U1096 ( n1182, n1184, n1187 );
nand U1097 ( n1185, n1184, n1178 );
nand U1098 ( n84, n1188, n1189 );
nand U1099 ( n1189, n1190, n1109 );
nand U1100 ( n1188, n1191, n1183 );
nand U1101 ( n79, n1192, n1193 );
nand U1102 ( n1193, n1190, n1113 );
nand U1103 ( n1190, n1191, n1187 );
nand U1104 ( n1192, n1191, n1178 );
nand U1105 ( n74, n1194, n1195 );
nand U1106 ( n1195, n1196, n1110 );
nand U1107 ( n1194, n1197, n1183 );
nand U1108 ( n69, n1198, n1199 );
nand U1109 ( n1199, n1196, n1114 );
nand U1110 ( n1196, n1197, n1187 );
nand U1111 ( n1198, n1197, n1178 );
nand U1112 ( n64, n1200, n1201 );
nand U1113 ( n1201, n1202, n1108 );
nand U1114 ( n1200, n1203, n1183 );
nand U1115 ( n616, n1204, n1205 );
nor U1116 ( n1205, n1206, n1207 );
nand U1117 ( n1207, n1208, n1209 );
nor U1118 ( n1206, n1210, n1211 );
nand U1119 ( n1211, n1212, n1213 );
nor U1120 ( n1204, n1214, n1215 );
nand U1121 ( n1215, n1216, n1217 );
nand U1122 ( n1217, n1218, n1219 );
nand U1123 ( n1218, n1220, n1221 );
nor U1124 ( n1221, n1222, n1223 );
nor U1125 ( n1223, n1224, n1225 );
nand U1126 ( n1225, n1226, n1227 );
nand U1127 ( n1227, n1228, n1090 );
nand U1128 ( n1228, n1229, n1230 );
nor U1129 ( n1229, n1231, n1232 );
nor U1130 ( n1232, K_2_, n1233 );
nor U1131 ( n1233, n2151, n1234 );
nor U1132 ( n1231, n2151, n1235 );
nand U1133 ( n1226, n1236, n2150 );
nand U1134 ( n1236, n1237, n1238 );
nand U1135 ( n1238, n2151, n1239 );
nand U1136 ( n1237, n1240, n1083 );
nand U1137 ( n1240, K_1_, n1239 );
nor U1138 ( n1220, n1241, n1242 );
nand U1139 ( n1216, n1243, n1244 );
nand U1140 ( n1244, n1245, n1246 );
nor U1141 ( n1245, n1247, n1248 );
nand U1142 ( n611, n1249, n1250 );
nor U1143 ( n1250, n1251, n1252 );
nand U1144 ( n1252, n1253, n1254 );
nand U1145 ( n1251, n1255, n1256 );
nor U1146 ( n1249, n1257, n1258 );
nand U1147 ( n1258, n1259, n1260 );
nand U1148 ( n1260, n1261, n1262 );
not U1149 ( n1259, n1214 );
nand U1150 ( n1214, n1263, n1264 );
or U1151 ( n1264, n1265, n1266 );
nor U1152 ( n1263, n1267, n1268 );
nor U1153 ( n1268, n1269, n1270 );
nand U1154 ( n1257, n1271, n1272 );
nand U1155 ( n1272, n1212, n1273 );
nand U1156 ( n1271, n1274, n1275 );
nand U1157 ( n606, n1276, n1277 );
nor U1158 ( n1277, n1278, n1279 );
nand U1159 ( n1279, n1280, n1281 );
nand U1160 ( n1281, n1282, n1283 );
nand U1161 ( n1280, n1284, n1285 );
nand U1162 ( n1278, n1286, n1209 );
nand U1163 ( n1209, n1287, n1288 );
nor U1164 ( n1287, n1289, n1213 );
nor U1165 ( n1286, n1222, n1267 );
not U1166 ( n1267, n1290 );
nor U1167 ( n1276, n1291, n1292 );
nand U1168 ( n1292, n1293, n1294 );
not U1169 ( n1294, n1248 );
nand U1170 ( n1248, n1295, n1296 );
nand U1171 ( n1295, n1212, n1297 );
nand U1172 ( n1291, n1298, n1299 );
or U1173 ( n1299, n1270, n1243 );
nand U1174 ( n1298, n1300, n1213 );
nand U1175 ( n601, n1301, n1302 );
nor U1176 ( n1302, n1303, n1304 );
nand U1177 ( n1304, n1305, n1253 );
nand U1178 ( n1305, n1306, n1307 );
nor U1179 ( n1306, n1297, n1308 );
and U1180 ( n1308, n1309, n1310 );
nand U1181 ( n1303, n1290, n1311 );
nand U1182 ( n1290, n1312, n1313 );
nand U1183 ( n1313, n1265, n1314 );
nand U1184 ( n1314, n1300, n1219 );
nor U1185 ( n1301, n1315, n1316 );
nand U1186 ( n1316, n1296, n1317 );
nand U1187 ( n1317, n1318, n1319 );
nand U1188 ( n1319, n1269, n1320 );
nand U1189 ( n1296, n1312, n1285 );
nor U1190 ( n1315, n1270, n1321 );
nand U1191 ( n596, n1322, n1323 );
and U1192 ( n1323, n1324, n1210 );
nor U1193 ( n1322, n1325, n1326 );
nor U1194 ( n1326, n1219, n1224 );
nor U1195 ( n1325, n1327, n1328 );
nand U1196 ( n591, n1329, n1330 );
nor U1197 ( n1330, n1331, n1332 );
nand U1198 ( n1332, n1333, n1334 );
nor U1199 ( n1334, n1335, n1336 );
nand U1200 ( n1336, n1337, n1338 );
nand U1201 ( n1338, n1339, n1130 );
nand U1202 ( n1337, n1340, n1122 );
nand U1203 ( n1335, n1341, n1342 );
nand U1204 ( n1342, n1343, n1126 );
nand U1205 ( n1341, n1344, n1128 );
nor U1206 ( n1333, n1345, n1346 );
nand U1207 ( n1346, n1347, n1348 );
nand U1208 ( n1348, n1349, n1137 );
nand U1209 ( n1347, n1350, n1139 );
nand U1210 ( n1345, n1351, n1352 );
nand U1211 ( n1352, n1353, n1132 );
nand U1212 ( n1351, n1354, n1135 );
nand U1213 ( n1331, n1355, n1356 );
nor U1214 ( n1356, n1357, n1358 );
nand U1215 ( n1358, n1359, n1360 );
nand U1216 ( n1360, n1203, n1108 );
nand U1217 ( n1359, n1191, n1109 );
nand U1218 ( n1357, n1361, n1362 );
nand U1219 ( n1362, n1197, n1110 );
nand U1220 ( n1361, n1184, n1111 );
nor U1221 ( n1355, n1363, n1364 );
nand U1222 ( n1364, n1365, n1366 );
nand U1223 ( n1366, n1367, n1121 );
nand U1224 ( n1365, n1368, n1124 );
nand U1225 ( n1363, n1369, n1370 );
nand U1226 ( n1370, n1371, n1117 );
nand U1227 ( n1369, n1372, n1119 );
nor U1228 ( n1329, n1373, n1374 );
nand U1229 ( n1374, n1375, n1376 );
nor U1230 ( n1376, n1377, n1378 );
nand U1231 ( n1378, n1379, n1380 );
nand U1232 ( n1380, n1381, n1161 );
nand U1233 ( n1379, n1382, n1163 );
nand U1234 ( n1377, n1383, n1384 );
nand U1235 ( n1384, n1385, n1157 );
nand U1236 ( n1383, n1386, n1159 );
nor U1237 ( n1375, n1387, n1388 );
nand U1238 ( n1388, n1389, n1390 );
nand U1239 ( n1390, n1391, n1169 );
nand U1240 ( n1389, n1179, n1171 );
nand U1241 ( n1387, n1392, n1393 );
nand U1242 ( n1393, n1394, n1165 );
nand U1243 ( n1392, n1395, n1167 );
nand U1244 ( n1373, n1396, n1397 );
nor U1245 ( n1397, n1398, n1399 );
nand U1246 ( n1399, n1400, n1401 );
nand U1247 ( n1401, n1402, n1145 );
nand U1248 ( n1400, n1403, n1147 );
nand U1249 ( n1398, n1404, n1405 );
nand U1250 ( n1405, n1406, n1141 );
nand U1251 ( n1404, n1407, n1143 );
nor U1252 ( n1396, n1408, n1409 );
nand U1253 ( n1409, n1410, n1411 );
nand U1254 ( n1411, n1412, n1153 );
nand U1255 ( n1410, n1413, n1155 );
nand U1256 ( n1408, n1414, n1415 );
nand U1257 ( n1415, n1416, n1149 );
nand U1258 ( n1414, n1417, n1151 );
nand U1259 ( n59, n1418, n1419 );
nand U1260 ( n1419, n1202, n1112 );
nand U1261 ( n1202, n1203, n1187 );
nand U1262 ( n1418, n1203, n1178 );
nand U1263 ( n586, n1420, n1421 );
nor U1264 ( n1421, n1422, n1423 );
nand U1265 ( n1423, n1424, n1425 );
nor U1266 ( n1425, n1426, n1427 );
nand U1267 ( n1427, n1428, n1429 );
nand U1268 ( n1429, n1339, n1131 );
nand U1269 ( n1428, n1340, n1133 );
nand U1270 ( n1426, n1430, n1431 );
nand U1271 ( n1431, n1343, n1127 );
nand U1272 ( n1430, n1344, n1129 );
nor U1273 ( n1424, n1432, n1433 );
nand U1274 ( n1433, n1434, n1435 );
nand U1275 ( n1435, n1349, n1138 );
nand U1276 ( n1434, n1350, n1140 );
nand U1277 ( n1432, n1436, n1437 );
nand U1278 ( n1437, n1353, n1134 );
nand U1279 ( n1436, n1354, n1136 );
nand U1280 ( n1422, n1438, n1439 );
nor U1281 ( n1439, n1440, n1441 );
nand U1282 ( n1441, n1442, n1443 );
nand U1283 ( n1443, n1203, n1112 );
and U1284 ( n1203, n1444, n1445 );
nand U1285 ( n1442, n1191, n1113 );
and U1286 ( n1191, n1446, n1447 );
nand U1287 ( n1440, n1448, n1449 );
nand U1288 ( n1449, n1197, n1114 );
and U1289 ( n1197, n1446, n1450 );
nand U1290 ( n1448, n1184, n1115 );
and U1291 ( n1184, n1450, n1445 );
nor U1292 ( n1438, n1451, n1452 );
nand U1293 ( n1452, n1453, n1454 );
nand U1294 ( n1454, n1367, n1123 );
nand U1295 ( n1453, n1368, n1125 );
nand U1296 ( n1451, n1455, n1456 );
nand U1297 ( n1456, n1371, n1118 );
nand U1298 ( n1455, n1372, n1120 );
nor U1299 ( n1420, n1457, n1458 );
nand U1300 ( n1458, n1459, n1460 );
nor U1301 ( n1460, n1461, n1462 );
nand U1302 ( n1462, n1463, n1464 );
nand U1303 ( n1464, n1381, n1162 );
nand U1304 ( n1463, n1382, n1164 );
nand U1305 ( n1461, n1465, n1466 );
nand U1306 ( n1466, n1385, n1158 );
nand U1307 ( n1465, n1386, n1160 );
nor U1308 ( n1459, n1467, n1468 );
nand U1309 ( n1468, n1469, n1470 );
nand U1310 ( n1470, n1391, n1170 );
nand U1311 ( n1469, n1179, n1116 );
nand U1312 ( n1467, n1471, n1472 );
nand U1313 ( n1472, n1394, n1166 );
nand U1314 ( n1471, n1395, n1168 );
nand U1315 ( n1457, n1473, n1474 );
nor U1316 ( n1474, n1475, n1476 );
nand U1317 ( n1476, n1477, n1478 );
nand U1318 ( n1478, n1402, n1146 );
nand U1319 ( n1477, n1403, n1148 );
nand U1320 ( n1475, n1479, n1480 );
nand U1321 ( n1480, n1406, n1142 );
nand U1322 ( n1479, n1407, n1144 );
nor U1323 ( n1473, n1481, n1482 );
nand U1324 ( n1482, n1483, n1484 );
nand U1325 ( n1484, n1412, n1154 );
nand U1326 ( n1483, n1413, n1156 );
nand U1327 ( n1481, n1485, n1486 );
nand U1328 ( n1486, n1416, n1150 );
nand U1329 ( n1485, n1417, n1152 );
xor U1330 ( n573, n2106, n1 );
nand U1331 ( n563, n1487, n1488 );
nand U1332 ( n1488, n568, n1101 );
and U1333 ( n568, n1489, n2149 );
nand U1334 ( n1487, n1490, n2109 );
nor U1335 ( n1490, n2149, n1491 );
nor U1336 ( n558, n1492, n1491 );
not U1337 ( n1491, n1489 );
nor U1338 ( n1489, n1493, n1494 );
or U1339 ( n1493, n2148, n1495 );
nor U1340 ( n1495, n2143, n2144 );
nor U1341 ( n1492, n1496, n1172 );
nor U1342 ( n1496, n2109, n2149 );
nand U1343 ( n553, n1497, n1498 );
nand U1344 ( n1498, n1499, n1187 );
nand U1345 ( n1499, n1500, n1275 );
nor U1346 ( n1500, n1501, n1307 );
nand U1347 ( n549, n1502, n1503 );
nand U1348 ( n1503, n1504, n1505 );
nor U1349 ( n1504, n2107, n2148 );
nand U1350 ( n545, n1506, n1507 );
nand U1351 ( n1507, n1508, NLOSS_REG );
not U1352 ( n1508, n1509 );
nand U1353 ( n1506, n1307, n1509 );
nand U1354 ( n1509, n1510, n1511 );
nand U1355 ( n1511, n1512, n1513 );
or U1356 ( n1513, n1283, n1243 );
nand U1357 ( n1283, n1514, n1515 );
nor U1358 ( n1515, n1516, n1517 );
nor U1359 ( n1517, n2151, n1239 );
not U1360 ( n1239, K_0_ );
nor U1361 ( n1516, K_0_, n1518 );
nand U1362 ( n1518, n2151, K_1_ );
nor U1363 ( n1514, n1519, n1520 );
nor U1364 ( n1520, n1521, n1522 );
not U1365 ( n1522, n1230 );
nor U1366 ( n1521, n1523, n1524 );
nand U1367 ( n1524, n1525, n1526 );
nand U1368 ( n1526, n1527, n1235 );
nor U1369 ( n1527, n1083, n1234 );
not U1370 ( n1234, K_3_ );
nand U1371 ( n1525, K_2_, n1083 );
nor U1372 ( n1523, n1528, n1090 );
nor U1373 ( n1519, n2150, n1230 );
nand U1374 ( n540, n1529, n1530 );
or U1375 ( n1530, n1531, n2148 );
nand U1376 ( n1529, n1532, n1531 );
nand U1377 ( n1531, n1533, n1534 );
nor U1378 ( n1534, n1535, n1536 );
nor U1379 ( n1536, n1310, n1328 );
nor U1380 ( n1310, n1300, n1285 );
nor U1381 ( n1535, n1537, n1538 );
nand U1382 ( n1538, n1212, n1539 );
nor U1383 ( n1533, n1540, n1541 );
nand U1384 ( n1532, n1542, n1543 );
nand U1385 ( n1543, n1544, n1210 );
nand U1386 ( n1544, n1224, n1545 );
nor U1387 ( n1542, n1546, n1547 );
nor U1388 ( n1547, n1307, n1548 );
nor U1389 ( n1548, n1549, n1300 );
nor U1390 ( n1549, n1501, n1213 );
nor U1391 ( n1546, n1311, n1550 );
nand U1392 ( n1550, n1274, n1213 );
nand U1393 ( n54, n1551, n1552 );
nand U1394 ( n1552, n1553, n1117 );
nand U1395 ( n1551, n1371, n1183 );
nand U1396 ( n535, n1502, n1554 );
or U1397 ( n1554, n1555, n2108 );
nand U1398 ( n1502, n2108, n1555 );
nor U1399 ( n1555, n1505, n2148 );
nand U1400 ( n1505, n1494, n1556 );
nand U1401 ( n1556, n1086, n1097 );
nand U1402 ( n1494, n1557, n1558 );
nand U1403 ( n1558, n1559, n1560 );
nor U1404 ( n1560, n1561, n1562 );
nor U1405 ( n1562, n1563, n1097 );
nor U1406 ( n1563, n2149, n1094 );
nor U1407 ( n1559, n2109, n1086 );
nand U1408 ( n1557, n1564, n1172 );
nand U1409 ( n1564, n1565, n1566 );
nand U1410 ( n1566, n1567, n1101 );
nand U1411 ( n1567, n2149, n2144 );
nor U1412 ( n1565, n1568, n1569 );
nor U1413 ( n1569, n2144, n1570 );
or U1414 ( n1570, n1094, n2149 );
nor U1415 ( n1568, n1561, n1086 );
nor U1416 ( n1561, n2143, n1094 );
nand U1417 ( n530, n1571, n1572 );
nand U1418 ( n1572, n1573, NUM_REG_0_ );
or U1419 ( n1571, n1573, n2122 );
nand U1420 ( n525, n1574, n1575 );
nand U1421 ( n1575, n1573, NUM_REG_1_ );
or U1422 ( n1574, n1573, n2118 );
not U1423 ( n1573, n1497 );
nand U1424 ( n520, n1576, n1577 );
nand U1425 ( n1577, n1578, n1096 );
nor U1426 ( n1576, n1579, n1580 );
nor U1427 ( n1580, n2132, n1581 );
nor U1428 ( n1579, n2127, n1582 );
nand U1429 ( n515, n1583, n1584 );
nand U1430 ( n1584, n1578, n1085 );
nor U1431 ( n1583, n1585, n1586 );
nor U1432 ( n1586, n2131, n1581 );
nor U1433 ( n1585, n2126, n1582 );
nand U1434 ( n510, n1587, n1588 );
nand U1435 ( n1588, n1578, n1087 );
nor U1436 ( n1587, n1589, n1590 );
nor U1437 ( n1590, n2130, n1581 );
nor U1438 ( n1589, n2125, n1582 );
nand U1439 ( n505, n1591, n1592 );
nand U1440 ( n1592, n1578, n1092 );
not U1441 ( n1578, n1593 );
nor U1442 ( n1591, n1594, n1595 );
nor U1443 ( n1595, n2129, n1581 );
nor U1444 ( n1594, n2124, n1582 );
nand U1445 ( n500, n1596, n1597 );
or U1446 ( n1597, n1593, n2145 );
nor U1447 ( n1596, n1598, n1599 );
nor U1448 ( n1599, n2128, n1581 );
nand U1449 ( n1581, n1593, n1600 );
nand U1450 ( n1600, n1309, n1265 );
nor U1451 ( n1598, n2123, n1582 );
nand U1452 ( n1582, n1593, n1601 );
nand U1453 ( n1601, n1539, n1327 );
nand U1454 ( n1593, n1602, n1603 );
nand U1455 ( n1603, n1604, n1210 );
nor U1456 ( n1602, n1605, n1606 );
nor U1457 ( n1606, n1309, n1607 );
not U1458 ( n1605, n1208 );
nand U1459 ( n1208, n1608, n1275 );
nor U1460 ( n1608, n1539, n1609 );
nand U1461 ( n495, n1610, n1611 );
nand U1462 ( n1611, n1612, n1094 );
nand U1463 ( n1610, n1613, n1614 );
nand U1464 ( n1613, n1615, n1616 );
nand U1465 ( n1616, n1539, n1083 );
nor U1466 ( n1615, n1284, n1617 );
nor U1467 ( n1617, n1273, n1618 );
or U1468 ( n1618, n1619, K_0_ );
nand U1469 ( n490, n1620, n1621 );
nand U1470 ( n1621, n1612, n1086 );
nand U1471 ( n1620, n1622, n1614 );
nand U1472 ( n1622, n1623, n1624 );
nand U1473 ( n1624, n1625, n1090 );
nand U1474 ( n1625, n1626, n1627 );
nand U1475 ( n1623, n1230, n1275 );
nand U1476 ( n49, n1628, n1629 );
nand U1477 ( n1629, n1553, n1118 );
nand U1478 ( n1553, n1371, n1187 );
nand U1479 ( n1628, n1371, n1178 );
and U1480 ( n1371, n1630, n1445 );
nand U1481 ( n485, n1631, n1632 );
nand U1482 ( n1632, n1612, n1097 );
nand U1483 ( n1631, n1633, n1614 );
not U1484 ( n1614, n1612 );
nor U1485 ( n1612, n1634, n1540 );
nand U1486 ( n1540, n1635, n1636 );
and U1487 ( n1636, n1255, n1637 );
nor U1488 ( n1635, n1638, n1639 );
nor U1489 ( n1639, n1545, n1640 );
nand U1490 ( n1640, n1641, n1269 );
nand U1491 ( n1545, n1274, n1297 );
or U1492 ( n1634, n1642, n1643 );
nor U1493 ( n1643, n1644, n1219 );
nor U1494 ( n1644, n1241, n1645 );
nor U1495 ( n1645, n1327, n1210 );
nor U1496 ( n1241, n1501, n1311 );
nand U1497 ( n1633, n1646, n1647 );
nand U1498 ( n1647, n1648, n1266 );
nand U1499 ( n480, n1649, n1650 );
nor U1500 ( n1649, n1651, n1652 );
nor U1501 ( n1652, n1653, n1654 );
nor U1502 ( n1654, n1655, n1656 );
nor U1503 ( n1656, n1657, n1658 );
nor U1504 ( n1655, n2139, n1659 );
nor U1505 ( n1651, n2116, n1660 );
nand U1506 ( n475, n1661, n1662 );
or U1507 ( n1662, n1660, n2142 );
nor U1508 ( n1661, n1663, n1664 );
nor U1509 ( n1664, n1665, n1666 );
not U1510 ( n1665, n1667 );
nor U1511 ( n1663, n2138, n1668 );
nand U1512 ( n470, n1669, n1670 );
or U1513 ( n1670, n1660, n2141 );
nor U1514 ( n1669, n1671, n1672 );
nor U1515 ( n1672, n1673, n1666 );
not U1516 ( n1673, n1674 );
nor U1517 ( n1671, n2137, n1668 );
nand U1518 ( n465, n1675, n1676 );
nand U1519 ( n1676, n1653, n1103 );
nand U1520 ( n1675, n1677, n1660 );
nand U1521 ( n1677, n1678, n1679 );
nand U1522 ( n1679, n1680, n1681 );
nor U1523 ( n1678, n1682, n1683 );
nor U1524 ( n1683, n2136, n1684 );
nor U1525 ( n1684, n1685, n1686 );
nand U1526 ( n1686, n1537, n1627 );
nor U1527 ( n1682, n1687, n1219 );
nor U1528 ( n1687, n1688, n1689 );
nor U1529 ( n1688, n1690, n1262 );
nand U1530 ( n460, n1691, n1692 );
nand U1531 ( n1692, n1653, n1102 );
nor U1532 ( n1691, n1693, n1694 );
nor U1533 ( n1694, n1666, n1695 );
not U1534 ( n1695, n1696 );
nand U1535 ( n1666, n1681, n1660 );
nand U1536 ( n1681, n1697, n1698 );
nand U1537 ( n1698, n1699, n1289 );
nor U1538 ( n1697, n1700, n1701 );
nor U1539 ( n1701, n1213, n1702 );
nand U1540 ( n1702, n1219, n1309 );
nor U1541 ( n1693, n2135, n1668 );
nand U1542 ( n1668, n1703, n1660 );
or U1543 ( n1703, n1685, n1704 );
or U1544 ( n1685, n1705, n1706 );
or U1545 ( n1705, n1707, n1708 );
nor U1546 ( n1708, n1690, n1709 );
nand U1547 ( n1709, n1275, n1710 );
nand U1548 ( n455, n1711, n1650 );
nand U1549 ( n1650, n1712, n1275 );
nor U1550 ( n1712, n1289, n1653 );
nor U1551 ( n1711, n1713, n1714 );
nor U1552 ( n1714, n1653, n1715 );
nor U1553 ( n1715, n1716, n1717 );
nor U1554 ( n1717, n2134, n1659 );
and U1555 ( n1659, n1718, n1719 );
nor U1556 ( n1719, n1720, n1721 );
and U1557 ( n1720, n1710, n1275 );
nor U1558 ( n1718, n1704, n1706 );
nand U1559 ( n1706, n1722, n1723 );
or U1560 ( n1723, n1328, n1690 );
nand U1561 ( n1722, n1243, n1288 );
nand U1562 ( n1704, n1627, n1724 );
or U1563 ( n1724, n1537, n1609 );
not U1564 ( n1627, n1604 );
nor U1565 ( n1604, n1266, n1690 );
nor U1566 ( n1716, n1657, n1725 );
not U1567 ( n1725, n1726 );
and U1568 ( n1657, n1727, n1728 );
nand U1569 ( n1728, n1219, n1729 );
nand U1570 ( n1729, n1730, n1609 );
nand U1571 ( n1730, n1289, n1297 );
nor U1572 ( n1727, n1700, n1699 );
nor U1573 ( n1699, n1710, n1273 );
and U1574 ( n1700, n1731, n1219 );
nand U1575 ( n1731, n1732, n1733 );
nand U1576 ( n1733, n1501, n1539 );
not U1577 ( n1732, n1689 );
nand U1578 ( n1689, n1311, n1734 );
nand U1579 ( n1734, n1274, n1735 );
not U1580 ( n1653, n1660 );
nor U1581 ( n1713, n2140, n1660 );
nand U1582 ( n1660, n1736, n1737 );
nor U1583 ( n1737, n1738, n1739 );
nand U1584 ( n1739, n1637, n1324 );
nand U1585 ( n1324, n1740, n1641 );
and U1586 ( n1740, n1269, n1318 );
nand U1587 ( n1637, n1741, n1300 );
nor U1588 ( n1738, n1262, n1742 );
nand U1589 ( n1742, n1539, n1309 );
nor U1590 ( n1736, n1743, n1744 );
nand U1591 ( n1744, n1293, n1745 );
nand U1592 ( n1745, n1746, n1210 );
nand U1593 ( n1746, n1747, n1748 );
nand U1594 ( n1748, n1300, n1749 );
nand U1595 ( n1749, n1646, n1750 );
nand U1596 ( n1750, n1297, n1219 );
nand U1597 ( n1747, n1285, n1307 );
and U1598 ( n1293, n1751, n1752 );
nand U1599 ( n1752, n1242, n1219 );
or U1600 ( n1242, n1318, n1753 );
nor U1601 ( n1751, n1754, n1642 );
and U1602 ( n1642, n1755, n1261 );
nor U1603 ( n1755, n1648, n1213 );
not U1604 ( n1754, n1255 );
nand U1605 ( n1255, n1269, n1753 );
nand U1606 ( n1743, n1756, n1757 );
nand U1607 ( n1757, n1758, n1213 );
nand U1608 ( n1758, n1759, n1760 );
nand U1609 ( n1760, n1761, n1690 );
nor U1610 ( n1759, n1762, n1247 );
nor U1611 ( n1247, n1609, n1210 );
nor U1612 ( n1762, n1539, n1763 );
nand U1613 ( n1763, n1501, n1219 );
nand U1614 ( n1756, n1764, n1297 );
nor U1615 ( n1764, n1765, n1690 );
nand U1616 ( n450, n1766, n1767 );
nand U1617 ( n1767, n1768, n1106 );
nand U1618 ( n1766, n1769, n1770 );
nand U1619 ( n1769, n1307, n1658 );
nand U1620 ( n445, n1771, n1772 );
nand U1621 ( n1772, n1773, n1667 );
nand U1622 ( n1667, n1774, n1775 );
nand U1623 ( n1775, n1776, n1658 );
nand U1624 ( n1771, n1768, n1107 );
nand U1625 ( n440, n1777, n1778 );
nand U1626 ( n1778, n1773, n1674 );
nand U1627 ( n1674, n1779, n1780 );
nand U1628 ( n1780, n1781, n1774 );
nand U1629 ( n1777, n1768, n1105 );
nand U1630 ( n44, n1782, n1783 );
nand U1631 ( n1783, n1784, n1119 );
nand U1632 ( n1782, n1372, n1183 );
nand U1633 ( n435, n1785, n1786 );
nand U1634 ( n1786, n1773, n1680 );
nand U1635 ( n1680, n1787, n1788 );
nand U1636 ( n1788, n1789, n1779 );
nand U1637 ( n1785, n1768, n1104 );
nand U1638 ( n430, n1790, n1791 );
nand U1639 ( n1791, n1773, n1696 );
xor U1640 ( n1696, n1787, n1792 );
nor U1641 ( n1792, n1793, n1102 );
not U1642 ( n1787, n1794 );
nor U1643 ( n1773, n1539, n1768 );
or U1644 ( n1790, n1770, n2135 );
nand U1645 ( n425, n1795, n1796 );
nand U1646 ( n1796, n1793, n1095 );
nor U1647 ( n1793, n1219, n2135 );
nor U1648 ( n1795, n1797, n1798 );
nor U1649 ( n1798, n1768, n1799 );
nor U1650 ( n1799, n1539, n1726 );
nand U1651 ( n1726, n1800, n1801 );
nand U1652 ( n1801, n1802, n1803 );
nand U1653 ( n1802, n2140, n1804 );
nand U1654 ( n1804, n1243, n1095 );
nand U1655 ( n1800, n1805, n1806 );
not U1656 ( n1806, n1803 );
nand U1657 ( n1803, n1794, n2115 );
nor U1658 ( n1794, n1779, n1789 );
nand U1659 ( n1789, n2114, n1807 );
nand U1660 ( n1807, n1243, n1104 );
or U1661 ( n1779, n1774, n1781 );
nand U1662 ( n1781, n2141, n1808 );
nand U1663 ( n1808, n1243, n1105 );
or U1664 ( n1774, n1776, n1658 );
nand U1665 ( n1658, n2116, n1809 );
nand U1666 ( n1809, n1243, n1106 );
nand U1667 ( n1776, n2142, n1810 );
nand U1668 ( n1810, n1243, n1107 );
nor U1669 ( n1805, n1095, n1811 );
nand U1670 ( n1811, n2135, n2140 );
nor U1671 ( n1797, n2134, n1770 );
nand U1672 ( n420, n1812, n1813 );
nand U1673 ( n1813, n1814, n1091 );
nand U1674 ( n1812, n1815, n1638 );
nor U1675 ( n1815, K_0_, n1619 );
nor U1676 ( n1619, n1235, K_1_ );
not U1677 ( n1235, K_2_ );
nand U1678 ( n415, n1816, n1817 );
nand U1679 ( n1817, n1638, n1230 );
not U1680 ( n1638, n1814 );
nand U1681 ( n1816, n1814, n1084 );
nand U1682 ( n1814, n1282, n1710 );
nand U1683 ( n1710, n1528, n1230 );
nor U1684 ( n1230, K_0_, K_1_ );
nor U1685 ( n1528, K_3_, K_2_ );
not U1686 ( n1282, n1253 );
nand U1687 ( n1253, n1512, n1219 );
not U1688 ( n1512, n1224 );
nand U1689 ( n410, n1818, n1819 );
or U1690 ( n1819, n1820, n2132 );
nand U1691 ( n405, n1821, n1822 );
or U1692 ( n1822, n1823, n2131 );
nand U1693 ( n1821, n1824, n2131 );
nor U1694 ( n1824, n2132, n1825 );
nand U1695 ( n400, n1826, n1827 );
or U1696 ( n1827, n1828, n1093 );
nand U1697 ( n1826, n1829, n1093 );
nand U1698 ( n395, n1830, n1831 );
or U1699 ( n1831, n1832, n2129 );
nand U1700 ( n1830, n1833, n2129 );
nor U1701 ( n1833, n2130, n1828 );
nand U1702 ( n390, n1834, n1835 );
nand U1703 ( n1835, n1836, n1100 );
nand U1704 ( n1836, n1832, n1837 );
nand U1705 ( n1837, n1838, n2129 );
nor U1706 ( n1832, n1829, n1839 );
nor U1707 ( n1839, n1825, n1093 );
nand U1708 ( n1829, n1823, n1840 );
nand U1709 ( n1840, n1838, n2131 );
and U1710 ( n1823, n1820, n1818 );
nand U1711 ( n1818, n1838, n2132 );
nand U1712 ( n1834, n1841, n2128 );
nor U1713 ( n1841, n1828, n1842 );
nand U1714 ( n1842, n1093, n1089 );
nand U1715 ( n1828, n1843, n1838 );
not U1716 ( n1838, n1825 );
nand U1717 ( n1825, n1297, n1820 );
nand U1718 ( n1820, n1768, n1844 );
nand U1719 ( n1844, n1243, n1845 );
nand U1720 ( n1845, n1246, n1846 );
nand U1721 ( n1846, n1741, n1285 );
not U1722 ( n1285, n1609 );
nand U1723 ( n1609, n1501, n1690 );
and U1724 ( n1246, n1224, n1847 );
nand U1725 ( n1847, n1753, n1848 );
nor U1726 ( n1753, n1309, n1262 );
nand U1727 ( n1224, n1849, n1212 );
nor U1728 ( n1849, n1297, n1539 );
not U1729 ( n1768, n1770 );
nand U1730 ( n1770, n1254, n1510 );
nand U1731 ( n1510, n1261, n1275 );
nand U1732 ( n1254, n1850, n1318 );
nor U1733 ( n1850, n1641, n1321 );
not U1734 ( n1641, n1320 );
nand U1735 ( n1320, n1843, n1851 );
nor U1736 ( n1851, n2130, n1852 );
nand U1737 ( n1852, n1089, n1100 );
nor U1738 ( n1843, n2131, n2132 );
nand U1739 ( n39, n1853, n1854 );
nand U1740 ( n1854, n1784, n1120 );
nand U1741 ( n1784, n1372, n1187 );
nand U1742 ( n1853, n1372, n1178 );
and U1743 ( n1372, n1444, n1446 );
nand U1744 ( n385, n1855, n1856 );
or U1745 ( n1856, n1857, n2127 );
nand U1746 ( n380, n1858, n1859 );
nand U1747 ( n1859, n1860, n1099 );
nand U1748 ( n1858, n1861, n2126 );
nor U1749 ( n1861, n2127, n1862 );
nand U1750 ( n375, n1863, n1864 );
or U1751 ( n1864, n1865, n1088 );
or U1752 ( n1863, n1866, n2125 );
nand U1753 ( n370, n1867, n1868 );
nand U1754 ( n1868, n1869, n1098 );
nand U1755 ( n1867, n1870, n2124 );
nor U1756 ( n1870, n2125, n1865 );
nand U1757 ( n365, n1871, n1872 );
nand U1758 ( n1872, n1873, n1173 );
nand U1759 ( n1873, n1874, n1875 );
nand U1760 ( n1875, n1876, n2124 );
not U1761 ( n1874, n1869 );
nand U1762 ( n1869, n1866, n1877 );
nand U1763 ( n1877, n1876, n2125 );
nor U1764 ( n1866, n1860, n1878 );
nor U1765 ( n1878, n1862, n1099 );
nand U1766 ( n1860, n1857, n1855 );
nand U1767 ( n1855, n1876, n2127 );
nand U1768 ( n1871, n1879, n2123 );
nor U1769 ( n1879, n1865, n1880 );
nand U1770 ( n1880, n1088, n1098 );
nand U1771 ( n1865, n1881, n1876 );
not U1772 ( n1876, n1862 );
nand U1773 ( n1862, n1882, n1297 );
and U1774 ( n1882, n1848, n1857 );
nand U1775 ( n1857, n1497, n1883 );
nand U1776 ( n1883, n1243, n1884 );
nand U1777 ( n1884, n1270, n1885 );
nand U1778 ( n1885, n1318, n1848 );
nor U1779 ( n1318, n1309, n1646 );
nand U1780 ( n1270, n1886, n1300 );
nor U1781 ( n1886, n1735, n1213 );
nand U1782 ( n1497, n1887, n1289 );
nor U1783 ( n1887, n1297, n1765 );
not U1784 ( n1765, n1288 );
nor U1785 ( n1288, n1888, n1735 );
nor U1786 ( n1881, n2126, n2127 );
nand U1787 ( n361, n1889, n1890 );
nor U1788 ( n1890, n1891, n1892 );
nor U1789 ( n1892, n1893, n1894 );
nand U1790 ( n1894, n2150, n2151 );
nor U1791 ( n1889, n1895, n1896 );
nor U1792 ( n1896, n2110, n1897 );
nor U1793 ( n1895, n1084, n1898 );
nand U1794 ( n1898, n2133, n1899 );
nand U1795 ( n357, n1900, n1901 );
nor U1796 ( n1901, n1891, n1902 );
nor U1797 ( n1902, n1893, n1903 );
nand U1798 ( n1903, n2150, n1083 );
nor U1799 ( n1900, n1904, n1905 );
nor U1800 ( n1905, n2111, n1897 );
nor U1801 ( n1904, n1084, n1906 );
nand U1802 ( n1906, n1899, n1091 );
nand U1803 ( n353, n1907, n1908 );
nor U1804 ( n1908, n1891, n1909 );
nor U1805 ( n1909, n1893, n1910 );
nand U1806 ( n1910, n2151, n1090 );
nor U1807 ( n1907, n1911, n1912 );
nor U1808 ( n1912, n2112, n1897 );
nor U1809 ( n1911, n1091, n1913 );
nand U1810 ( n1913, n1899, n1084 );
not U1811 ( n1899, n1914 );
nand U1812 ( n349, n1915, n1916 );
nor U1813 ( n1916, n1891, n1917 );
nor U1814 ( n1917, n1893, n1918 );
nand U1815 ( n1918, n1083, n1090 );
nand U1816 ( n1893, n1919, n1920 );
nand U1817 ( n1920, n1921, n1922 );
nand U1818 ( n1922, n1648, n1923 );
nor U1819 ( n1921, n1707, n1222 );
not U1820 ( n1222, n1256 );
not U1821 ( n1707, n1626 );
and U1822 ( n1891, n1924, n1761 );
not U1823 ( n1761, n1311 );
nand U1824 ( n1311, n1648, n1307 );
nor U1825 ( n1924, n1925, n1888 );
nor U1826 ( n1915, n1926, n1927 );
nor U1827 ( n1927, n2113, n1897 );
and U1828 ( n1897, n1928, n1929 );
nor U1829 ( n1929, n1925, n1930 );
nand U1830 ( n1930, n1256, n1626 );
nand U1831 ( n1626, n1721, n1297 );
nor U1832 ( n1721, n1289, n1735 );
nand U1833 ( n1735, n1210, n1539 );
nand U1834 ( n1256, n1284, n1300 );
not U1835 ( n1284, n1262 );
nand U1836 ( n1262, n1648, n1297 );
nor U1837 ( n1928, n1931, n1932 );
nand U1838 ( n1932, n1933, n1934 );
nand U1839 ( n1934, n1261, n1648 );
nand U1840 ( n1933, n1212, n1307 );
nor U1841 ( n1926, n1914, n1935 );
nand U1842 ( n1935, n1091, n1084 );
nand U1843 ( n1914, n1936, n1307 );
nor U1844 ( n1936, n1925, n1937 );
nor U1845 ( n1937, n1212, n1275 );
not U1846 ( n1925, n1919 );
nand U1847 ( n1919, n1938, n1939 );
nor U1848 ( n1939, n1940, n1941 );
nand U1849 ( n1941, n1942, n1943 );
nand U1850 ( n1943, n1944, n1261 );
nor U1851 ( n1944, n1213, n1321 );
not U1852 ( n1321, n1269 );
nor U1853 ( n1269, n1219, n1848 );
nand U1854 ( n1848, n1945, n1946 );
nor U1855 ( n1946, n1947, n1948 );
nand U1856 ( n1948, n1949, n1950 );
xor U1857 ( n1950, n1088, n2130 );
xnor U1858 ( n1949, n2127, n2132 );
xor U1859 ( n1947, n2126, n2131 );
nor U1860 ( n1945, n1951, n1952 );
xor U1861 ( n1952, n2123, n2128 );
xor U1862 ( n1951, n2124, n2129 );
nand U1863 ( n1942, n1212, n1953 );
nand U1864 ( n1953, n1537, n1954 );
nand U1865 ( n1954, n1312, n1210 );
nand U1866 ( n1537, n1243, n1297 );
not U1867 ( n1212, n1265 );
nand U1868 ( n1265, n1289, n1501 );
not U1869 ( n1501, n1888 );
nor U1870 ( n1940, n1274, n1328 );
nand U1871 ( n1328, n1243, n1312 );
not U1872 ( n1312, n1646 );
nand U1873 ( n1646, n1307, n1297 );
not U1874 ( n1297, n1213 );
not U1875 ( n1243, n1219 );
nor U1876 ( n1938, n1955, n1541 );
nand U1877 ( n1541, n1956, n1957 );
nand U1878 ( n1957, n1261, n1210 );
not U1879 ( n1261, n1958 );
nand U1880 ( n1956, n1959, n1648 );
not U1881 ( n1648, n1210 );
nor U1882 ( n1959, n1219, n1923 );
nand U1883 ( n1923, n1266, n1958 );
nand U1884 ( n1958, n1274, n1539 );
not U1885 ( n1274, n1309 );
nand U1886 ( n1309, n1690, n1888 );
nand U1887 ( n1219, n1960, n1961 );
nor U1888 ( n1961, n1174, n1962 );
nand U1889 ( n1962, n2141, n2142 );
nor U1890 ( n1960, n1103, n1963 );
nand U1891 ( n1963, n2115, n2116 );
and U1892 ( n1955, n1931, n1300 );
not U1893 ( n1300, n1327 );
nand U1894 ( n1327, n1289, n1888 );
nand U1895 ( n1888, n2117, n1964 );
not U1896 ( n1289, n1690 );
nand U1897 ( n1690, GAMMA_REG_1_, n1964 );
nand U1898 ( n1931, n1607, n1965 );
nand U1899 ( n1965, n1275, n1307 );
not U1900 ( n1307, n1539 );
not U1901 ( n1275, n1273 );
nand U1902 ( n1273, n1213, n1210 );
not U1903 ( n1607, n1741 );
nor U1904 ( n1741, n1210, n1266 );
nand U1905 ( n1266, n1539, n1213 );
nand U1906 ( n1213, GAMMA_REG_2_, n1964 );
nand U1907 ( n1539, GAMMA_REG_3_, n1964 );
nand U1908 ( n1210, GAMMA_REG_4_, n1964 );
not U1909 ( n1964, START );
nand U1910 ( n344, n1966, n1967 );
nand U1911 ( n1967, n1968, n1121 );
nand U1912 ( n1966, n1367, n1183 );
nand U1913 ( n34, n1969, n1970 );
nand U1914 ( n1970, n1971, n1122 );
nand U1915 ( n1969, n1340, n1183 );
nand U1916 ( n339, n1972, n1973 );
nand U1917 ( n1973, n1968, n1123 );
nand U1918 ( n1968, n1367, n1187 );
nand U1919 ( n1972, n1367, n1178 );
and U1920 ( n1367, n1974, n1447 );
nand U1921 ( n334, n1975, n1976 );
nand U1922 ( n1976, n1977, n1124 );
nand U1923 ( n1975, n1368, n1183 );
nand U1924 ( n329, n1978, n1979 );
nand U1925 ( n1979, n1977, n1125 );
nand U1926 ( n1977, n1368, n1187 );
nand U1927 ( n1978, n1368, n1178 );
and U1928 ( n1368, n1974, n1450 );
nand U1929 ( n324, n1980, n1981 );
nand U1930 ( n1981, n1982, n1126 );
nand U1931 ( n1980, n1343, n1183 );
nand U1932 ( n319, n1983, n1984 );
nand U1933 ( n1984, n1982, n1127 );
nand U1934 ( n1982, n1343, n1187 );
nand U1935 ( n1983, n1343, n1178 );
and U1936 ( n1343, n1985, n1447 );
nand U1937 ( n314, n1986, n1987 );
nand U1938 ( n1987, n1988, n1128 );
nand U1939 ( n1986, n1344, n1183 );
nand U1940 ( n309, n1989, n1990 );
nand U1941 ( n1990, n1988, n1129 );
nand U1942 ( n1988, n1344, n1187 );
nand U1943 ( n1989, n1344, n1178 );
and U1944 ( n1344, n1985, n1450 );
nand U1945 ( n304, n1991, n1992 );
nand U1946 ( n1992, n1993, n1130 );
nand U1947 ( n1991, n1339, n1183 );
nand U1948 ( n299, n1994, n1995 );
nand U1949 ( n1995, n1993, n1131 );
nand U1950 ( n1993, n1339, n1187 );
nand U1951 ( n1994, n1339, n1178 );
and U1952 ( n1339, n1974, n1444 );
nand U1953 ( n294, n1996, n1997 );
nand U1954 ( n1997, n1998, n1132 );
nand U1955 ( n1996, n1353, n1183 );
nand U1956 ( n29, n1999, n2000 );
nand U1957 ( n2000, n1971, n1133 );
nand U1958 ( n1971, n1340, n1187 );
nand U1959 ( n1999, n1340, n1178 );
and U1960 ( n1340, n1630, n1446 );
and U1961 ( n1446, n2001, n1092 );
nand U1962 ( n289, n2002, n2003 );
nand U1963 ( n2003, n1998, n1134 );
nand U1964 ( n1998, n1353, n1187 );
nand U1965 ( n2002, n1353, n1178 );
and U1966 ( n1353, n1974, n1630 );
and U1967 ( n1974, n2004, n2145 );
nor U1968 ( n2004, n1085, n1092 );
nand U1969 ( n284, n2005, n2006 );
nand U1970 ( n2006, n2007, n1135 );
nand U1971 ( n2005, n1354, n1183 );
nand U1972 ( n279, n2008, n2009 );
nand U1973 ( n2009, n2007, n1136 );
nand U1974 ( n2007, n1354, n1187 );
nand U1975 ( n2008, n1354, n1178 );
and U1976 ( n1354, n1985, n1444 );
nand U1977 ( n274, n2010, n2011 );
nand U1978 ( n2011, n2012, n1137 );
nand U1979 ( n2010, n1349, n1183 );
nand U1980 ( n269, n2013, n2014 );
nand U1981 ( n2014, n2012, n1138 );
nand U1982 ( n2012, n1349, n1187 );
nand U1983 ( n2013, n1349, n1178 );
and U1984 ( n1349, n1985, n1630 );
and U1985 ( n1985, n2015, n2145 );
nor U1986 ( n2015, n2119, n1092 );
nand U1987 ( n264, n2016, n2017 );
nand U1988 ( n2017, n2018, n1139 );
nand U1989 ( n2016, n1350, n1183 );
nand U1990 ( n259, n2019, n2020 );
nand U1991 ( n2020, n2018, n1140 );
nand U1992 ( n2018, n1350, n1187 );
nand U1993 ( n2019, n1350, n1178 );
and U1994 ( n1350, n2021, n1447 );
nand U1995 ( n254, n2022, n2023 );
nand U1996 ( n2023, n2024, n1141 );
nand U1997 ( n2022, n1406, n1183 );
nand U1998 ( n249, n2025, n2026 );
nand U1999 ( n2026, n2024, n1142 );
nand U2000 ( n2024, n1406, n1187 );
nand U2001 ( n2025, n1406, n1178 );
and U2002 ( n1406, n2021, n1450 );
nand U2003 ( n244, n2027, n2028 );
nand U2004 ( n2028, n2029, n1143 );
nand U2005 ( n2027, n1407, n1183 );
nand U2006 ( n239, n2030, n2031 );
nand U2007 ( n2031, n2029, n1144 );
nand U2008 ( n2029, n1407, n1187 );
nand U2009 ( n2030, n1407, n1178 );
and U2010 ( n1407, n2032, n1447 );
nand U2011 ( n234, n2033, n2034 );
nand U2012 ( n2034, n2035, n1145 );
nand U2013 ( n2033, n1402, n1183 );
nand U2014 ( n229, n2036, n2037 );
nand U2015 ( n2037, n2035, n1146 );
nand U2016 ( n2035, n1402, n1187 );
nand U2017 ( n2036, n1402, n1178 );
and U2018 ( n1402, n2032, n1450 );
nand U2019 ( n224, n2038, n2039 );
nand U2020 ( n2039, n2040, n1147 );
nand U2021 ( n2038, n1403, n1183 );
nand U2022 ( n219, n2041, n2042 );
nand U2023 ( n2042, n2040, n1148 );
nand U2024 ( n2040, n1403, n1187 );
nand U2025 ( n2041, n1403, n1178 );
and U2026 ( n1403, n2021, n1444 );
nand U2027 ( n214, n2043, n2044 );
nand U2028 ( n2044, n2045, n1149 );
nand U2029 ( n2043, n1416, n1183 );
nand U2030 ( n209, n2046, n2047 );
nand U2031 ( n2047, n2045, n1150 );
nand U2032 ( n2045, n1416, n1187 );
nand U2033 ( n2046, n1416, n1178 );
and U2034 ( n1416, n2021, n1630 );
and U2035 ( n2021, n2048, n2145 );
nor U2036 ( n2048, n2146, n1085 );
nand U2037 ( n204, n2049, n2050 );
nand U2038 ( n2050, n2051, n1151 );
nand U2039 ( n2049, n1417, n1183 );
nand U2040 ( n199, n2052, n2053 );
nand U2041 ( n2053, n2051, n1152 );
nand U2042 ( n2051, n1417, n1187 );
nand U2043 ( n2052, n1417, n1178 );
and U2044 ( n1417, n2032, n1444 );
nand U2045 ( n194, n2054, n2055 );
nand U2046 ( n2055, n2056, n1153 );
nand U2047 ( n2054, n1412, n1183 );
nand U2048 ( n189, n2057, n2058 );
nand U2049 ( n2058, n2056, n1154 );
nand U2050 ( n2056, n1412, n1187 );
nand U2051 ( n2057, n1412, n1178 );
and U2052 ( n1412, n2032, n1630 );
and U2053 ( n2032, n2059, n2145 );
nor U2054 ( n2059, n2119, n2146 );
nand U2055 ( n184, n2060, n2061 );
nand U2056 ( n2061, n2062, n1155 );
nand U2057 ( n2060, n1413, n1183 );
nand U2058 ( n179, n2063, n2064 );
nand U2059 ( n2064, n2062, n1156 );
nand U2060 ( n2062, n1413, n1187 );
nand U2061 ( n2063, n1413, n1178 );
and U2062 ( n1413, n2065, n1447 );
nand U2063 ( n174, n2066, n2067 );
nand U2064 ( n2067, n2068, n1157 );
nand U2065 ( n2066, n1385, n1183 );
nand U2066 ( n169, n2069, n2070 );
nand U2067 ( n2070, n2068, n1158 );
nand U2068 ( n2068, n1385, n1187 );
nand U2069 ( n2069, n1385, n1178 );
and U2070 ( n1385, n2065, n1450 );
nand U2071 ( n164, n2071, n2072 );
nand U2072 ( n2072, n2073, n1159 );
nand U2073 ( n2071, n1386, n1183 );
nand U2074 ( n159, n2074, n2075 );
nand U2075 ( n2075, n2073, n1160 );
nand U2076 ( n2073, n1386, n1187 );
nand U2077 ( n2074, n1386, n1178 );
and U2078 ( n1386, n2076, n1447 );
nand U2079 ( n154, n2077, n2078 );
nand U2080 ( n2078, n2079, n1161 );
nand U2081 ( n2077, n1381, n1183 );
nand U2082 ( n149, n2080, n2081 );
nand U2083 ( n2081, n2079, n1162 );
nand U2084 ( n2079, n1381, n1187 );
nand U2085 ( n2080, n1381, n1178 );
and U2086 ( n1381, n2076, n1450 );
nor U2087 ( n1450, n1087, n2147 );
nand U2088 ( n144, n2082, n2083 );
nand U2089 ( n2083, n2084, n1163 );
nand U2090 ( n2082, n1382, n1183 );
nand U2091 ( n139, n2085, n2086 );
nand U2092 ( n2086, n2084, n1164 );
nand U2093 ( n2084, n1382, n1187 );
nand U2094 ( n2085, n1382, n1178 );
and U2095 ( n1382, n2065, n1444 );
nand U2096 ( n134, n2087, n2088 );
nand U2097 ( n2088, n2089, n1165 );
nand U2098 ( n2087, n1394, n1183 );
nand U2099 ( n129, n2090, n2091 );
nand U2100 ( n2091, n2089, n1166 );
nand U2101 ( n2089, n1394, n1187 );
nand U2102 ( n2090, n1394, n1178 );
and U2103 ( n1394, n2065, n1630 );
and U2104 ( n2065, n2092, n2146 );
nor U2105 ( n2092, n2145, n1085 );
nand U2106 ( n124, n2093, n2094 );
nand U2107 ( n2094, n2095, n1167 );
nand U2108 ( n2093, n1395, n1183 );
nand U2109 ( n119, n2096, n2097 );
nand U2110 ( n2097, n2095, n1168 );
nand U2111 ( n2095, n1395, n1187 );
nand U2112 ( n2096, n1395, n1178 );
and U2113 ( n1395, n2076, n1444 );
nor U2114 ( n1444, n1096, n2120 );
nand U2115 ( n114, n2098, n2099 );
nand U2116 ( n2099, n2100, n1169 );
nand U2117 ( n2098, n1391, n1183 );
nand U2118 ( n109, n2101, n2102 );
nand U2119 ( n2102, n2100, n1170 );
nand U2120 ( n2100, n1391, n1187 );
nand U2121 ( n2101, n1391, n1178 );
and U2122 ( n1391, n2076, n1630 );
nor U2123 ( n1630, n2147, n2120 );
and U2124 ( n2076, n2001, n2146 );
nor U2125 ( n2001, n2119, n2145 );
nand U2126 ( n104, n2103, n2104 );
nand U2127 ( n2104, n1177, n1171 );
nand U2128 ( n1177, n1179, n1187 );
nand U2129 ( n2103, n1183, n1179 );
and U2130 ( n1179, n1447, n1445 );
and U2131 ( n1445, n2105, n2119 );
nor U2132 ( n2105, n2145, n2146 );
nor U2133 ( n1447, n1087, n1096 );
endmodule

