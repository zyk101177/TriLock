
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule

module b20_ori ( clk, reset, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_,
SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_,
SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_,
SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, ADD_1068_U4,
ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59,
ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47,
ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52,
ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123 );
input clk, reset, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_,
SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_,
SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_,
SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_;
output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
U126, U123;
wire P2_WR_REG, P1_WR_REG, P2_RD_REG, P1_RD_REG, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, ex_wire30, ex_wire31, ex_wire32, ex_wire33, ex_wire34, ex_wire35, ex_wire36, ex_wire37, ex_wire38, ex_wire39, ex_wire40, ex_wire41, ex_wire42, ex_wire43, P2_ADDR_REG_19_,
P1_ADDR_REG_19_, P1_DATAO_REG_9_, P1_DATAO_REG_8_, P1_DATAO_REG_7_,
P1_DATAO_REG_6_, P1_DATAO_REG_5_, P1_DATAO_REG_4_, P1_DATAO_REG_3_,
P1_DATAO_REG_31_, P1_DATAO_REG_30_, P1_DATAO_REG_2_, P1_DATAO_REG_29_,
P1_DATAO_REG_28_, P1_DATAO_REG_27_, P1_DATAO_REG_26_,
P1_DATAO_REG_25_, P1_DATAO_REG_24_, P1_DATAO_REG_23_,
P1_DATAO_REG_22_, P1_DATAO_REG_21_, P1_DATAO_REG_20_, P1_DATAO_REG_1_,
P1_DATAO_REG_19_, P1_DATAO_REG_18_, P1_DATAO_REG_17_,
P1_DATAO_REG_16_, P1_DATAO_REG_15_, P1_DATAO_REG_14_,
P1_DATAO_REG_13_, P1_DATAO_REG_12_, P1_DATAO_REG_11_,
P1_DATAO_REG_10_, P1_DATAO_REG_0_, P2_DATAO_REG_9_, P2_DATAO_REG_8_,
P2_DATAO_REG_7_, P2_DATAO_REG_6_, P2_DATAO_REG_5_, P2_DATAO_REG_4_,
P2_DATAO_REG_3_, P2_DATAO_REG_31_, P2_DATAO_REG_30_, P2_DATAO_REG_2_,
P2_DATAO_REG_29_, P2_DATAO_REG_28_, P2_DATAO_REG_27_,
P2_DATAO_REG_26_, P2_DATAO_REG_25_, P2_DATAO_REG_24_,
P2_DATAO_REG_23_, P2_DATAO_REG_22_, P2_DATAO_REG_21_,
P2_DATAO_REG_20_, P2_DATAO_REG_1_, P2_DATAO_REG_19_, P2_DATAO_REG_18_,
P2_DATAO_REG_17_, P2_DATAO_REG_16_, P2_DATAO_REG_15_,
P2_DATAO_REG_14_, P2_DATAO_REG_13_, P2_DATAO_REG_12_,
P2_DATAO_REG_11_, P2_DATAO_REG_10_, P2_DATAO_REG_0_, P1_STATE_REG,
n1325, n1315, n1310, n1305, n1300, n1295, n1290, n1285, n1280, n1275,
n1270, n1265, n1260, n1255, n1250, n1245, n1240, n1235, n1230, n1225,
n1220, n1215, n1210, n1205, n1200, n1195, n1190, n1185, n1180, n1175,
n1170, n1005, n1000, n995, n990, n985, n980, n975, n970, n965, n960,
n955, n950, n945, n940, n935, n930, n925, n920, n915, n910, n905,
n900, n890, n885, n880, n875, n870, n865, n860, n855, n850, n845,
n840, n835, n830, n825, n820, n815, n810, n805, n800, n795, n790,
n785, n780, n775, n770, n765, n760, n755, n750, P1_D_REG_31_, n425,
P1_D_REG_30_, n420, P1_D_REG_29_, n415, P1_D_REG_28_, n410,
P1_D_REG_27_, n405, P1_D_REG_26_, n400, P1_D_REG_25_, n395,
P1_D_REG_24_, n390, P1_D_REG_23_, n385, n380, P1_D_REG_21_, n375,
P1_D_REG_20_, n370, P1_D_REG_19_, n365, P1_D_REG_18_, n360,
P1_D_REG_17_, n355, P1_D_REG_16_, n350, P1_D_REG_15_, n345,
P1_D_REG_14_, n340, P1_D_REG_13_, n335, P1_D_REG_12_, n330,
P1_D_REG_11_, n325, P1_D_REG_10_, n320, P1_D_REG_9_, n315,
P1_D_REG_8_, n310, n305, P1_D_REG_6_, n300, P1_D_REG_5_, n295,
P1_D_REG_4_, n290, P1_D_REG_3_, n285, P1_D_REG_2_, n280, n265, n260,
n255, n250, n245, n240, n235, n230, n225, n220, n215, n210, n205,
n200, n195, n190, n185, n180, n175, n170, n165, n160, n155, n150,
n145, n140, n135, n130, n125, n120, n115, n110, n895, P1_B_REG,
P1_REG2_REG_0_, n270, n275, n430, n435, n440, n445, n450, n455, n460,
n465, n470, n475, n480, n485, n490, n495, n500, n505, n510, n515,
n520, n525, n530, n535, n540, n545, n550, n555, n560, n565, n570,
n575, n580, n585, n590, n595, n600, n605, n610, n615, n620, n625,
n630, n635, n640, n645, n650, n655, n660, n665, n670, n675, n680,
n685, n690, n695, n700, n705, n710, n715, n720, n725, n730, n735,
n740, n745, n1010, n1015, n1020, n1025, n1030, n1035, n1040, n1045,
n1050, n1055, n1060, n1065, n1070, n1075, n1080, n1085, n1090, n1095,
n1100, n1105, n1110, n1115, n1120, n1125, n1130, n1135, n1140, n1145,
n1150, n1155, n1160, n1165, P1_IR_REG_31_, P1_IR_REG_0_, P1_IR_REG_1_,
P1_IR_REG_2_, P1_IR_REG_3_, P1_IR_REG_4_, P1_IR_REG_5_, P1_IR_REG_6_,
P1_IR_REG_7_, P1_IR_REG_8_, P1_IR_REG_9_, P1_IR_REG_10_,
P1_IR_REG_11_, P1_IR_REG_12_, P1_IR_REG_13_, P1_IR_REG_14_,
P1_IR_REG_15_, P1_IR_REG_16_, P1_IR_REG_17_, P1_IR_REG_18_,
P1_IR_REG_19_, P1_IR_REG_20_, P1_IR_REG_21_, P1_IR_REG_22_,
P1_IR_REG_23_, P1_IR_REG_24_, P1_IR_REG_25_, P1_IR_REG_26_,
P1_IR_REG_27_, P1_IR_REG_28_, P1_IR_REG_29_, P1_IR_REG_30_,
P1_REG2_REG_1_, P1_REG1_REG_1_, P1_REG0_REG_1_, P1_REG3_REG_1_,
P1_REG2_REG_2_, P1_REG1_REG_2_, P1_REG0_REG_2_, P1_REG3_REG_2_,
P1_REG0_REG_0_, P1_REG1_REG_0_, P1_REG2_REG_3_, P1_REG1_REG_3_,
P1_REG0_REG_3_, P1_REG2_REG_4_, P1_REG1_REG_4_, P1_REG0_REG_4_,
P1_REG2_REG_5_, P1_REG1_REG_5_, P1_REG0_REG_5_, P1_REG2_REG_6_,
P1_REG1_REG_6_, P1_REG0_REG_6_, P1_REG2_REG_7_, P1_REG1_REG_7_,
P1_REG0_REG_7_, P1_REG2_REG_8_, P1_REG1_REG_8_, P1_REG0_REG_8_,
P1_REG2_REG_9_, P1_REG1_REG_9_, P1_REG0_REG_9_, P1_REG2_REG_10_,
P1_REG1_REG_10_, P1_REG0_REG_10_, P1_REG2_REG_11_, P1_REG1_REG_11_,
P1_REG0_REG_11_, P1_REG2_REG_12_, P1_REG1_REG_12_, P1_REG0_REG_12_,
P1_REG2_REG_13_, P1_REG1_REG_13_, P1_REG0_REG_13_, P1_REG2_REG_14_,
P1_REG1_REG_14_, P1_REG0_REG_14_, P1_REG2_REG_15_, P1_REG1_REG_15_,
P1_REG0_REG_15_, P1_REG2_REG_16_, P1_REG1_REG_16_, P1_REG0_REG_16_,
P1_REG2_REG_17_, P1_REG1_REG_17_, P1_REG0_REG_17_, P1_REG2_REG_18_,
P1_REG1_REG_18_, P1_REG0_REG_18_, P1_REG1_REG_19_, P1_REG0_REG_19_,
P1_REG1_REG_20_, P1_REG0_REG_20_, P1_REG1_REG_21_, P1_REG0_REG_21_,
P1_REG1_REG_22_, P1_REG0_REG_22_, P1_REG1_REG_23_, P1_REG0_REG_23_,
P1_REG1_REG_24_, P1_REG0_REG_24_, P1_REG1_REG_25_, P1_REG0_REG_25_,
P1_REG1_REG_26_, P1_REG0_REG_26_, P1_REG1_REG_27_, P1_REG0_REG_27_,
P1_REG1_REG_28_, P1_REG0_REG_28_, P1_REG1_REG_29_, P1_REG0_REG_29_,
P1_REG1_REG_30_, P1_REG0_REG_30_, P1_REG1_REG_31_, P1_REG0_REG_31_,
P1_REG3_REG_18_, P1_ADDR_REG_18_, P1_ADDR_REG_17_, P1_REG3_REG_16_,
P1_ADDR_REG_16_, P1_ADDR_REG_15_, P1_REG3_REG_14_, P1_ADDR_REG_14_,
P1_ADDR_REG_13_, P1_REG3_REG_12_, P1_ADDR_REG_12_, P1_ADDR_REG_11_,
P1_REG3_REG_10_, P1_ADDR_REG_10_, P1_ADDR_REG_9_, P1_REG3_REG_8_,
P1_ADDR_REG_8_, P1_ADDR_REG_7_, P1_REG3_REG_6_, P1_ADDR_REG_6_,
P1_ADDR_REG_5_, P1_REG3_REG_4_, P1_ADDR_REG_4_, P1_REG3_REG_3_,
P1_ADDR_REG_3_, P1_ADDR_REG_2_, P1_ADDR_REG_0_, P1_REG3_REG_26_,
P1_REG3_REG_22_, P1_REG3_REG_20_, P1_REG3_REG_24_, P1_REG3_REG_28_,
P1_D_REG_0_, P1_D_REG_1_, P2_STATE_REG, n2550, n2540, n2535, n2530,
n2525, n2520, n2515, n2510, n2505, n2500, n2495, n2490, n2485, n2480,
n2475, n2470, n2465, n2460, n2455, n2450, n2445, n2440, n2435, n2430,
n2425, n2420, n2415, n2410, n2405, n2400, n2230, n2225, n2220, n2215,
n2210, n2205, n2200, n2195, n2190, n2185, n2180, n2175, n2170, n2165,
n2160, n2155, n2150, n2145, n2140, n2135, n2130, n2125, n2120, n2115,
n2110, n2105, n2100, n2095, n2090, n2085, n2080, n2075, n2070, n2065,
n2060, n2055, n2050, n2045, n2040, n2035, n2030, n2025, n2020, n2015,
n2010, n2005, n2000, n1995, n1990, n1985, n1980, n1975, P2_D_REG_31_,
n1650, P2_D_REG_30_, n1645, P2_D_REG_29_, n1640, P2_D_REG_28_, n1635,
P2_D_REG_27_, n1630, P2_D_REG_26_, n1625, P2_D_REG_25_, n1620,
P2_D_REG_24_, n1615, P2_D_REG_23_, n1610, n1605, P2_D_REG_21_, n1600,
P2_D_REG_20_, n1595, P2_D_REG_19_, n1590, P2_D_REG_18_, n1585,
P2_D_REG_17_, n1580, P2_D_REG_16_, n1575, P2_D_REG_15_, n1570,
P2_D_REG_14_, n1565, P2_D_REG_13_, n1560, P2_D_REG_12_, n1555,
P2_D_REG_11_, n1550, P2_D_REG_10_, n1545, P2_D_REG_9_, n1540,
P2_D_REG_8_, n1535, n1530, P2_D_REG_6_, n1525, P2_D_REG_5_, n1520,
P2_D_REG_4_, n1515, P2_D_REG_3_, n1510, P2_D_REG_2_, n1505, n1490,
n1485, n1480, n1475, n1470, n1465, n1460, n1455, n1450, n1445, n1440,
n1435, n1430, n1425, n1420, n1415, n1410, n1405, n1400, n1395, n1390,
n1385, n1380, n1375, n1370, n1365, n1360, n1355, n1350, n1345, n1340,
n1335, n2395, P2_B_REG, n1495, n1500, n1655, n1660, n1665, n1670,
n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720,
n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770,
n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820,
n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870,
n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1910, n1915, n1920,
n1925, n1930, n1935, n1940, n1945, n1950, n1955, n1960, n1965, n1970,
n2235, n2240, n2245, n2250, n2255, n2260, n2265, n2270, n2275, n2280,
n2285, n2290, n2295, n2300, n2305, n2310, n2315, n2320, n2325, n2330,
n2335, n2340, n2345, n2350, n2355, n2360, n2365, n2370, n2375, n2380,
n2385, n2390, P2_IR_REG_31_, P2_IR_REG_0_, P2_IR_REG_1_, P2_IR_REG_2_,
P2_IR_REG_3_, P2_IR_REG_4_, P2_IR_REG_5_, P2_IR_REG_6_, P2_IR_REG_7_,
P2_IR_REG_8_, P2_IR_REG_9_, P2_IR_REG_10_, P2_IR_REG_11_,
P2_IR_REG_12_, P2_IR_REG_13_, P2_IR_REG_14_, P2_IR_REG_15_,
P2_IR_REG_16_, P2_IR_REG_17_, P2_IR_REG_18_, P2_IR_REG_19_,
P2_IR_REG_20_, P2_IR_REG_21_, P2_IR_REG_22_, P2_IR_REG_23_,
P2_IR_REG_24_, P2_IR_REG_25_, P2_IR_REG_26_, P2_IR_REG_27_,
P2_IR_REG_28_, P2_IR_REG_29_, P2_IR_REG_30_, P2_REG0_REG_1_,
P2_REG1_REG_1_, P2_REG2_REG_1_, P2_REG3_REG_1_, P2_REG0_REG_2_,
P2_REG1_REG_2_, P2_REG2_REG_2_, P2_REG3_REG_2_, P2_REG0_REG_0_,
P2_REG1_REG_0_, P2_REG2_REG_0_, P2_REG3_REG_0_, P2_REG0_REG_3_,
P2_REG1_REG_3_, P2_REG2_REG_3_, P2_REG0_REG_4_, P2_REG1_REG_4_,
P2_REG2_REG_4_, P2_REG0_REG_5_, P2_REG1_REG_5_, P2_REG2_REG_5_,
P2_REG0_REG_6_, P2_REG1_REG_6_, P2_REG2_REG_6_, P2_REG0_REG_7_,
P2_REG1_REG_7_, P2_REG2_REG_7_, P2_REG0_REG_8_, P2_REG1_REG_8_,
P2_REG2_REG_8_, P2_REG0_REG_9_, P2_REG1_REG_9_, P2_REG2_REG_9_,
P2_REG0_REG_10_, P2_REG1_REG_10_, P2_REG2_REG_10_, P2_REG0_REG_11_,
P2_REG1_REG_11_, P2_REG2_REG_11_, P2_REG0_REG_12_, P2_REG1_REG_12_,
P2_REG2_REG_12_, P2_REG0_REG_13_, P2_REG1_REG_13_, P2_REG2_REG_13_,
P2_REG0_REG_14_, P2_REG1_REG_14_, P2_REG2_REG_14_, P2_REG0_REG_15_,
P2_REG1_REG_15_, P2_REG2_REG_15_, P2_REG0_REG_16_, P2_REG1_REG_16_,
P2_REG2_REG_16_, P2_REG0_REG_17_, P2_REG1_REG_17_, P2_REG2_REG_17_,
P2_REG0_REG_18_, P2_REG1_REG_18_, P2_REG2_REG_18_, P2_REG0_REG_19_,
P2_REG1_REG_19_, P2_REG1_REG_20_, P2_REG0_REG_20_, P2_REG1_REG_21_,
P2_REG0_REG_21_, P2_REG1_REG_22_, P2_REG0_REG_22_, P2_REG1_REG_23_,
P2_REG0_REG_23_, P2_REG1_REG_24_, P2_REG0_REG_24_, P2_REG1_REG_25_,
P2_REG0_REG_25_, P2_REG1_REG_26_, P2_REG0_REG_26_, P2_REG1_REG_27_,
P2_REG0_REG_27_, P2_REG1_REG_28_, P2_REG0_REG_28_, P2_REG1_REG_29_,
P2_REG0_REG_29_, P2_REG1_REG_30_, P2_REG0_REG_30_, P2_REG1_REG_31_,
P2_REG0_REG_31_, P2_REG3_REG_19_, P2_REG3_REG_18_, P2_ADDR_REG_18_,
P2_REG3_REG_17_, P2_ADDR_REG_17_, P2_REG3_REG_16_, P2_ADDR_REG_16_,
P2_REG3_REG_15_, P2_ADDR_REG_15_, P2_REG3_REG_14_, P2_ADDR_REG_14_,
P2_REG3_REG_13_, P2_ADDR_REG_13_, P2_REG3_REG_12_, P2_ADDR_REG_12_,
P2_REG3_REG_11_, P2_ADDR_REG_11_, P2_REG3_REG_10_, P2_ADDR_REG_10_,
P2_REG3_REG_9_, P2_ADDR_REG_9_, P2_REG3_REG_8_, P2_ADDR_REG_8_,
P2_REG3_REG_7_, P2_ADDR_REG_7_, P2_REG3_REG_6_, P2_ADDR_REG_6_,
P2_REG3_REG_5_, P2_ADDR_REG_5_, P2_REG3_REG_4_, P2_ADDR_REG_4_,
P2_REG3_REG_3_, P2_ADDR_REG_3_, P2_ADDR_REG_2_, P2_ADDR_REG_1_,
P2_ADDR_REG_0_, P2_REG3_REG_26_, P2_REG3_REG_22_, P2_REG3_REG_20_,
P2_REG3_REG_24_, P2_REG3_REG_25_, P2_REG3_REG_21_, P2_REG3_REG_28_,
P2_REG3_REG_23_, P2_REG3_REG_27_, P2_D_REG_0_, P2_D_REG_1_, n1, n2,
n3, n4, n5, n6, n7, n8, n9, n10, n14, n15, n17, n18, n19, n20, n21,
n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n50,
n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
n65, n66, n67, n69, n70, n71, n73, n74, n75, n76, n77, n78, n81, n82,
n83, n84, n87, n88, n89, n90, n92, n93, n94, n95, n96, n97, n98, n99,
n101, n102, n103, n104, n105, n106, n107, n108, n109, n111, n112,
n113, n114, n116, n117, n118, n119, n121, n122, n123, n124, n126,
n128, n129, n131, n132, n133, n134, n136, n137, n138, n139, n141,
n142, n143, n144, n146, n147, n148, n149, n151, n152, n153, n154,
n156, n157, n158, n159, n161, n162, n163, n164, n166, n168, n171,
n172, n173, n174, n176, n177, n178, n179, n182, n183, n184, n186,
n187, n188, n191, n192, n193, n194, n196, n197, n198, n199, n201,
n202, n203, n204, n206, n207, n208, n209, n211, n212, n213, n214,
n216, n217, n218, n219, n221, n222, n224, n226, n227, n228, n229,
n231, n232, n233, n234, n236, n237, n238, n239, n241, n242, n243,
n244, n246, n247, n248, n249, n251, n252, n253, n254, n256, n257,
n258, n259, n261, n262, n263, n264, n266, n267, n268, n269, n271,
n272, n273, n274, n276, n277, n278, n279, n281, n282, n283, n284,
n286, n287, n288, n289, n291, n292, n293, n294, n296, n297, n298,
n299, n301, n302, n303, n304, n306, n307, n308, n309, n311, n312,
n313, n314, n316, n317, n318, n319, n321, n322, n323, n324, n326,
n327, n328, n329, n331, n332, n333, n334, n336, n337, n338, n339,
n341, n344, n346, n348, n349, n351, n352, n353, n354, n356, n357,
n358, n359, n361, n363, n364, n366, n367, n369, n371, n372, n373,
n374, n376, n377, n378, n379, n381, n382, n383, n384, n386, n387,
n388, n389, n391, n392, n393, n394, n396, n398, n399, n401, n402,
n403, n404, n406, n407, n408, n409, n411, n419, n421, n504, n506,
n507, n508, n509, n511, n512, n513, n514, n516, n517, n518, n519,
n521, n522, n523, n524, n526, n527, n528, n529, n531, n532, n533,
n534, n536, n537, n538, n539, n541, n542, n543, n544, n546, n547,
n548, n549, n551, n552, n553, n554, n556, n557, n558, n559, n561,
n562, n563, n564, n567, n568, n569, n571, n572, n573, n574, n576,
n578, n579, n581, n582, n583, n584, n586, n587, n588, n589, n591,
n592, n593, n594, n596, n597, n598, n599, n601, n602, n603, n604,
n606, n607, n608, n609, n611, n612, n613, n614, n616, n617, n618,
n619, n622, n624, n626, n627, n628, n629, n631, n632, n633, n634,
n636, n637, n638, n639, n641, n642, n644, n646, n647, n648, n649,
n651, n652, n654, n656, n657, n658, n659, n661, n662, n663, n664,
n666, n667, n668, n669, n672, n673, n674, n677, n678, n679, n681,
n683, n684, n687, n688, n689, n691, n692, n693, n694, n696, n697,
n698, n699, n701, n702, n703, n704, n706, n707, n708, n709, n711,
n712, n714, n716, n717, n719, n721, n722, n723, n724, n726, n727,
n728, n729, n731, n732, n733, n734, n736, n737, n739, n741, n742,
n743, n744, n746, n747, n748, n749, n751, n752, n753, n754, n756,
n757, n759, n761, n762, n763, n764, n766, n767, n768, n769, n771,
n772, n773, n774, n776, n777, n781, n783, n787, n788, n789, n791,
n792, n793, n794, n796, n797, n798, n799, n801, n802, n803, n807,
n808, n809, n811, n812, n813, n814, n816, n817, n827, n828, n849,
n851, n853, n854, n856, n857, n858, n859, n861, n862, n863, n864,
n866, n867, n868, n871, n872, n873, n874, n876, n877, n878, n879,
n882, n883, n884, n886, n887, n888, n889, n891, n893, n894, n896,
n897, n898, n902, n903, n904, n906, n907, n909, n911, n912, n914,
n916, n917, n918, n919, n921, n922, n923, n924, n926, n927, n928,
n929, n932, n933, n934, n936, n937, n938, n939, n941, n942, n944,
n946, n947, n948, n949, n951, n952, n953, n954, n956, n957, n959,
n961, n962, n963, n964, n966, n967, n968, n969, n971, n972, n973,
n974, n976, n977, n978, n979, n981, n982, n983, n984, n986, n987,
n988, n989, n991, n992, n993, n994, n996, n997, n998, n999, n1001,
n1002, n1003, n1004, n1007, n1008, n1009, n1011, n1013, n1021, n1022,
n1149, n1176, n1177, n1178, n1179, n1181, n1182, n1183, n1184, n1186,
n1187, n1188, n1189, n1191, n1192, n1193, n1194, n1196, n1197, n1198,
n1199, n1201, n1202, n1203, n1204, n1206, n1207, n1208, n1209, n1211,
n1212, n1213, n1214, n1217, n1218, n1219, n1221, n1222, n1223, n1224,
n1226, n1227, n1228, n1229, n1231, n1232, n1233, n1234, n1236, n1237,
n1238, n1239, n1241, n1242, n1243, n1244, n1246, n1247, n1248, n1249,
n1251, n1253, n1254, n1256, n1257, n1258, n1259, n1261, n1262, n1263,
n1264, n1266, n1267, n1268, n1269, n1271, n1272, n1273, n1274, n1276,
n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1286, n1287, n1288,
n1289, n1291, n1292, n1293, n1294, n1296, n1297, n1298, n1299, n1301,
n1302, n1303, n1304, n1306, n1307, n1308, n1309, n1311, n1312, n1313,
n1314, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1336,
n1337, n1338, n1339, n1341, n1342, n1343, n1344, n1346, n1347, n1348,
n1349, n1351, n1352, n1353, n1354, n1356, n1357, n1358, n1359, n1361,
n1362, n1363, n1364, n1367, n1368, n1369, n1371, n1372, n1373, n1374,
n1376, n1377, n1378, n1379, n1381, n1382, n1383, n1384, n1386, n1387,
n1388, n1389, n1391, n1392, n1393, n1394, n1396, n1397, n1398, n1399,
n1401, n1402, n1403, n1404, n1406, n1407, n1408, n1409, n1411, n1412,
n1413, n1414, n1416, n1417, n1418, n1419, n1421, n1422, n1423, n1424,
n1426, n1427, n1428, n1429, n1431, n1432, n1433, n1434, n1436, n1437,
n1438, n1439, n1441, n1442, n1443, n1444, n1446, n1447, n1448, n1449,
n1451, n1452, n1453, n1454, n1456, n1457, n1458, n1459, n1461, n1462,
n1463, n1464, n1466, n1467, n1468, n1469, n1471, n1472, n1473, n1474,
n1476, n1477, n1478, n1479, n1481, n1482, n1483, n1484, n1486, n1487,
n1488, n1489, n1491, n1492, n1493, n1494, n1496, n1497, n1498, n1499,
n1501, n1502, n1503, n1504, n1506, n1507, n1508, n1509, n1511, n1512,
n1513, n1514, n1516, n1517, n1518, n1519, n1521, n1522, n1523, n1524,
n1526, n1527, n1528, n1529, n1531, n1532, n1533, n1534, n1536, n1537,
n1538, n1539, n1541, n1542, n1543, n1544, n1546, n1547, n1548, n1549,
n1551, n1552, n1553, n1554, n1556, n1557, n1558, n1559, n1561, n1562,
n1563, n1564, n1566, n1567, n1568, n1569, n1571, n1572, n1573, n1574,
n1576, n1577, n1578, n1579, n1581, n1582, n1583, n1584, n1586, n1587,
n1588, n1589, n1591, n1592, n1593, n1594, n1596, n1597, n1598, n1599,
n1601, n1602, n1603, n1604, n1606, n1607, n1608, n1609, n1611, n1612,
n1613, n1614, n1616, n1617, n1618, n1619, n1621, n1622, n1623, n1624,
n1627, n1628, n1629, n1631, n1632, n1633, n1634, n1636, n1637, n1638,
n1639, n1641, n1642, n1643, n1644, n1646, n1647, n1648, n1649, n1651,
n1652, n1653, n1654, n1656, n1657, n1658, n1659, n1661, n1662, n1663,
n1664, n1666, n1667, n1668, n1669, n1671, n1672, n1673, n1674, n1676,
n1677, n1678, n1679, n1681, n1682, n1683, n1684, n1686, n1687, n1688,
n1689, n1691, n1692, n1693, n1694, n1696, n1697, n1698, n1699, n1701,
n1702, n1703, n1704, n1706, n1707, n1708, n1709, n1711, n1712, n1713,
n1714, n1716, n1717, n1718, n1719, n1721, n1722, n1723, n1724, n1726,
n1727, n1728, n1729, n1731, n1732, n1733, n1734, n1736, n1737, n1738,
n1739, n1741, n1742, n1743, n1744, n1746, n1747, n1748, n1749, n1751,
n1752, n1753, n1754, n1756, n1757, n1758, n1759, n1761, n1762, n1763,
n1764, n1766, n1767, n1768, n1769, n1771, n1772, n1773, n1774, n1776,
n1777, n1778, n1779, n1781, n1782, n1783, n1784, n1786, n1787, n1788,
n1789, n1791, n1792, n1793, n1794, n1796, n1797, n1798, n1799, n1801,
n1802, n1803, n1804, n1806, n1807, n1808, n1809, n1811, n1812, n1813,
n1814, n1816, n1817, n1818, n1819, n1821, n1822, n1823, n1824, n1826,
n1827, n1828, n1829, n1831, n1832, n1833, n1834, n1836, n1837, n1838,
n1839, n1841, n1842, n1843, n1844, n1846, n1847, n1848, n1849, n1851,
n1852, n1853, n1854, n1856, n1857, n1858, n1859, n1861, n1862, n1863,
n1864, n1866, n1867, n1868, n1869, n1871, n1872, n1873, n1874, n1876,
n1877, n1878, n1879, n1881, n1882, n1883, n1884, n1886, n1887, n1888,
n1889, n1891, n1893, n1894, n1896, n1897, n1898, n1899, n1901, n1902,
n1903, n1904, n1906, n1907, n1908, n1909, n1912, n1913, n1914, n1916,
n1917, n1918, n1919, n1921, n1922, n1923, n1924, n1926, n1927, n1928,
n1929, n1931, n1932, n1933, n1934, n1936, n1937, n1938, n1939, n1941,
n1942, n1943, n1944, n1946, n1947, n1948, n1949, n1951, n1952, n1953,
n1954, n1956, n1957, n1958, n1959, n1961, n1962, n1963, n1964, n1966,
n1967, n1968, n1969, n1971, n1972, n1973, n1974, n1976, n1977, n1978,
n1979, n1981, n1982, n1983, n1984, n1986, n1987, n1988, n1989, n1991,
n1992, n1993, n1994, n1996, n1997, n1998, n1999, n2001, n2002, n2003,
n2004, n2006, n2007, n2008, n2009, n2011, n2012, n2013, n2014, n2016,
n2017, n2018, n2019, n2021, n2022, n2023, n2024, n2026, n2027, n2028,
n2029, n2031, n2032, n2033, n2034, n2036, n2037, n2038, n2039, n2041,
n2042, n2043, n2044, n2046, n2047, n2048, n2049, n2051, n2052, n2053,
n2054, n2056, n2057, n2058, n2059, n2061, n2062, n2063, n2064, n2066,
n2067, n2068, n2069, n2071, n2072, n2073, n2074, n2076, n2077, n2078,
n2079, n2081, n2082, n2083, n2084, n2086, n2087, n2088, n2089, n2091,
n2092, n2093, n2094, n2096, n2097, n2098, n2099, n2101, n2102, n2103,
n2104, n2106, n2107, n2108, n2109, n2111, n2112, n2113, n2114, n2116,
n2117, n2118, n2119, n2121, n2122, n2123, n2124, n2126, n2127, n2128,
n2129, n2131, n2132, n2133, n2134, n2136, n2137, n2138, n2139, n2141,
n2142, n2143, n2144, n2146, n2147, n2148, n2149, n2151, n2152, n2153,
n2154, n2156, n2157, n2158, n2159, n2161, n2162, n2163, n2164, n2166,
n2167, n2168, n2169, n2171, n2172, n2173, n2174, n2176, n2177, n2178,
n2179, n2181, n2182, n2183, n2184, n2186, n2187, n2188, n2189, n2191,
n2192, n2193, n2194, n2196, n2197, n2198, n2199, n2201, n2202, n2203,
n2204, n2206, n2207, n2208, n2209, n2211, n2212, n2213, n2214, n2216,
n2217, n2218, n2219, n2221, n2222, n2223, n2224, n2226, n2227, n2228,
n2229, n2231, n2232, n2233, n2234, n2236, n2237, n2238, n2239, n2241,
n2242, n2243, n2244, n2246, n2247, n2248, n2249, n2251, n2252, n2253,
n2254, n2256, n2257, n2258, n2259, n2261, n2262, n2263, n2264, n2266,
n2267, n2268, n2269, n2271, n2272, n2273, n2274, n2276, n2277, n2278,
n2279, n2281, n2282, n2283, n2284, n2286, n2287, n2288, n2289, n2291,
n2292, n2293, n2294, n2296, n2297, n2298, n2299, n2301, n2302, n2303,
n2304, n2306, n2307, n2308, n2309, n2311, n2312, n2313, n2314, n2316,
n2317, n2318, n2319, n2321, n2322, n2323, n2324, n2326, n2327, n2328,
n2329, n2331, n2332, n2333, n2334, n2336, n2337, n2338, n2339, n2341,
n2342, n2343, n2344, n2346, n2347, n2348, n2349, n2351, n2352, n2353,
n2354, n2356, n2357, n2358, n2359, n2361, n2362, n2363, n2364, n2366,
n2367, n2368, n2369, n2371, n2372, n2373, n2374, n2376, n2377, n2378,
n2379, n2381, n2382, n2383, n2384, n2386, n2387, n2388, n2389, n2391,
n2392, n2393, n2394, n2396, n2397, n2398, n2399, n2401, n2402, n2403,
n2404, n2406, n2407, n2408, n2409, n2411, n2412, n2413, n2414, n2416,
n2417, n2418, n2419, n2421, n2422, n2423, n2424, n2426, n2427, n2428,
n2429, n2431, n2432, n2433, n2434, n2436, n2437, n2438, n2439, n2441,
n2442, n2443, n2444, n2446, n2447, n2448, n2449, n2451, n2452, n2453,
n2454, n2456, n2457, n2458, n2459, n2461, n2462, n2463, n2464, n2466,
n2467, n2468, n2469, n2471, n2472, n2473, n2474, n2476, n2477, n2478,
n2479, n2481, n2482, n2483, n2484, n2486, n2487, n2488, n2489, n2491,
n2492, n2493, n2494, n2496, n2497, n2498, n2499, n2501, n2502, n2503,
n2504, n2506, n2507, n2508, n2509, n2511, n2512, n2513, n2514, n2516,
n2517, n2518, n2519, n2521, n2522, n2523, n2524, n2526, n2527, n2528,
n2529, n2531, n2532, n2533, n2534, n2536, n2537, n2538, n2539, n2541,
n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2551, n2552,
n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
n2673, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
n2704, n2705, n2706, n2707, n2710, n2711, n2712, n2713, n2714, n2715,
n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
n2736, n2737, n2738, n2739, n2740, n2741, n2743, n2744, n2745, n2746,
n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2756, n2757,
n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2838, n2839,
n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
n3050, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3161, n3162, n3163,
n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
n3304, n3305, n3306, n3307, n3308, n3309, n3312, n3313, n3314, n3315,
n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
n3326, n3327, n3328, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
n3368, n3369, n3370, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
n3519, n3520, n3521, n3522, n3523, n3524, n3526, n3527, n3528, n3529,
n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3589, n3590, n3591,
n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3650, n3651, n3652,
n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3861, n3862, n3863,
n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
n3904, n3905, n3906, n3907, n3909, n3910, n3911, n3912, n3913, n3914,
n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
n4005, n4006, n4007, n4008, n4009, n4011, n4012, n4013, n4014, n4015,
n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4134, n4135, n4136,
n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
n4357, n4358, n4359, n4360, n4361, n4362, n4364, n4365, n4366, n4367,
n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
n4868, n4869, n4870, n4871, n4872, n4874, n4875, n4876, n4877, n4878,
n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4977, n4978, n4979,
n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
n5260, n5261, n5262, n5263, n5264, n5265, n5267, n5268, n5269, n5270,
n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
n5301, n5302, n5303, n5304, n5305, n5306, n5308, n5309, n5310, n5311,
n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
n5552, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5681, n5682, n5683,
n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
n5784, n5785, n5786, n5787, n5788, n5790, n5791, n5792, n5793, n5794,
n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5915,
n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
n6096, n6097, n6098, n6099, n6100, n6102, n6103, n6104, n6105, n6106,
n6107, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
n6820, n6821, n6822, n6823, n6824, n6825, n6828, n6829, n6830, n6831,
n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
n7004, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
n7026, n7027, n7028, n7029, n7030, n7032, n7033, n7034, n7035, n7036,
n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
n7079, n7080, n7081, n7082, n7083, n7084, n7086, n7087, n7088, n7089,
n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
n7220, n7221, n7222, n7223, n7224, n7226, n7227, n7228, n7229, n7230,
n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
n7271, n7272, n7273, n7274, n7276, n7277, n7278, n7279, n7280, n7281,
n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
n7302, n7303, n7304, n7305, n7308, n7309, n7310, n7311, n7312, n7313,
n7314, n7317, n7318, n7319, n7321, n7322, n7323, n7324, n7325, n7326,
n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
n7417, n7418, n7419, n7420, n7421, n7424, n7425, n7426, n7427, n7428,
n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
n7639, n7640, n7641, n7642, n7643, n7644, n7646, n7647, n7648, n7649,
n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
n8290, n8291, n8292, n8293, n8296, n8297, n8298, n8299, n8300, n8301,
n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8701, n8702, n8703,
n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
n8904, n8905, n8906, n8907, n8908, n8909, n8911, n8912, n8913, n8914,
n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
n9865, n9866, n9867, n9868, n9869, n9870, n9872, n9873, n9874, n9875,
n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9884, n9885, n9886,
n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
n9977, n9978, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
n10392, n10393, n10394, n10397, n10398, n10399, n10400, n10401,
n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
n10834, n10835, n10836, n10837, n10838, n10839, n10842, n10843,
n10844, n10845, n10846, n10847, n10848, n10849, n10851, n10852,
n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
n11533, n11534, n11535, n11536, n11537;

dff P1_STATE_REG_reg ( clk, reset, P1_STATE_REG, n11535 );
not U_inv0 ( n10956, P1_STATE_REG );
dff P2_STATE_REG_reg ( clk, reset, P2_STATE_REG, n11530 );
dff P2_RD_REG_reg ( clk, reset, P2_RD_REG, n2550 );
dff P1_IR_REG_0__reg ( clk, reset, P1_IR_REG_0_, n110 );
not U_inv1 ( n10957, P1_IR_REG_0_ );
dff P1_B_REG_reg ( clk, reset, P1_B_REG, n1170 );
not U_inv2 ( n11111, P1_B_REG );
dff P1_REG0_REG_29__reg ( clk, reset, P1_REG0_REG_29_, n575 );
dff P1_DATAO_REG_29__reg ( clk, reset, P1_DATAO_REG_29_, n1155 );
dff P1_REG0_REG_30__reg ( clk, reset, P1_REG0_REG_30_, n580 );
dff P1_DATAO_REG_30__reg ( clk, reset, P1_DATAO_REG_30_, n1160 );
dff P1_REG0_REG_31__reg ( clk, reset, P1_REG0_REG_31_, n585 );
dff P1_DATAO_REG_31__reg ( clk, reset, P1_DATAO_REG_31_, n1165 );
dff P2_IR_REG_0__reg ( clk, reset, P2_IR_REG_0_, n1335 );
not U_inv3 ( n10960, P2_IR_REG_0_ );
dff P2_IR_REG_2__reg ( clk, reset, P2_IR_REG_2_, n1345 );
dff P2_IR_REG_3__reg ( clk, reset, P2_IR_REG_3_, n1350 );
dff P2_IR_REG_4__reg ( clk, reset, P2_IR_REG_4_, n1355 );
dff P2_IR_REG_6__reg ( clk, reset, P2_IR_REG_6_, n1365 );
dff P2_REG0_REG_6__reg ( clk, reset, P2_REG0_REG_6_, n1685 );
not U_inv4 ( n11001, P2_REG0_REG_6_ );
dff P2_REG0_REG_7__reg ( clk, reset, P2_REG0_REG_7_, n1690 );
not U_inv5 ( n11006, P2_REG0_REG_7_ );
dff P2_REG0_REG_8__reg ( clk, reset, P2_REG0_REG_8_, n1695 );
not U_inv6 ( n11021, P2_REG0_REG_8_ );
dff P2_B_REG_reg ( clk, reset, P2_B_REG, n2395 );
not U_inv7 ( n11157, P2_B_REG );
dff P2_REG3_REG_15__reg ( clk, reset, P2_REG3_REG_15_, n2400 );
not U_inv8 ( n11180, P2_REG3_REG_15_ );
dff P2_REG0_REG_16__reg ( clk, reset, P2_REG0_REG_16_, n1735 );
not U_inv9 ( n11062, P2_REG0_REG_16_ );
dff P2_REG0_REG_17__reg ( clk, reset, P2_REG0_REG_17_, n1740 );
not U_inv10 ( n11065, P2_REG0_REG_17_ );
dff P2_REG0_REG_18__reg ( clk, reset, P2_REG0_REG_18_, n1745 );
not U_inv11 ( n11073, P2_REG0_REG_18_ );
dff P2_REG0_REG_22__reg ( clk, reset, P2_REG0_REG_22_, n1765 );
not U_inv12 ( n11098, P2_REG0_REG_22_ );
dff P2_REG0_REG_23__reg ( clk, reset, P2_REG0_REG_23_, n1770 );
not U_inv13 ( n11102, P2_REG0_REG_23_ );
dff P2_REG0_REG_24__reg ( clk, reset, P2_REG0_REG_24_, n1775 );
not U_inv14 ( n11119, P2_REG0_REG_24_ );
dff P2_REG0_REG_25__reg ( clk, reset, P2_REG0_REG_25_, n1780 );
not U_inv15 ( n11113, P2_REG0_REG_25_ );
dff P2_REG0_REG_26__reg ( clk, reset, P2_REG0_REG_26_, n1785 );
not U_inv16 ( n11116, P2_REG0_REG_26_ );
dff P2_REG0_REG_27__reg ( clk, reset, P2_REG0_REG_27_, n1790 );
not U_inv17 ( n11140, P2_REG0_REG_27_ );
dff P2_REG0_REG_29__reg ( clk, reset, P2_REG0_REG_29_, n1800 );
not U_inv18 ( n11149, P2_REG0_REG_29_ );
dff P2_REG2_REG_28__reg ( clk, reset, ex_wire0, n2115 );
not U_inv19 ( n11144, ex_wire0 );
dff P2_DATAO_REG_28__reg ( clk, reset, P2_DATAO_REG_28_, n2375 );
dff P1_REG0_REG_28__reg ( clk, reset, P1_REG0_REG_28_, n570 );
dff P1_DATAO_REG_28__reg ( clk, reset, P1_DATAO_REG_28_, n1150 );
dff P2_IR_REG_28__reg ( clk, reset, P2_IR_REG_28_, n1475 );
dff P2_REG0_REG_0__reg ( clk, reset, P2_REG0_REG_0_, n1655 );
not U_inv20 ( n10969, P2_REG0_REG_0_ );
dff P2_REG0_REG_1__reg ( clk, reset, P2_REG0_REG_1_, n1660 );
not U_inv21 ( n10994, P2_REG0_REG_1_ );
dff P2_REG0_REG_2__reg ( clk, reset, P2_REG0_REG_2_, n1665 );
not U_inv22 ( n10997, P2_REG0_REG_2_ );
dff P2_REG0_REG_4__reg ( clk, reset, P2_REG0_REG_4_, n1675 );
not U_inv23 ( n10999, P2_REG0_REG_4_ );
dff P2_REG0_REG_5__reg ( clk, reset, P2_REG0_REG_5_, n1680 );
not U_inv24 ( n10990, P2_REG0_REG_5_ );
dff P2_REG2_REG_9__reg ( clk, reset, P2_REG2_REG_9_, n2020 );
not U_inv25 ( n11016, P2_REG2_REG_9_ );
dff P2_REG0_REG_10__reg ( clk, reset, P2_REG0_REG_10_, n1705 );
not U_inv26 ( n11019, P2_REG0_REG_10_ );
dff P2_REG0_REG_11__reg ( clk, reset, P2_REG0_REG_11_, n1710 );
not U_inv27 ( n11029, P2_REG0_REG_11_ );
dff P2_REG0_REG_12__reg ( clk, reset, P2_REG0_REG_12_, n1715 );
not U_inv28 ( n11035, P2_REG0_REG_12_ );
dff P2_REG2_REG_13__reg ( clk, reset, P2_REG2_REG_13_, n2040 );
not U_inv29 ( n11036, P2_REG2_REG_13_ );
dff P2_REG0_REG_14__reg ( clk, reset, P2_REG0_REG_14_, n1725 );
not U_inv30 ( n11054, P2_REG0_REG_14_ );
dff P2_REG0_REG_19__reg ( clk, reset, P2_REG0_REG_19_, n1750 );
not U_inv31 ( n11083, P2_REG0_REG_19_ );
dff P2_REG0_REG_20__reg ( clk, reset, P2_REG0_REG_20_, n1755 );
not U_inv32 ( n11081, P2_REG0_REG_20_ );
dff P2_REG0_REG_21__reg ( clk, reset, P2_REG0_REG_21_, n1760 );
not U_inv33 ( n11095, P2_REG0_REG_21_ );
dff P2_DATAO_REG_21__reg ( clk, reset, P2_DATAO_REG_21_, n2340 );
dff P1_REG3_REG_27__reg ( clk, reset, ex_wire1, n1310 );
not U_inv34 ( n11121, ex_wire1 );
dff P1_REG2_REG_27__reg ( clk, reset, ex_wire2, n885 );
not U_inv35 ( n11136, ex_wire2 );
dff P1_DATAO_REG_27__reg ( clk, reset, P1_DATAO_REG_27_, n1145 );
dff P1_IR_REG_30__reg ( clk, reset, P1_IR_REG_30_, n260 );
dff P1_DATAO_REG_0__reg ( clk, reset, P1_DATAO_REG_0_, n1010 );
dff P2_REG2_REG_3__reg ( clk, reset, P2_REG2_REG_3_, n1990 );
not U_inv36 ( n10983, P2_REG2_REG_3_ );
dff P2_DATAO_REG_3__reg ( clk, reset, P2_DATAO_REG_3_, n2250 );
dff P1_REG0_REG_12__reg ( clk, reset, P1_REG0_REG_12_, n490 );
dff P1_DATAO_REG_12__reg ( clk, reset, P1_DATAO_REG_12_, n1070 );
dff P1_REG0_REG_21__reg ( clk, reset, P1_REG0_REG_21_, n535 );
dff P1_DATAO_REG_21__reg ( clk, reset, P1_DATAO_REG_21_, n1115 );
dff P2_IR_REG_21__reg ( clk, reset, P2_IR_REG_21_, n1440 );
dff P2_IR_REG_22__reg ( clk, reset, P2_IR_REG_22_, n1445 );
dff P2_IR_REG_23__reg ( clk, reset, P2_IR_REG_23_, n1450 );
dff P2_IR_REG_24__reg ( clk, reset, P2_IR_REG_24_, n1455 );
dff P2_IR_REG_27__reg ( clk, reset, P2_IR_REG_27_, n1470 );
dff P2_IR_REG_29__reg ( clk, reset, P2_IR_REG_29_, n1480 );
dff P2_IR_REG_30__reg ( clk, reset, P2_IR_REG_30_, n1485 );
dff P2_IR_REG_26__reg ( clk, reset, P2_IR_REG_26_, n1465 );
dff P2_D_REG_31__reg ( clk, reset, P2_D_REG_31_, n1650 );
dff P2_D_REG_30__reg ( clk, reset, P2_D_REG_30_, n1645 );
dff P2_D_REG_29__reg ( clk, reset, P2_D_REG_29_, n1640 );
dff P2_D_REG_28__reg ( clk, reset, P2_D_REG_28_, n1635 );
dff P2_D_REG_27__reg ( clk, reset, P2_D_REG_27_, n1630 );
dff P2_D_REG_26__reg ( clk, reset, P2_D_REG_26_, n1625 );
dff P2_D_REG_25__reg ( clk, reset, P2_D_REG_25_, n1620 );
dff P2_D_REG_24__reg ( clk, reset, P2_D_REG_24_, n1615 );
dff P2_D_REG_23__reg ( clk, reset, P2_D_REG_23_, n1610 );
dff P2_D_REG_21__reg ( clk, reset, P2_D_REG_21_, n1600 );
dff P2_D_REG_20__reg ( clk, reset, P2_D_REG_20_, n1595 );
dff P2_D_REG_19__reg ( clk, reset, P2_D_REG_19_, n1590 );
dff P2_D_REG_18__reg ( clk, reset, P2_D_REG_18_, n1585 );
dff P2_D_REG_17__reg ( clk, reset, P2_D_REG_17_, n1580 );
dff P2_D_REG_16__reg ( clk, reset, P2_D_REG_16_, n1575 );
dff P2_D_REG_15__reg ( clk, reset, P2_D_REG_15_, n1570 );
dff P2_D_REG_14__reg ( clk, reset, P2_D_REG_14_, n1565 );
dff P2_D_REG_13__reg ( clk, reset, P2_D_REG_13_, n1560 );
dff P2_D_REG_12__reg ( clk, reset, P2_D_REG_12_, n1555 );
dff P2_D_REG_11__reg ( clk, reset, P2_D_REG_11_, n1550 );
dff P2_D_REG_10__reg ( clk, reset, P2_D_REG_10_, n1545 );
dff P2_D_REG_9__reg ( clk, reset, P2_D_REG_9_, n1540 );
dff P2_D_REG_8__reg ( clk, reset, P2_D_REG_8_, n1535 );
dff P2_D_REG_6__reg ( clk, reset, P2_D_REG_6_, n1525 );
dff P2_D_REG_5__reg ( clk, reset, P2_D_REG_5_, n1520 );
dff P2_D_REG_4__reg ( clk, reset, P2_D_REG_4_, n1515 );
dff P2_D_REG_3__reg ( clk, reset, P2_D_REG_3_, n1510 );
dff P2_D_REG_2__reg ( clk, reset, P2_D_REG_2_, n1505 );
dff P2_D_REG_22__reg ( clk, reset, ex_wire3, n1605 );
not U_inv37 ( n11135, ex_wire3 );
dff P2_D_REG_7__reg ( clk, reset, ex_wire4, n1530 );
not U_inv38 ( n11134, ex_wire4 );
dff P2_D_REG_0__reg ( clk, reset, P2_D_REG_0_, n1495 );
dff P2_DATAO_REG_29__reg ( clk, reset, P2_DATAO_REG_29_, n2380 );
dff P2_DATAO_REG_27__reg ( clk, reset, P2_DATAO_REG_27_, n2370 );
dff P2_DATAO_REG_26__reg ( clk, reset, P2_DATAO_REG_26_, n2365 );
dff P2_DATAO_REG_25__reg ( clk, reset, P2_DATAO_REG_25_, n2360 );
dff P2_DATAO_REG_24__reg ( clk, reset, P2_DATAO_REG_24_, n2355 );
dff P2_DATAO_REG_23__reg ( clk, reset, P2_DATAO_REG_23_, n2350 );
dff P2_DATAO_REG_22__reg ( clk, reset, P2_DATAO_REG_22_, n2345 );
dff P2_DATAO_REG_20__reg ( clk, reset, P2_DATAO_REG_20_, n2335 );
dff P2_DATAO_REG_19__reg ( clk, reset, P2_DATAO_REG_19_, n2330 );
dff P2_DATAO_REG_18__reg ( clk, reset, P2_DATAO_REG_18_, n2325 );
dff P2_DATAO_REG_17__reg ( clk, reset, P2_DATAO_REG_17_, n2320 );
dff P2_DATAO_REG_16__reg ( clk, reset, P2_DATAO_REG_16_, n2315 );
dff P2_DATAO_REG_15__reg ( clk, reset, P2_DATAO_REG_15_, n2310 );
dff P2_DATAO_REG_14__reg ( clk, reset, P2_DATAO_REG_14_, n2305 );
dff P2_DATAO_REG_13__reg ( clk, reset, P2_DATAO_REG_13_, n2300 );
dff P2_DATAO_REG_12__reg ( clk, reset, P2_DATAO_REG_12_, n2295 );
dff P2_DATAO_REG_11__reg ( clk, reset, P2_DATAO_REG_11_, n2290 );
dff P2_DATAO_REG_10__reg ( clk, reset, P2_DATAO_REG_10_, n2285 );
dff P2_DATAO_REG_9__reg ( clk, reset, P2_DATAO_REG_9_, n2280 );
dff P2_DATAO_REG_8__reg ( clk, reset, P2_DATAO_REG_8_, n2275 );
dff P2_DATAO_REG_7__reg ( clk, reset, P2_DATAO_REG_7_, n2270 );
dff P2_DATAO_REG_6__reg ( clk, reset, P2_DATAO_REG_6_, n2265 );
dff P2_DATAO_REG_5__reg ( clk, reset, P2_DATAO_REG_5_, n2260 );
dff P2_DATAO_REG_4__reg ( clk, reset, P2_DATAO_REG_4_, n2255 );
dff P2_DATAO_REG_2__reg ( clk, reset, P2_DATAO_REG_2_, n2245 );
dff P2_DATAO_REG_1__reg ( clk, reset, P2_DATAO_REG_1_, n2240 );
dff P1_IR_REG_1__reg ( clk, reset, P1_IR_REG_1_, n115 );
dff P1_REG0_REG_16__reg ( clk, reset, P1_REG0_REG_16_, n510 );
dff P1_REG0_REG_17__reg ( clk, reset, P1_REG0_REG_17_, n515 );
dff P1_DATAO_REG_17__reg ( clk, reset, P1_DATAO_REG_17_, n1095 );
dff P1_REG0_REG_18__reg ( clk, reset, P1_REG0_REG_18_, n520 );
dff P1_DATAO_REG_18__reg ( clk, reset, P1_DATAO_REG_18_, n1100 );
dff P1_REG0_REG_20__reg ( clk, reset, P1_REG0_REG_20_, n530 );
dff P1_DATAO_REG_20__reg ( clk, reset, P1_DATAO_REG_20_, n1110 );
dff P1_REG0_REG_22__reg ( clk, reset, P1_REG0_REG_22_, n540 );
dff P1_DATAO_REG_22__reg ( clk, reset, P1_DATAO_REG_22_, n1120 );
dff P1_REG0_REG_23__reg ( clk, reset, P1_REG0_REG_23_, n545 );
dff P1_DATAO_REG_23__reg ( clk, reset, P1_DATAO_REG_23_, n1125 );
dff P1_REG0_REG_24__reg ( clk, reset, P1_REG0_REG_24_, n550 );
dff P1_DATAO_REG_24__reg ( clk, reset, P1_DATAO_REG_24_, n1130 );
dff P1_REG0_REG_25__reg ( clk, reset, P1_REG0_REG_25_, n555 );
dff P1_DATAO_REG_25__reg ( clk, reset, P1_DATAO_REG_25_, n1135 );
dff P2_IR_REG_25__reg ( clk, reset, P2_IR_REG_25_, n1460 );
dff P2_D_REG_1__reg ( clk, reset, P2_D_REG_1_, n1500 );
dff P1_REG0_REG_26__reg ( clk, reset, P1_REG0_REG_26_, n560 );
dff P1_DATAO_REG_26__reg ( clk, reset, P1_DATAO_REG_26_, n1140 );
dff P1_IR_REG_26__reg ( clk, reset, P1_IR_REG_26_, n240 );
dff P1_WR_REG_reg ( clk, reset, P1_WR_REG, n11448 );
dff P1_DATAO_REG_1__reg ( clk, reset, P1_DATAO_REG_1_, n1015 );
dff P1_REG0_REG_3__reg ( clk, reset, P1_REG0_REG_3_, n445 );
dff P1_REG3_REG_15__reg ( clk, reset, ex_wire5, n1175 );
not U_inv39 ( n11059, ex_wire5 );
dff P1_REG2_REG_15__reg ( clk, reset, P1_REG2_REG_15_, n825 );
not U_inv40 ( n11067, P1_REG2_REG_15_ );
dff P1_DATAO_REG_15__reg ( clk, reset, P1_DATAO_REG_15_, n1085 );
dff P1_REG3_REG_19__reg ( clk, reset, ex_wire6, n1285 );
not U_inv41 ( n11072, ex_wire6 );
dff P1_REG2_REG_19__reg ( clk, reset, ex_wire7, n845 );
not U_inv42 ( n11086, ex_wire7 );
dff P1_DATAO_REG_19__reg ( clk, reset, P1_DATAO_REG_19_, n1105 );
dff P1_IR_REG_19__reg ( clk, reset, P1_IR_REG_19_, n205 );
dff P1_IR_REG_27__reg ( clk, reset, P1_IR_REG_27_, n245 );
not U_inv43 ( n10961, P1_IR_REG_27_ );
dff P1_IR_REG_25__reg ( clk, reset, P1_IR_REG_25_, n235 );
dff P1_IR_REG_24__reg ( clk, reset, P1_IR_REG_24_, n230 );
dff P1_IR_REG_23__reg ( clk, reset, P1_IR_REG_23_, n225 );
dff P1_IR_REG_21__reg ( clk, reset, P1_IR_REG_21_, n215 );
dff P1_IR_REG_22__reg ( clk, reset, P1_IR_REG_22_, n220 );
dff P1_IR_REG_20__reg ( clk, reset, P1_IR_REG_20_, n210 );
dff P1_IR_REG_17__reg ( clk, reset, P1_IR_REG_17_, n195 );
dff P1_IR_REG_18__reg ( clk, reset, P1_IR_REG_18_, n200 );
dff P1_IR_REG_15__reg ( clk, reset, P1_IR_REG_15_, n185 );
not U_inv44 ( n11055, P1_IR_REG_15_ );
dff P1_IR_REG_3__reg ( clk, reset, P1_IR_REG_3_, n125 );
not U_inv45 ( n10971, P1_IR_REG_3_ );
dff P1_D_REG_31__reg ( clk, reset, P1_D_REG_31_, n425 );
dff P1_D_REG_30__reg ( clk, reset, P1_D_REG_30_, n420 );
dff P1_D_REG_29__reg ( clk, reset, P1_D_REG_29_, n415 );
dff P1_D_REG_28__reg ( clk, reset, P1_D_REG_28_, n410 );
dff P1_D_REG_27__reg ( clk, reset, P1_D_REG_27_, n405 );
dff P1_D_REG_26__reg ( clk, reset, P1_D_REG_26_, n400 );
dff P1_D_REG_25__reg ( clk, reset, P1_D_REG_25_, n395 );
dff P1_D_REG_24__reg ( clk, reset, P1_D_REG_24_, n390 );
dff P1_D_REG_23__reg ( clk, reset, P1_D_REG_23_, n385 );
dff P1_D_REG_21__reg ( clk, reset, P1_D_REG_21_, n375 );
dff P1_D_REG_20__reg ( clk, reset, P1_D_REG_20_, n370 );
dff P1_D_REG_19__reg ( clk, reset, P1_D_REG_19_, n365 );
dff P1_D_REG_18__reg ( clk, reset, P1_D_REG_18_, n360 );
dff P1_D_REG_17__reg ( clk, reset, P1_D_REG_17_, n355 );
dff P1_D_REG_16__reg ( clk, reset, P1_D_REG_16_, n350 );
dff P1_D_REG_15__reg ( clk, reset, P1_D_REG_15_, n345 );
dff P1_D_REG_14__reg ( clk, reset, P1_D_REG_14_, n340 );
dff P1_D_REG_13__reg ( clk, reset, P1_D_REG_13_, n335 );
dff P1_D_REG_12__reg ( clk, reset, P1_D_REG_12_, n330 );
dff P1_D_REG_11__reg ( clk, reset, P1_D_REG_11_, n325 );
dff P1_D_REG_10__reg ( clk, reset, P1_D_REG_10_, n320 );
dff P1_D_REG_9__reg ( clk, reset, P1_D_REG_9_, n315 );
dff P1_D_REG_8__reg ( clk, reset, P1_D_REG_8_, n310 );
dff P1_D_REG_6__reg ( clk, reset, P1_D_REG_6_, n300 );
dff P1_D_REG_5__reg ( clk, reset, P1_D_REG_5_, n295 );
dff P1_D_REG_4__reg ( clk, reset, P1_D_REG_4_, n290 );
dff P1_D_REG_3__reg ( clk, reset, P1_D_REG_3_, n285 );
dff P1_D_REG_2__reg ( clk, reset, P1_D_REG_2_, n280 );
dff P1_D_REG_22__reg ( clk, reset, ex_wire8, n380 );
not U_inv46 ( n11129, ex_wire8 );
dff P1_D_REG_7__reg ( clk, reset, ex_wire9, n305 );
not U_inv47 ( n11128, ex_wire9 );
dff P1_D_REG_1__reg ( clk, reset, P1_D_REG_1_, n275 );
dff P1_D_REG_0__reg ( clk, reset, P1_D_REG_0_, n270 );
dff P1_REG1_REG_31__reg ( clk, reset, P1_REG1_REG_31_, n745 );
not U_inv48 ( n11130, P1_REG1_REG_31_ );
dff P1_REG1_REG_30__reg ( clk, reset, P1_REG1_REG_30_, n740 );
not U_inv49 ( n11132, P1_REG1_REG_30_ );
dff P1_REG1_REG_29__reg ( clk, reset, P1_REG1_REG_29_, n735 );
not U_inv50 ( n11147, P1_REG1_REG_29_ );
dff P1_REG1_REG_28__reg ( clk, reset, P1_REG1_REG_28_, n730 );
not U_inv51 ( n11142, P1_REG1_REG_28_ );
dff P1_REG1_REG_26__reg ( clk, reset, P1_REG1_REG_26_, n720 );
not U_inv52 ( n11127, P1_REG1_REG_26_ );
dff P1_REG1_REG_25__reg ( clk, reset, P1_REG1_REG_25_, n715 );
not U_inv53 ( n11125, P1_REG1_REG_25_ );
dff P1_REG1_REG_24__reg ( clk, reset, P1_REG1_REG_24_, n710 );
not U_inv54 ( n11124, P1_REG1_REG_24_ );
dff P1_REG1_REG_23__reg ( clk, reset, P1_REG1_REG_23_, n705 );
not U_inv55 ( n11109, P1_REG1_REG_23_ );
dff P1_REG1_REG_22__reg ( clk, reset, P1_REG1_REG_22_, n700 );
not U_inv56 ( n11105, P1_REG1_REG_22_ );
dff P1_REG1_REG_21__reg ( clk, reset, P1_REG1_REG_21_, n695 );
not U_inv57 ( n11089, P1_REG1_REG_21_ );
dff P1_REG1_REG_20__reg ( clk, reset, P1_REG1_REG_20_, n690 );
not U_inv58 ( n11091, P1_REG1_REG_20_ );
dff P1_REG1_REG_18__reg ( clk, reset, P1_REG1_REG_18_, n680 );
not U_inv59 ( n11093, P1_REG1_REG_18_ );
dff P1_REG1_REG_17__reg ( clk, reset, P1_REG1_REG_17_, n675 );
not U_inv60 ( n11085, P1_REG1_REG_17_ );
dff P1_REG1_REG_16__reg ( clk, reset, P1_REG1_REG_16_, n670 );
not U_inv61 ( n11076, P1_REG1_REG_16_ );
dff P1_REG1_REG_12__reg ( clk, reset, P1_REG1_REG_12_, n650 );
not U_inv62 ( n11051, P1_REG1_REG_12_ );
dff P1_REG1_REG_3__reg ( clk, reset, P1_REG1_REG_3_, n605 );
not U_inv63 ( n10982, P1_REG1_REG_3_ );
dff P1_IR_REG_29__reg ( clk, reset, P1_IR_REG_29_, n255 );
dff P1_IR_REG_28__reg ( clk, reset, P1_IR_REG_28_, n250 );
dff P1_RD_REG_reg ( clk, reset, P1_RD_REG, n1325 );
dff P1_REG2_REG_31__reg ( clk, reset, ex_wire10, n905 );
not U_inv64 ( n11131, ex_wire10 );
dff P1_REG1_REG_1__reg ( clk, reset, P1_REG1_REG_1_, n595 );
not U_inv65 ( n10973, P1_REG1_REG_1_ );
dff P1_REG0_REG_1__reg ( clk, reset, P1_REG0_REG_1_, n435 );
dff P1_REG1_REG_0__reg ( clk, reset, P1_REG1_REG_0_, n590 );
not U_inv66 ( n10963, P1_REG1_REG_0_ );
dff P1_REG0_REG_0__reg ( clk, reset, P1_REG0_REG_0_, n430 );
dff P1_REG3_REG_0__reg ( clk, reset, ex_wire11, n1220 );
not U_inv67 ( n10965, ex_wire11 );
dff P1_REG2_REG_0__reg ( clk, reset, P1_REG2_REG_0_, n750 );
not U_inv68 ( n10964, P1_REG2_REG_0_ );
dff P1_REG1_REG_2__reg ( clk, reset, P1_REG1_REG_2_, n600 );
not U_inv69 ( n10977, P1_REG1_REG_2_ );
dff P1_REG0_REG_2__reg ( clk, reset, P1_REG0_REG_2_, n440 );
dff P1_REG3_REG_1__reg ( clk, reset, P1_REG3_REG_1_, n1270 );
not U_inv70 ( n10972, P1_REG3_REG_1_ );
dff P1_REG2_REG_1__reg ( clk, reset, P1_REG2_REG_1_, n755 );
not U_inv71 ( n10974, P1_REG2_REG_1_ );
dff P1_REG3_REG_2__reg ( clk, reset, P1_REG3_REG_2_, n1195 );
not U_inv72 ( n10976, P1_REG3_REG_2_ );
dff P1_REG2_REG_2__reg ( clk, reset, P1_REG2_REG_2_, n760 );
not U_inv73 ( n10975, P1_REG2_REG_2_ );
dff P1_DATAO_REG_2__reg ( clk, reset, P1_DATAO_REG_2_, n1020 );
dff P1_REG1_REG_10__reg ( clk, reset, P1_REG1_REG_10_, n640 );
not U_inv74 ( n11043, P1_REG1_REG_10_ );
dff P1_REG0_REG_10__reg ( clk, reset, P1_REG0_REG_10_, n480 );
dff P1_REG2_REG_9__reg ( clk, reset, P1_REG2_REG_9_, n795 );
not U_inv75 ( n11044, P1_REG2_REG_9_ );
dff P1_REG2_REG_8__reg ( clk, reset, P1_REG2_REG_8_, n790 );
not U_inv76 ( n11032, P1_REG2_REG_8_ );
dff P1_REG2_REG_7__reg ( clk, reset, P1_REG2_REG_7_, n785 );
not U_inv77 ( n11024, P1_REG2_REG_7_ );
dff P1_REG2_REG_6__reg ( clk, reset, P1_REG2_REG_6_, n780 );
not U_inv78 ( n11020, P1_REG2_REG_6_ );
dff P1_REG2_REG_5__reg ( clk, reset, P1_REG2_REG_5_, n775 );
not U_inv79 ( n11011, P1_REG2_REG_5_ );
dff P1_REG2_REG_4__reg ( clk, reset, P1_REG2_REG_4_, n770 );
not U_inv80 ( n11007, P1_REG2_REG_4_ );
dff P1_REG3_REG_3__reg ( clk, reset, P1_REG3_REG_3_, n1290 );
not U_inv81 ( n11002, P1_REG3_REG_3_ );
dff P1_REG2_REG_3__reg ( clk, reset, P1_REG2_REG_3_, n765 );
not U_inv82 ( n10981, P1_REG2_REG_3_ );
dff P1_DATAO_REG_4__reg ( clk, reset, P1_DATAO_REG_4_, n1030 );
dff P1_IR_REG_4__reg ( clk, reset, P1_IR_REG_4_, n130 );
dff P1_REG3_REG_4__reg ( clk, reset, P1_REG3_REG_4_, n1230 );
not U_inv83 ( n11165, P1_REG3_REG_4_ );
dff P1_REG1_REG_4__reg ( clk, reset, P1_REG1_REG_4_, n610 );
not U_inv84 ( n11009, P1_REG1_REG_4_ );
dff P1_REG0_REG_4__reg ( clk, reset, P1_REG0_REG_4_, n450 );
dff P1_DATAO_REG_5__reg ( clk, reset, P1_DATAO_REG_5_, n1035 );
dff P2_IR_REG_5__reg ( clk, reset, P2_IR_REG_5_, n1360 );
dff P1_IR_REG_5__reg ( clk, reset, P1_IR_REG_5_, n135 );
dff P1_REG3_REG_5__reg ( clk, reset, ex_wire12, n1245 );
not U_inv85 ( n11003, ex_wire12 );
dff P1_REG1_REG_5__reg ( clk, reset, P1_REG1_REG_5_, n615 );
not U_inv86 ( n11012, P1_REG1_REG_5_ );
dff P1_REG0_REG_5__reg ( clk, reset, P1_REG0_REG_5_, n455 );
dff P1_DATAO_REG_6__reg ( clk, reset, P1_DATAO_REG_6_, n1040 );
dff P1_IR_REG_6__reg ( clk, reset, P1_IR_REG_6_, n140 );
dff P1_REG3_REG_6__reg ( clk, reset, P1_REG3_REG_6_, n1185 );
not U_inv87 ( n11164, P1_REG3_REG_6_ );
dff P1_REG1_REG_6__reg ( clk, reset, P1_REG1_REG_6_, n620 );
not U_inv88 ( n11023, P1_REG1_REG_6_ );
dff P1_REG0_REG_6__reg ( clk, reset, P1_REG0_REG_6_, n460 );
dff P1_DATAO_REG_7__reg ( clk, reset, P1_DATAO_REG_7_, n1045 );
dff P2_IR_REG_7__reg ( clk, reset, P2_IR_REG_7_, n1370 );
not U_inv89 ( n10978, P2_IR_REG_7_ );
dff P1_IR_REG_7__reg ( clk, reset, P1_IR_REG_7_, n145 );
not U_inv90 ( n11008, P1_IR_REG_7_ );
dff P1_REG3_REG_7__reg ( clk, reset, ex_wire13, n1315 );
not U_inv91 ( n10955, ex_wire13 );
dff P1_REG1_REG_7__reg ( clk, reset, P1_REG1_REG_7_, n625 );
not U_inv92 ( n11025, P1_REG1_REG_7_ );
dff P1_REG0_REG_7__reg ( clk, reset, P1_REG0_REG_7_, n465 );
dff P1_DATAO_REG_8__reg ( clk, reset, P1_DATAO_REG_8_, n1050 );
dff P2_IR_REG_8__reg ( clk, reset, P2_IR_REG_8_, n1375 );
dff P1_IR_REG_8__reg ( clk, reset, P1_IR_REG_8_, n150 );
dff P1_REG3_REG_8__reg ( clk, reset, P1_REG3_REG_8_, n1275 );
not U_inv93 ( n11163, P1_REG3_REG_8_ );
dff P1_REG1_REG_8__reg ( clk, reset, P1_REG1_REG_8_, n630 );
not U_inv94 ( n11034, P1_REG1_REG_8_ );
dff P1_REG0_REG_8__reg ( clk, reset, P1_REG0_REG_8_, n470 );
dff P1_DATAO_REG_9__reg ( clk, reset, P1_DATAO_REG_9_, n1055 );
dff P2_IR_REG_9__reg ( clk, reset, P2_IR_REG_9_, n1380 );
dff P1_IR_REG_9__reg ( clk, reset, P1_IR_REG_9_, n155 );
dff P1_REG3_REG_9__reg ( clk, reset, ex_wire14, n1225 );
not U_inv95 ( n11026, ex_wire14 );
dff P1_REG1_REG_9__reg ( clk, reset, P1_REG1_REG_9_, n635 );
not U_inv96 ( n11045, P1_REG1_REG_9_ );
dff P1_REG0_REG_9__reg ( clk, reset, P1_REG0_REG_9_, n475 );
dff P1_REG1_REG_11__reg ( clk, reset, P1_REG1_REG_11_, n645 );
not U_inv97 ( n11053, P1_REG1_REG_11_ );
dff P1_REG0_REG_11__reg ( clk, reset, P1_REG0_REG_11_, n485 );
dff P1_REG3_REG_10__reg ( clk, reset, P1_REG3_REG_10_, n1295 );
not U_inv98 ( n11162, P1_REG3_REG_10_ );
dff P1_REG2_REG_10__reg ( clk, reset, P1_REG2_REG_10_, n800 );
not U_inv99 ( n11041, P1_REG2_REG_10_ );
dff P1_DATAO_REG_11__reg ( clk, reset, P1_DATAO_REG_11_, n1065 );
dff P1_IR_REG_11__reg ( clk, reset, P1_IR_REG_11_, n165 );
not U_inv100 ( n11037, P1_IR_REG_11_ );
dff P1_IR_REG_12__reg ( clk, reset, P1_IR_REG_12_, n170 );
dff P1_REG3_REG_11__reg ( clk, reset, ex_wire15, n1200 );
not U_inv101 ( n11030, ex_wire15 );
dff P1_REG2_REG_11__reg ( clk, reset, P1_REG2_REG_11_, n805 );
not U_inv102 ( n11052, P1_REG2_REG_11_ );
dff P1_IR_REG_13__reg ( clk, reset, P1_IR_REG_13_, n175 );
dff P1_REG1_REG_13__reg ( clk, reset, P1_REG1_REG_13_, n655 );
not U_inv103 ( n11047, P1_REG1_REG_13_ );
dff P1_REG0_REG_13__reg ( clk, reset, P1_REG0_REG_13_, n495 );
dff P1_REG3_REG_12__reg ( clk, reset, P1_REG3_REG_12_, n1260 );
not U_inv104 ( n11161, P1_REG3_REG_12_ );
dff P1_REG2_REG_12__reg ( clk, reset, P1_REG2_REG_12_, n810 );
not U_inv105 ( n11049, P1_REG2_REG_12_ );
dff P1_DATAO_REG_13__reg ( clk, reset, P1_DATAO_REG_13_, n1075 );
dff P1_IR_REG_14__reg ( clk, reset, P1_IR_REG_14_, n180 );
dff P1_REG1_REG_14__reg ( clk, reset, P1_REG1_REG_14_, n660 );
not U_inv106 ( n11074, P1_REG1_REG_14_ );
dff P1_REG0_REG_14__reg ( clk, reset, P1_REG0_REG_14_, n500 );
dff P1_REG3_REG_13__reg ( clk, reset, ex_wire16, n1210 );
not U_inv107 ( n11042, ex_wire16 );
dff P1_REG2_REG_13__reg ( clk, reset, P1_REG2_REG_13_, n815 );
not U_inv108 ( n11046, P1_REG2_REG_13_ );
dff P1_REG3_REG_14__reg ( clk, reset, P1_REG3_REG_14_, n1305 );
not U_inv109 ( n11160, P1_REG3_REG_14_ );
dff P1_REG2_REG_16__reg ( clk, reset, P1_REG2_REG_16_, n830 );
not U_inv110 ( n11075, P1_REG2_REG_16_ );
dff P1_REG3_REG_16__reg ( clk, reset, P1_REG3_REG_16_, n1250 );
not U_inv111 ( n11159, P1_REG3_REG_16_ );
dff P1_REG3_REG_17__reg ( clk, reset, ex_wire17, n1240 );
not U_inv112 ( n11066, ex_wire17 );
dff P1_REG3_REG_18__reg ( clk, reset, P1_REG3_REG_18_, n1190 );
not U_inv113 ( n11158, P1_REG3_REG_18_ );
dff P1_REG2_REG_14__reg ( clk, reset, P1_REG2_REG_14_, n820 );
not U_inv114 ( n11071, P1_REG2_REG_14_ );
dff P1_DATAO_REG_14__reg ( clk, reset, P1_DATAO_REG_14_, n1080 );
dff P1_DATAO_REG_10__reg ( clk, reset, P1_DATAO_REG_10_, n1060 );
dff P2_IR_REG_10__reg ( clk, reset, P2_IR_REG_10_, n1385 );
dff P2_IR_REG_11__reg ( clk, reset, P2_IR_REG_11_, n1390 );
not U_inv115 ( n11010, P2_IR_REG_11_ );
dff P2_IR_REG_13__reg ( clk, reset, P2_IR_REG_13_, n1400 );
dff P2_IR_REG_14__reg ( clk, reset, P2_IR_REG_14_, n1405 );
dff P2_IR_REG_15__reg ( clk, reset, P2_IR_REG_15_, n1410 );
not U_inv116 ( n11038, P2_IR_REG_15_ );
dff P2_IR_REG_12__reg ( clk, reset, P2_IR_REG_12_, n1395 );
dff P1_IR_REG_10__reg ( clk, reset, P1_IR_REG_10_, n160 );
dff P1_REG1_REG_19__reg ( clk, reset, P1_REG1_REG_19_, n685 );
not U_inv117 ( n11087, P1_REG1_REG_19_ );
dff P1_REG0_REG_19__reg ( clk, reset, P1_REG0_REG_19_, n525 );
dff P1_REG3_REG_20__reg ( clk, reset, P1_REG3_REG_20_, n1215 );
dff P1_REG2_REG_21__reg ( clk, reset, ex_wire18, n855 );
not U_inv118 ( n11088, ex_wire18 );
dff P1_REG3_REG_21__reg ( clk, reset, ex_wire19, n1265 );
not U_inv119 ( n11077, ex_wire19 );
dff P1_REG3_REG_22__reg ( clk, reset, P1_REG3_REG_22_, n1205 );
dff P1_REG3_REG_23__reg ( clk, reset, ex_wire20, n1300 );
not U_inv120 ( n11100, ex_wire20 );
dff P1_REG3_REG_24__reg ( clk, reset, P1_REG3_REG_24_, n1235 );
dff P1_REG3_REG_25__reg ( clk, reset, ex_wire21, n1255 );
not U_inv121 ( n11108, ex_wire21 );
dff P1_REG1_REG_15__reg ( clk, reset, P1_REG1_REG_15_, n665 );
not U_inv122 ( n11068, P1_REG1_REG_15_ );
dff P1_REG0_REG_15__reg ( clk, reset, P1_REG0_REG_15_, n505 );
dff P1_DATAO_REG_3__reg ( clk, reset, P1_DATAO_REG_3_, n1025 );
dff P2_IR_REG_1__reg ( clk, reset, P2_IR_REG_1_, n1340 );
dff P1_ADDR_REG_2__reg ( clk, reset, P1_ADDR_REG_2_, n995 );
dff P1_ADDR_REG_3__reg ( clk, reset, P1_ADDR_REG_3_, n990 );
dff P1_ADDR_REG_4__reg ( clk, reset, P1_ADDR_REG_4_, n985 );
dff P1_ADDR_REG_5__reg ( clk, reset, P1_ADDR_REG_5_, n980 );
dff P1_ADDR_REG_6__reg ( clk, reset, P1_ADDR_REG_6_, n975 );
dff P1_ADDR_REG_7__reg ( clk, reset, P1_ADDR_REG_7_, n970 );
dff P1_ADDR_REG_8__reg ( clk, reset, P1_ADDR_REG_8_, n965 );
dff P1_ADDR_REG_9__reg ( clk, reset, P1_ADDR_REG_9_, n960 );
dff P1_ADDR_REG_10__reg ( clk, reset, P1_ADDR_REG_10_, n955 );
dff P1_ADDR_REG_11__reg ( clk, reset, P1_ADDR_REG_11_, n950 );
dff P1_ADDR_REG_12__reg ( clk, reset, P1_ADDR_REG_12_, n945 );
dff P1_ADDR_REG_13__reg ( clk, reset, P1_ADDR_REG_13_, n940 );
dff P1_ADDR_REG_14__reg ( clk, reset, P1_ADDR_REG_14_, n935 );
dff P1_ADDR_REG_15__reg ( clk, reset, P1_ADDR_REG_15_, n930 );
dff P1_ADDR_REG_16__reg ( clk, reset, P1_ADDR_REG_16_, n925 );
dff P1_REG3_REG_26__reg ( clk, reset, P1_REG3_REG_26_, n1180 );
dff P1_REG1_REG_27__reg ( clk, reset, P1_REG1_REG_27_, n725 );
not U_inv123 ( n11137, P1_REG1_REG_27_ );
dff P1_REG0_REG_27__reg ( clk, reset, P1_REG0_REG_27_, n565 );
dff P1_REG2_REG_26__reg ( clk, reset, ex_wire22, n880 );
not U_inv124 ( n11126, ex_wire22 );
dff P1_REG2_REG_25__reg ( clk, reset, ex_wire23, n875 );
not U_inv125 ( n11123, ex_wire23 );
dff P1_REG2_REG_24__reg ( clk, reset, ex_wire24, n870 );
not U_inv126 ( n11122, ex_wire24 );
dff P1_REG2_REG_23__reg ( clk, reset, ex_wire25, n865 );
not U_inv127 ( n11107, ex_wire25 );
dff P1_REG2_REG_22__reg ( clk, reset, ex_wire26, n860 );
not U_inv128 ( n11104, ex_wire26 );
dff P1_REG2_REG_20__reg ( clk, reset, ex_wire27, n850 );
not U_inv129 ( n11090, ex_wire27 );
dff P1_REG2_REG_18__reg ( clk, reset, P1_REG2_REG_18_, n840 );
not U_inv130 ( n11092, P1_REG2_REG_18_ );
dff P1_REG2_REG_17__reg ( clk, reset, P1_REG2_REG_17_, n835 );
not U_inv131 ( n11084, P1_REG2_REG_17_ );
dff P1_ADDR_REG_17__reg ( clk, reset, P1_ADDR_REG_17_, n920 );
dff P1_ADDR_REG_18__reg ( clk, reset, P1_ADDR_REG_18_, n915 );
not U_inv132 ( n11106, P1_ADDR_REG_18_ );
dff P1_ADDR_REG_19__reg ( clk, reset, P1_ADDR_REG_19_, n910 );
not U_inv133 ( n10959, P1_ADDR_REG_19_ );
dff P1_DATAO_REG_16__reg ( clk, reset, P1_DATAO_REG_16_, n1090 );
dff P2_IR_REG_16__reg ( clk, reset, P2_IR_REG_16_, n1415 );
dff P2_IR_REG_17__reg ( clk, reset, P2_IR_REG_17_, n1420 );
dff P2_IR_REG_18__reg ( clk, reset, P2_IR_REG_18_, n1425 );
dff P2_IR_REG_19__reg ( clk, reset, P2_IR_REG_19_, n1430 );
not U_inv134 ( n10996, P2_IR_REG_19_ );
dff P2_IR_REG_20__reg ( clk, reset, P2_IR_REG_20_, n1435 );
dff P1_IR_REG_16__reg ( clk, reset, P1_IR_REG_16_, n190 );
dff P1_IR_REG_2__reg ( clk, reset, P1_IR_REG_2_, n120 );
dff P2_DATAO_REG_0__reg ( clk, reset, P2_DATAO_REG_0_, n2235 );
dff P2_REG1_REG_29__reg ( clk, reset, P2_REG1_REG_29_, n1960 );
not U_inv135 ( n11150, P2_REG1_REG_29_ );
dff P2_REG1_REG_27__reg ( clk, reset, P2_REG1_REG_27_, n1950 );
not U_inv136 ( n11141, P2_REG1_REG_27_ );
dff P2_REG1_REG_26__reg ( clk, reset, P2_REG1_REG_26_, n1945 );
not U_inv137 ( n11117, P2_REG1_REG_26_ );
dff P2_REG1_REG_25__reg ( clk, reset, P2_REG1_REG_25_, n1940 );
not U_inv138 ( n11114, P2_REG1_REG_25_ );
dff P2_REG1_REG_24__reg ( clk, reset, P2_REG1_REG_24_, n1935 );
not U_inv139 ( n11120, P2_REG1_REG_24_ );
dff P2_REG1_REG_23__reg ( clk, reset, P2_REG1_REG_23_, n1930 );
not U_inv140 ( n11103, P2_REG1_REG_23_ );
dff P2_REG1_REG_22__reg ( clk, reset, P2_REG1_REG_22_, n1925 );
not U_inv141 ( n11099, P2_REG1_REG_22_ );
dff P2_REG1_REG_21__reg ( clk, reset, P2_REG1_REG_21_, n1920 );
not U_inv142 ( n11096, P2_REG1_REG_21_ );
dff P2_REG1_REG_20__reg ( clk, reset, P2_REG1_REG_20_, n1915 );
not U_inv143 ( n11082, P2_REG1_REG_20_ );
dff P2_REG1_REG_19__reg ( clk, reset, P2_REG1_REG_19_, n1910 );
not U_inv144 ( n11078, P2_REG1_REG_19_ );
dff P2_REG1_REG_18__reg ( clk, reset, P2_REG1_REG_18_, n1905 );
not U_inv145 ( n11070, P2_REG1_REG_18_ );
dff P2_REG1_REG_17__reg ( clk, reset, P2_REG1_REG_17_, n1900 );
not U_inv146 ( n11064, P2_REG1_REG_17_ );
dff P2_REG1_REG_16__reg ( clk, reset, P2_REG1_REG_16_, n1895 );
not U_inv147 ( n11061, P2_REG1_REG_16_ );
dff P2_REG1_REG_14__reg ( clk, reset, P2_REG1_REG_14_, n1885 );
not U_inv148 ( n11050, P2_REG1_REG_14_ );
dff P2_REG1_REG_12__reg ( clk, reset, P2_REG1_REG_12_, n1875 );
not U_inv149 ( n11033, P2_REG1_REG_12_ );
dff P2_REG1_REG_11__reg ( clk, reset, P2_REG1_REG_11_, n1870 );
not U_inv150 ( n11028, P2_REG1_REG_11_ );
dff P2_REG1_REG_10__reg ( clk, reset, P2_REG1_REG_10_, n1865 );
not U_inv151 ( n11015, P2_REG1_REG_10_ );
dff P2_REG1_REG_8__reg ( clk, reset, P2_REG1_REG_8_, n1855 );
not U_inv152 ( n11017, P2_REG1_REG_8_ );
dff P2_REG1_REG_7__reg ( clk, reset, P2_REG1_REG_7_, n1850 );
not U_inv153 ( n11005, P2_REG1_REG_7_ );
dff P2_REG1_REG_6__reg ( clk, reset, P2_REG1_REG_6_, n1845 );
not U_inv154 ( n11000, P2_REG1_REG_6_ );
dff P2_REG1_REG_5__reg ( clk, reset, P2_REG1_REG_5_, n1840 );
not U_inv155 ( n10980, P2_REG1_REG_5_ );
dff P2_REG1_REG_4__reg ( clk, reset, P2_REG1_REG_4_, n1835 );
not U_inv156 ( n10995, P2_REG1_REG_4_ );
dff P2_REG1_REG_2__reg ( clk, reset, P2_REG1_REG_2_, n1825 );
not U_inv157 ( n10991, P2_REG1_REG_2_ );
dff P2_REG1_REG_1__reg ( clk, reset, P2_REG1_REG_1_, n1820 );
not U_inv158 ( n10986, P2_REG1_REG_1_ );
dff P2_REG1_REG_0__reg ( clk, reset, P2_REG1_REG_0_, n1815 );
not U_inv159 ( n10967, P2_REG1_REG_0_ );
dff P2_REG3_REG_3__reg ( clk, reset, P2_REG3_REG_3_, n2515 );
not U_inv160 ( n10958, P2_REG3_REG_3_ );
dff P2_REG3_REG_1__reg ( clk, reset, P2_REG3_REG_1_, n2495 );
not U_inv161 ( n10987, P2_REG3_REG_1_ );
dff P2_REG3_REG_16__reg ( clk, reset, P2_REG3_REG_16_, n2475 );
not U_inv162 ( n11179, P2_REG3_REG_16_ );
dff P2_REG3_REG_17__reg ( clk, reset, P2_REG3_REG_17_, n2465 );
not U_inv163 ( n11178, P2_REG3_REG_17_ );
dff P2_REG2_REG_17__reg ( clk, reset, P2_REG2_REG_17_, n2060 );
not U_inv164 ( n11063, P2_REG2_REG_17_ );
dff P2_REG3_REG_4__reg ( clk, reset, P2_REG3_REG_4_, n2455 );
not U_inv165 ( n10970, P2_REG3_REG_4_ );
dff P2_REG3_REG_5__reg ( clk, reset, P2_REG3_REG_5_, n2470 );
not U_inv166 ( n11177, P2_REG3_REG_5_ );
dff P2_REG3_REG_2__reg ( clk, reset, P2_REG3_REG_2_, n2420 );
not U_inv167 ( n10992, P2_REG3_REG_2_ );
dff P2_REG3_REG_18__reg ( clk, reset, P2_REG3_REG_18_, n2415 );
not U_inv168 ( n11176, P2_REG3_REG_18_ );
dff P2_REG3_REG_19__reg ( clk, reset, P2_REG3_REG_19_, n2510 );
not U_inv169 ( n11175, P2_REG3_REG_19_ );
dff P2_REG2_REG_18__reg ( clk, reset, P2_REG2_REG_18_, n2065 );
not U_inv170 ( n11069, P2_REG2_REG_18_ );
dff P2_REG3_REG_6__reg ( clk, reset, P2_REG3_REG_6_, n2410 );
not U_inv171 ( n11174, P2_REG3_REG_6_ );
dff P2_REG3_REG_14__reg ( clk, reset, P2_REG3_REG_14_, n2530 );
not U_inv172 ( n11173, P2_REG3_REG_14_ );
dff P2_REG3_REG_13__reg ( clk, reset, P2_REG3_REG_13_, n2435 );
not U_inv173 ( n11172, P2_REG3_REG_13_ );
dff P2_REG3_REG_12__reg ( clk, reset, P2_REG3_REG_12_, n2485 );
not U_inv174 ( n11171, P2_REG3_REG_12_ );
dff P2_REG2_REG_12__reg ( clk, reset, P2_REG2_REG_12_, n2035 );
not U_inv175 ( n11031, P2_REG2_REG_12_ );
dff P2_REG3_REG_11__reg ( clk, reset, P2_REG3_REG_11_, n2425 );
not U_inv176 ( n11170, P2_REG3_REG_11_ );
dff P2_REG3_REG_10__reg ( clk, reset, P2_REG3_REG_10_, n2520 );
not U_inv177 ( n11169, P2_REG3_REG_10_ );
dff P2_REG2_REG_10__reg ( clk, reset, P2_REG2_REG_10_, n2025 );
not U_inv178 ( n11013, P2_REG2_REG_10_ );
dff P2_REG3_REG_9__reg ( clk, reset, P2_REG3_REG_9_, n2450 );
not U_inv179 ( n11168, P2_REG3_REG_9_ );
dff P2_REG3_REG_8__reg ( clk, reset, P2_REG3_REG_8_, n2500 );
not U_inv180 ( n11167, P2_REG3_REG_8_ );
dff P2_REG3_REG_7__reg ( clk, reset, P2_REG3_REG_7_, n2540 );
not U_inv181 ( n11166, P2_REG3_REG_7_ );
dff P2_REG2_REG_7__reg ( clk, reset, P2_REG2_REG_7_, n2010 );
not U_inv182 ( n11004, P2_REG2_REG_7_ );
dff P2_REG3_REG_0__reg ( clk, reset, P2_REG3_REG_0_, n2445 );
not U_inv183 ( n10968, P2_REG3_REG_0_ );
dff P2_REG3_REG_20__reg ( clk, reset, P2_REG3_REG_20_, n2440 );
dff P2_REG3_REG_21__reg ( clk, reset, P2_REG3_REG_21_, n2490 );
dff P2_REG3_REG_22__reg ( clk, reset, P2_REG3_REG_22_, n2430 );
dff P2_REG3_REG_25__reg ( clk, reset, P2_REG3_REG_25_, n2480 );
dff P2_REG3_REG_24__reg ( clk, reset, P2_REG3_REG_24_, n2460 );
dff P2_REG3_REG_23__reg ( clk, reset, P2_REG3_REG_23_, n2525 );
dff P2_REG3_REG_26__reg ( clk, reset, P2_REG3_REG_26_, n2405 );
dff P2_REG3_REG_28__reg ( clk, reset, P2_REG3_REG_28_, n2505 );
dff P2_REG3_REG_27__reg ( clk, reset, P2_REG3_REG_27_, n2535 );
dff P2_REG2_REG_15__reg ( clk, reset, P2_REG2_REG_15_, n2050 );
not U_inv184 ( n11056, P2_REG2_REG_15_ );
dff P2_REG1_REG_15__reg ( clk, reset, P2_REG1_REG_15_, n1890 );
not U_inv185 ( n11057, P2_REG1_REG_15_ );
dff P2_REG1_REG_13__reg ( clk, reset, P2_REG1_REG_13_, n1880 );
not U_inv186 ( n11039, P2_REG1_REG_13_ );
dff P2_REG0_REG_31__reg ( clk, reset, P2_REG0_REG_31_, n1810 );
not U_inv187 ( n11152, P2_REG0_REG_31_ );
dff P2_REG2_REG_31__reg ( clk, reset, ex_wire28, n2130 );
not U_inv188 ( n11151, ex_wire28 );
dff P2_REG2_REG_30__reg ( clk, reset, ex_wire29, n2125 );
not U_inv189 ( n11154, ex_wire29 );
dff P2_REG1_REG_31__reg ( clk, reset, P2_REG1_REG_31_, n1970 );
not U_inv190 ( n11153, P2_REG1_REG_31_ );
dff P2_REG1_REG_30__reg ( clk, reset, P2_REG1_REG_30_, n1965 );
not U_inv191 ( n11156, P2_REG1_REG_30_ );
dff P2_DATAO_REG_31__reg ( clk, reset, P2_DATAO_REG_31_, n2390 );
dff P2_REG0_REG_30__reg ( clk, reset, P2_REG0_REG_30_, n1805 );
not U_inv192 ( n11155, P2_REG0_REG_30_ );
dff P2_DATAO_REG_30__reg ( clk, reset, P2_DATAO_REG_30_, n2385 );
dff P2_REG0_REG_15__reg ( clk, reset, P2_REG0_REG_15_, n1730 );
not U_inv193 ( n11058, P2_REG0_REG_15_ );
dff P2_REG0_REG_13__reg ( clk, reset, P2_REG0_REG_13_, n1720 );
not U_inv194 ( n11040, P2_REG0_REG_13_ );
dff P2_REG1_REG_9__reg ( clk, reset, P2_REG1_REG_9_, n1860 );
not U_inv195 ( n11018, P2_REG1_REG_9_ );
dff P2_REG0_REG_9__reg ( clk, reset, P2_REG0_REG_9_, n1700 );
not U_inv196 ( n11022, P2_REG0_REG_9_ );
dff P2_REG1_REG_3__reg ( clk, reset, P2_REG1_REG_3_, n1830 );
not U_inv197 ( n10985, P2_REG1_REG_3_ );
dff P2_REG0_REG_3__reg ( clk, reset, P2_REG0_REG_3_, n1670 );
not U_inv198 ( n10993, P2_REG0_REG_3_ );
dff P1_REG2_REG_30__reg ( clk, reset, ex_wire30, n900 );
not U_inv199 ( n11133, ex_wire30 );
dff P1_REG3_REG_28__reg ( clk, reset, P1_REG3_REG_28_, n1280 );
dff P1_REG2_REG_28__reg ( clk, reset, ex_wire31, n890 );
not U_inv200 ( n11138, ex_wire31 );
dff P2_REG1_REG_28__reg ( clk, reset, P2_REG1_REG_28_, n1955 );
not U_inv201 ( n11146, P2_REG1_REG_28_ );
dff P2_REG0_REG_28__reg ( clk, reset, P2_REG0_REG_28_, n1795 );
not U_inv202 ( n11145, P2_REG0_REG_28_ );
dff P2_REG2_REG_21__reg ( clk, reset, ex_wire32, n2080 );
not U_inv203 ( n11094, ex_wire32 );
dff P2_REG2_REG_20__reg ( clk, reset, ex_wire33, n2075 );
not U_inv204 ( n11080, ex_wire33 );
dff P2_REG2_REG_19__reg ( clk, reset, ex_wire34, n2070 );
not U_inv205 ( n11079, ex_wire34 );
dff P2_REG2_REG_14__reg ( clk, reset, P2_REG2_REG_14_, n2045 );
not U_inv206 ( n11048, P2_REG2_REG_14_ );
dff P2_REG2_REG_11__reg ( clk, reset, P2_REG2_REG_11_, n2030 );
not U_inv207 ( n11027, P2_REG2_REG_11_ );
dff P2_REG2_REG_5__reg ( clk, reset, P2_REG2_REG_5_, n2000 );
not U_inv208 ( n10979, P2_REG2_REG_5_ );
dff P2_REG2_REG_6__reg ( clk, reset, P2_REG2_REG_6_, n2005 );
not U_inv209 ( n10998, P2_REG2_REG_6_ );
dff P2_REG2_REG_4__reg ( clk, reset, P2_REG2_REG_4_, n1995 );
not U_inv210 ( n10988, P2_REG2_REG_4_ );
dff P2_REG2_REG_2__reg ( clk, reset, P2_REG2_REG_2_, n1985 );
not U_inv211 ( n10989, P2_REG2_REG_2_ );
dff P2_REG2_REG_1__reg ( clk, reset, P2_REG2_REG_1_, n1980 );
not U_inv212 ( n10984, P2_REG2_REG_1_ );
dff P2_REG2_REG_0__reg ( clk, reset, P2_REG2_REG_0_, n1975 );
not U_inv213 ( n10966, P2_REG2_REG_0_ );
dff P2_ADDR_REG_1__reg ( clk, reset, P2_ADDR_REG_1_, n2225 );
dff P2_ADDR_REG_2__reg ( clk, reset, P2_ADDR_REG_2_, n2220 );
dff P2_ADDR_REG_3__reg ( clk, reset, P2_ADDR_REG_3_, n2215 );
dff P2_ADDR_REG_4__reg ( clk, reset, P2_ADDR_REG_4_, n2210 );
dff P2_ADDR_REG_5__reg ( clk, reset, P2_ADDR_REG_5_, n2205 );
dff P2_ADDR_REG_6__reg ( clk, reset, P2_ADDR_REG_6_, n2200 );
dff P2_ADDR_REG_7__reg ( clk, reset, P2_ADDR_REG_7_, n2195 );
dff P2_ADDR_REG_0__reg ( clk, reset, P2_ADDR_REG_0_, n2230 );
dff P2_REG2_REG_29__reg ( clk, reset, ex_wire35, n2120 );
not U_inv214 ( n11148, ex_wire35 );
dff P2_REG2_REG_27__reg ( clk, reset, ex_wire36, n2110 );
not U_inv215 ( n11139, ex_wire36 );
dff P2_REG2_REG_26__reg ( clk, reset, ex_wire37, n2105 );
not U_inv216 ( n11115, ex_wire37 );
dff P2_REG2_REG_25__reg ( clk, reset, ex_wire38, n2100 );
not U_inv217 ( n11112, ex_wire38 );
dff P2_REG2_REG_24__reg ( clk, reset, ex_wire39, n2095 );
not U_inv218 ( n11118, ex_wire39 );
dff P2_REG2_REG_23__reg ( clk, reset, ex_wire40, n2090 );
not U_inv219 ( n11101, ex_wire40 );
dff P2_REG2_REG_22__reg ( clk, reset, ex_wire41, n2085 );
not U_inv220 ( n11097, ex_wire41 );
dff P2_REG2_REG_16__reg ( clk, reset, P2_REG2_REG_16_, n2055 );
not U_inv221 ( n11060, P2_REG2_REG_16_ );
dff P2_REG2_REG_8__reg ( clk, reset, P2_REG2_REG_8_, n2015 );
not U_inv222 ( n11014, P2_REG2_REG_8_ );
dff P2_ADDR_REG_8__reg ( clk, reset, P2_ADDR_REG_8_, n2190 );
dff P2_ADDR_REG_12__reg ( clk, reset, P2_ADDR_REG_12_, n2170 );
dff P2_ADDR_REG_13__reg ( clk, reset, P2_ADDR_REG_13_, n2165 );
dff P2_ADDR_REG_14__reg ( clk, reset, P2_ADDR_REG_14_, n2160 );
dff P2_ADDR_REG_17__reg ( clk, reset, P2_ADDR_REG_17_, n2145 );
dff P2_ADDR_REG_18__reg ( clk, reset, P2_ADDR_REG_18_, n2140 );
not U_inv223 ( n11110, P2_ADDR_REG_18_ );
dff P2_ADDR_REG_19__reg ( clk, reset, P2_ADDR_REG_19_, n2135 );
dff P2_ADDR_REG_15__reg ( clk, reset, P2_ADDR_REG_15_, n2155 );
dff P2_ADDR_REG_16__reg ( clk, reset, P2_ADDR_REG_16_, n2150 );
dff P2_ADDR_REG_9__reg ( clk, reset, P2_ADDR_REG_9_, n2185 );
dff P2_ADDR_REG_10__reg ( clk, reset, P2_ADDR_REG_10_, n2180 );
dff P2_ADDR_REG_11__reg ( clk, reset, P2_ADDR_REG_11_, n2175 );
dff P1_REG2_REG_29__reg ( clk, reset, ex_wire42, n895 );
not U_inv224 ( n11143, ex_wire42 );
dff P1_ADDR_REG_0__reg ( clk, reset, P1_ADDR_REG_0_, n1005 );
dff P1_ADDR_REG_1__reg ( clk, reset, ex_wire43, n1000 );
not U_inv225 ( n10962, ex_wire43 );
dff P2_WR_REG_reg ( clk, reset, P2_WR_REG, n11388 );
dff P2_IR_REG_31__reg ( clk, reset, P2_IR_REG_31_, n1490 );
dff P1_IR_REG_31__reg ( clk, reset, P1_IR_REG_31_, n265 );
not U10979 ( n344, n2719 );
nand U10980 ( n6777, n8146, n929 );
nand U10981 ( n6776, n8145, n4769 );
nor U10982 ( n2719, n348, n9387 );
nand U10983 ( n2774, n9385, n9384 );
nand U10984 ( n2775, n9386, n353 );
nand U10985 ( n2906, n9392, n359 );
nand U10986 ( n4739, n6515, n4743 );
nand U10987 ( n6780, n8144, n4769 );
nand U10988 ( n2713, n9357, n3970 );
not U10989 ( n352, n2906 );
nor U10990 ( n3515, n332, n338 );
not U10991 ( n283, n2728 );
not U10992 ( n339, n9149 );
not U10993 ( n107, n9152 );
nand U10994 ( n8749, n9364, n9302 );
nand U10995 ( n6677, n11403, n4713 );
nand U10996 ( n2769, n9392, n9384 );
nor U10997 ( n5408, n11386, n5314 );
nand U10998 ( n5187, n8144, n907 );
buf U10999 ( n11496, n103 );
buf U11000 ( n11516, n78 );
buf U11001 ( n11475, n909 );
buf U11002 ( n11444, n11226 );
buf U11003 ( n11436, n11227 );
or U11004 ( n6496, n11406, n4715 );
buf U11005 ( n11357, n11358 );
buf U11006 ( n11356, n11358 );
not U11007 ( n11258, n11316 );
buf U11008 ( n11405, n11235 );
buf U11009 ( n11406, n11235 );
buf U11010 ( n11438, n1908 );
buf U11011 ( n11428, n11429 );
buf U11012 ( n11366, n6133 );
buf U11013 ( n11427, n11429 );
buf U11014 ( n11374, n6112 );
buf U11015 ( n11447, n11238 );
buf U11016 ( n11431, n11430 );
buf U11017 ( n11361, n11362 );
buf U11018 ( n11387, n11389 );
buf U11019 ( n11360, n11362 );
buf U11020 ( n11432, n11430 );
not U11021 ( n11415, n11416 );
not U11022 ( n11414, n11416 );
nor U11023 ( n2736, n321, n1923 );
buf U11024 ( n11420, n11242 );
buf U11025 ( n11330, n11335 );
nor U11026 ( n6789, n4056, n629 );
nor U11027 ( n5303, n998, n4640 );
nor U11028 ( n5276, n4096, n652 );
buf U11029 ( n11347, n6665 );
nor U11030 ( n7032, n4513, n993 );
nor U11031 ( n3012, n266, n2074 );
buf U11032 ( n11384, n11243 );
nor U11033 ( n3013, n313, n2058 );
buf U11034 ( n11331, n11334 );
nor U11035 ( n5247, n4211, n736 );
nor U11036 ( n3011, n312, n2069 );
nor U11037 ( n5261, n4046, n974 );
nor U11038 ( n3784, n2459, n291 );
nor U11039 ( n3735, n2409, n184 );
nor U11040 ( n3416, n2226, n197 );
nor U11041 ( n3628, n2342, n133 );
nor U11042 ( n3601, n2327, n298 );
buf U11043 ( n11329, n11335 );
buf U11044 ( n11332, n11334 );
buf U11045 ( n11317, n11314 );
buf U11046 ( n11316, n11314 );
buf U11047 ( n11396, n11390 );
buf U11048 ( n11412, n11244 );
buf U11049 ( n11378, n6106 );
nand U11050 ( n2778, n3982, n9376 );
nor U11051 ( n3166, n2719, n333 );
buf U11052 ( n11319, n11318 );
buf U11053 ( n11320, n11318 );
buf U11054 ( n11424, n11425 );
buf U11055 ( n11423, n11425 );
nand U11056 ( n6859, n6515, n6642 );
buf U11057 ( n11430, n2538 );
buf U11058 ( n11398, n4039 );
buf U11059 ( n11416, n11248 );
buf U11060 ( n11341, n11339 );
buf U11061 ( n11340, n11339 );
nor U11062 ( n2665, n11418, n4006 );
nor U11063 ( n1898, n11418, n4015 );
nor U11064 ( n4199, n6792, n11382 );
nor U11065 ( n4640, n6924, n11382 );
nor U11066 ( n1923, n11418, n4223 );
nor U11067 ( n1934, n11418, n4432 );
nor U11068 ( n4063, n6861, n11382 );
nor U11069 ( n1968, n11418, n4755 );
buf U11070 ( n11306, n10471 );
or U11071 ( n10472, n10769, n326 );
buf U11072 ( n11299, n10485 );
buf U11073 ( n11310, n10468 );
buf U11074 ( n11335, n11336 );
nor U11075 ( n1979, n11418, n5340 );
nor U11076 ( n2024, n11418, n5392 );
nor U11077 ( n2069, n11418, n5810 );
nor U11078 ( n2013, n11418, n5365 );
nand U11079 ( n9149, n9354, n9355 );
buf U11080 ( n11343, n6666 );
nor U11081 ( n2058, n11418, n5574 );
nor U11082 ( n4468, n7277, n11382 );
buf U11083 ( n11351, n6662 );
nor U11084 ( n4268, n7227, n11383 );
nor U11085 ( n2103, n11418, n6180 );
buf U11086 ( n11334, n11336 );
nand U11087 ( n2426, n10040, n10041 );
buf U11088 ( n11481, n11483 );
buf U11089 ( n11452, n11454 );
buf U11090 ( n11314, n9727 );
buf U11091 ( n11373, n6122 );
buf U11092 ( n11318, n8614 );
nand U11093 ( n6692, n8142, n6495 );
buf U11094 ( n11339, n6718 );
buf U11095 ( n11534, n11536 );
buf U11096 ( n11528, n11531 );
nand U11097 ( n9356, n10826, n10827 );
nand U11098 ( n4769, n8187, n8188 );
buf U11099 ( n11531, n11532 );
buf U11100 ( n11536, n11537 );
nor U11101 ( n7564, n7685, n509 );
nand U11102 ( n2297, n11443, n2298 );
nor U11103 ( n8755, n8756, n8734 );
nor U11104 ( n8756, n1, n8740 );
buf U11105 ( n11500, n11496 );
nand U11106 ( n9660, n249, n224 );
not U11107 ( n93, n8740 );
not U11108 ( n263, n3007 );
not U11109 ( n97, n8808 );
nand U11110 ( n2866, n244, n2892 );
nand U11111 ( n2892, n32, n252 );
nand U11112 ( n2889, n2866, n2867 );
not U11113 ( n666, n7154 );
and U11114 ( n1957, n2866, n2867 );
nor U11115 ( n3171, n30, n3132 );
nor U11116 ( n3147, n214, n3171 );
not U11117 ( n17, n2958 );
not U11118 ( n221, n3132 );
nand U11119 ( n7185, n7189, n7154 );
not U11120 ( n517, n7189 );
nor U11121 ( n7197, n7154, n516 );
not U11122 ( n89, n8999 );
buf U11123 ( n11499, n11496 );
or U11124 ( n3168, n3171, n214 );
not U11125 ( n663, n4253 );
nand U11126 ( n3210, n30, n216 );
not U11127 ( n14, n3237 );
xnor U11128 ( n6261, n679, n588 );
buf U11129 ( n11513, n11516 );
nor U11130 ( n7488, n559, n7359 );
nor U11131 ( n7521, n7685, n511 );
not U11132 ( n213, n3208 );
not U11133 ( n509, n7525 );
and U11134 ( n7527, n7505, n7488 );
not U11135 ( n11442, n11444 );
not U11136 ( n11434, n11436 );
not U11137 ( n11435, n11436 );
not U11138 ( n11443, n11444 );
nor U11139 ( n7600, n7604, n7605 );
nor U11140 ( n7604, n7575, n7610 );
nand U11141 ( n7605, n7606, n6682 );
nand U11142 ( n7610, n7611, n716 );
not U11143 ( n25, n3663 );
not U11144 ( n556, n6329 );
nor U11145 ( n3698, n171, n3699 );
nand U11146 ( n3699, n26, n331 );
xnor U11147 ( n2298, n142, n35 );
nor U11148 ( n7688, n593, n7359 );
buf U11149 ( n11498, n11496 );
buf U11150 ( n11514, n11516 );
not U11151 ( n123, n3350 );
buf U11152 ( n11511, n11517 );
buf U11153 ( n11512, n11517 );
buf U11154 ( n11515, n11516 );
nor U11155 ( n7728, n7731, n7732 );
nand U11156 ( n7732, n7733, n6682 );
nor U11157 ( n7731, n7697, n7737 );
nand U11158 ( n7733, n7734, n7735 );
and U11159 ( n7739, n7716, n7688 );
buf U11160 ( n11479, n11475 );
not U11161 ( n10, n3737 );
nor U11162 ( n7832, n549, n7359 );
not U11163 ( n9, n3827 );
and U11164 ( n7988, n7965, n7932 );
and U11165 ( n7886, n7871, n7832 );
nor U11166 ( n8016, n7359, n543 );
not U11167 ( n543, n6445 );
buf U11168 ( n11363, n6496 );
nor U11169 ( n7925, n506, n7933 );
nand U11170 ( n7933, n6682, n739 );
not U11171 ( n20, n3922 );
nor U11172 ( n8050, n7359, n597 );
buf U11173 ( n11478, n11475 );
buf U11174 ( n11477, n11475 );
nand U11175 ( n6472, n11480, n6474 );
and U11176 ( n7734, n727, n4826 );
nor U11177 ( n8090, n7359, n542 );
buf U11178 ( n11364, n6496 );
buf U11179 ( n11365, n6496 );
not U11180 ( n11355, n11356 );
buf U11181 ( n11272, n11357 );
buf U11182 ( n11270, n11357 );
buf U11183 ( n11271, n11357 );
buf U11184 ( n11502, n84 );
buf U11185 ( n11503, n84 );
buf U11186 ( n11504, n84 );
not U11187 ( n241, n10243 );
nand U11188 ( n8778, n8605, n9256 );
nand U11189 ( n9256, n8611, n8608 );
nand U11190 ( n8644, n9235, n9236 );
nand U11191 ( n9235, n9330, n9331 );
nand U11192 ( n9236, n9237, n89 );
nand U11193 ( n9330, n9332, n9001 );
nand U11194 ( n9027, n9133, n9134 );
nand U11195 ( n9133, n9169, n9170 );
nand U11196 ( n9134, n9135, n97 );
nand U11197 ( n9169, n9171, n8810 );
not U11198 ( n1, n8853 );
nand U11199 ( n8911, n8872, n8874 );
nor U11200 ( n9135, n8715, n8983 );
nand U11201 ( n8611, n8607, n9257 );
nand U11202 ( n9257, n8609, n9094 );
nand U11203 ( n8726, n8744, n106 );
not U11204 ( n106, n8729 );
nor U11205 ( n8744, n8754, n8732 );
nor U11206 ( n8754, n8730, n8755 );
and U11207 ( n9237, n9010, n9009 );
nand U11208 ( n8727, n8728, n8729 );
nor U11209 ( n8728, n8730, n8731 );
nor U11210 ( n8731, n8732, n8629 );
or U11211 ( n8629, n8733, n8734 );
or U11212 ( n8733, n8735, n8736 );
nor U11213 ( n8736, n104, n8737 );
nor U11214 ( n8735, n8740, n8741 );
or U11215 ( n4872, n11181, n4844 );
nand U11216 ( n11181, n4835, n4853 );
not U11217 ( n238, n2684 );
nor U11218 ( n2715, n2716, n2717 );
nand U11219 ( n2717, n333, n232 );
not U11220 ( n232, n2712 );
not U11221 ( n574, n6788 );
not U11222 ( n589, n7545 );
not U11223 ( n588, n7360 );
nor U11224 ( n7640, n5250, n591 );
not U11225 ( n591, n7742 );
nand U11226 ( n6832, n6833, n6834 );
nand U11227 ( n6833, n522, n902 );
nand U11228 ( n6834, n6835, n628 );
nand U11229 ( n6835, n573, n6836 );
not U11230 ( n573, n6838 );
nor U11231 ( n9107, n8853, n9110 );
nand U11232 ( n9110, n9109, n94 );
nor U11233 ( n4770, n4800, n4801 );
nand U11234 ( n4800, n4817, n4818 );
nand U11235 ( n4801, n4802, n4803 );
nor U11236 ( n4817, n4824, n4825 );
nor U11237 ( n2710, n238, n2690 );
nor U11238 ( n2737, n19, n2741 );
nand U11239 ( n2741, n231, n238 );
nand U11240 ( n2730, n336, n2703 );
not U11241 ( n576, n6715 );
nand U11242 ( n8847, n8852, n8853 );
nand U11243 ( n8852, n94, n8854 );
nand U11244 ( n9669, n2761, n2684 );
and U11245 ( n6843, n6845, n6846 );
not U11246 ( n50, n8699 );
nor U11247 ( n2738, n2739, n2740 );
nand U11248 ( n2740, n2684, n229 );
nand U11249 ( n9462, n9464, n9465 );
nor U11250 ( n9464, n9469, n9470 );
nor U11251 ( n9465, n9466, n9467 );
nor U11252 ( n9470, n9471, n9472 );
not U11253 ( n614, n6711 );
not U11254 ( n19, n2739 );
not U11255 ( n11337, n11338 );
nand U11256 ( n9472, n251, n2825 );
not U11257 ( n251, n9473 );
and U11258 ( n6766, n6764, n903 );
and U11259 ( n6762, n6764, n902 );
nor U11260 ( n6756, n6757, n6758 );
nand U11261 ( n6757, n6767, n6768 );
nand U11262 ( n6758, n6680, n6759 );
nand U11263 ( n6767, n576, n917 );
nor U11264 ( n6710, n576, n6711 );
not U11265 ( n633, n6893 );
nand U11266 ( n6163, n6882, n6883 );
nor U11267 ( n6883, n6884, n6885 );
nor U11268 ( n6882, n6909, n6910 );
nand U11269 ( n6885, n6886, n6887 );
and U11270 ( n2848, n2893, n2888 );
not U11271 ( n586, n6123 );
not U11272 ( n224, n2839 );
nand U11273 ( n9657, n9658, n9659 );
nor U11274 ( n9658, n9662, n9663 );
nor U11275 ( n9659, n9660, n9661 );
or U11276 ( n9663, n211, n3229 );
nand U11277 ( n6723, n614, n6722 );
nor U11278 ( n6697, n6680, n618 );
nand U11279 ( n8740, n8854, n9111 );
nand U11280 ( n2783, n352, n19 );
and U11281 ( n1891, n2682, n2683 );
nand U11282 ( n2683, n2684, n2685 );
nand U11283 ( n2682, n2688, n238 );
nand U11284 ( n2685, n233, n2686 );
nor U11285 ( n9556, n9466, n9469 );
nand U11286 ( n2766, n352, n2739 );
nand U11287 ( n8734, n8757, n8758 );
nand U11288 ( n8758, n8759, n93 );
not U11289 ( n35, n3617 );
not U11290 ( n34, n3487 );
nand U11291 ( n3821, n3900, n3901 );
nand U11292 ( n7646, n7690, n7691 );
nand U11293 ( n7691, n7692, n7693 );
nor U11294 ( n7690, n7694, n7695 );
nor U11295 ( n7695, n7696, n7697 );
nand U11296 ( n7525, n7568, n7569 );
nand U11297 ( n7569, n7570, n7571 );
nor U11298 ( n7568, n7572, n7573 );
nor U11299 ( n7573, n7574, n7575 );
not U11300 ( n526, n8025 );
nand U11301 ( n2958, n3004, n3005 );
nand U11302 ( n3004, n3008, n271 );
nand U11303 ( n3005, n263, n3006 );
nand U11304 ( n3008, n3009, n3010 );
nand U11305 ( n3526, n138, n3573 );
nand U11306 ( n3573, n3574, n136 );
nand U11307 ( n3710, n182, n3731 );
nand U11308 ( n3731, n183, n3732 );
nand U11309 ( n3192, n218, n3236 );
nand U11310 ( n3236, n3237, n212 );
nand U11311 ( n3237, n206, n3281 );
nand U11312 ( n3281, n3282, n203 );
not U11313 ( n252, n2887 );
not U11314 ( n569, n7044 );
nand U11315 ( n7073, n7074, n7075 );
nand U11316 ( n7074, n519, n902 );
nand U11317 ( n7075, n7076, n649 );
nand U11318 ( n7076, n7077, n7078 );
nand U11319 ( n3007, n9554, n276 );
nand U11320 ( n2820, n2823, n2824 );
nand U11321 ( n2824, n2825, n2826 );
nand U11322 ( n2823, n2827, n2828 );
nand U11323 ( n2826, n2793, n246 );
not U11324 ( n522, n6783 );
nor U11325 ( n1883, n1891, n11444 );
nand U11326 ( n2688, n236, n2689 );
nand U11327 ( n2689, n33, n233 );
not U11328 ( n228, n2761 );
nor U11329 ( n8807, n8808, n8809 );
nand U11330 ( n8809, n8810, n8811 );
nand U11331 ( n8811, n2, n96 );
not U11332 ( n2, n8815 );
xnor U11333 ( n1917, n228, n33 );
nor U11334 ( n8806, n8812, n8813 );
xnor U11335 ( n8812, n8817, n99 );
nand U11336 ( n8813, n8814, n96 );
nand U11337 ( n8814, n8815, n8816 );
not U11338 ( n233, n2690 );
nand U11339 ( n8808, n8816, n9170 );
nand U11340 ( n9170, n99, n105 );
not U11341 ( n105, n8817 );
not U11342 ( n587, n6722 );
not U11343 ( n32, n2882 );
not U11344 ( n612, n4806 );
nand U11345 ( n9644, n267, n274 );
nand U11346 ( n9606, n9597, n9607 );
nand U11347 ( n9607, n3384, n9608 );
nand U11348 ( n9608, n9609, n9501 );
nor U11349 ( n9609, n9610, n9611 );
nor U11350 ( n4818, n4819, n4820 );
nand U11351 ( n4819, n4823, n739 );
nand U11352 ( n4820, n4821, n4822 );
nand U11353 ( n6146, n6799, n6800 );
nand U11354 ( n6799, n6803, n6804 );
nand U11355 ( n6800, n6801, n604 );
nand U11356 ( n6804, n6745, n628 );
xnor U11357 ( n6134, n4806, n6722 );
xnor U11358 ( n1938, n2803, n224 );
not U11359 ( n18, n2793 );
nand U11360 ( n8975, n8980, n8815 );
nand U11361 ( n8980, n96, n8816 );
nand U11362 ( n7154, n7214, n7259 );
nand U11363 ( n2828, n18, n248 );
nor U11364 ( n2876, n2879, n2880 );
nor U11365 ( n2879, n2882, n2883 );
nor U11366 ( n2880, n32, n2881 );
nand U11367 ( n2883, n2884, n252 );
not U11368 ( n521, n6894 );
and U11369 ( n7940, n7943, n7944 );
not U11370 ( n604, n4822 );
nand U11371 ( n2877, n2885, n2886 );
or U11372 ( n2885, n2888, n243 );
nand U11373 ( n2886, n2887, n244 );
not U11374 ( n244, n2881 );
nand U11375 ( n9666, n171, n2884 );
nand U11376 ( n3103, n274, n3111 );
nand U11377 ( n3111, n3006, n276 );
nand U11378 ( n6887, n6888, n903 );
nand U11379 ( n6886, n6888, n902 );
nor U11380 ( n6905, n521, n6892 );
nor U11381 ( n7115, n7077, n7103 );
nand U11382 ( n9109, n9111, n8757 );
not U11383 ( n243, n2884 );
nor U11384 ( n9108, n95, n8854 );
not U11385 ( n95, n9109 );
nand U11386 ( n6158, n6876, n6877 );
nand U11387 ( n6877, n6878, n6745 );
nand U11388 ( n6876, n582, n4794 );
not U11389 ( n582, n6745 );
not U11390 ( n529, n4301 );
nor U11391 ( n4789, n4790, n4791 );
nand U11392 ( n4791, n4792, n4793 );
nand U11393 ( n4790, n632, n4794 );
nand U11394 ( n4174, n4175, n609 );
not U11395 ( n609, n4176 );
nand U11396 ( n6896, n633, n4794 );
nor U11397 ( n6904, n6894, n6896 );
not U11398 ( n249, n2926 );
and U11399 ( n3074, n274, n3111 );
nand U11400 ( n2867, n2890, n2891 );
nand U11401 ( n2891, n2882, n2888 );
nor U11402 ( n2890, n2887, n243 );
not U11403 ( n30, n3146 );
nand U11404 ( n2082, n3150, n3151 );
nor U11405 ( n3151, n3152, n3153 );
nor U11406 ( n3150, n3172, n3173 );
nor U11407 ( n3152, n3168, n3169 );
nand U11408 ( n3170, n3147, n3148 );
not U11409 ( n15, n3060 );
and U11410 ( n3122, n3124, n221 );
and U11411 ( n3124, n3125, n3126 );
nor U11412 ( n6891, n6893, n6894 );
nand U11413 ( n6964, n521, n903 );
xnor U11414 ( n1983, n2926, n32 );
and U11415 ( n2941, n2916, n336 );
nand U11416 ( n4175, n4185, n4186 );
not U11417 ( n632, n6931 );
and U11418 ( n7093, n649, n7044 );
nand U11419 ( n6951, n903, n6894 );
nand U11420 ( n3132, n3185, n222 );
not U11421 ( n151, n9519 );
not U11422 ( n94, n8759 );
nand U11423 ( n7046, n7044, n649 );
nor U11424 ( n3153, n3148, n3154 );
nor U11425 ( n3154, n3155, n3156 );
nand U11426 ( n3156, n3157, n3158 );
nand U11427 ( n3155, n3161, n3162 );
nand U11428 ( n2936, n352, n2916 );
xor U11429 ( n6170, n6931, n6880 );
not U11430 ( n104, n8739 );
nand U11431 ( n2898, n248, n246 );
not U11432 ( n257, n2997 );
nand U11433 ( n9661, n3047, n257 );
not U11434 ( n216, n3211 );
not U11435 ( n567, n7029 );
nor U11436 ( n4910, n4911, n4912 );
nor U11437 ( n4912, n4913, n4914 );
nor U11438 ( n4911, n4921, n4922 );
nor U11439 ( n4913, n4915, n4916 );
nand U11440 ( n6213, n7101, n7102 );
or U11441 ( n7101, n7044, n647 );
nand U11442 ( n7102, n648, n7044 );
not U11443 ( n648, n7103 );
nand U11444 ( n7223, n917, n7029 );
nor U11445 ( n2981, n2996, n2997 );
nor U11446 ( n2996, n2998, n2999 );
nand U11447 ( n2998, n3002, n3003 );
nand U11448 ( n2999, n3000, n3001 );
nand U11449 ( n3003, n17, n336 );
nand U11450 ( n7188, n7206, n7207 );
nor U11451 ( n7206, n659, n667 );
nand U11452 ( n7207, n666, n7208 );
nand U11453 ( n7189, n7202, n7203 );
nand U11454 ( n7203, n903, n7188 );
nor U11455 ( n7202, n7204, n7205 );
and U11456 ( n7204, n7188, n902 );
xor U11457 ( n6189, n637, n6933 );
nor U11458 ( n3220, n3224, n3225 );
nor U11459 ( n3225, n3226, n3212 );
nor U11460 ( n3224, n3228, n213 );
nor U11461 ( n3226, n3211, n3146 );
nor U11462 ( n8906, n8907, n8908 );
nand U11463 ( n8908, n8909, n8874 );
nand U11464 ( n8909, n3, n8873 );
not U11465 ( n3, n8872 );
not U11466 ( n516, n7208 );
and U11467 ( n8905, n8907, n11182 );
and U11468 ( n11182, n8911, n8873 );
not U11469 ( n642, n4385 );
nand U11470 ( n7000, n903, n6844 );
nand U11471 ( n3110, n3074, n352 );
nor U11472 ( n2073, n3142, n3143 );
and U11473 ( n3143, n273, n3144 );
and U11474 ( n3142, n3147, n3148 );
nand U11475 ( n3144, n3145, n3130 );
nand U11476 ( n2987, n352, n2958 );
nand U11477 ( n4253, n4635, n4261 );
nand U11478 ( n8999, n8836, n9331 );
and U11479 ( n7255, n7266, n7267 );
nand U11480 ( n7267, n7208, n7259 );
nor U11481 ( n5221, n5223, n651 );
nor U11482 ( n5223, n5225, n5226 );
not U11483 ( n651, n5224 );
nand U11484 ( n5226, n707, n697 );
not U11485 ( n519, n7023 );
nor U11486 ( n7261, n7268, n7269 );
nor U11487 ( n7268, n7255, n514 );
nor U11488 ( n7269, n7255, n513 );
not U11489 ( n514, n7192 );
nand U11490 ( n6225, n7166, n7167 );
or U11491 ( n7166, n7029, n659 );
nand U11492 ( n7167, n654, n7029 );
not U11493 ( n654, n7168 );
nand U11494 ( n7258, n7266, n7267 );
xor U11495 ( n6237, n7226, n4809 );
not U11496 ( n641, n4382 );
not U11497 ( n512, n7195 );
nand U11498 ( n3104, n31, n333 );
nand U11499 ( n7191, n7192, n7188 );
nand U11500 ( n8866, n8871, n8872 );
nand U11501 ( n8871, n8873, n8874 );
not U11502 ( n661, n4953 );
nand U11503 ( n3158, n352, n3006 );
nand U11504 ( n3162, n336, n3006 );
and U11505 ( n2092, n3206, n3207 );
nand U11506 ( n3207, n3208, n3209 );
nand U11507 ( n3206, n219, n3210 );
nand U11508 ( n3209, n3146, n222 );
nor U11509 ( n9853, n9859, n9860 );
nand U11510 ( n9860, n9861, n9862 );
nand U11511 ( n9859, n9869, n9870 );
nor U11512 ( n9861, n9863, n9864 );
nand U11513 ( n2113, n3246, n3247 );
nand U11514 ( n3246, n30, n211 );
or U11515 ( n3247, n3248, n30 );
nand U11516 ( n3145, n221, n3146 );
not U11517 ( n532, n4260 );
nor U11518 ( n7116, n7117, n4821 );
nor U11519 ( n7117, n7118, n7119 );
nand U11520 ( n7118, n7122, n7123 );
nand U11521 ( n7119, n7120, n7121 );
nand U11522 ( n7123, n518, n902 );
not U11523 ( n269, n3047 );
nand U11524 ( n9941, n156, n9942 );
not U11525 ( n156, n9943 );
nand U11526 ( n9662, n3148, n3092 );
nand U11527 ( n7697, n7693, n7736 );
nor U11528 ( n7355, n7357, n7358 );
and U11529 ( n7358, n7144, n902 );
nor U11530 ( n7357, n7359, n588 );
nor U11531 ( n7349, n679, n7350 );
nor U11532 ( n7350, n7351, n7352 );
nand U11533 ( n7352, n7353, n7354 );
nand U11534 ( n7351, n7355, n7356 );
nand U11535 ( n3257, n14, n352 );
not U11536 ( n637, n4793 );
nand U11537 ( n7575, n7609, n7571 );
nor U11538 ( n8998, n8999, n9000 );
nand U11539 ( n9000, n9001, n9002 );
nand U11540 ( n9002, n4, n88 );
not U11541 ( n4, n8835 );
nand U11542 ( n3260, n14, n336 );
nand U11543 ( n2167, n2168, n2169 );
nand U11544 ( n2169, n11522, n2171 );
nand U11545 ( n2168, n11514, n2172 );
xor U11546 ( n6249, n7276, n4799 );
xnor U11547 ( n3221, n3229, n3192 );
not U11548 ( n102, n8873 );
and U11549 ( n3447, n192, n3479 );
nand U11550 ( n3468, n192, n3479 );
not U11551 ( n644, n4792 );
not U11552 ( n199, n9742 );
and U11553 ( n7425, n7415, n903 );
not U11554 ( n202, n9548 );
nand U11555 ( n4454, n4458, n4260 );
nand U11556 ( n4458, n668, n4261 );
not U11557 ( n122, n3339 );
nor U11558 ( n4696, n722, n4478 );
nand U11559 ( n7353, n903, n7144 );
nand U11560 ( n7417, n902, n7415 );
nand U11561 ( n8829, n8834, n8835 );
nand U11562 ( n8834, n88, n8836 );
nand U11563 ( n3305, n352, n3282 );
nand U11564 ( n4633, n4076, n704 );
nor U11565 ( n9517, n157, n149 );
nand U11566 ( n9626, n9517, n183 );
nor U11567 ( n9621, n9624, n9625 );
nand U11568 ( n9625, n9626, n174 );
not U11569 ( n667, n7152 );
nand U11570 ( n3353, n29, n122 );
nand U11571 ( n3345, n3346, n3347 );
nand U11572 ( n3346, n11491, n2171 );
nand U11573 ( n3347, n2158, n11410 );
nor U11574 ( n3460, n3472, n194 );
nor U11575 ( n3472, n3473, n3474 );
nand U11576 ( n3474, n3475, n3476 );
nand U11577 ( n3473, n3477, n3478 );
not U11578 ( n262, n3092 );
buf U11579 ( n11501, n11497 );
buf U11580 ( n11497, n103 );
buf U11581 ( n11522, n76 );
buf U11582 ( n11521, n76 );
nand U11583 ( n2257, n2258, n2259 );
nand U11584 ( n2258, n11514, n2262 );
nand U11585 ( n2259, n11522, n2261 );
nand U11586 ( n2346, n2347, n2348 );
nand U11587 ( n2347, n11514, n2351 );
nand U11588 ( n2348, n11522, n2349 );
nand U11589 ( n2302, n2303, n2304 );
nand U11590 ( n2303, n11514, n2307 );
nand U11591 ( n2304, n11522, n2306 );
nand U11592 ( n2433, n2434, n2436 );
nand U11593 ( n2434, n11514, n2438 );
nand U11594 ( n2436, n11522, n2437 );
buf U11595 ( n11518, n77 );
buf U11596 ( n11519, n77 );
nand U11597 ( n2389, n2391, n2392 );
nand U11598 ( n2391, n11514, n2394 );
nand U11599 ( n2392, n11523, n2393 );
buf U11600 ( n11523, n76 );
not U11601 ( n559, n7456 );
nor U11602 ( n7486, n7487, n7488 );
nor U11603 ( n7487, n7359, n697 );
buf U11604 ( n11520, n77 );
not U11605 ( n647, n4821 );
not U11606 ( n214, n3130 );
nand U11607 ( n3475, n3447, n352 );
nand U11608 ( n2178, n11443, n2182 );
nor U11609 ( n7518, n694, n7519 );
not U11610 ( n694, n4784 );
nor U11611 ( n7519, n7520, n7521 );
nor U11612 ( n7520, n7359, n7456 );
not U11613 ( n511, n7482 );
xnor U11614 ( n3362, n3327, n3373 );
not U11615 ( n27, n3566 );
and U11616 ( n2248, n3557, n3558 );
nand U11617 ( n3557, n3563, n3531 );
nand U11618 ( n3558, n3559, n3560 );
nor U11619 ( n3563, n3564, n3565 );
not U11620 ( n273, n3148 );
nor U11621 ( n3208, n3229, n3211 );
nand U11622 ( n9488, n9489, n212 );
nand U11623 ( n9489, n9490, n9491 );
nor U11624 ( n9490, n9546, n9547 );
nor U11625 ( n9491, n9492, n9493 );
not U11626 ( n96, n8985 );
nor U11627 ( n3506, n3507, n3508 );
nand U11628 ( n3508, n3509, n3510 );
nand U11629 ( n3507, n3511, n3512 );
nand U11630 ( n3509, n352, n3385 );
nor U11631 ( n3511, n3513, n3514 );
nor U11632 ( n3513, n3515, n3487 );
and U11633 ( n3514, n3385, n336 );
not U11634 ( n534, n4281 );
nor U11635 ( n3564, n3537, n3566 );
not U11636 ( n211, n3267 );
nand U11637 ( n6322, n7555, n7556 );
nor U11638 ( n7556, n7557, n7558 );
nor U11639 ( n7555, n7561, n7562 );
nor U11640 ( n7558, n7544, n7559 );
nor U11641 ( n7561, n703, n7563 );
not U11642 ( n703, n4779 );
nor U11643 ( n7563, n7564, n7565 );
nor U11644 ( n7565, n7359, n7545 );
nor U11645 ( n7517, n4784, n7522 );
nand U11646 ( n7522, n511, n6682 );
nand U11647 ( n3453, n3454, n3455 );
nand U11648 ( n3454, n11492, n2216 );
nand U11649 ( n3455, n11411, n2208 );
nand U11650 ( n9493, n206, n218 );
buf U11651 ( n11296, n11289 );
nand U11652 ( n3545, n3546, n3547 );
nand U11653 ( n3547, n11491, n2261 );
nand U11654 ( n3546, n2248, n11410 );
nor U11655 ( n4663, n536, n4633 );
nor U11656 ( n3594, n3515, n3605 );
nor U11657 ( n3605, n3606, n3607 );
nor U11658 ( n3607, n3590, n3566 );
nor U11659 ( n3606, n27, n3589 );
not U11660 ( n722, n4526 );
nor U11661 ( n7557, n4779, n7560 );
nand U11662 ( n7560, n509, n6682 );
not U11663 ( n219, n3212 );
buf U11664 ( n11295, n11289 );
nand U11665 ( n2207, n11443, n2208 );
not U11666 ( n668, n4462 );
buf U11667 ( n11297, n11289 );
nand U11668 ( n6297, n7503, n7504 );
nand U11669 ( n7504, n7505, n7456 );
nand U11670 ( n7503, n559, n4784 );
nand U11671 ( n2542, n2543, n2544 );
nand U11672 ( n2543, n2546, n11513 );
nand U11673 ( n2544, n11442, n8 );
xor U11674 ( n3567, n3560, n3526 );
not U11675 ( n923, n4193 );
buf U11676 ( n11293, n11288 );
xnor U11677 ( n2232, n3500, n34 );
not U11678 ( n26, n3678 );
nor U11679 ( n3668, n3515, n3663 );
nand U11680 ( n3663, n3669, n3670 );
nand U11681 ( n3669, n3675, n3638 );
nand U11682 ( n3670, n3671, n3672 );
nor U11683 ( n3675, n3676, n3677 );
or U11684 ( n2272, n11183, n11184 );
nor U11685 ( n11183, n3566, n3590 );
nor U11686 ( n11184, n3589, n27 );
not U11687 ( n743, n7779 );
buf U11688 ( n11298, n4193 );
nor U11689 ( n4788, n4795, n4796 );
nand U11690 ( n4796, n729, n4797 );
nand U11691 ( n4795, n4798, n4799 );
nand U11692 ( n7606, n7607, n7608 );
and U11693 ( n7607, n698, n4778 );
nand U11694 ( n7608, n508, n7609 );
not U11695 ( n508, n7574 );
nand U11696 ( n5050, n732, n4973 );
not U11697 ( n732, n4979 );
nand U11698 ( n9682, n208, n3295 );
nand U11699 ( n9672, n9680, n9681 );
nor U11700 ( n9680, n9684, n9685 );
nor U11701 ( n9681, n9682, n9683 );
nand U11702 ( n9685, n3625, n3590 );
nand U11703 ( n7611, n7574, n698 );
nor U11704 ( n3676, n3645, n3678 );
nand U11705 ( n4969, n4970, n4971 );
nand U11706 ( n4971, n4972, n4973 );
nand U11707 ( n4970, n4982, n4983 );
nand U11708 ( n4972, n4974, n4975 );
nor U11709 ( n7635, n7685, n7644 );
xnor U11710 ( n7644, n4823, n7574 );
nand U11711 ( n3650, n3627, n3626 );
nand U11712 ( n2307, n3619, n3620 );
nor U11713 ( n3620, n3621, n3622 );
nor U11714 ( n3619, n3630, n3631 );
nor U11715 ( n3622, n3623, n3624 );
and U11716 ( n3648, n11185, n3650 );
or U11717 ( n11185, n334, n134 );
nand U11718 ( n2351, n3695, n3696 );
nor U11719 ( n3696, n3697, n3698 );
nor U11720 ( n3695, n3703, n3704 );
nor U11721 ( n3697, n3700, n3701 );
nor U11722 ( n3703, n3693, n3705 );
nor U11723 ( n3705, n3706, n3707 );
nor U11724 ( n3706, n334, n3683 );
nor U11725 ( n3707, n3515, n26 );
nand U11726 ( n6317, n7542, n7543 );
nand U11727 ( n7543, n589, n4779 );
or U11728 ( n7542, n7544, n589 );
xor U11729 ( n6329, n4778, n7567 );
nand U11730 ( n7559, n6837, n7545 );
xnor U11731 ( n3597, n3590, n3574 );
not U11732 ( n5, n9094 );
nor U11733 ( n8602, n8603, n8604 );
nand U11734 ( n8603, n8608, n8609 );
nand U11735 ( n8604, n8605, n8606 );
nand U11736 ( n8606, n5, n8607 );
nand U11737 ( n3614, n3615, n3616 );
nand U11738 ( n3615, n11492, n2306 );
nand U11739 ( n3616, n11411, n2298 );
not U11740 ( n593, n7668 );
nor U11741 ( n7686, n7687, n7688 );
nor U11742 ( n7687, n7359, n724 );
nor U11743 ( n3621, n142, n3629 );
nand U11744 ( n3629, n331, n3617 );
not U11745 ( n208, n3373 );
xnor U11746 ( n6341, n4823, n7603 );
xnor U11747 ( n2337, n26, n3693 );
nand U11748 ( n3690, n3691, n3692 );
nand U11749 ( n3692, n11492, n2349 );
nand U11750 ( n3691, n2337, n11410 );
nand U11751 ( n3623, n3600, n134 );
nand U11752 ( n9089, n9095, n9094 );
nand U11753 ( n9095, n8607, n8609 );
nor U11754 ( n7680, n7685, n7689 );
nand U11755 ( n7689, n7646, n4828 );
nor U11756 ( n3350, n3373, n3339 );
buf U11757 ( n11517, n78 );
nand U11758 ( n2373, n3725, n3726 );
nor U11759 ( n3726, n3727, n3728 );
nor U11760 ( n3725, n3739, n3740 );
nor U11761 ( n3728, n3710, n3729 );
and U11762 ( n3739, n331, n2366 );
not U11763 ( n201, n3295 );
buf U11764 ( n11294, n11289 );
nor U11765 ( n3680, n3672, n3650 );
nor U11766 ( n3763, n3515, n3758 );
buf U11767 ( n11437, n11227 );
not U11768 ( n679, n4798 );
nand U11769 ( n7737, n7738, n721 );
nand U11770 ( n7738, n7696, n727 );
nand U11771 ( n7735, n507, n7736 );
not U11772 ( n507, n7696 );
nor U11773 ( n3667, n3627, n3679 );
nand U11774 ( n3679, n3672, n3626 );
or U11775 ( n9683, n194, n3405 );
not U11776 ( n11403, n11405 );
nand U11777 ( n3755, n3756, n3757 );
nand U11778 ( n3757, n11492, n2393 );
nand U11779 ( n3756, n23, n11410 );
not U11780 ( n23, n3758 );
nor U11781 ( n7767, n7685, n7781 );
xnor U11782 ( n7781, n4797, n7696 );
nand U11783 ( n3701, n3683, n3626 );
buf U11784 ( n11292, n11288 );
nand U11785 ( n3771, n24, n152 );
nor U11786 ( n4774, n4782, n4783 );
nand U11787 ( n4783, n4784, n4785 );
nand U11788 ( n4782, n4786, n4787 );
nor U11789 ( n7698, n7359, n7663 );
buf U11790 ( n11439, n11438 );
buf U11791 ( n11440, n11438 );
not U11792 ( n194, n3456 );
buf U11793 ( n11441, n11438 );
not U11794 ( n553, n6377 );
nand U11795 ( n6365, n7714, n7715 );
nand U11796 ( n7715, n7716, n7668 );
nand U11797 ( n7714, n593, n4826 );
and U11798 ( n3803, n331, n2404 );
not U11799 ( n11402, n11405 );
not U11800 ( n11404, n11406 );
nand U11801 ( n3737, n3732, n3626 );
buf U11802 ( n11525, n75 );
buf U11803 ( n11524, n75 );
not U11804 ( n689, n4787 );
nor U11805 ( n7932, n546, n7359 );
not U11806 ( n549, n7812 );
not U11807 ( n552, n7778 );
nor U11808 ( n7830, n7831, n7832 );
nor U11809 ( n7831, n7359, n737 );
nor U11810 ( n7930, n7931, n7932 );
nor U11811 ( n7931, n7359, n748 );
nor U11812 ( n7729, n7668, n7730 );
nand U11813 ( n7730, n6837, n4826 );
buf U11814 ( n11526, n75 );
nand U11815 ( n3827, n3833, n3626 );
not U11816 ( n191, n3500 );
nand U11817 ( n9684, n3560, n191 );
buf U11818 ( n11480, n11476 );
buf U11819 ( n11476, n909 );
nor U11820 ( n3847, n3515, n3842 );
nor U11821 ( n3773, n3767, n3737 );
nand U11822 ( n3404, n122, n126 );
nor U11823 ( n3432, n334, n198 );
not U11824 ( n506, n7842 );
nor U11825 ( n3762, n3732, n3772 );
nand U11826 ( n3772, n3767, n3626 );
nor U11827 ( n7875, n7878, n7879 );
nor U11828 ( n7878, n4812, n7884 );
nand U11829 ( n7879, n7880, n6682 );
nand U11830 ( n7884, n7885, n742 );
nor U11831 ( n7824, n524, n7833 );
nand U11832 ( n7833, n6682, n729 );
nor U11833 ( n3858, n3854, n3827 );
nand U11834 ( n4777, n4778, n4779 );
nor U11835 ( n8694, n8695, n8696 );
nand U11836 ( n8696, n8697, n8698 );
nand U11837 ( n8697, n6, n8699 );
and U11838 ( n8693, n8695, n11186 );
and U11839 ( n11186, n8701, n8699 );
nand U11840 ( n3839, n3840, n3841 );
nand U11841 ( n3841, n11492, n2437 );
nand U11842 ( n3840, n22, n11410 );
not U11843 ( n22, n3842 );
nor U11844 ( n3846, n3833, n3857 );
nand U11845 ( n3857, n3854, n3626 );
nor U11846 ( n9675, n9676, n9677 );
nand U11847 ( n9676, n3730, n3672 );
nand U11848 ( n9677, n3825, n3767 );
nand U11849 ( n3851, n3852, n163 );
nor U11850 ( n3877, n334, n3883 );
xnor U11851 ( n3883, n3879, n3779 );
not U11852 ( n171, n3693 );
nand U11853 ( n4823, n7609, n698 );
not U11854 ( n698, n7570 );
or U11855 ( n7885, n7842, n7836 );
xor U11856 ( n2453, n3879, n3852 );
nand U11857 ( n6430, n7975, n7976 );
nor U11858 ( n7976, n7977, n7978 );
nor U11859 ( n7975, n7988, n7989 );
nor U11860 ( n7977, n7980, n7981 );
nand U11861 ( n4778, n7571, n716 );
not U11862 ( n716, n7572 );
nand U11863 ( n3879, n163, n166 );
not U11864 ( n163, n3809 );
nor U11865 ( n3898, n334, n3902 );
nor U11866 ( n3902, n3903, n3904 );
nor U11867 ( n3904, n3905, n3906 );
nor U11868 ( n3903, n3907, n3885 );
nor U11869 ( n7945, n7359, n7907 );
nor U11870 ( n7843, n7359, n7807 );
xor U11871 ( n6445, n4827, n552 );
not U11872 ( n159, n3907 );
nand U11873 ( n6401, n7869, n7870 );
nand U11874 ( n7870, n7871, n7812 );
nand U11875 ( n7869, n549, n4812 );
nand U11876 ( n7505, n693, n697 );
buf U11877 ( n11368, n11366 );
buf U11878 ( n11367, n11366 );
xnor U11879 ( n2469, n159, n3882 );
buf U11880 ( n11369, n11366 );
nor U11881 ( n7876, n7812, n7877 );
nand U11882 ( n7877, n4812, n6837 );
not U11883 ( n88, n9006 );
not U11884 ( n21, n3900 );
nand U11885 ( n3922, n3939, n3940 );
or U11886 ( n3939, n3931, n21 );
nand U11887 ( n3940, n21, n3933 );
buf U11888 ( n11290, n11288 );
nand U11889 ( n4824, n4828, n4829 );
nand U11890 ( n3892, n3893, n3894 );
nand U11891 ( n3894, n11492, n2481 );
nand U11892 ( n3893, n11411, n2469 );
not U11893 ( n739, n7910 );
nand U11894 ( n3906, n3907, n48 );
xor U11895 ( n8023, n4827, n7985 );
not U11896 ( n597, n6457 );
not U11897 ( n729, n7810 );
nand U11898 ( n4826, n7693, n721 );
nand U11899 ( n4825, n4826, n4827 );
not U11900 ( n721, n7694 );
not U11901 ( n147, n3825 );
nand U11902 ( n4797, n7736, n727 );
not U11903 ( n727, n7692 );
not U11904 ( n152, n3743 );
not U11905 ( n709, n4828 );
nand U11906 ( n3624, n3625, n3626 );
not U11907 ( n142, n3625 );
nand U11908 ( n3729, n3730, n3626 );
xnor U11909 ( n8057, n4829, n526 );
and U11910 ( n3958, n331, n2511 );
not U11911 ( n754, n4829 );
not U11912 ( n542, n6469 );
nand U11913 ( n6474, n8081, n8082 );
nor U11914 ( n8082, n8083, n8084 );
nor U11915 ( n8081, n8090, n8091 );
nor U11916 ( n8083, n7785, n8085 );
xor U11917 ( n8085, n4785, n8060 );
nor U11918 ( n8084, n7786, n8085 );
and U11919 ( n2546, n3971, n8 );
nand U11920 ( n3971, n334, n3515 );
nor U11921 ( n8123, n7359, n541 );
nand U11922 ( n7871, n737, n733 );
buf U11923 ( n11291, n11288 );
not U11924 ( n936, n5419 );
nand U11925 ( n7716, n719, n724 );
not U11926 ( n934, n5418 );
nand U11927 ( n7965, n746, n748 );
buf U11928 ( n11375, n11374 );
buf U11929 ( n11376, n11374 );
buf U11930 ( n11377, n11374 );
not U11931 ( n11445, n11447 );
not U11932 ( n11426, n11427 );
not U11933 ( n11386, n11387 );
nand U11934 ( n10802, n81, n71 );
not U11935 ( n11446, n11447 );
not U11936 ( n906, n4440 );
buf U11937 ( n11281, n11428 );
buf U11938 ( n11280, n11428 );
buf U11939 ( n11279, n11428 );
buf U11940 ( n11509, n82 );
buf U11941 ( n11508, n82 );
buf U11942 ( n11510, n82 );
not U11943 ( n11359, n11360 );
buf U11944 ( n11506, n83 );
buf U11945 ( n11505, n83 );
buf U11946 ( n11507, n83 );
buf U11947 ( n11473, n912 );
buf U11948 ( n11472, n912 );
buf U11949 ( n11275, n11361 );
buf U11950 ( n11274, n11361 );
buf U11951 ( n11273, n11361 );
buf U11952 ( n11474, n912 );
not U11953 ( n334, n3626 );
buf U11954 ( n11464, n922 );
buf U11955 ( n11465, n922 );
buf U11956 ( n11469, n916 );
buf U11957 ( n11470, n916 );
buf U11958 ( n11471, n916 );
not U11959 ( n84, n3987 );
nand U11960 ( n6682, n7785, n7786 );
nor U11961 ( n7785, n902, n903 );
not U11962 ( n331, n3515 );
buf U11963 ( n11461, n941 );
buf U11964 ( n11491, n346 );
buf U11965 ( n11462, n941 );
buf U11966 ( n11450, n1022 );
buf U11967 ( n11463, n941 );
buf U11968 ( n11449, n1022 );
buf U11969 ( n11451, n1022 );
and U11970 ( n7685, n7785, n7786 );
buf U11971 ( n11492, n346 );
buf U11972 ( n11466, n919 );
buf U11973 ( n11468, n919 );
buf U11974 ( n11490, n419 );
buf U11975 ( n11467, n919 );
not U11976 ( n911, n4712 );
buf U11977 ( n11489, n419 );
buf U11978 ( n11488, n419 );
nand U11979 ( n10189, n10205, n117 );
nor U11980 ( n10205, n10207, n10208 );
not U11981 ( n117, n10206 );
nor U11982 ( n10207, n10211, n10212 );
nand U11983 ( n10206, n10246, n10247 );
nor U11984 ( n10247, n241, n10248 );
nor U11985 ( n10246, n10259, n10236 );
nor U11986 ( n10248, n10249, n10250 );
nand U11987 ( n9648, n9687, n9688 );
nor U11988 ( n9687, n10233, n10234 );
nor U11989 ( n9688, n9689, n9690 );
nor U11990 ( n10234, n10235, n10236 );
nor U11991 ( n9695, n10189, n10190 );
nand U11992 ( n10190, n10191, n10192 );
or U11993 ( n10192, n10181, n10180 );
nand U11994 ( n10191, n10202, n10203 );
not U11995 ( n11325, n11330 );
nor U11996 ( n9689, n10204, n10189 );
nor U11997 ( n10204, n10213, n10214 );
nor U11998 ( n10214, n10202, n10203 );
and U11999 ( n10213, n10212, n10211 );
not U12000 ( n11326, n11330 );
nand U12001 ( n10243, n10239, n10240 );
nand U12002 ( n8743, n9123, n9124 );
nand U12003 ( n9123, n8656, n8658 );
nand U12004 ( n9124, n9125, n8659 );
or U12005 ( n9125, n8658, n8656 );
nand U12006 ( n8938, n9271, n9272 );
nand U12007 ( n9272, n50, n8702 );
nor U12008 ( n9271, n9273, n9274 );
nor U12009 ( n9274, n92, n9275 );
nand U12010 ( n8952, n9251, n9252 );
nand U12011 ( n9251, n8776, n8778 );
nand U12012 ( n9252, n9253, n8779 );
or U12013 ( n9253, n8778, n8776 );
nand U12014 ( n9077, n9141, n9142 );
nand U12015 ( n9142, n102, n8912 );
nor U12016 ( n9141, n9143, n9144 );
nor U12017 ( n9144, n101, n9145 );
nand U12018 ( n8893, n9263, n9264 );
nand U12019 ( n9263, n8938, n8937 );
nand U12020 ( n9264, n8935, n9265 );
or U12021 ( n9265, n8937, n8938 );
nand U12022 ( n8681, n9243, n9244 );
nand U12023 ( n9243, n8952, n8951 );
nand U12024 ( n9244, n8949, n9245 );
or U12025 ( n9245, n8951, n8952 );
nand U12026 ( n8872, n9155, n9156 );
nand U12027 ( n9155, n9160, n9159 );
nand U12028 ( n9156, n9157, n9158 );
or U12029 ( n9157, n9159, n9160 );
nand U12030 ( n8701, n9064, n8698 );
nor U12031 ( n9273, n9277, n8701 );
nor U12032 ( n9277, n8702, n9276 );
nor U12033 ( n9143, n9147, n8911 );
nor U12034 ( n9147, n8912, n9146 );
nand U12035 ( n9094, n9258, n9259 );
nand U12036 ( n9258, n8891, n8893 );
nand U12037 ( n9259, n9260, n8894 );
or U12038 ( n9260, n8893, n8891 );
not U12039 ( n11419, n11420 );
nand U12040 ( n8853, n9118, n9119 );
nand U12041 ( n9118, n8739, n8743 );
nand U12042 ( n9119, n9120, n8738 );
or U12043 ( n9120, n8743, n8739 );
nand U12044 ( n8658, n9128, n9129 );
nand U12045 ( n9128, n9025, n9027 );
nand U12046 ( n9129, n9130, n9028 );
or U12047 ( n9130, n9027, n9025 );
nand U12048 ( n9010, n9238, n9239 );
nand U12049 ( n9238, n8679, n8681 );
nand U12050 ( n9239, n9240, n8682 );
or U12051 ( n9240, n8681, n8679 );
nand U12052 ( n9158, n9230, n9231 );
nand U12053 ( n9230, n8642, n8644 );
nand U12054 ( n9231, n9232, n8645 );
or U12055 ( n9232, n8644, n8642 );
and U12056 ( n8715, n9136, n9137 );
nand U12057 ( n9136, n9075, n9077 );
nand U12058 ( n9137, n9138, n9078 );
or U12059 ( n9138, n9077, n9075 );
nor U12060 ( n10233, n10245, n10206 );
nor U12061 ( n10245, n10303, n10304 );
and U12062 ( n10303, n10210, n10209 );
and U12063 ( n10304, n10250, n10249 );
nor U12064 ( n5203, n624, n1004 );
nor U12065 ( n5196, n5308, n5203 );
nor U12066 ( n5308, n626, n5202 );
nand U12067 ( n5188, n5189, n5190 );
nor U12068 ( n5190, n5191, n5192 );
nor U12069 ( n5189, n5206, n5207 );
nand U12070 ( n5192, n5193, n5194 );
and U12071 ( n5205, n5197, n5304 );
nor U12072 ( n5304, n5305, n5306 );
nor U12073 ( n5186, n5187, n5188 );
nand U12074 ( n5207, n5208, n5209 );
nand U12075 ( n5208, n5303, n5205 );
nand U12076 ( n5209, n5210, n5211 );
nor U12077 ( n5211, n5212, n5213 );
and U12078 ( n5210, n5302, n5205 );
and U12079 ( n5185, n5188, n926 );
nand U12080 ( n8741, n8742, n8743 );
or U12081 ( n8742, n8738, n8739 );
nor U12082 ( n9571, n9572, n9573 );
nor U12083 ( n9573, n9574, n242 );
nor U12084 ( n9572, n9575, n9576 );
nand U12085 ( n9576, n9577, n9578 );
nand U12086 ( n9577, n9581, n9582 );
nor U12087 ( n9581, n2735, n9583 );
nor U12088 ( n9582, n9580, n9552 );
nor U12089 ( n9583, n2736, n9584 );
xor U12090 ( n8627, n8628, n8629 );
nand U12091 ( n9653, n9654, n9655 );
nor U12092 ( n9654, n9672, n9673 );
nor U12093 ( n9655, n9656, n9657 );
nand U12094 ( n9673, n9674, n9675 );
nand U12095 ( n4835, n4869, n4870 );
nor U12096 ( n4833, n4867, n4868 );
nor U12097 ( n4868, n4869, n4870 );
nor U12098 ( n4867, n4871, n4872 );
nand U12099 ( n4871, n4909, n4910 );
nor U12100 ( n10235, n10237, n10238 );
nor U12101 ( n10238, n10239, n10240 );
nor U12102 ( n10237, n10241, n10242 );
nand U12103 ( n10242, n10243, n10244 );
nor U12104 ( n9105, n9112, n9113 );
nor U12105 ( n9112, n8740, n9114 );
nand U12106 ( n9114, n9115, n8757 );
nand U12107 ( n9115, n1, n94 );
nand U12108 ( n5193, n5197, n5198 );
nor U12109 ( n10259, n237, n10244 );
not U12110 ( n237, n10241 );
nand U12111 ( n4844, n4874, n4866 );
nand U12112 ( n4874, n622, n4863 );
not U12113 ( n622, n4865 );
nor U12114 ( n4842, n4843, n4844 );
nor U12115 ( n4843, n4845, n4846 );
nor U12116 ( n4845, n4861, n4862 );
nand U12117 ( n4846, n4847, n4848 );
nand U12118 ( n4834, n4835, n4836 );
nand U12119 ( n4836, n4837, n4838 );
nand U12120 ( n4838, n4839, n4840 );
nor U12121 ( n4837, n4841, n4842 );
or U12122 ( n4866, n4840, n4839 );
nor U12123 ( n2684, n9552, n9460 );
nand U12124 ( n2562, n2678, n2679 );
nor U12125 ( n2679, n2680, n2681 );
nor U12126 ( n2678, n2692, n1889 );
nor U12127 ( n2680, n2658, n1899 );
nand U12128 ( n2712, n2720, n2721 );
nand U12129 ( n2721, n2684, n2691 );
nand U12130 ( n2720, n2690, n238 );
nand U12131 ( n6788, n5298, n6922 );
nand U12132 ( n6922, n6923, n5302 );
nand U12133 ( n7009, n6982, n5300 );
or U12134 ( n7029, n5283, n11187 );
and U12135 ( n11187, n7226, n5271 );
nand U12136 ( n7545, n5232, n7566 );
nand U12137 ( n7566, n7567, n5229 );
nor U12138 ( n7360, n5289, n7380 );
nor U12139 ( n7380, n7381, n5295 );
nor U12140 ( n7778, n5255, n8017 );
and U12141 ( n8017, n8018, n5265 );
nor U12142 ( n8018, n596, n8019 );
or U12143 ( n7226, n5294, n11188 );
and U12144 ( n11188, n7276, n5292 );
nor U12145 ( n6916, n574, n6859 );
nand U12146 ( n6151, n6815, n6816 );
nor U12147 ( n6815, n6853, n6854 );
nor U12148 ( n6816, n6817, n6818 );
nor U12149 ( n6853, n998, n6677 );
nor U12150 ( n7603, n7637, n5235 );
and U12151 ( n7637, n7638, n5241 );
nor U12152 ( n7638, n7640, n7641 );
nor U12153 ( n7641, n7642, n5267 );
nor U12154 ( n7435, n7436, n7437 );
nor U12155 ( n7437, n7438, n7439 );
nor U12156 ( n7439, n5238, n589 );
nor U12157 ( n7775, n7776, n7777 );
and U12158 ( n7776, n5259, n7780 );
nor U12159 ( n7777, n7778, n7779 );
not U12160 ( n596, n8055 );
nand U12161 ( n7567, n5242, n7602 );
nand U12162 ( n7602, n7603, n699 );
not U12163 ( n699, n5231 );
nand U12164 ( n6531, n6795, n6796 );
nor U12165 ( n6796, n6797, n6798 );
nor U12166 ( n6795, n6814, n6151 );
nor U12167 ( n6797, n1001, n11363 );
nand U12168 ( n6838, n6913, n6914 );
nand U12169 ( n6914, n927, n6788 );
nor U12170 ( n6913, n6915, n6916 );
and U12171 ( n6915, n6788, n914 );
nand U12172 ( n6818, n6819, n6820 );
nand U12173 ( n6820, n6821, n4822 );
nand U12174 ( n6819, n604, n6828 );
nand U12175 ( n6821, n6822, n6823 );
nand U12176 ( n6982, n7027, n7028 );
nor U12177 ( n7027, n5275, n7030 );
nand U12178 ( n7028, n5224, n7029 );
nor U12179 ( n7030, n658, n5276 );
nand U12180 ( n6923, n5299, n6974 );
nand U12181 ( n6974, n6933, n5301 );
or U12182 ( n7276, n5296, n11189 );
and U12183 ( n11189, n588, n5293 );
not U12184 ( n11383, n11384 );
nor U12185 ( n7742, n7772, n5248 );
and U12186 ( n7772, n7773, n5268 );
nor U12187 ( n7773, n5261, n7774 );
nor U12188 ( n7774, n5247, n7775 );
nor U12189 ( n4841, n4863, n4864 );
nand U12190 ( n4864, n4865, n4866 );
nand U12191 ( n8848, n1, n8849 );
xor U12192 ( n8849, n8850, n8851 );
nor U12193 ( n4802, n4810, n4811 );
nand U12194 ( n4811, n4812, n4813 );
nand U12195 ( n4810, n4814, n4815 );
xnor U12196 ( n4814, n626, n1003 );
nand U12197 ( n2716, n2722, n2723 );
nand U12198 ( n2723, n2711, n2687 );
nand U12199 ( n2722, n33, n2710 );
nand U12200 ( n2703, n2731, n2732 );
and U12201 ( n2732, n2733, n2734 );
nor U12202 ( n2731, n2737, n2738 );
nand U12203 ( n2734, n2735, n2684 );
nand U12204 ( n2729, n337, n2703 );
nand U12205 ( n6715, n6742, n6787 );
nand U12206 ( n6787, n6744, n6788 );
nor U12207 ( n6124, n6126, n6111 );
nor U12208 ( n2711, n2691, n2684 );
nand U12209 ( n6764, n6781, n6782 );
nand U12210 ( n6782, n6783, n6784 );
nand U12211 ( n6783, n6841, n6842 );
and U12212 ( n6841, n6847, n6848 );
nand U12213 ( n6842, n6843, n6844 );
nand U12214 ( n6848, n6845, n6849 );
nor U12215 ( n6845, n6897, n627 );
not U12216 ( n627, n6908 );
nand U12217 ( n6908, n998, n629 );
nor U12218 ( n6779, n5187, n6764 );
nand U12219 ( n8699, n9063, n9062 );
nor U12220 ( n9275, n50, n8702 );
nand U12221 ( n6525, n6669, n6126 );
nor U12222 ( n6669, n6716, n6717 );
nor U12223 ( n6717, n11466, n619 );
nor U12224 ( n6716, n586, n11342 );
nand U12225 ( n6691, n6785, n6786 );
nand U12226 ( n6785, n917, n6715 );
nand U12227 ( n6786, n914, n6715 );
nor U12228 ( n6774, n6777, n6764 );
and U12229 ( n2707, n11190, n11191 );
nand U12230 ( n11190, n2687, n2711 );
nand U12231 ( n11191, n2710, n33 );
and U12232 ( n4851, n4861, n4862 );
and U12233 ( n4853, n4888, n4889 );
or U12234 ( n4889, n4860, n4859 );
nor U12235 ( n4888, n4894, n4851 );
nor U12236 ( n4894, n4850, n4852 );
nand U12237 ( n4847, n4853, n4854 );
nand U12238 ( n4854, n4855, n4856 );
nand U12239 ( n4856, n4857, n4858 );
nand U12240 ( n4855, n4859, n4860 );
nand U12241 ( n7780, n7890, n5253 );
and U12242 ( n7890, n748, n5260 );
nand U12243 ( n5260, n7891, n752 );
nor U12244 ( n7891, n971, n7892 );
nand U12245 ( n2733, n2736, n238 );
or U12246 ( n8698, n9062, n9063 );
nand U12247 ( n2839, n2796, n226 );
nor U12248 ( n2825, n2839, n2798 );
nor U12249 ( n9468, n9559, n2917 );
nand U12250 ( n9559, n229, n2825 );
not U12251 ( n226, n2794 );
or U12252 ( n9467, n9468, n2735 );
xnor U12253 ( n8923, n8743, n8738 );
nand U12254 ( n4848, n4849, n4850 );
nor U12255 ( n4849, n608, n4851 );
not U12256 ( n608, n4852 );
nand U12257 ( n7779, n7893, n7894 );
and U12258 ( n7893, n746, n5259 );
not U12259 ( n746, n7892 );
nor U12260 ( n6754, n6769, n4806 );
nor U12261 ( n6769, n6691, n6770 );
nand U12262 ( n6770, n523, n6771 );
nand U12263 ( n6771, n927, n6715 );
not U12264 ( n229, n2736 );
nand U12265 ( n6528, n6738, n6739 );
nor U12266 ( n6739, n6740, n6741 );
nor U12267 ( n6738, n6751, n6139 );
nor U12268 ( n6740, n1002, n11363 );
not U12269 ( n523, n6686 );
not U12270 ( n618, n4807 );
nand U12271 ( n6711, n6726, n6727 );
nand U12272 ( n6726, n5306, n4807 );
nand U12273 ( n6727, n5198, n618 );
nand U12274 ( n6706, n6707, n6708 );
nand U12275 ( n6707, n6709, n917 );
nand U12276 ( n6708, n6709, n914 );
nor U12277 ( n6709, n613, n6710 );
not U12278 ( n613, n6712 );
nand U12279 ( n2739, n2790, n2791 );
nand U12280 ( n2791, n2792, n2793 );
and U12281 ( n2790, n2796, n2797 );
nor U12282 ( n2792, n2794, n2795 );
nor U12283 ( n2760, n2761, n2762 );
nor U12284 ( n2762, n2763, n2764 );
nand U12285 ( n2763, n2770, n2771 );
nand U12286 ( n2764, n2765, n2766 );
nand U12287 ( n2565, n2745, n2746 );
nor U12288 ( n2746, n2747, n2748 );
nor U12289 ( n2745, n2756, n1924 );
nor U12290 ( n2747, n322, n11431 );
nand U12291 ( n2797, n2798, n226 );
nor U12292 ( n2761, n2736, n2735 );
not U12293 ( n748, n7912 );
and U12294 ( n6680, n6760, n6761 );
nor U12295 ( n6760, n6765, n6766 );
nor U12296 ( n6761, n6762, n6763 );
and U12297 ( n6765, n6764, n926 );
and U12298 ( n6763, n6764, n924 );
nor U12299 ( n9584, n2794, n9585 );
nor U12300 ( n9585, n9586, n9587 );
nor U12301 ( n9586, n9588, n9589 );
nand U12302 ( n9587, n248, n2796 );
nand U12303 ( n9471, n9474, n229 );
nand U12304 ( n9474, n9475, n3013 );
and U12305 ( n9475, n271, n2959 );
nor U12306 ( n6744, n6789, n5305 );
nand U12307 ( n6784, n999, n607 );
nand U12308 ( n6768, n576, n914 );
nand U12309 ( n6759, n576, n927 );
not U12310 ( n246, n2795 );
nand U12311 ( n9589, n2917, n246 );
nand U12312 ( n6713, n6714, n6712 );
nand U12313 ( n6714, n614, n6715 );
and U12314 ( n9469, n9560, n2795 );
nor U12315 ( n9560, n2736, n2839 );
not U12316 ( n231, n2735 );
nor U12317 ( n6893, n636, n997 );
nand U12318 ( n6849, n633, n6850 );
nand U12319 ( n6540, n6864, n6865 );
nor U12320 ( n6865, n6866, n6867 );
nor U12321 ( n6864, n6881, n6163 );
nor U12322 ( n6867, n999, n11363 );
nand U12323 ( n6910, n6911, n6912 );
nand U12324 ( n6911, n6917, n4794 );
nand U12325 ( n6912, n6878, n6838 );
nand U12326 ( n6917, n6918, n6919 );
nor U12327 ( n4803, n4804, n4805 );
nand U12328 ( n4804, n4808, n4809 );
nand U12329 ( n4805, n4806, n4807 );
nand U12330 ( n2803, n2844, n2845 );
nand U12331 ( n2845, n2846, n2847 );
and U12332 ( n2844, n2850, n2851 );
and U12333 ( n2846, n2848, n2849 );
not U12334 ( n33, n2687 );
nand U12335 ( n2893, n318, n247 );
nor U12336 ( n2779, n2780, n2781 );
nand U12337 ( n2780, n2786, n2787 );
nand U12338 ( n2781, n2782, n2783 );
nor U12339 ( n2787, n2788, n2789 );
nand U12340 ( n2851, n2848, n2852 );
nand U12341 ( n2852, n252, n2853 );
nand U12342 ( n6123, n6719, n6720 );
nand U12343 ( n6720, n6721, n618 );
nand U12344 ( n6719, n6723, n6712 );
nor U12345 ( n6721, n5306, n587 );
not U12346 ( n103, n8749 );
not U12347 ( n92, n9276 );
nor U12348 ( n9466, n226, n2736 );
nor U12349 ( n9557, n9468, n9558 );
nand U12350 ( n9558, n231, n2959 );
nor U12351 ( n2690, n234, n321 );
xnor U12352 ( n4806, n1001, n617 );
nand U12353 ( n8737, n93, n8738 );
xor U12354 ( n9116, n339, n9199 );
nor U12355 ( n9199, n9200, n9201 );
nor U12356 ( n9201, n318, n8749 );
nor U12357 ( n9200, n107, n247 );
or U12358 ( n9111, n9117, n9116 );
nor U12359 ( n2681, n1891, n11413 );
xnor U12360 ( n8657, n8658, n8659 );
nor U12361 ( n2788, n2739, n2775 );
nor U12362 ( n6858, n6789, n574 );
nor U12363 ( n6857, n6858, n6859 );
nand U12364 ( n6119, n6120, n6121 );
or U12365 ( n6120, n11381, n619 );
nand U12366 ( n6121, n11370, n6123 );
buf U12367 ( n11338, n11233 );
nand U12368 ( n3617, n3635, n3636 );
nand U12369 ( n3635, n3641, n3642 );
nand U12370 ( n3636, n3637, n3638 );
nand U12371 ( n3641, n3643, n3644 );
nand U12372 ( n3900, n3941, n3942 );
nand U12373 ( n3942, n3943, n3944 );
nand U12374 ( n3487, n3528, n3529 );
nand U12375 ( n3528, n3533, n3534 );
nand U12376 ( n3529, n3530, n3531 );
nand U12377 ( n3533, n3535, n3536 );
nor U12378 ( n3530, n3532, n35 );
nor U12379 ( n3637, n3639, n3640 );
nor U12380 ( n1862, n1863, n1864 );
nand U12381 ( n9473, n9591, n9592 );
nand U12382 ( n9592, n3014, n2959 );
and U12383 ( n9591, n2956, n2914 );
nor U12384 ( n9588, n9590, n9473 );
nor U12385 ( n9590, n9593, n9594 );
nand U12386 ( n9593, n9554, n2959 );
nand U12387 ( n9594, n9595, n9596 );
nand U12388 ( n7023, n7081, n7082 );
nand U12389 ( n7082, n7083, n7084 );
nand U12390 ( n7373, n7480, n7481 );
nand U12391 ( n7481, n7482, n7483 );
and U12392 ( n7574, n7648, n11192 );
nand U12393 ( n11192, n7646, n7647 );
nand U12394 ( n7144, n7370, n7371 );
and U12395 ( n7370, n7375, n7376 );
nand U12396 ( n7371, n7372, n7373 );
or U12397 ( n7375, n7378, n683 );
nand U12398 ( n7842, n7934, n7935 );
nand U12399 ( n7935, n7936, n7937 );
nand U12400 ( n7936, n7938, n7939 );
nand U12401 ( n7939, n7940, n7941 );
not U12402 ( n524, n7829 );
nand U12403 ( n6844, n7021, n7022 );
nand U12404 ( n7022, n7023, n7024 );
nor U12405 ( n7696, n7782, n7783 );
nor U12406 ( n7783, n524, n7784 );
nand U12407 ( n8060, n8086, n8087 );
nand U12408 ( n8087, n8088, n8089 );
nand U12409 ( n8025, n8058, n8059 );
nand U12410 ( n8059, n8060, n8061 );
nand U12411 ( n7482, n7523, n7524 );
nand U12412 ( n7524, n7525, n7526 );
nand U12413 ( n7941, n526, n7942 );
not U12414 ( n248, n2798 );
nand U12415 ( n3282, n3325, n3326 );
nand U12416 ( n3326, n3327, n3328 );
nand U12417 ( n2916, n2956, n2957 );
nand U12418 ( n2957, n2958, n2959 );
nand U12419 ( n2793, n2914, n2915 );
nand U12420 ( n2915, n2916, n2917 );
nand U12421 ( n3006, n278, n3191 );
nand U12422 ( n3191, n3192, n3193 );
or U12423 ( n3385, n3527, n11193 );
and U12424 ( n11193, n186, n3526 );
nand U12425 ( n3732, n3775, n3776 );
nand U12426 ( n3775, n3780, n3781 );
nand U12427 ( n3776, n3777, n151 );
nand U12428 ( n3780, n3782, n3783 );
nand U12429 ( n3627, n174, n3682 );
nand U12430 ( n3682, n3683, n172 );
not U12431 ( n172, n3684 );
nand U12432 ( n3683, n177, n3709 );
nand U12433 ( n3709, n3710, n178 );
not U12434 ( n178, n3711 );
nand U12435 ( n3779, n161, n3884 );
nand U12436 ( n3884, n3885, n3886 );
nand U12437 ( n3600, n3627, n129 );
not U12438 ( n129, n3628 );
or U12439 ( n3885, n11194, n3909 );
and U12440 ( n11194, n3910, n48 );
and U12441 ( n3574, n3598, n143 );
nand U12442 ( n3598, n3599, n3600 );
nor U12443 ( n3599, n3601, n3602 );
and U12444 ( n3327, n3380, n3381 );
nand U12445 ( n3380, n3382, n3383 );
and U12446 ( n3382, n3386, n3387 );
nand U12447 ( n3383, n3384, n3385 );
and U12448 ( n3777, n3778, n3779 );
not U12449 ( n348, n9394 );
nand U12450 ( n3944, n287, n168 );
nor U12451 ( n2887, n253, n317 );
nand U12452 ( n7044, n658, n7158 );
nand U12453 ( n7158, n7029, n656 );
not U12454 ( n656, n5280 );
nor U12455 ( n7127, n569, n6859 );
nand U12456 ( n6206, n7056, n7057 );
nor U12457 ( n7056, n7086, n7087 );
nor U12458 ( n7057, n7058, n7059 );
nor U12459 ( n7086, n993, n6677 );
nand U12460 ( n6549, n7036, n7037 );
nor U12461 ( n7037, n7038, n7039 );
nor U12462 ( n7036, n7055, n6206 );
nor U12463 ( n7038, n996, n11363 );
nand U12464 ( n7059, n7060, n7061 );
nand U12465 ( n7061, n7062, n4792 );
nand U12466 ( n7060, n644, n7069 );
nand U12467 ( n7062, n7063, n7064 );
and U12468 ( n7077, n7124, n7125 );
nand U12469 ( n7125, n927, n7044 );
nor U12470 ( n7124, n7126, n7127 );
and U12471 ( n7126, n7044, n914 );
nor U12472 ( n10208, n10209, n10210 );
nor U12473 ( n9554, n9476, n3012 );
nand U12474 ( n1947, n2814, n2815 );
nor U12475 ( n2814, n2829, n2830 );
nor U12476 ( n2815, n2816, n2817 );
nor U12477 ( n2829, n318, n283 );
nand U12478 ( n2817, n2818, n2819 );
nand U12479 ( n2818, n336, n2820 );
nand U12480 ( n2819, n351, n2820 );
nor U12481 ( n2827, n224, n2795 );
nand U12482 ( n2568, n2807, n2808 );
nor U12483 ( n2808, n2809, n2810 );
nor U12484 ( n2807, n2813, n1947 );
nor U12485 ( n2809, n321, n11431 );
nand U12486 ( n2816, n2821, n2822 );
nand U12487 ( n2821, n352, n2820 );
nand U12488 ( n2822, n337, n2820 );
nand U12489 ( n6919, n574, n927 );
buf U12490 ( n11264, n11331 );
nand U12491 ( n1942, n1943, n1944 );
nand U12492 ( n1944, n1946, n11522 );
nand U12493 ( n1943, n11513, n1947 );
nand U12494 ( n2888, n317, n253 );
nand U12495 ( n8815, n8981, n8982 );
nand U12496 ( n8981, n8984, n8714 );
or U12497 ( n8982, n8983, n8715 );
xnor U12498 ( n8729, n8745, n8746 );
nor U12499 ( n8746, n8747, n8748 );
xnor U12500 ( n8745, n339, n8750 );
nor U12501 ( n8748, n321, n8749 );
nor U12502 ( n1873, n1864, n1876 );
nor U12503 ( n6823, n6824, n6825 );
and U12504 ( n6825, n6783, n924 );
nor U12505 ( n6824, n522, n6777 );
nand U12506 ( n8089, n966, n601 );
nor U12507 ( n6946, n6931, n6947 );
nor U12508 ( n6947, n6948, n6949 );
nand U12509 ( n6949, n6950, n6951 );
nand U12510 ( n6948, n6954, n6955 );
nand U12511 ( n6543, n6927, n6928 );
nor U12512 ( n6928, n6929, n6930 );
nor U12513 ( n6927, n6942, n6175 );
nor U12514 ( n6929, n998, n11363 );
buf U12515 ( n11348, n11347 );
nand U12516 ( n2748, n2749, n2750 );
nand U12517 ( n2750, n1916, n11491 );
nand U12518 ( n2749, n11411, n1917 );
nor U12519 ( n6960, n6961, n6962 );
nand U12520 ( n6961, n6967, n6968 );
nand U12521 ( n6962, n6963, n6964 );
nor U12522 ( n6968, n6969, n6970 );
and U12523 ( n6967, n11195, n11196 );
nand U12524 ( n11195, n6923, n914 );
nand U12525 ( n11196, n6923, n917 );
nor U12526 ( n6840, n5187, n6783 );
nor U12527 ( n5224, n5280, n5276 );
nor U12528 ( n6817, n603, n6851 );
not U12529 ( n603, n6803 );
nand U12530 ( n6851, n914, n6852 );
nand U12531 ( n6852, n6788, n628 );
xnor U12532 ( n9026, n9027, n9028 );
xnor U12533 ( n8850, n339, n9204 );
nor U12534 ( n9204, n9205, n9206 );
nor U12535 ( n9206, n317, n8749 );
nor U12536 ( n9205, n107, n253 );
nand U12537 ( n8854, n8851, n8850 );
xor U12538 ( n8817, n339, n9177 );
nor U12539 ( n9177, n9178, n9179 );
nor U12540 ( n9179, n312, n8749 );
nor U12541 ( n9178, n107, n277 );
nor U12542 ( n9171, n8985, n9173 );
nor U12543 ( n9173, n98, n9174 );
nand U12544 ( n9174, n97, n8714 );
nand U12545 ( n6722, n6742, n6743 );
nand U12546 ( n6743, n6744, n6745 );
nor U12547 ( n2843, n2778, n2803 );
nand U12548 ( n2686, n236, n2687 );
nand U12549 ( n2830, n2831, n2832 );
nand U12550 ( n2832, n224, n2833 );
nand U12551 ( n2831, n2838, n2839 );
nand U12552 ( n2833, n2834, n2835 );
and U12553 ( n6822, n11197, n11198 );
nand U12554 ( n11197, n6783, n926 );
nand U12555 ( n11198, n6783, n903 );
nand U12556 ( n6745, n5298, n6879 );
nand U12557 ( n6879, n6880, n5302 );
nand U12558 ( n6880, n5299, n6932 );
nand U12559 ( n6932, n6933, n5301 );
and U12560 ( n6933, n6982, n5300 );
not U12561 ( n48, n9524 );
nor U12562 ( n8732, n8628, n8626 );
xnor U12563 ( n8626, n339, n8760 );
nor U12564 ( n8760, n8761, n8762 );
nor U12565 ( n8762, n319, n8749 );
nor U12566 ( n8761, n107, n227 );
nor U12567 ( n8747, n107, n234 );
nand U12568 ( n3901, n288, n49 );
not U12569 ( n271, n9476 );
nor U12570 ( n2930, n2945, n2926 );
nor U12571 ( n2945, n2946, n2947 );
nand U12572 ( n2946, n2952, n2953 );
nand U12573 ( n2947, n2948, n2949 );
nand U12574 ( n2574, n2920, n2921 );
nor U12575 ( n2921, n2922, n2923 );
nor U12576 ( n2920, n2927, n1992 );
nor U12577 ( n2922, n318, n11431 );
nand U12578 ( n2882, n2853, n2962 );
nand U12579 ( n2962, n2849, n2847 );
nand U12580 ( n8061, n968, n762 );
not U12581 ( n267, n3013 );
nor U12582 ( n9595, n9602, n9603 );
nor U12583 ( n9603, n3013, n9604 );
nor U12584 ( n9602, n9605, n9606 );
nor U12585 ( n9604, n9483, n9555 );
and U12586 ( n9597, n9642, n9643 );
nor U12587 ( n9642, n9549, n9645 );
nor U12588 ( n9643, n9494, n9644 );
nor U12589 ( n9645, n9601, n9646 );
nor U12590 ( n3009, n3013, n3014 );
nand U12591 ( n1987, n1988, n1989 );
nand U12592 ( n1989, n1991, n11522 );
nand U12593 ( n1988, n11514, n1992 );
nand U12594 ( n6846, n996, n638 );
and U12595 ( n8730, n8628, n8626 );
nor U12596 ( n1874, n1867, n242 );
nand U12597 ( n4822, n6784, n6781 );
nand U12598 ( n1903, n1913, n1914 );
nand U12599 ( n1914, n1916, n11521 );
nand U12600 ( n1913, n11443, n1917 );
nor U12601 ( n6801, n6789, n6802 );
nor U12602 ( n6802, n5303, n6745 );
nor U12603 ( n6798, n583, n11342 );
not U12604 ( n583, n6146 );
nand U12605 ( n8757, n9116, n9117 );
and U12606 ( n2834, n11199, n11200 );
nand U12607 ( n11199, n2803, n338 );
nand U12608 ( n11200, n2803, n333 );
not U12609 ( n236, n2691 );
nand U12610 ( n8976, n2, n8977 );
xor U12611 ( n8977, n8978, n8979 );
nor U12612 ( n6741, n6134, n11342 );
nand U12613 ( n3010, n3011, n264 );
not U12614 ( n264, n3012 );
nand U12615 ( n2810, n2811, n2812 );
nand U12616 ( n2811, n1946, n11491 );
nand U12617 ( n2812, n11411, n1938 );
nand U12618 ( n2571, n2856, n2857 );
nor U12619 ( n2857, n2858, n2859 );
nor U12620 ( n2856, n2868, n1969 );
nor U12621 ( n2858, n319, n11431 );
nand U12622 ( n2895, n2896, n2897 );
nand U12623 ( n2896, n2907, n2884 );
nand U12624 ( n2897, n2898, n2899 );
nand U12625 ( n2907, n2908, n2909 );
nor U12626 ( n2902, n18, n2775 );
nor U12627 ( n2905, n18, n2906 );
nand U12628 ( n7214, n991, n669 );
nand U12629 ( n7151, n7152, n7153 );
or U12630 ( n7153, n7154, n7155 );
nand U12631 ( n6892, n6845, n6847 );
nand U12632 ( n6902, n6906, n6907 );
nand U12633 ( n6906, n6897, n4794 );
or U12634 ( n6907, n633, n6892 );
nor U12635 ( n2932, n2933, n2934 );
nand U12636 ( n2933, n2939, n2940 );
nand U12637 ( n2934, n2935, n2936 );
nor U12638 ( n2940, n2941, n2942 );
nor U12639 ( n2935, n2937, n2938 );
and U12640 ( n2938, n2916, n351 );
nor U12641 ( n2937, n344, n2882 );
nand U12642 ( n6884, n6898, n6899 );
nand U12643 ( n6898, n6903, n6901 );
nand U12644 ( n6899, n6900, n6901 );
nor U12645 ( n6901, n6904, n6905 );
nand U12646 ( n2872, n2873, n2874 );
nand U12647 ( n2873, n2878, n2876 );
nand U12648 ( n2874, n2875, n2876 );
nor U12649 ( n2878, n2778, n2877 );
nor U12650 ( n6995, n637, n6996 );
nor U12651 ( n6996, n6997, n6998 );
nand U12652 ( n6998, n6999, n7000 );
nand U12653 ( n6997, n7003, n7004 );
nand U12654 ( n6546, n6978, n6979 );
nor U12655 ( n6979, n6980, n6981 );
nor U12656 ( n6978, n6991, n6194 );
nor U12657 ( n6980, n997, n11363 );
nand U12658 ( n6894, n6850, n6971 );
nand U12659 ( n6971, n6844, n6846 );
nand U12660 ( n7944, n971, n752 );
nor U12661 ( n6803, n5303, n604 );
nand U12662 ( n2881, n2848, n2850 );
nor U12663 ( n2875, n344, n2877 );
nand U12664 ( n2884, n2893, n2850 );
nand U12665 ( n7024, n994, n646 );
nand U12666 ( n5250, n7643, n719 );
not U12667 ( n719, n7642 );
nand U12668 ( n2037, n3035, n3036 );
nor U12669 ( n3035, n3067, n3068 );
nor U12670 ( n3036, n3037, n3038 );
nor U12671 ( n3067, n313, n283 );
nand U12672 ( n3060, n3097, n3098 );
nor U12673 ( n3097, n3101, n3102 );
nor U12674 ( n3098, n3099, n3100 );
nor U12675 ( n3102, n3074, n2906 );
nor U12676 ( n3056, n3012, n3058 );
nor U12677 ( n3058, n3059, n3060 );
nor U12678 ( n3059, n334, n267 );
nand U12679 ( n2580, n3028, n3029 );
nor U12680 ( n3029, n3030, n3031 );
nor U12681 ( n3028, n3034, n2037 );
nor U12682 ( n3030, n316, n11431 );
nand U12683 ( n3037, n3045, n3046 );
nand U12684 ( n3046, n3047, n3048 );
nand U12685 ( n3045, n3053, n269 );
nand U12686 ( n3048, n3049, n3050 );
nand U12687 ( n3053, n3054, n3055 );
nor U12688 ( n3054, n3061, n3062 );
nor U12689 ( n3055, n3056, n3057 );
nor U12690 ( n3061, n2778, n3024 );
nor U12691 ( n3099, n3074, n2775 );
nand U12692 ( n7084, n993, n652 );
xnor U12693 ( n8713, n8714, n8715 );
nor U12694 ( n6888, n6889, n6890 );
nor U12695 ( n6889, n6895, n6896 );
nor U12696 ( n6890, n6891, n6892 );
nor U12697 ( n6895, n6897, n521 );
not U12698 ( n628, n6789 );
nand U12699 ( n2032, n2033, n2034 );
nand U12700 ( n2034, n2036, n11522 );
nand U12701 ( n2033, n11514, n2037 );
xor U12702 ( n4170, n4180, n617 );
xnor U12703 ( n4180, n1001, n923 );
nand U12704 ( n4168, n4169, n616 );
nor U12705 ( n4169, n4171, n4172 );
not U12706 ( n616, n4170 );
nor U12707 ( n4172, n4173, n4174 );
nand U12708 ( n7943, n969, n756 );
nor U12709 ( n7010, n7011, n7012 );
nand U12710 ( n7012, n7013, n7014 );
nand U12711 ( n7011, n7017, n7018 );
or U12712 ( n7014, n6844, n5187 );
nand U12713 ( n6218, n7113, n7114 );
nor U12714 ( n7113, n7128, n7129 );
nor U12715 ( n7114, n7115, n7116 );
nor U12716 ( n7129, n992, n6677 );
nand U12717 ( n6552, n7097, n7098 );
nor U12718 ( n7098, n7099, n7100 );
nor U12719 ( n7097, n7112, n6218 );
nor U12720 ( n7099, n994, n11363 );
nand U12721 ( n5213, n5214, n628 );
nand U12722 ( n5214, n5215, n5216 );
nor U12723 ( n5215, n5274, n5275 );
nor U12724 ( n5216, n5217, n5218 );
nand U12725 ( n2849, n316, n259 );
nand U12726 ( n9596, n9597, n9598 );
nand U12727 ( n9598, n9599, n202 );
and U12728 ( n9599, n3381, n212 );
nor U12729 ( n2692, n239, n11415 );
nand U12730 ( n7152, n7214, n7215 );
nand U12731 ( n7215, n7216, n7217 );
nand U12732 ( n4167, n4179, n4170 );
nor U12733 ( n4179, n4176, n4181 );
nor U12734 ( n4181, n4055, n4171 );
nor U12735 ( n7128, n647, n7130 );
nor U12736 ( n7130, n7131, n7132 );
nand U12737 ( n7132, n7133, n7134 );
nand U12738 ( n7131, n7137, n7138 );
nor U12739 ( n8759, n8850, n8851 );
nor U12740 ( n6866, n581, n11342 );
not U12741 ( n581, n6158 );
nor U12742 ( n3809, n291, n164 );
not U12743 ( n536, n4077 );
nand U12744 ( n4210, n4672, n4029 );
nor U12745 ( n4672, n4673, n4674 );
nor U12746 ( n4674, n4675, n4031 );
nor U12747 ( n4673, n4676, n4027 );
nand U12748 ( n4403, n4682, n4683 );
nand U12749 ( n4683, n761, n4135 );
nor U12750 ( n4682, n4684, n4685 );
nor U12751 ( n4685, n969, n4686 );
nand U12752 ( n4557, n4618, n4619 );
nand U12753 ( n4619, n687, n4365 );
nor U12754 ( n4618, n4620, n4621 );
nor U12755 ( n4621, n987, n4622 );
nand U12756 ( n4134, n4543, n4131 );
nand U12757 ( n4364, n4324, n4326 );
nand U12758 ( n4301, n641, n4605 );
nand U12759 ( n4605, n4187, n4385 );
nor U12760 ( n4614, n4152, n4461 );
and U12761 ( n4506, n4612, n4613 );
nand U12762 ( n4612, n4634, n4635 );
nand U12763 ( n4613, n4614, n663 );
nand U12764 ( n4634, n4636, n4255 );
nand U12765 ( n4626, n4629, n4630 );
nand U12766 ( n4630, n4631, n704 );
or U12767 ( n4629, n4633, n536 );
nand U12768 ( n4631, n4074, n4632 );
and U12769 ( n4603, n4302, n529 );
or U12770 ( n4236, n4446, n11297 );
nand U12771 ( n4191, n4598, n634 );
nand U12772 ( n4178, n4187, n4188 );
nand U12773 ( n4188, n4189, n4190 );
or U12774 ( n4189, n4192, n642 );
or U12775 ( n4190, n4191, n642 );
and U12776 ( n4055, n4184, n4175 );
and U12777 ( n4184, n4178, n4177 );
xor U12778 ( n4304, n636, n923 );
not U12779 ( n634, n4599 );
or U12780 ( n8609, n9092, n9093 );
nand U12781 ( n4794, n6908, n6847 );
nor U12782 ( n4771, n4772, n4773 );
nand U12783 ( n4773, n4774, n4775 );
nand U12784 ( n4772, n4788, n4789 );
nor U12785 ( n4775, n4776, n4777 );
not U12786 ( n658, n5279 );
nor U12787 ( n4176, n4183, n999 );
nand U12788 ( n8816, n8979, n8978 );
xnor U12789 ( n8978, n339, n9187 );
nor U12790 ( n9187, n9188, n9189 );
nor U12791 ( n9189, n311, n8749 );
nor U12792 ( n9188, n107, n279 );
nand U12793 ( n2926, n2917, n2914 );
not U12794 ( n274, n3011 );
not U12795 ( n161, n9542 );
not U12796 ( n166, n3853 );
nand U12797 ( n6836, n5303, n6837 );
not U12798 ( n611, n4183 );
nand U12799 ( n2859, n2860, n2861 );
nand U12800 ( n2861, n1961, n11491 );
nand U12801 ( n2860, n1957, n11410 );
nor U12802 ( n7090, n7091, n6859 );
nor U12803 ( n7091, n5276, n569 );
not U12804 ( n99, n9172 );
nor U12805 ( n2982, n257, n2983 );
nor U12806 ( n2983, n2984, n2985 );
nand U12807 ( n2984, n2990, n2991 );
nand U12808 ( n2985, n2986, n2987 );
nand U12809 ( n2577, n2965, n2966 );
nor U12810 ( n2966, n2967, n2968 );
nor U12811 ( n2965, n2978, n2014 );
nor U12812 ( n2967, n317, n11432 );
nand U12813 ( n2014, n2979, n2980 );
nor U12814 ( n2979, n3015, n3016 );
nor U12815 ( n2980, n2981, n2982 );
nor U12816 ( n3016, n314, n283 );
nand U12817 ( n3146, n3133, n3278 );
nand U12818 ( n3278, n3126, n3123 );
nor U12819 ( n3172, n3174, n273 );
nor U12820 ( n3174, n3175, n3176 );
nand U12821 ( n3175, n3181, n3182 );
nand U12822 ( n3176, n3177, n3178 );
nor U12823 ( n3091, n3092, n3093 );
nor U12824 ( n3093, n3094, n3095 );
nand U12825 ( n3094, n3104, n3105 );
nand U12826 ( n3095, n15, n3096 );
nand U12827 ( n2586, n3136, n3137 );
nor U12828 ( n3137, n3138, n3139 );
nor U12829 ( n3136, n3149, n2082 );
nor U12830 ( n3138, n313, n11431 );
nand U12831 ( n2583, n3077, n3078 );
nor U12832 ( n3078, n3079, n3080 );
nor U12833 ( n3077, n3087, n2059 );
nor U12834 ( n3079, n314, n11431 );
nand U12835 ( n3125, n312, n277 );
nand U12836 ( n4238, n4446, n11298 );
nand U12837 ( n2077, n2078, n2079 );
nand U12838 ( n2079, n2081, n11521 );
nand U12839 ( n2078, n11514, n2082 );
xnor U12840 ( n4054, n4055, n999 );
nor U12841 ( n6969, n6777, n6894 );
nor U12842 ( n7043, n7032, n7044 );
nor U12843 ( n7039, n572, n11341 );
not U12844 ( n572, n6201 );
nand U12845 ( n6201, n7040, n7041 );
nand U12846 ( n7040, n7045, n7046 );
nand U12847 ( n7041, n7042, n644 );
nor U12848 ( n7042, n5276, n7043 );
xor U12849 ( n8739, n339, n9196 );
nor U12850 ( n9196, n9197, n9198 );
nor U12851 ( n9198, n316, n8749 );
nor U12852 ( n9197, n107, n259 );
nand U12853 ( n8607, n9093, n9092 );
not U12854 ( n724, n7667 );
nand U12855 ( n4173, n4177, n4178 );
nor U12856 ( n3782, n3785, n3786 );
and U12857 ( n2942, n2916, n337 );
nand U12858 ( n7259, n989, n674 );
nand U12859 ( n2923, n2924, n2925 );
nand U12860 ( n2924, n1991, n11491 );
nand U12861 ( n2925, n11411, n1983 );
not U12862 ( n276, n9555 );
nand U12863 ( n7937, n972, n747 );
or U12864 ( n8608, n8612, n8613 );
nand U12865 ( n3783, n3784, n3778 );
not U12866 ( n531, n4187 );
nor U12867 ( n4595, n4596, n4597 );
nand U12868 ( n4597, n4186, n4177 );
nor U12869 ( n4596, n4600, n4185 );
nor U12870 ( n4600, n642, n531 );
xor U12871 ( n8656, n339, n9193 );
nor U12872 ( n9193, n9194, n9195 );
nor U12873 ( n9195, n314, n8749 );
nor U12874 ( n9194, n107, n272 );
nor U12875 ( n7836, n973, n741 );
nand U12876 ( n4186, n4192, n4191 );
xor U12877 ( n9025, n339, n9190 );
nor U12878 ( n9190, n9191, n9192 );
nor U12879 ( n9192, n313, n8749 );
nor U12880 ( n9191, n107, n266 );
nor U12881 ( n6931, n6897, n6893 );
nand U12882 ( n8810, n8817, n9172 );
xnor U12883 ( n4239, n601, n11295 );
nand U12884 ( n3128, n3129, n3125 );
nand U12885 ( n3129, n3130, n3131 );
or U12886 ( n3131, n3132, n3133 );
nor U12887 ( n6751, n11466, n617 );
nor U12888 ( n2756, n234, n11414 );
xnor U12889 ( n9076, n9077, n9078 );
nand U12890 ( n3185, n311, n279 );
nand U12891 ( n9519, n3781, n3861 );
or U12892 ( n2949, n2916, n2906 );
nand U12893 ( n5218, n5298, n5299 );
and U12894 ( n7058, n7045, n11201 );
and U12895 ( n11201, n914, n7046 );
xnor U12896 ( n4544, n762, n11293 );
nor U12897 ( n4686, n761, n4135 );
not U12898 ( n761, n4132 );
nand U12899 ( n10160, n10166, n10170 );
nand U12900 ( n10170, n10165, n10164 );
nand U12901 ( n10166, n10180, n10181 );
nor U12902 ( n9701, n10159, n10160 );
nor U12903 ( n10159, n261, n10161 );
not U12904 ( n261, n10162 );
nand U12905 ( n9698, n9699, n9700 );
nand U12906 ( n9699, n10163, n268 );
nand U12907 ( n9700, n9701, n9702 );
not U12908 ( n268, n10164 );
nand U12909 ( n6230, n7178, n7179 );
nor U12910 ( n7178, n7218, n7219 );
nor U12911 ( n7179, n7180, n7181 );
nor U12912 ( n7219, n991, n6677 );
nand U12913 ( n6555, n7162, n7163 );
nor U12914 ( n7163, n7164, n7165 );
nor U12915 ( n7162, n7177, n6230 );
nor U12916 ( n7164, n993, n11363 );
nor U12917 ( n7180, n7198, n659 );
nor U12918 ( n7198, n7199, n7200 );
nand U12919 ( n7200, n517, n7201 );
nand U12920 ( n7199, n7209, n7210 );
nor U12921 ( n9697, n10162, n10167 );
nand U12922 ( n10167, n254, n10161 );
not U12923 ( n254, n10160 );
nor U12924 ( n3043, n3012, n3074 );
nor U12925 ( n3041, n3043, n2775 );
nor U12926 ( n3161, n3163, n3164 );
nor U12927 ( n3163, n3166, n3167 );
nor U12928 ( n3164, n214, n3165 );
nand U12929 ( n3167, n3130, n3132 );
nand U12930 ( n3068, n3069, n3070 );
nand U12931 ( n3069, n3072, n3042 );
nand U12932 ( n3070, n3071, n3042 );
nor U12933 ( n3072, n3073, n2906 );
not U12934 ( n183, n3735 );
nor U12935 ( n4380, n4383, n4384 );
nor U12936 ( n4383, n4386, n4187 );
nor U12937 ( n4384, n531, n4385 );
xnor U12938 ( n4386, n4387, n996 );
nor U12939 ( n6930, n6170, n11342 );
nor U12940 ( n9483, n3011, n3193 );
nor U12941 ( n10163, n10165, n256 );
not U12942 ( n256, n10166 );
nand U12943 ( n8605, n8613, n8612 );
nand U12944 ( n3019, n3020, n3021 );
nand U12945 ( n3020, n333, n2847 );
nand U12946 ( n3021, n338, n2847 );
nor U12947 ( n3106, n3107, n3108 );
nand U12948 ( n3107, n3114, n3115 );
nand U12949 ( n3108, n3109, n3110 );
nor U12950 ( n3114, n3118, n3119 );
nand U12951 ( n3130, n3185, n3186 );
nand U12952 ( n3186, n3187, n216 );
or U12953 ( n6878, n5303, n6789 );
nand U12954 ( n2997, n2959, n2956 );
nor U12955 ( n3211, n309, n217 );
not U12956 ( n742, n7883 );
nand U12957 ( n4298, n529, n4303 );
xnor U12958 ( n4303, n997, n4304 );
nand U12959 ( n7201, n567, n927 );
and U12960 ( n7004, n11202, n11203 );
nand U12961 ( n11202, n6844, n902 );
nand U12962 ( n11203, n6844, n924 );
nand U12963 ( n4914, n4924, n4925 );
nand U12964 ( n4925, n4917, n4918 );
nand U12965 ( n4924, n4930, n4931 );
nand U12966 ( n4922, n4923, n639 );
nor U12967 ( n4923, n4932, n4933 );
not U12968 ( n639, n4914 );
nor U12969 ( n4932, n4938, n4939 );
nand U12970 ( n4299, n4300, n4301 );
nand U12971 ( n4300, n4302, n634 );
nor U12972 ( n7100, n571, n11341 );
not U12973 ( n571, n6213 );
nand U12974 ( n7224, n914, n7029 );
nor U12975 ( n8985, n8978, n8979 );
nor U12976 ( n5212, n5297, n5218 );
and U12977 ( n5297, n5300, n5301 );
nor U12978 ( n3743, n293, n153 );
nand U12979 ( n3001, n17, n351 );
nand U12980 ( n4185, n4302, n641 );
not U12981 ( n631, n4177 );
nor U12982 ( n4909, n5175, n5176 );
nor U12983 ( n5175, n4930, n4931 );
nor U12984 ( n5176, n4857, n4858 );
or U12985 ( n7210, n7029, n6859 );
nand U12986 ( n3169, n338, n3170 );
nand U12987 ( n3002, n17, n337 );
nand U12988 ( n7208, n7155, n7321 );
nand U12989 ( n7321, n7144, n681 );
nor U12990 ( n7181, n667, n7182 );
nor U12991 ( n7182, n7183, n7184 );
nand U12992 ( n7183, n7190, n7191 );
nand U12993 ( n7184, n7185, n7186 );
and U12994 ( n7205, n7188, n924 );
nor U12995 ( n6981, n6189, n11342 );
nand U12996 ( n2104, n3214, n3215 );
nor U12997 ( n3214, n3230, n3231 );
nor U12998 ( n3215, n3216, n3217 );
nand U12999 ( n3230, n3234, n3235 );
nor U13000 ( n3228, n3227, n30 );
nand U13001 ( n2589, n3196, n3197 );
nor U13002 ( n3197, n3198, n3199 );
nor U13003 ( n3196, n3213, n2104 );
nor U13004 ( n3198, n312, n11431 );
nand U13005 ( n3217, n3218, n3219 );
nand U13006 ( n3218, n3221, n336 );
nand U13007 ( n3219, n3220, n338 );
not U13008 ( n154, n3769 );
nor U13009 ( n3638, n132, n3674 );
not U13010 ( n132, n3642 );
nand U13011 ( n3642, n298, n133 );
nor U13012 ( n3643, n3645, n3646 );
nor U13013 ( n3646, n131, n3647 );
not U13014 ( n131, n3638 );
not U13015 ( n222, n3227 );
buf U13016 ( n11494, n108 );
not U13017 ( n182, n3738 );
nor U13018 ( n3062, n344, n3024 );
nand U13019 ( n4385, n996, n4387 );
nor U13020 ( n3073, n3012, n3074 );
nand U13021 ( n2127, n3250, n3251 );
nor U13022 ( n3251, n3252, n3253 );
nor U13023 ( n3250, n3265, n3266 );
nor U13024 ( n3253, n3254, n211 );
not U13025 ( n212, n9601 );
nor U13026 ( n3265, n3267, n3268 );
nor U13027 ( n3268, n3269, n3270 );
nand U13028 ( n3269, n3276, n3277 );
nand U13029 ( n3270, n3271, n3165 );
nand U13030 ( n2592, n3240, n3241 );
nor U13031 ( n3241, n3242, n3243 );
nor U13032 ( n3240, n3249, n2127 );
nor U13033 ( n3242, n311, n11431 );
nor U13034 ( n3182, n3183, n3184 );
nor U13035 ( n3184, n3166, n3130 );
and U13036 ( n3183, n3188, n221 );
and U13037 ( n3049, n11204, n11205 );
nand U13038 ( n11204, n3024, n338 );
nand U13039 ( n11205, n3024, n333 );
or U13040 ( n3000, n2958, n2906 );
not U13041 ( n31, n3065 );
nand U13042 ( n2122, n2123, n2124 );
nand U13043 ( n2124, n11522, n2126 );
nand U13044 ( n2123, n11514, n2127 );
nor U13045 ( n3119, n31, n2778 );
nand U13046 ( n4381, n4382, n4187 );
nand U13047 ( n3139, n3140, n3141 );
nand U13048 ( n3140, n2081, n11491 );
nand U13049 ( n3141, n2073, n11410 );
not U13050 ( n278, n9549 );
nor U13051 ( n2813, n227, n11415 );
nand U13052 ( n2002, n2975, n2976 );
nand U13053 ( n2976, n2977, n2847 );
or U13054 ( n2975, n2847, n257 );
nand U13055 ( n2968, n2969, n2970 );
nand U13056 ( n2970, n2006, n11491 );
nand U13057 ( n2969, n11411, n2002 );
nand U13058 ( n4635, n992, n4637 );
nor U13059 ( n4636, n4462, n4638 );
nor U13060 ( n4638, n4253, n4459 );
nand U13061 ( n8836, n8832, n8833 );
nor U13062 ( n9332, n9006, n9333 );
nor U13063 ( n9333, n90, n9334 );
not U13064 ( n90, n9011 );
nand U13065 ( n9334, n89, n9012 );
nand U13066 ( n6242, n7243, n7244 );
nor U13067 ( n7243, n7271, n7272 );
nor U13068 ( n7244, n7245, n7246 );
nor U13069 ( n7271, n989, n6677 );
nand U13070 ( n6558, n7230, n7231 );
nor U13071 ( n7231, n7232, n7233 );
nor U13072 ( n7230, n7242, n6242 );
nor U13073 ( n7232, n992, n11363 );
nand U13074 ( n7246, n7247, n7248 );
nand U13075 ( n7247, n7260, n7217 );
nand U13076 ( n7248, n7249, n7250 );
nand U13077 ( n7260, n7261, n7262 );
nand U13078 ( n7250, n7251, n7252 );
nor U13079 ( n7251, n7256, n7257 );
nor U13080 ( n7252, n7253, n7254 );
and U13081 ( n7256, n7258, n926 );
nor U13082 ( n5217, n5219, n5220 );
nand U13083 ( n5219, n5269, n5270 );
nand U13084 ( n5220, n5221, n5222 );
and U13085 ( n5269, n5272, n5273 );
nor U13086 ( n6814, n11466, n607 );
nor U13087 ( n7257, n7255, n5187 );
nor U13088 ( n7064, n7065, n7066 );
and U13089 ( n7066, n7023, n924 );
nor U13090 ( n7065, n519, n6777 );
nor U13091 ( n7253, n7255, n6777 );
nor U13092 ( n7262, n7263, n7264 );
nor U13093 ( n7263, n7208, n7265 );
nor U13094 ( n7264, n7255, n512 );
nand U13095 ( n7265, n926, n7258 );
nand U13096 ( n4793, n6846, n6850 );
nand U13097 ( n3277, n30, n338 );
and U13098 ( n3157, n11206, n11207 );
nand U13099 ( n11206, n3006, n337 );
nand U13100 ( n11207, n3006, n351 );
nor U13101 ( n7165, n568, n11341 );
not U13102 ( n568, n6225 );
or U13103 ( n9331, n9013, n9014 );
nand U13104 ( n7272, n7273, n7274 );
nand U13105 ( n7273, n927, n6237 );
nand U13106 ( n7274, n917, n6237 );
nor U13107 ( n7296, n673, n7297 );
not U13108 ( n673, n4799 );
nor U13109 ( n7297, n7298, n7299 );
nand U13110 ( n7298, n7304, n7305 );
nand U13111 ( n6561, n7280, n7281 );
nor U13112 ( n7281, n7282, n7283 );
nor U13113 ( n7280, n7292, n6254 );
nor U13114 ( n7282, n991, n11363 );
nor U13115 ( n4382, n4387, n996 );
not U13116 ( n203, n9600 );
not U13117 ( n177, n9529 );
nor U13118 ( n7310, n7311, n7312 );
nand U13119 ( n7311, n7317, n7318 );
nand U13120 ( n7312, n7313, n7314 );
nor U13121 ( n7318, n7187, n7192 );
and U13122 ( n7313, n11208, n11209 );
nand U13123 ( n11208, n7276, n917 );
nand U13124 ( n11209, n7276, n927 );
xnor U13125 ( n4457, n923, n669 );
nand U13126 ( n4261, n991, n4457 );
nor U13127 ( n7317, n7195, n7319 );
and U13128 ( n7319, n7276, n914 );
nor U13129 ( n9547, n9600, n3325 );
nor U13130 ( n9646, n9547, n9495 );
nor U13131 ( n3531, n187, n3562 );
not U13132 ( n187, n3534 );
nand U13133 ( n3534, n302, n188 );
nor U13134 ( n3535, n3537, n3538 );
nor U13135 ( n3538, n139, n3539 );
not U13136 ( n139, n3531 );
not U13137 ( n518, n7083 );
nand U13138 ( n8867, n3, n8868 );
xor U13139 ( n8868, n8869, n8870 );
and U13140 ( n7063, n11210, n11211 );
nand U13141 ( n11210, n7023, n926 );
nand U13142 ( n11211, n7023, n903 );
nor U13143 ( n7195, n7208, n5187 );
nand U13144 ( n3105, n31, n338 );
nor U13145 ( n7080, n5187, n7023 );
or U13146 ( n3178, n3006, n2906 );
nand U13147 ( n7186, n7187, n7188 );
not U13148 ( n513, n7187 );
nor U13149 ( n7192, n7208, n6777 );
nor U13150 ( n3047, n9476, n3014 );
xor U13151 ( n9227, n9158, n9159 );
nor U13152 ( n3645, n297, n173 );
nand U13153 ( n4947, n5137, n5138 );
nand U13154 ( n5138, n672, n5139 );
not U13155 ( n672, n5140 );
nor U13156 ( n4942, n4948, n4949 );
nand U13157 ( n4948, n4954, n4955 );
nand U13158 ( n4949, n661, n4950 );
nand U13159 ( n4954, n5115, n5116 );
nand U13160 ( n5137, n4938, n4939 );
nand U13161 ( n4921, n4940, n4941 );
nor U13162 ( n4940, n5117, n5118 );
nor U13163 ( n4941, n4942, n4943 );
nor U13164 ( n5117, n5139, n5166 );
nand U13165 ( n4953, n5120, n5121 );
nor U13166 ( n5121, n5122, n5123 );
nor U13167 ( n5120, n5136, n4947 );
nor U13168 ( n5122, n5131, n5130 );
nand U13169 ( n1959, n1961, n11522 );
not U13170 ( n218, n9494 );
nor U13171 ( n4916, n4917, n4918 );
xor U13172 ( n2028, n269, n3024 );
nand U13173 ( n3031, n3032, n3033 );
nand U13174 ( n3032, n2036, n11491 );
nand U13175 ( n3033, n11411, n2028 );
not U13176 ( n136, n9545 );
and U13177 ( n3386, n198, n3389 );
xnor U13178 ( n4505, n923, n652 );
nor U13179 ( n3300, n3295, n3301 );
nor U13180 ( n3301, n3302, n3303 );
nand U13181 ( n3302, n3308, n3309 );
nand U13182 ( n3303, n3304, n3305 );
nand U13183 ( n2595, n3285, n3286 );
nor U13184 ( n3286, n3287, n3288 );
nor U13185 ( n3285, n3296, n2149 );
nor U13186 ( n3287, n309, n11431 );
nor U13187 ( n3304, n3306, n3307 );
and U13188 ( n3307, n3282, n351 );
nor U13189 ( n3306, n344, n3123 );
and U13190 ( n7305, n11212, n11213 );
nand U13191 ( n11212, n7208, n902 );
nand U13192 ( n11213, n7208, n924 );
nand U13193 ( n3199, n3200, n3201 );
nand U13194 ( n3201, n2096, n11491 );
nand U13195 ( n3200, n2092, n11410 );
not U13196 ( n174, n3702 );
nand U13197 ( n9832, n9851, n9852 );
nor U13198 ( n9851, n10070, n10071 );
nor U13199 ( n9852, n9853, n9854 );
nor U13200 ( n10071, n10072, n10073 );
nor U13201 ( n9937, n9938, n9939 );
nor U13202 ( n9939, n9940, n9941 );
nor U13203 ( n9938, n9956, n9943 );
nand U13204 ( n9940, n9944, n9945 );
nand U13205 ( n9881, n9934, n9935 );
nand U13206 ( n9934, n10034, n10035 );
nand U13207 ( n9935, n9936, n9937 );
nor U13208 ( n9936, n10032, n10033 );
nor U13209 ( n9956, n9963, n9964 );
nor U13210 ( n9963, n10002, n10003 );
nand U13211 ( n9964, n9965, n9966 );
or U13212 ( n9965, n9962, n9961 );
nor U13213 ( n9869, n9875, n9876 );
nor U13214 ( n9876, n9877, n9878 );
nor U13215 ( n9875, n9881, n9882 );
nand U13216 ( n9878, n9879, n9880 );
nand U13217 ( n9966, n9942, n9967 );
nand U13218 ( n9967, n9968, n9969 );
nand U13219 ( n9969, n9970, n9971 );
or U13220 ( n9968, n9947, n9946 );
nor U13221 ( n9942, n11214, n11215 );
and U13222 ( n11214, n10002, n10003 );
nor U13223 ( n11215, n9971, n9970 );
nor U13224 ( n9743, n9749, n9750 );
nand U13225 ( n9750, n199, n9751 );
nand U13226 ( n9749, n9783, n9784 );
nand U13227 ( n9751, n9752, n9753 );
nor U13228 ( n9702, n9703, n9704 );
nor U13229 ( n9704, n9705, n9706 );
nor U13230 ( n9703, n9707, n9708 );
and U13231 ( n9707, n9706, n9705 );
nand U13232 ( n9801, n9805, n9806 );
or U13233 ( n9806, n9804, n9803 );
nor U13234 ( n9805, n9829, n9830 );
and U13235 ( n9830, n9831, n9832 );
nand U13236 ( n9719, n9737, n9738 );
nand U13237 ( n9738, n9739, n121 );
nor U13238 ( n9737, n9743, n9744 );
not U13239 ( n121, n9740 );
nor U13240 ( n9711, n9715, n9716 );
nor U13241 ( n9716, n9717, n9718 );
nor U13242 ( n9715, n9719, n9720 );
nand U13243 ( n9720, n9721, n9722 );
nand U13244 ( n9708, n9709, n9710 );
nand U13245 ( n9709, n9717, n9718 );
nand U13246 ( n9710, n9711, n9712 );
nand U13247 ( n9712, n9713, n9714 );
nand U13248 ( n9784, n9785, n9786 );
or U13249 ( n9786, n9753, n9752 );
nand U13250 ( n9785, n9801, n9802 );
nand U13251 ( n9802, n9803, n9804 );
nand U13252 ( n3243, n3244, n3245 );
nand U13253 ( n3244, n11492, n2126 );
nand U13254 ( n3245, n11411, n2113 );
not U13255 ( n664, n4637 );
nor U13256 ( n2868, n247, n11415 );
nor U13257 ( n7233, n7270, n11341 );
not U13258 ( n98, n8984 );
nor U13259 ( n5118, n5119, n4953 );
nor U13260 ( n5119, n5135, n5145 );
nand U13261 ( n5145, n5146, n5147 );
or U13262 ( n5147, n5116, n5115 );
xnor U13263 ( n4401, n752, n11294 );
nor U13264 ( n6881, n11466, n629 );
nand U13265 ( n4260, n4459, n4460 );
or U13266 ( n4460, n4461, n4152 );
nor U13267 ( n4252, n4253, n4254 );
nand U13268 ( n4254, n4255, n4256 );
nand U13269 ( n4256, n532, n668 );
not U13270 ( n206, n9495 );
nor U13271 ( n3314, n3315, n3316 );
nand U13272 ( n3315, n3321, n3322 );
nand U13273 ( n3316, n3317, n3318 );
nor U13274 ( n3322, n3323, n3324 );
nor U13275 ( n7782, n731, n976 );
and U13276 ( n3321, n11216, n11217 );
nand U13277 ( n11216, n3123, n338 );
nand U13278 ( n11217, n3123, n333 );
nand U13279 ( n7314, n516, n926 );
not U13280 ( n196, n3416 );
and U13281 ( n3384, n3482, n196 );
and U13282 ( n7372, n691, n7374 );
nand U13283 ( n7374, n987, n683 );
nand U13284 ( n3387, n3388, n196 );
nand U13285 ( n7121, n518, n926 );
nor U13286 ( n3042, n269, n3013 );
nor U13287 ( n9006, n8833, n8832 );
nand U13288 ( n7122, n518, n924 );
nor U13289 ( n4462, n4457, n991 );
nand U13290 ( n9943, n9957, n9958 );
nand U13291 ( n9957, n9961, n9962 );
nand U13292 ( n9958, n9959, n9960 );
nor U13293 ( n3092, n3012, n3013 );
nand U13294 ( n7736, n977, n728 );
nor U13295 ( n4251, n4257, n4258 );
xnor U13296 ( n4257, n992, n664 );
nand U13297 ( n4258, n4259, n668 );
nand U13298 ( n4259, n4260, n4261 );
nand U13299 ( n7693, n978, n723 );
nor U13300 ( n4943, n4944, n4945 );
nand U13301 ( n4945, n662, n4946 );
not U13302 ( n662, n4947 );
not U13303 ( n143, n9508 );
nand U13304 ( n6564, n7333, n7334 );
nor U13305 ( n7334, n7335, n7336 );
nor U13306 ( n7333, n7345, n6266 );
nor U13307 ( n7335, n989, n11363 );
nor U13308 ( n3537, n301, n137 );
nor U13309 ( n5274, n5276, n5277 );
nor U13310 ( n5277, n5278, n5279 );
nor U13311 ( n5278, n5280, n5281 );
nor U13312 ( n5281, n5282, n5283 );
xnor U13313 ( n4504, n4506, n993 );
nand U13314 ( n3126, n308, n204 );
nand U13315 ( n3258, n14, n351 );
nor U13316 ( n3254, n3255, n3256 );
nand U13317 ( n3255, n3259, n3260 );
nand U13318 ( n3256, n3257, n3258 );
nand U13319 ( n3259, n14, n337 );
nor U13320 ( n9145, n102, n8912 );
nor U13321 ( n8983, n8714, n8984 );
xor U13322 ( n4341, n747, n923 );
nand U13323 ( n7609, n981, n702 );
nand U13324 ( n8835, n9007, n9008 );
nand U13325 ( n9007, n9011, n9012 );
nand U13326 ( n9008, n9009, n9010 );
and U13327 ( n4933, n4920, n4919 );
nand U13328 ( n2977, n2849, n2853 );
not U13329 ( n29, n3334 );
nand U13330 ( n2172, n3355, n3356 );
nor U13331 ( n3355, n3374, n3375 );
nor U13332 ( n3356, n3357, n3358 );
nand U13333 ( n3374, n3378, n3379 );
nor U13334 ( n3361, n3365, n3366 );
nor U13335 ( n3365, n3367, n123 );
nor U13336 ( n3367, n3368, n29 );
nand U13337 ( n2598, n3342, n3343 );
nor U13338 ( n3343, n3344, n3345 );
nor U13339 ( n3342, n3354, n2172 );
nor U13340 ( n3344, n308, n11432 );
nand U13341 ( n3358, n3359, n3360 );
nand U13342 ( n3359, n336, n3362 );
nand U13343 ( n3360, n3361, n338 );
xnor U13344 ( n4279, n702, n11294 );
nand U13345 ( n4478, n4699, n4283 );
and U13346 ( n4074, n4694, n4695 );
nand U13347 ( n4695, n4696, n4697 );
nand U13348 ( n4694, n4698, n4699 );
nor U13349 ( n4697, n978, n4488 );
nand U13350 ( n4698, n4700, n4480 );
nor U13351 ( n4700, n701, n4701 );
not U13352 ( n701, n4282 );
nor U13353 ( n4701, n4478, n4485 );
nand U13354 ( n4792, n7024, n7021 );
nand U13355 ( n7134, n903, n7083 );
xnor U13356 ( n4037, n736, n11292 );
nand U13357 ( n4027, n734, n4035 );
not U13358 ( n734, n4675 );
nor U13359 ( n8997, n9003, n9004 );
xor U13360 ( n9003, n9013, n9014 );
nand U13361 ( n9004, n9005, n88 );
nand U13362 ( n9005, n8835, n8836 );
not U13363 ( n138, n9509 );
nor U13364 ( n7283, n564, n11341 );
not U13365 ( n564, n6249 );
or U13366 ( n7120, n7083, n5187 );
nor U13367 ( n7361, n7362, n7363 );
nand U13368 ( n7363, n7364, n7365 );
nand U13369 ( n7362, n7366, n7367 );
or U13370 ( n7364, n7144, n5187 );
nor U13371 ( n7366, n7368, n7369 );
nor U13372 ( n7369, n6777, n7144 );
nor U13373 ( n7368, n7360, n7359 );
nor U13374 ( n3425, n29, n2778 );
nand U13375 ( n2194, n3407, n3408 );
nor U13376 ( n3407, n3440, n3441 );
nor U13377 ( n3408, n3409, n3410 );
nor U13378 ( n3440, n304, n283 );
nand U13379 ( n2601, n3392, n3393 );
nor U13380 ( n3393, n3394, n3395 );
nor U13381 ( n3392, n3406, n2194 );
nor U13382 ( n3394, n307, n11432 );
nand U13383 ( n3409, n3419, n3420 );
nand U13384 ( n3419, n3426, n3405 );
nand U13385 ( n3420, n3421, n3404 );
nand U13386 ( n3426, n3427, n3428 );
xnor U13387 ( n8643, n8644, n8645 );
nand U13388 ( n8873, n8870, n8869 );
nand U13389 ( n3235, n3221, n337 );
nor U13390 ( n4915, n4919, n4920 );
nand U13391 ( n3234, n3221, n351 );
xor U13392 ( n2052, n262, n3065 );
nand U13393 ( n3080, n3081, n3082 );
nand U13394 ( n3082, n2051, n11491 );
nand U13395 ( n3081, n11411, n2052 );
not U13396 ( n186, n9612 );
not U13397 ( n198, n3446 );
nand U13398 ( n7571, n982, n717 );
nand U13399 ( n3479, n3385, n3482 );
nor U13400 ( n3466, n3447, n2775 );
and U13401 ( n3366, n11218, n3352 );
or U13402 ( n11218, n3339, n3334 );
nor U13403 ( n3470, n3447, n2906 );
nand U13404 ( n5166, n5137, n5140 );
not U13405 ( n649, n5276 );
nor U13406 ( n7694, n723, n978 );
nor U13407 ( n7045, n644, n7032 );
and U13408 ( n3333, n126, n3335 );
nand U13409 ( n3335, n307, n209 );
xnor U13410 ( n4489, n717, n11295 );
nor U13411 ( n3323, n2775, n3282 );
or U13412 ( n8874, n8869, n8870 );
nand U13413 ( n9945, n9946, n9947 );
not U13414 ( n691, n7410 );
nand U13415 ( n7415, n7426, n7427 );
and U13416 ( n7426, n4813, n7378 );
nand U13417 ( n7427, n7373, n691 );
nand U13418 ( n6278, n7404, n7405 );
nor U13419 ( n7404, n7428, n7429 );
nor U13420 ( n7405, n7406, n7407 );
nor U13421 ( n7429, n986, n6677 );
nor U13422 ( n7406, n7373, n7418 );
nand U13423 ( n7418, n7419, n7378 );
nand U13424 ( n7419, n7420, n7421 );
nor U13425 ( n7420, n7424, n7425 );
nand U13426 ( n6567, n7391, n7392 );
nor U13427 ( n7392, n7393, n7394 );
nor U13428 ( n7391, n7403, n6278 );
nor U13429 ( n7393, n988, n11364 );
and U13430 ( n7421, n11219, n11220 );
nand U13431 ( n11219, n7415, n902 );
nand U13432 ( n11220, n7415, n924 );
nand U13433 ( n9742, n9747, n9754 );
nand U13434 ( n9754, n207, n9745 );
not U13435 ( n207, n9748 );
or U13436 ( n9747, n9724, n9723 );
nand U13437 ( n7647, n979, n712 );
nor U13438 ( n7692, n728, n977 );
xnor U13439 ( n4575, n741, n11298 );
nor U13440 ( n2927, n253, n11414 );
nand U13441 ( n9548, n203, n3328 );
nand U13442 ( n9001, n9014, n9013 );
not U13443 ( n659, n4808 );
and U13444 ( n7424, n7415, n926 );
nor U13445 ( n3339, n306, n124 );
not U13446 ( n101, n9146 );
nand U13447 ( n7354, n926, n7144 );
nor U13448 ( n3427, n3434, n3435 );
nor U13449 ( n3434, n2778, n3334 );
nor U13450 ( n3435, n344, n3334 );
or U13451 ( n9009, n9012, n9011 );
nor U13452 ( n7407, n7408, n7409 );
nor U13453 ( n7409, n7410, n4813 );
nor U13454 ( n7408, n7411, n7412 );
nand U13455 ( n7411, n7416, n7417 );
nand U13456 ( n7412, n7413, n7414 );
nand U13457 ( n7413, n903, n7415 );
nand U13458 ( n7414, n926, n7415 );
and U13459 ( n3309, n11221, n11222 );
nand U13460 ( n11221, n3282, n336 );
nand U13461 ( n11222, n3282, n337 );
xor U13462 ( n4149, n674, n923 );
nor U13463 ( n3370, n3372, n123 );
and U13464 ( n3372, n126, n3334 );
nand U13465 ( n7356, n924, n7144 );
nor U13466 ( n7570, n702, n981 );
not U13467 ( n11328, n11329 );
nand U13468 ( n8830, n4, n8831 );
xor U13469 ( n8831, n8832, n8833 );
nor U13470 ( n6942, n11466, n636 );
nand U13471 ( n7416, n924, n7415 );
nand U13472 ( n4821, n7084, n7081 );
nor U13473 ( n10032, n9959, n9960 );
nand U13474 ( n2041, n2048, n2049 );
nand U13475 ( n2049, n2051, n11522 );
nand U13476 ( n2048, n11443, n2052 );
nand U13477 ( n7526, n983, n706 );
nor U13478 ( n10033, n10034, n10035 );
nor U13479 ( n9744, n9745, n9746 );
nand U13480 ( n9746, n9747, n9748 );
or U13481 ( n3318, n3282, n2906 );
nor U13482 ( n7572, n717, n982 );
xnor U13483 ( n2142, n3123, n3295 );
nand U13484 ( n3288, n3289, n3290 );
nand U13485 ( n3290, n2141, n11491 );
nand U13486 ( n3289, n11411, n2142 );
nor U13487 ( n3148, n3011, n9555 );
xnor U13488 ( n9040, n9010, n9012 );
nor U13489 ( n9739, n9741, n9742 );
nand U13490 ( n7078, n7032, n6837 );
or U13491 ( n9721, n9714, n9713 );
not U13492 ( n126, n3368 );
nor U13493 ( n5282, n5284, n5285 );
nand U13494 ( n5285, n5222, n5286 );
nand U13495 ( n5284, n5272, n5271 );
nand U13496 ( n5286, n5287, n5288 );
nand U13497 ( n9874, n9879, n9898 );
nand U13498 ( n9898, n176, n9877 );
not U13499 ( n176, n9880 );
or U13500 ( n9882, n9874, n11223 );
and U13501 ( n11223, n9873, n9872 );
nand U13502 ( n9879, n9865, n9866 );
nor U13503 ( n4076, n4665, n4478 );
or U13504 ( n4665, n4525, n4488 );
nor U13505 ( n7336, n563, n11341 );
not U13506 ( n563, n6261 );
not U13507 ( n157, n3785 );
nor U13508 ( n9610, n9613, n9614 );
nand U13509 ( n9614, n186, n136 );
nor U13510 ( n9613, n9615, n3602 );
nor U13511 ( n9615, n9616, n9617 );
nand U13512 ( n9617, n9618, n9619 );
nand U13513 ( n9618, n3905, n9620 );
nand U13514 ( n9619, n9524, n9620 );
and U13515 ( n9620, n9621, n9622 );
nand U13516 ( n9632, n9633, n9634 );
nor U13517 ( n9633, n3684, n3711 );
nand U13518 ( n9634, n148, n9635 );
not U13519 ( n148, n9624 );
nand U13520 ( n9635, n9636, n3778 );
nand U13521 ( n9636, n9637, n9626 );
nand U13522 ( n9637, n9638, n151 );
nor U13523 ( n9638, n3735, n9639 );
nand U13524 ( n9616, n9629, n9630 );
nor U13525 ( n9629, n9508, n3628 );
nand U13526 ( n9630, n9631, n9632 );
nor U13527 ( n9631, n3601, n3702 );
nand U13528 ( n2004, n2006, n11522 );
and U13529 ( n2158, n3348, n3349 );
nand U13530 ( n3349, n3350, n3351 );
nand U13531 ( n3348, n3352, n3353 );
nand U13532 ( n3351, n3334, n126 );
nor U13533 ( n5132, n5134, n5135 );
nand U13534 ( n5135, n5156, n5157 );
nand U13535 ( n5157, n5128, n5127 );
nand U13536 ( n5156, n5131, n5130 );
nand U13537 ( n5123, n5124, n5125 );
nand U13538 ( n5125, n5126, n684 );
nand U13539 ( n5124, n5132, n692 );
not U13540 ( n684, n5127 );
xnor U13541 ( n4071, n706, n11293 );
not U13542 ( n704, n4664 );
nand U13543 ( n2604, n3450, n3451 );
nor U13544 ( n3451, n3452, n3453 );
nor U13545 ( n3450, n3457, n2217 );
nor U13546 ( n3452, n306, n11432 );
nor U13547 ( n3477, n3480, n3481 );
nor U13548 ( n3481, n2775, n3468 );
nor U13549 ( n3480, n28, n3471 );
not U13550 ( n28, n3439 );
nor U13551 ( n5288, n5294, n5296 );
and U13552 ( n5222, n5291, n5292 );
or U13553 ( n5291, n5293, n5294 );
nand U13554 ( n9624, n9640, n9641 );
nor U13555 ( n9640, n9529, n3738 );
nand U13556 ( n9641, n3786, n183 );
nand U13557 ( n2212, n2213, n2214 );
nand U13558 ( n2214, n11522, n2216 );
nand U13559 ( n2213, n11514, n2217 );
nand U13560 ( n5272, n5288, n5295 );
nor U13561 ( n9639, n3784, n3886 );
nand U13562 ( n7483, n984, n696 );
xnor U13563 ( n4322, n688, n11291 );
nor U13564 ( n4622, n687, n4365 );
not U13565 ( n687, n4325 );
nor U13566 ( n3462, n3463, n3433 );
nor U13567 ( n3463, n3471, n3439 );
nor U13568 ( n5126, n5128, n5129 );
and U13569 ( n5129, n5130, n5131 );
nor U13570 ( n5136, n677, n4946 );
not U13571 ( n677, n4944 );
buf U13572 ( n11266, n11331 );
nor U13573 ( n7103, n5276, n7032 );
not U13574 ( n149, n3781 );
nand U13575 ( n9857, n10072, n10073 );
and U13576 ( n9862, n9857, n10077 );
nand U13577 ( n10077, n141, n9855 );
not U13578 ( n141, n9858 );
xnor U13579 ( n4555, n678, n11290 );
nand U13580 ( n2182, n3402, n3403 );
nand U13581 ( n3403, n3404, n3334 );
nand U13582 ( n3402, n29, n3405 );
nand U13583 ( n3395, n3396, n3397 );
nand U13584 ( n3397, n2186, n11491 );
nand U13585 ( n3396, n11411, n2182 );
nor U13586 ( n3905, n3909, n3910 );
nor U13587 ( n10070, n9868, n10074 );
nand U13588 ( n10074, n9862, n9867 );
buf U13589 ( n11267, n11332 );
xor U13590 ( n6273, n4813, n7381 );
nor U13591 ( n7428, n7430, n6273 );
nor U13592 ( n2978, n259, n11415 );
buf U13593 ( n11268, n11332 );
xnor U13594 ( n4521, n712, n11296 );
nand U13595 ( n2131, n2138, n2139 );
nand U13596 ( n2139, n2141, n11521 );
nand U13597 ( n2138, n11443, n2142 );
nor U13598 ( n3418, n3416, n3447 );
nand U13599 ( n3441, n3442, n3443 );
nand U13600 ( n3442, n3445, n3414 );
nand U13601 ( n3443, n3444, n3414 );
nor U13602 ( n3445, n3418, n2906 );
nand U13603 ( n3410, n3411, n3412 );
nand U13604 ( n3412, n3413, n3414 );
nand U13605 ( n3411, n3417, n3414 );
nor U13606 ( n3413, n3415, n2775 );
or U13607 ( n9870, n11224, n9872 );
or U13608 ( n11224, n9873, n9874 );
xnor U13609 ( n4556, n988, n4557 );
not U13610 ( n76, n1864 );
not U13611 ( n78, n1878 );
not U13612 ( n11410, n11412 );
nor U13613 ( n6991, n11466, n638 );
nand U13614 ( n2221, n2228, n2229 );
nand U13615 ( n2228, n11443, n2232 );
nand U13616 ( n2229, n2231, n11521 );
nand U13617 ( n2311, n2318, n2319 );
nand U13618 ( n2318, n25, n11442 );
nand U13619 ( n2319, n2321, n11521 );
nand U13620 ( n2442, n2449, n2451 );
nand U13621 ( n2449, n2453, n11442 );
nand U13622 ( n2451, n2452, n11521 );
nand U13623 ( n2354, n2362, n2363 );
nand U13624 ( n2362, n11443, n2366 );
nand U13625 ( n2363, n2364, n11521 );
nand U13626 ( n2094, n2096, n11521 );
not U13627 ( n77, n1867 );
nor U13628 ( n9854, n9855, n9856 );
nand U13629 ( n9856, n9857, n9858 );
nor U13630 ( n3415, n3416, n3447 );
nor U13631 ( n9487, n3011, n9549 );
buf U13632 ( n11265, n11331 );
nor U13633 ( n7475, n7477, n4787 );
nor U13634 ( n7477, n7478, n7479 );
nor U13635 ( n7478, n7436, n7486 );
nor U13636 ( n7479, n7473, n7373 );
nand U13637 ( n6578, n7448, n7449 );
nor U13638 ( n7449, n7450, n7451 );
nor U13639 ( n7448, n7465, n6290 );
nor U13640 ( n7450, n987, n11364 );
nand U13641 ( n6290, n7466, n7467 );
nor U13642 ( n7467, n7468, n7469 );
nor U13643 ( n7466, n7475, n7476 );
nor U13644 ( n7469, n7430, n7452 );
nand U13645 ( n2518, n2519, n2521 );
nand U13646 ( n2519, n11514, n2523 );
nand U13647 ( n2521, n11523, n2522 );
nand U13648 ( n2477, n2478, n2479 );
nand U13649 ( n2478, n11515, n2482 );
nand U13650 ( n2479, n11523, n2481 );
nand U13651 ( n7456, n707, n7529 );
or U13652 ( n7529, n589, n5238 );
not U13653 ( n134, n3601 );
nor U13654 ( n9622, n3784, n9623 );
nand U13655 ( n9623, n161, n134 );
not U13656 ( n11327, n11329 );
nand U13657 ( n3229, n3193, n278 );
nand U13658 ( n3476, n3447, n351 );
nand U13659 ( n4809, n7214, n7216 );
and U13660 ( n7266, n7217, n4809 );
xnor U13661 ( n8680, n8681, n8682 );
nand U13662 ( n6581, n7499, n7500 );
nor U13663 ( n7500, n7501, n7502 );
nor U13664 ( n7499, n7514, n6302 );
nor U13665 ( n7501, n986, n11364 );
nand U13666 ( n6302, n7515, n7516 );
nor U13667 ( n7515, n7527, n7528 );
nor U13668 ( n7516, n7517, n7518 );
nor U13669 ( n7528, n983, n6677 );
nand U13670 ( n9722, n9723, n9724 );
nand U13671 ( n3478, n3447, n337 );
buf U13672 ( n11349, n11347 );
nor U13673 ( n9863, n128, n9867 );
not U13674 ( n128, n9868 );
nor U13675 ( n9864, n9865, n9866 );
nor U13676 ( n7394, n6273, n11341 );
nor U13677 ( n3504, n3516, n3500 );
nor U13678 ( n3516, n3517, n3518 );
nand U13679 ( n3518, n3519, n3520 );
nand U13680 ( n3517, n3521, n3522 );
nand U13681 ( n2607, n3490, n3491 );
nor U13682 ( n3491, n3492, n3493 );
nor U13683 ( n3490, n3501, n2239 );
nor U13684 ( n3492, n304, n11432 );
nor U13685 ( n3521, n3523, n3524 );
nor U13686 ( n3523, n34, n3515 );
nor U13687 ( n3524, n2775, n3385 );
nand U13688 ( n3379, n337, n3362 );
nand U13689 ( n3378, n351, n3362 );
nand U13690 ( n3566, n3539, n3608 );
or U13691 ( n3608, n35, n3532 );
nand U13692 ( n2262, n3549, n3550 );
nor U13693 ( n3549, n3569, n3570 );
nor U13694 ( n3550, n3551, n3552 );
nor U13695 ( n3569, n301, n283 );
nand U13696 ( n2610, n3542, n3543 );
nor U13697 ( n3543, n3544, n3545 );
nor U13698 ( n3542, n3548, n2262 );
nor U13699 ( n3544, n303, n11432 );
nand U13700 ( n3552, n3553, n3554 );
nand U13701 ( n3553, n3567, n336 );
nand U13702 ( n3554, n2248, n3555 );
nand U13703 ( n3555, n3556, n2778 );
nor U13704 ( n3559, n3537, n3561 );
nor U13705 ( n3561, n3562, n27 );
nor U13706 ( n7468, n7473, n7474 );
nand U13707 ( n7474, n7373, n4787 );
and U13708 ( n5270, n693, n5271 );
xor U13709 ( n4207, n731, n923 );
xnor U13710 ( n4628, n696, n11292 );
nand U13711 ( n3212, n221, n3187 );
nor U13712 ( n9492, n9496, n9497 );
nand U13713 ( n9496, n196, n3381 );
nand U13714 ( n9497, n202, n9498 );
nand U13715 ( n9498, n9499, n198 );
nor U13716 ( n3034, n272, n11415 );
nand U13717 ( n4281, n4485, n4486 );
nand U13718 ( n4486, n4487, n711 );
not U13719 ( n711, n4488 );
nor U13720 ( n4477, n4478, n4479 );
nand U13721 ( n4479, n4480, n4481 );
nand U13722 ( n4481, n534, n4282 );
nor U13723 ( n3267, n9601, n9494 );
nor U13724 ( n7168, n5280, n5279 );
nand U13725 ( n6584, n7538, n7539 );
nor U13726 ( n7539, n7540, n7541 );
nor U13727 ( n7538, n7554, n6322 );
nor U13728 ( n7540, n984, n11364 );
not U13729 ( n533, n4324 );
nor U13730 ( n4359, n4360, n4361 );
nand U13731 ( n4361, n4362, n4326 );
nand U13732 ( n4362, n533, n4325 );
xor U13733 ( n8950, n8951, n8952 );
and U13734 ( n4358, n4360, n11225 );
and U13735 ( n11225, n4364, n4325 );
or U13736 ( n3519, n3385, n2906 );
nor U13737 ( n4476, n4482, n4483 );
xnor U13738 ( n4482, n982, n4489 );
nand U13739 ( n4483, n4484, n4282 );
nand U13740 ( n4484, n4281, n4283 );
nor U13741 ( n7055, n11466, n646 );
xnor U13742 ( n2208, n3439, n3456 );
nand U13743 ( n6285, n7452, n7453 );
nand U13744 ( n7453, n7454, n689 );
nor U13745 ( n7454, n7436, n7455 );
nor U13746 ( n7455, n7434, n7456 );
nor U13747 ( n7451, n561, n11341 );
not U13748 ( n561, n6285 );
nand U13749 ( n3510, n351, n3385 );
nor U13750 ( n9504, n9509, n9510 );
nor U13751 ( n9510, n9511, n9512 );
nand U13752 ( n9511, n9543, n9544 );
nand U13753 ( n9512, n9513, n9514 );
nor U13754 ( n9513, n9525, n9526 );
nor U13755 ( n9526, n9527, n9528 );
nor U13756 ( n9525, n9530, n9531 );
nand U13757 ( n9528, n177, n174 );
nand U13758 ( n9499, n3482, n9500 );
nand U13759 ( n9500, n9501, n9502 );
nand U13760 ( n9502, n186, n9503 );
nand U13761 ( n9503, n9504, n9505 );
nand U13762 ( n3512, n337, n3385 );
not U13763 ( n681, n7146 );
nand U13764 ( n11289, n4702, n4703 );
buf U13765 ( n11269, n11332 );
nor U13766 ( n9546, n9548, n3389 );
xnor U13767 ( n4658, n984, n4659 );
nand U13768 ( n4659, n4660, n4632 );
nor U13769 ( n4660, n4662, n4663 );
nor U13770 ( n4662, n4664, n4074 );
nand U13771 ( n9605, n3389, n198 );
nand U13772 ( n2613, n3577, n3578 );
nor U13773 ( n3578, n3579, n3580 );
nor U13774 ( n3577, n3591, n2284 );
nor U13775 ( n3579, n302, n11432 );
nand U13776 ( n9783, n9741, n9740 );
not U13777 ( n11418, n11420 );
xnor U13778 ( n4526, n723, n11297 );
nand U13779 ( n7452, n7470, n7471 );
nor U13780 ( n7470, n7434, n689 );
nand U13781 ( n7471, n7456, n693 );
xnor U13782 ( n4418, n728, n11290 );
nand U13783 ( n4277, n4278, n534 );
xnor U13784 ( n4278, n981, n4279 );
nand U13785 ( n4320, n4321, n533 );
xnor U13786 ( n4321, n986, n4322 );
nand U13787 ( n5014, n5021, n4982 );
nor U13788 ( n5021, n757, n5061 );
nor U13789 ( n5061, n763, n4993 );
not U13790 ( n757, n4992 );
nand U13791 ( n4995, n5041, n5042 );
nand U13792 ( n5042, n5034, n5033 );
nand U13793 ( n5041, n5037, n5036 );
nor U13794 ( n4961, n4962, n4963 );
nor U13795 ( n4962, n5092, n5093 );
nand U13796 ( n4963, n4964, n4965 );
nand U13797 ( n4964, n5083, n726 );
and U13798 ( n4982, n5022, n5023 );
nor U13799 ( n5022, n5049, n5050 );
nor U13800 ( n5023, n5024, n5025 );
nor U13801 ( n5049, n5037, n5036 );
nor U13802 ( n5000, n5013, n5014 );
nor U13803 ( n5013, n5015, n5016 );
and U13804 ( n4951, n4958, n4959 );
nand U13805 ( n4958, n5096, n5097 );
nand U13806 ( n4959, n4960, n4961 );
nor U13807 ( n4960, n5094, n5095 );
nand U13808 ( n4965, n4966, n4967 );
nor U13809 ( n4966, n5073, n5074 );
nor U13810 ( n4967, n4968, n4969 );
nand U13811 ( n5074, n5075, n5076 );
nor U13812 ( n5024, n4997, n5038 );
nand U13813 ( n5038, n744, n4996 );
not U13814 ( n744, n4995 );
nand U13815 ( n9514, n9515, n9516 );
nor U13816 ( n9515, n9517, n9518 );
nor U13817 ( n9518, n9519, n9520 );
nand U13818 ( n9520, n9521, n3778 );
nand U13819 ( n9521, n9522, n9523 );
nand U13820 ( n9523, n48, n3886 );
nor U13821 ( n7502, n558, n11341 );
not U13822 ( n558, n6297 );
or U13823 ( n11226, n2545, n1878 );
nor U13824 ( n9611, n9612, n138 );
nand U13825 ( n4276, n4280, n4281 );
nand U13826 ( n4280, n4282, n4283 );
or U13827 ( n11227, n2539, n1878 );
nand U13828 ( n7249, n666, n7216 );
nor U13829 ( n3087, n266, n11415 );
nand U13830 ( n4319, n4323, n4324 );
nand U13831 ( n4323, n4325, n4326 );
nand U13832 ( n5025, n5026, n5027 );
nand U13833 ( n5027, n4978, n4977 );
nand U13834 ( n5026, n5032, n749 );
not U13835 ( n749, n5033 );
nor U13836 ( n5032, n5034, n5035 );
and U13837 ( n5035, n5036, n5037 );
nand U13838 ( n3570, n3571, n3572 );
nand U13839 ( n3571, n3567, n352 );
nand U13840 ( n3572, n3567, n351 );
nand U13841 ( n4193, n4702, n4703 );
nand U13842 ( n11288, n4702, n4703 );
nor U13843 ( n9501, n3527, n3388 );
nand U13844 ( n9530, n9541, n9522 );
nor U13845 ( n9541, n3909, n9517 );
nor U13846 ( n7112, n11466, n652 );
nand U13847 ( n3493, n3494, n3495 );
nand U13848 ( n3495, n2231, n11491 );
nand U13849 ( n3494, n11411, n2232 );
nand U13850 ( n2328, n3665, n3666 );
nor U13851 ( n3665, n3680, n3681 );
nor U13852 ( n3666, n3667, n3668 );
nor U13853 ( n3681, n297, n283 );
nand U13854 ( n3678, n3647, n3708 );
or U13855 ( n3708, n3640, n3639 );
nand U13856 ( n2619, n3653, n3654 );
nor U13857 ( n3654, n3655, n3656 );
nor U13858 ( n3653, n3664, n2328 );
nor U13859 ( n3655, n299, n11432 );
nor U13860 ( n3671, n3645, n3673 );
nor U13861 ( n3673, n3674, n26 );
nand U13862 ( n3580, n3581, n3582 );
nand U13863 ( n3582, n2276, n11491 );
nand U13864 ( n3581, n11411, n2272 );
nand U13865 ( n5244, n5245, n5246 );
nor U13866 ( n5246, n5247, n5248 );
nor U13867 ( n5245, n5249, n5250 );
nor U13868 ( n5249, n5251, n5252 );
nor U13869 ( n5262, n5263, n5264 );
nand U13870 ( n5264, n743, n5265 );
nor U13871 ( n5225, n5227, n5228 );
nand U13872 ( n5228, n5229, n5230 );
nand U13873 ( n5227, n5233, n5234 );
nand U13874 ( n5230, n5231, n5232 );
nand U13875 ( n5251, n5256, n5257 );
nand U13876 ( n5257, n5258, n5259 );
nor U13877 ( n5256, n5261, n5262 );
nand U13878 ( n5258, n5260, n748 );
nor U13879 ( n5233, n5237, n5238 );
nor U13880 ( n5237, n5239, n5240 );
nand U13881 ( n5240, n5236, n5241 );
nand U13882 ( n5239, n5243, n5244 );
nand U13883 ( n4799, n7217, n7259 );
nand U13884 ( n4950, n4951, n4952 );
not U13885 ( n11382, n11384 );
nor U13886 ( n9522, n9542, n3784 );
not U13887 ( n11315, n9727 );
nand U13888 ( n6587, n7585, n7586 );
nor U13889 ( n7586, n7587, n7588 );
nor U13890 ( n7585, n7597, n6334 );
nor U13891 ( n7588, n983, n11364 );
xnor U13892 ( n8777, n8778, n8779 );
nor U13893 ( n4979, n4981, n4980 );
nor U13894 ( n3295, n9600, n9495 );
xnor U13895 ( n4072, n983, n4073 );
nand U13896 ( n4073, n4074, n4075 );
nand U13897 ( n4075, n4076, n4077 );
and U13898 ( n9516, n9533, n9534 );
nor U13899 ( n9534, n3702, n9529 );
nor U13900 ( n9533, n3786, n3738 );
not U13901 ( n692, n5133 );
nor U13902 ( n9527, n3711, n3735 );
nand U13903 ( n3656, n3657, n3658 );
nand U13904 ( n3658, n2321, n11491 );
nand U13905 ( n3657, n25, n11410 );
nand U13906 ( n4973, n5051, n5052 );
not U13907 ( n44, n3205 );
nand U13908 ( n6590, n7620, n7621 );
nor U13909 ( n7621, n7622, n7623 );
nor U13910 ( n7620, n7632, n6346 );
nor U13911 ( n7622, n982, n11364 );
nor U13912 ( n3630, n3625, n3632 );
nor U13913 ( n3632, n3633, n3634 );
nor U13914 ( n3634, n3515, n3617 );
nor U13915 ( n3633, n3628, n3648 );
nand U13916 ( n2616, n3611, n3612 );
nor U13917 ( n3612, n3613, n3614 );
nor U13918 ( n3611, n3618, n2307 );
nor U13919 ( n3613, n301, n11432 );
nand U13920 ( n2622, n3687, n3688 );
nor U13921 ( n3688, n3689, n3690 );
nor U13922 ( n3687, n3694, n2351 );
nor U13923 ( n3689, n298, n11432 );
nor U13924 ( n7541, n557, n11341 );
not U13925 ( n557, n6317 );
nor U13926 ( n9544, n9545, n9508 );
nand U13927 ( n5073, n5086, n5087 );
nand U13928 ( n5087, n714, n5088 );
not U13929 ( n714, n5089 );
nand U13930 ( n5086, n5092, n5093 );
nor U13931 ( n5083, n5077, n5073 );
nand U13932 ( n5263, n759, n8055 );
not U13933 ( n759, n8019 );
nand U13934 ( n5252, n5253, n5254 );
nand U13935 ( n5254, n743, n5255 );
buf U13936 ( n11495, n108 );
nor U13937 ( n8601, n8610, n8611 );
xor U13938 ( n8610, n8612, n8613 );
nor U13939 ( n3149, n277, n11415 );
nor U13940 ( n7177, n11466, n657 );
nand U13941 ( n4798, n681, n7155 );
nand U13942 ( n4992, n4988, n4989 );
nor U13943 ( n4986, n4990, n4991 );
nand U13944 ( n4991, n4992, n4993 );
nand U13945 ( n4983, n4984, n4985 );
nor U13946 ( n4984, n4994, n4995 );
nor U13947 ( n4985, n4986, n4987 );
nor U13948 ( n4994, n753, n4996 );
nand U13949 ( n6358, n7678, n7679 );
nor U13950 ( n7678, n7698, n7699 );
nor U13951 ( n7679, n7680, n7681 );
nor U13952 ( n7699, n978, n6677 );
nor U13953 ( n7681, n7682, n4828 );
nor U13954 ( n7682, n7683, n7684 );
nor U13955 ( n7683, n7642, n7686 );
nor U13956 ( n7684, n7685, n7646 );
nand U13957 ( n6593, n7659, n7660 );
nor U13958 ( n7660, n7661, n7662 );
nor U13959 ( n7659, n7677, n6358 );
nor U13960 ( n7661, n981, n11364 );
not U13961 ( n763, n4990 );
nor U13962 ( n3248, n3211, n3227 );
nand U13963 ( n5146, n5134, n5133 );
buf U13964 ( n11260, n11317 );
nor U13965 ( n9543, n3628, n3684 );
not U13966 ( n43, n3294 );
or U13967 ( n4975, n11228, n4977 );
or U13968 ( n11228, n4978, n4979 );
nand U13969 ( n7668, n5267, n7741 );
nand U13970 ( n7741, n7742, n7643 );
buf U13971 ( n11261, n11317 );
nor U13972 ( n5094, n5088, n5098 );
nand U13973 ( n5098, n5086, n5089 );
nand U13974 ( n3373, n3328, n3325 );
nor U13975 ( n3352, n208, n3368 );
xnor U13976 ( n4813, n683, n987 );
not U13977 ( n753, n4997 );
nand U13978 ( n9505, n9506, n136 );
nand U13979 ( n9506, n146, n9507 );
not U13980 ( n146, n3602 );
nand U13981 ( n9507, n3601, n143 );
nor U13982 ( n7587, n556, n11341 );
nor U13983 ( n4987, n4988, n4989 );
nand U13984 ( n9090, n5, n9091 );
xor U13985 ( n9091, n9092, n9093 );
and U13986 ( n5236, n5232, n5242 );
nor U13987 ( n3213, n279, n11415 );
xor U13988 ( n2366, n3730, n3639 );
nand U13989 ( n2625, n3714, n3715 );
nor U13990 ( n3715, n3716, n3717 );
nor U13991 ( n3714, n3724, n2373 );
nor U13992 ( n3716, n297, n11432 );
not U13993 ( n853, n5588 );
buf U13994 ( n11459, n964 );
nor U13995 ( n7242, n11466, n669 );
not U13996 ( n42, n3401 );
xnor U13997 ( n2171, n3294, n209 );
not U13998 ( n24, n3749 );
nand U13999 ( n2394, n3760, n3761 );
nor U14000 ( n3760, n3773, n3774 );
nor U14001 ( n3761, n3762, n3763 );
nor U14002 ( n3774, n293, n283 );
nand U14003 ( n3758, n3764, n3765 );
nand U14004 ( n3764, n3770, n3771 );
nand U14005 ( n3765, n3766, n3767 );
nor U14006 ( n3770, n3769, n3767 );
nand U14007 ( n2628, n3752, n3753 );
nor U14008 ( n3753, n3754, n3755 );
nor U14009 ( n3752, n3759, n2394 );
nor U14010 ( n3754, n296, n11432 );
nor U14011 ( n3766, n3743, n3768 );
nor U14012 ( n3768, n3769, n24 );
nand U14013 ( n4974, n4980, n4981 );
not U14014 ( n11259, n11316 );
nor U14015 ( n5095, n5096, n5097 );
nand U14016 ( n6596, n7710, n7711 );
nor U14017 ( n7711, n7712, n7713 );
nor U14018 ( n7710, n7725, n6370 );
nor U14019 ( n7712, n979, n11364 );
nand U14020 ( n6370, n7726, n7727 );
nor U14021 ( n7726, n7739, n7740 );
nor U14022 ( n7727, n7728, n7729 );
nor U14023 ( n7740, n977, n6677 );
not U14024 ( n602, n5016 );
nor U14025 ( n7623, n6341, n11341 );
xnor U14026 ( n8892, n8893, n8894 );
or U14027 ( n5243, n5250, n11229 );
and U14028 ( n11229, n5267, n5268 );
nor U14029 ( n5113, n706, n11406 );
nand U14030 ( n5234, n5235, n5236 );
nand U14031 ( n6353, n7663, n7664 );
nand U14032 ( n7664, n7665, n709 );
nor U14033 ( n7665, n7642, n7666 );
nor U14034 ( n7666, n7667, n7668 );
nand U14035 ( n3717, n3718, n3719 );
nand U14036 ( n3719, n2364, n11491 );
nand U14037 ( n3718, n11411, n2366 );
nor U14038 ( n7662, n594, n11340 );
not U14039 ( n594, n6353 );
or U14040 ( n5075, n5052, n5051 );
not U14041 ( n697, n7434 );
nand U14042 ( n3405, n3381, n3389 );
nand U14043 ( n6599, n7752, n7753 );
nor U14044 ( n7753, n7754, n7755 );
nor U14045 ( n7752, n7764, n6382 );
nor U14046 ( n7754, n978, n11364 );
nand U14047 ( n5076, n5077, n5078 );
not U14048 ( n192, n3388 );
not U14049 ( n693, n7436 );
not U14050 ( n41, n3499 );
not U14051 ( n707, n7438 );
xnor U14052 ( n2216, n3401, n197 );
nand U14053 ( n4787, n7378, n691 );
nand U14054 ( n7663, n7700, n7701 );
nor U14055 ( n7700, n7667, n709 );
nand U14056 ( n7701, n7668, n719 );
nor U14057 ( n1908, n11431, n1878 );
nor U14058 ( n3456, n3416, n3446 );
nor U14059 ( n3249, n217, n11415 );
xor U14060 ( n8907, n101, n8912 );
nand U14061 ( n6377, n7769, n7770 );
nand U14062 ( n7770, n7742, n7771 );
nand U14063 ( n7769, n4797, n591 );
nand U14064 ( n7771, n7643, n5267 );
xor U14065 ( n8936, n8937, n8938 );
nor U14066 ( n7713, n592, n11340 );
not U14067 ( n592, n6365 );
nand U14068 ( n2404, n3804, n3805 );
nand U14069 ( n3805, n3806, n3749 );
nand U14070 ( n3804, n24, n147 );
nand U14071 ( n3806, n152, n154 );
nand U14072 ( n2631, n3789, n3790 );
nor U14073 ( n3790, n3791, n3792 );
nor U14074 ( n3789, n3799, n2417 );
nor U14075 ( n3791, n294, n11433 );
nand U14076 ( n2417, n3800, n3801 );
nor U14077 ( n3800, n3828, n3829 );
nor U14078 ( n3801, n3802, n3803 );
nor U14079 ( n3829, n292, n283 );
nor U14080 ( n7292, n674, n11466 );
not U14081 ( n909, n6111 );
nor U14082 ( n4026, n4027, n4028 );
nand U14083 ( n4028, n4029, n4030 );
nand U14084 ( n4030, n537, n4031 );
not U14085 ( n537, n4036 );
nor U14086 ( n3727, n3733, n3734 );
or U14087 ( n3734, n3730, n3735 );
nor U14088 ( n3733, n3736, n10 );
nor U14089 ( n3736, n334, n182 );
not U14090 ( n75, n8798 );
nand U14091 ( n6394, n7822, n7823 );
nor U14092 ( n7822, n7843, n7844 );
nor U14093 ( n7823, n7824, n7825 );
nor U14094 ( n7844, n974, n6677 );
nor U14095 ( n7825, n7826, n729 );
nor U14096 ( n7826, n7827, n7828 );
nor U14097 ( n7827, n5247, n7830 );
nor U14098 ( n7828, n7685, n7829 );
nand U14099 ( n6602, n7803, n7804 );
nor U14100 ( n7804, n7805, n7806 );
nor U14101 ( n7803, n7821, n6394 );
nor U14102 ( n7805, n977, n11364 );
nand U14103 ( n7812, n7888, n7889 );
nand U14104 ( n7889, n7780, n5259 );
nand U14105 ( n7888, n743, n552 );
not U14106 ( n546, n7913 );
nor U14107 ( n7926, n7927, n739 );
nor U14108 ( n7927, n7928, n7929 );
nor U14109 ( n7929, n7685, n7842 );
nor U14110 ( n7928, n7892, n7930 );
nand U14111 ( n6614, n7903, n7904 );
nor U14112 ( n7904, n7905, n7906 );
nor U14113 ( n7903, n7922, n6418 );
nor U14114 ( n7905, n974, n11364 );
nand U14115 ( n6418, n7923, n7924 );
nor U14116 ( n7923, n7945, n7946 );
nor U14117 ( n7924, n7925, n7926 );
nor U14118 ( n7946, n972, n6677 );
not U14119 ( n726, n5078 );
xnor U14120 ( n2261, n3499, n188 );
not U14121 ( n40, n3586 );
nor U14122 ( n4025, n4032, n4033 );
xnor U14123 ( n4032, n974, n4037 );
nand U14124 ( n4033, n4034, n4031 );
nand U14125 ( n4034, n4035, n4036 );
xor U14126 ( n4360, n987, n4365 );
nor U14127 ( n3802, n3823, n3824 );
nand U14128 ( n3824, n147, n3778 );
nor U14129 ( n3823, n3826, n9 );
nor U14130 ( n3826, n334, n157 );
or U14131 ( n3833, n3784, n11230 );
and U14132 ( n11230, n3861, n3779 );
nand U14133 ( n3500, n3482, n192 );
buf U14134 ( n11381, n11378 );
nand U14135 ( n3792, n3793, n3794 );
nand U14136 ( n3794, n2408, n11491 );
nand U14137 ( n3793, n11411, n2404 );
nor U14138 ( n3414, n3405, n3446 );
nor U14139 ( n6397, n736, n11381 );
nor U14140 ( n7755, n553, n11340 );
nor U14141 ( n6465, n762, n11381 );
nor U14142 ( n6477, n601, n11381 );
nor U14143 ( n6421, n747, n11381 );
nor U14144 ( n6409, n741, n11381 );
nor U14145 ( n6441, n752, n11381 );
nor U14146 ( n6453, n756, n11381 );
nor U14147 ( n6385, n731, n11380 );
buf U14148 ( n11380, n11378 );
buf U14149 ( n11379, n11378 );
nand U14150 ( n2438, n3844, n3845 );
nor U14151 ( n3844, n3858, n3859 );
nor U14152 ( n3845, n3846, n3847 );
nor U14153 ( n3859, n291, n283 );
nand U14154 ( n3882, n3822, n3821 );
nand U14155 ( n2634, n3836, n3837 );
nor U14156 ( n3837, n3838, n3839 );
nor U14157 ( n3836, n3843, n2438 );
nor U14158 ( n3838, n293, n11433 );
nor U14159 ( n3855, n3809, n3856 );
nor U14160 ( n3856, n3853, n3852 );
and U14161 ( n3852, n3817, n3880 );
nand U14162 ( n3880, n3881, n3882 );
nand U14163 ( n3881, n289, n162 );
nand U14164 ( n3842, n3848, n3849 );
nand U14165 ( n3849, n3850, n3851 );
nand U14166 ( n3848, n3855, n3854 );
nor U14167 ( n3850, n3853, n3854 );
buf U14168 ( n11262, n11317 );
nor U14169 ( n3296, n204, n11415 );
nor U14170 ( n3828, n3830, n3831 );
nand U14171 ( n3830, n3626, n157 );
nand U14172 ( n3831, n3825, n3832 );
nand U14173 ( n3832, n3833, n3778 );
nor U14174 ( n7345, n678, n11466 );
nand U14175 ( n4573, n4574, n537 );
xnor U14176 ( n4574, n973, n4575 );
nand U14177 ( n6406, n7873, n7874 );
nor U14178 ( n7873, n7886, n7887 );
nor U14179 ( n7874, n7875, n7876 );
nor U14180 ( n7887, n973, n6677 );
nand U14181 ( n7880, n7881, n4812 );
nor U14182 ( n7881, n7836, n7882 );
nor U14183 ( n7882, n7883, n506 );
nand U14184 ( n6605, n7857, n7858 );
nor U14185 ( n7858, n7859, n7860 );
nor U14186 ( n7857, n7872, n6406 );
nor U14187 ( n7860, n976, n11364 );
nor U14188 ( n3590, n9545, n9509 );
nand U14189 ( n4779, n7526, n7523 );
nand U14190 ( n4784, n7483, n7480 );
buf U14191 ( n11493, n108 );
not U14192 ( n6, n9064 );
not U14193 ( n39, n3662 );
xnor U14194 ( n2306, n3586, n144 );
nor U14195 ( n3560, n9612, n3527 );
nand U14196 ( n4572, n4576, n4036 );
nand U14197 ( n4576, n4031, n4035 );
nor U14198 ( n3767, n3738, n3735 );
nand U14199 ( n6389, n7807, n7808 );
nand U14200 ( n7808, n7809, n7810 );
nor U14201 ( n7809, n5247, n7811 );
nor U14202 ( n7811, n5261, n7812 );
nand U14203 ( n6413, n7907, n7908 );
nand U14204 ( n7908, n7909, n7910 );
nor U14205 ( n7909, n7892, n7911 );
nor U14206 ( n7911, n7912, n7913 );
nor U14207 ( n7806, n551, n11340 );
not U14208 ( n551, n6389 );
nor U14209 ( n7906, n547, n11340 );
not U14210 ( n547, n6413 );
nand U14211 ( n2637, n3864, n3865 );
nor U14212 ( n3865, n3866, n3867 );
nor U14213 ( n3864, n3874, n2461 );
nor U14214 ( n3866, n292, n11433 );
nor U14215 ( n3693, n3645, n3674 );
nor U14216 ( n9674, n9678, n9679 );
nand U14217 ( n9678, n159, n3854 );
nand U14218 ( n9679, n3972, n3933 );
xnor U14219 ( n4342, n4343, n972 );
nor U14220 ( n3933, n3909, n9524 );
nor U14221 ( n3672, n3628, n3601 );
nand U14222 ( n6617, n7959, n7960 );
nor U14223 ( n7960, n7961, n7962 );
nor U14224 ( n7959, n7974, n6430 );
nor U14225 ( n7961, n973, n11365 );
nor U14226 ( n3625, n9508, n3602 );
nor U14227 ( n3730, n9529, n3711 );
nand U14228 ( n2640, n3889, n3890 );
nor U14229 ( n3890, n3891, n3892 );
nor U14230 ( n3889, n3895, n2482 );
nor U14231 ( n3891, n291, n11433 );
nand U14232 ( n7907, n7947, n7948 );
nor U14233 ( n7947, n7912, n7910 );
nand U14234 ( n7948, n7913, n746 );
nand U14235 ( n7807, n7845, n7846 );
nor U14236 ( n7845, n5261, n7810 );
nand U14237 ( n7846, n7812, n733 );
and U14238 ( n3854, n3778, n157 );
nand U14239 ( n9060, n6, n9061 );
xor U14240 ( n9061, n9062, n9063 );
xnor U14241 ( n2349, n3662, n173 );
nor U14242 ( n7403, n683, n11467 );
not U14243 ( n38, n3723 );
nor U14244 ( n3354, n209, n11415 );
nand U14245 ( n3907, n161, n3886 );
nand U14246 ( n3959, n3941, n3944 );
nand U14247 ( n6620, n8000, n8001 );
nor U14248 ( n8001, n8002, n8003 );
nor U14249 ( n8000, n8012, n6450 );
nor U14250 ( n8003, n972, n11365 );
nor U14251 ( n3825, n3786, n149 );
nor U14252 ( n3589, n3537, n3562 );
nand U14253 ( n9059, n9065, n9064 );
nand U14254 ( n9065, n8699, n8698 );
nor U14255 ( n7859, n548, n11340 );
not U14256 ( n548, n6401 );
nor U14257 ( n7962, n544, n11340 );
not U14258 ( n544, n6425 );
nand U14259 ( n6425, n7963, n7964 );
nand U14260 ( n7964, n7965, n7913 );
nand U14261 ( n7963, n546, n4786 );
nand U14262 ( n3867, n3868, n3869 );
nand U14263 ( n3869, n2452, n11491 );
nand U14264 ( n3868, n2453, n11410 );
buf U14265 ( n11393, n11396 );
nor U14266 ( n4715, n11382, n6037 );
nor U14267 ( n6133, n11363, n6111 );
not U14268 ( n868, n5934 );
nor U14269 ( n7544, n5238, n7438 );
xnor U14270 ( n4402, n971, n4403 );
nor U14271 ( n7978, n7913, n7979 );
nand U14272 ( n7979, n6837, n4786 );
nand U14273 ( n2502, n3924, n3925 );
nor U14274 ( n3924, n3937, n3938 );
nor U14275 ( n3925, n3926, n3927 );
nor U14276 ( n3938, n287, n283 );
nor U14277 ( n3926, n3933, n3934 );
nor U14278 ( n3934, n3935, n3936 );
nor U14279 ( n3935, n3166, n3900 );
and U14280 ( n3936, n3626, n3910 );
nand U14281 ( n2643, n3913, n3914 );
nor U14282 ( n3914, n3915, n3916 );
nor U14283 ( n3913, n3923, n2502 );
nor U14284 ( n3915, n289, n11433 );
nand U14285 ( n7985, n7942, n8024 );
nand U14286 ( n8024, n8025, n7943 );
nor U14287 ( n7980, n4786, n7986 );
nand U14288 ( n7986, n7987, n7944 );
nand U14289 ( n7987, n527, n7938 );
not U14290 ( n527, n7985 );
nor U14291 ( n3932, n334, n3910 );
nand U14292 ( n3927, n3928, n3929 );
nand U14293 ( n3929, n3930, n3931 );
nand U14294 ( n3928, n3932, n3933 );
nor U14295 ( n3930, n21, n3166 );
nor U14296 ( n3565, n188, n302 );
xnor U14297 ( n2393, n3723, n184 );
not U14298 ( n37, n3798 );
nand U14299 ( n4828, n7647, n7648 );
nor U14300 ( n8002, n543, n11340 );
nor U14301 ( n7910, n7836, n7883 );
nor U14302 ( n7465, n688, n11467 );
nand U14303 ( n7981, n7982, n6682 );
nand U14304 ( n7982, n7983, n7984 );
and U14305 ( n7983, n4786, n7938 );
nand U14306 ( n7984, n7985, n7944 );
nand U14307 ( n3916, n3917, n3918 );
nand U14308 ( n3918, n2493, n11491 );
nand U14309 ( n3917, n20, n11410 );
nor U14310 ( n3406, n124, n11415 );
nor U14311 ( n8053, n8019, n8054 );
nor U14312 ( n8054, n8022, n8055 );
nand U14313 ( n6623, n8035, n8036 );
nor U14314 ( n8036, n8037, n8038 );
nor U14315 ( n8035, n8046, n6462 );
nor U14316 ( n8037, n971, n11365 );
nand U14317 ( n6457, n8051, n8052 );
nand U14318 ( n8051, n8056, n5263 );
nand U14319 ( n8052, n8053, n754 );
nor U14320 ( n8056, n8022, n754 );
buf U14321 ( n11394, n11396 );
nor U14322 ( n7810, n7784, n7782 );
not U14323 ( n737, n5261 );
nor U14324 ( n3677, n133, n298 );
buf U14325 ( n11350, n11347 );
xor U14326 ( n8695, n92, n8702 );
xnor U14327 ( n4812, n736, n974 );
not U14328 ( n538, n4543 );
nor U14329 ( n4127, n4128, n4129 );
nand U14330 ( n4129, n4130, n4131 );
nand U14331 ( n4130, n538, n4132 );
and U14332 ( n8965, n1247, n11505 );
xnor U14333 ( n2437, n3798, n158 );
not U14334 ( n36, n3873 );
and U14335 ( n4126, n4128, n11231 );
and U14336 ( n11231, n4134, n4132 );
xnor U14337 ( n2511, n3959, n3943 );
nand U14338 ( n2646, n3947, n3948 );
nor U14339 ( n3948, n3949, n3950 );
nor U14340 ( n3947, n3953, n2523 );
nor U14341 ( n3949, n288, n11433 );
buf U14342 ( n11392, n11397 );
nor U14343 ( n8797, n168, n8798 );
nand U14344 ( n4827, n7938, n7944 );
nor U14345 ( n9067, n49, n8798 );
nand U14346 ( n3931, n3901, n3822 );
nor U14347 ( n3700, n3702, n3684 );
nand U14348 ( n4786, n7937, n7934 );
nand U14349 ( n4829, n7943, n7942 );
nand U14350 ( n4785, n8061, n8058 );
nand U14351 ( n6502, n11480, n6504 );
nand U14352 ( n6484, n11480, n6486 );
nand U14353 ( n6626, n8070, n8071 );
nor U14354 ( n8071, n8072, n8073 );
nor U14355 ( n8070, n8080, n6474 );
nor U14356 ( n8073, n969, n11365 );
nand U14357 ( n6469, n8092, n8093 );
nand U14358 ( n8093, n8094, n8055 );
nand U14359 ( n8092, n596, n4785 );
or U14360 ( n8094, n8022, n8019 );
nand U14361 ( n4780, n8086, n8089 );
nor U14362 ( n8038, n597, n11340 );
nand U14363 ( n2649, n3965, n3966 );
nor U14364 ( n3965, n3975, n3976 );
nor U14365 ( n3966, n2546, n3967 );
nor U14366 ( n3975, n287, n11431 );
not U14367 ( n8, n3972 );
not U14368 ( n11411, n11412 );
nor U14369 ( n3457, n197, n11415 );
nand U14370 ( n3950, n3951, n3952 );
nand U14371 ( n3952, n11492, n2522 );
nand U14372 ( n3951, n11411, n2511 );
not U14373 ( n733, n5247 );
nor U14374 ( n7514, n696, n11467 );
nand U14375 ( n4541, n4542, n538 );
xnor U14376 ( n4542, n968, n4544 );
not U14377 ( n81, n2652 );
nor U14378 ( n3976, n3972, n11413 );
nor U14379 ( n7554, n706, n11467 );
xnor U14380 ( n2481, n3873, n162 );
nor U14381 ( n4439, n966, n11399 );
nor U14382 ( n3501, n193, n11415 );
buf U14383 ( n11399, n11398 );
not U14384 ( n541, n6481 );
nand U14385 ( n6629, n8109, n8110 );
nor U14386 ( n8110, n8111, n8112 );
nor U14387 ( n8109, n8119, n6486 );
nor U14388 ( n8111, n968, n11365 );
nor U14389 ( n4144, n991, n11400 );
nor U14390 ( n4413, n978, n11399 );
nor U14391 ( n4567, n974, n11399 );
buf U14392 ( n11400, n11398 );
nor U14393 ( n4314, n987, n11400 );
nand U14394 ( n5419, n11460, n5975 );
nor U14395 ( n4271, n982, n11400 );
nor U14396 ( n4121, n971, n11400 );
nor U14397 ( n4246, n993, n11400 );
nor U14398 ( n4202, n977, n11400 );
nor U14399 ( n4589, n999, n11399 );
nor U14400 ( n4396, n972, n11399 );
nor U14401 ( n4449, n992, n11399 );
nor U14402 ( n4375, n997, n11400 );
nor U14403 ( n4471, n983, n11399 );
nor U14404 ( n4653, n986, n11399 );
nor U14405 ( n4336, n973, n11400 );
nor U14406 ( n4550, n989, n11399 );
nor U14407 ( n4293, n998, n11400 );
nor U14408 ( n4516, n981, n11399 );
nor U14409 ( n4353, n988, n11400 );
nor U14410 ( n4162, n1002, n11400 );
nor U14411 ( n4499, n994, n11399 );
nand U14412 ( n4540, n4545, n4543 );
nand U14413 ( n4545, n4132, n4131 );
nor U14414 ( n4546, n969, n11399 );
nor U14415 ( n4241, n968, n11400 );
nor U14416 ( n4087, n996, n11401 );
nor U14417 ( n4066, n984, n11401 );
buf U14418 ( n11401, n11398 );
nor U14419 ( n4049, n1001, n11401 );
nor U14420 ( n4020, n976, n11401 );
nor U14421 ( n4105, n979, n11401 );
nor U14422 ( n8072, n542, n11340 );
nand U14423 ( n5418, n6037, n5975 );
xor U14424 ( n8124, n4780, n8088 );
nor U14425 ( n6112, n4748, n6111 );
nor U14426 ( n3591, n137, n11414 );
nor U14427 ( n7632, n702, n11467 );
nor U14428 ( n5202, n1003, n1004 );
nand U14429 ( n4232, n4233, n4234 );
nor U14430 ( n3548, n188, n11415 );
not U14431 ( n329, n2672 );
xor U14432 ( n4128, n969, n4135 );
nand U14433 ( n4231, n599, n4235 );
not U14434 ( n599, n4233 );
nand U14435 ( n4235, n4236, n4237 );
nand U14436 ( n4237, n967, n4238 );
nor U14437 ( n8112, n541, n11340 );
nor U14438 ( n7597, n717, n11467 );
not U14439 ( n879, n5907 );
xor U14440 ( n4233, n966, n4239 );
nor U14441 ( n8139, n966, n11365 );
nor U14442 ( n3953, n168, n11414 );
nand U14443 ( n2701, n2672, n11419 );
nor U14444 ( n3694, n173, n11414 );
nor U14445 ( n3759, n184, n11414 );
nor U14446 ( n3923, n49, n11414 );
nor U14447 ( n3895, n162, n11414 );
nor U14448 ( n3664, n133, n11414 );
nor U14449 ( n3618, n144, n11414 );
nor U14450 ( n3843, n158, n11414 );
nor U14451 ( n3724, n179, n11414 );
nor U14452 ( n3799, n153, n11414 );
nor U14453 ( n3874, n164, n11414 );
nor U14454 ( n7677, n712, n11467 );
nor U14455 ( n7989, n971, n6677 );
nor U14456 ( n7562, n982, n6677 );
nor U14457 ( n8135, n528, n11340 );
not U14458 ( n528, n6493 );
not U14459 ( n942, n4744 );
buf U14460 ( n11395, n11396 );
nor U14461 ( n7476, n984, n6677 );
not U14462 ( n11422, n11423 );
nor U14463 ( n6909, n997, n6677 );
nor U14464 ( n4441, n4443, n4444 );
xor U14465 ( n4443, n4445, n4446 );
xnor U14466 ( n4445, n967, n923 );
not U14467 ( n71, n1203 );
nand U14468 ( n10808, n10801, n10802 );
and U14469 ( n10800, n10801, n10802 );
nor U14470 ( n7872, n736, n11467 );
not U14471 ( n69, n1229 );
not U14472 ( n70, n1194 );
nand U14473 ( n1614, n1616, n1617 );
nand U14474 ( n1617, n1618, n11284 );
nand U14475 ( n1616, n1631, n70 );
nor U14476 ( n1618, n1619, n1621 );
nand U14477 ( n1354, n1356, n1357 );
nand U14478 ( n1357, n1358, n11284 );
nand U14479 ( n1356, n1371, n70 );
nor U14480 ( n1358, n1359, n1361 );
nand U14481 ( n1283, n1284, n1286 );
nand U14482 ( n1286, n1287, n11285 );
nand U14483 ( n1284, n1306, n70 );
nor U14484 ( n1287, n1288, n1289 );
nor U14485 ( n4440, n4044, n11282 );
nor U14486 ( n7725, n723, n11467 );
nor U14487 ( n7922, n741, n11467 );
nor U14488 ( n7974, n747, n11468 );
nor U14489 ( n8012, n752, n11468 );
nor U14490 ( n7821, n731, n11467 );
nor U14491 ( n8080, n762, n11468 );
nor U14492 ( n7764, n728, n11467 );
nor U14493 ( n8046, n756, n11468 );
nor U14494 ( n8119, n601, n11468 );
buf U14495 ( n11391, n11397 );
buf U14496 ( n11263, n11317 );
not U14497 ( n949, n4734 );
not U14498 ( n11358, n6651 );
nand U14499 ( n6651, n942, n8179 );
nand U14500 ( n8179, n8180, n8181 );
nand U14501 ( n8180, n948, n8184 );
nand U14502 ( n8181, n949, n8182 );
nand U14503 ( n8182, n5315, n918 );
buf U14504 ( n11278, n11424 );
buf U14505 ( n11277, n11424 );
buf U14506 ( n11276, n11424 );
not U14507 ( n109, n9225 );
not U14508 ( n82, n8795 );
nor U14509 ( n4242, n601, n4243 );
nor U14510 ( n8959, n287, n11319 );
nor U14511 ( n8091, n966, n6677 );
not U14512 ( n932, n6677 );
nor U14513 ( n8918, n317, n11320 );
nor U14514 ( n8708, n311, n11320 );
nor U14515 ( n8944, n298, n11319 );
nor U14516 ( n8886, n293, n11320 );
nor U14517 ( n8842, n318, n11320 );
nor U14518 ( n9020, n314, n11319 );
nor U14519 ( n8801, n313, n11320 );
nor U14520 ( n8930, n292, n11319 );
nor U14521 ( n9035, n301, n11319 );
nor U14522 ( n8771, n297, n11320 );
nor U14523 ( n9084, n294, n11319 );
nor U14524 ( n8900, n308, n11320 );
nor U14525 ( n8970, n312, n11319 );
nor U14526 ( n8824, n302, n11320 );
nor U14527 ( n8721, n322, n11320 );
nor U14528 ( n9070, n309, n11319 );
nor U14529 ( n8992, n303, n11319 );
nor U14530 ( n9101, n319, n11319 );
nor U14531 ( n9219, n306, n11319 );
nor U14532 ( n8861, n307, n11320 );
nor U14533 ( n8621, n321, n11321 );
nor U14534 ( n8637, n304, n11321 );
nor U14535 ( n8651, n316, n11321 );
nor U14536 ( n8596, n296, n11321 );
nor U14537 ( n8674, n299, n11321 );
buf U14538 ( n11460, n964 );
nor U14539 ( n3631, n298, n283 );
nor U14540 ( n3173, n311, n283 );
nor U14541 ( n3740, n294, n283 );
nor U14542 ( n2894, n317, n283 );
nor U14543 ( n3266, n308, n283 );
not U14544 ( n336, n2775 );
not U14545 ( n83, n9113 );
nor U14546 ( n3704, n296, n283 );
not U14547 ( n333, n2778 );
not U14548 ( n332, n3166 );
not U14549 ( n912, n4240 );
not U14550 ( n891, n5883 );
nand U14551 ( n3626, n3973, n3974 );
nor U14552 ( n3973, n336, n352 );
nor U14553 ( n3974, n351, n337 );
not U14554 ( n918, n4709 );
nor U14555 ( n9054, n287, n8795 );
nand U14556 ( n8963, n9366, n109 );
not U14557 ( n922, n4243 );
buf U14558 ( n11433, n11430 );
nor U14559 ( n8785, n286, n8795 );
not U14560 ( n916, n4444 );
nor U14561 ( n4535, n966, n4240 );
nand U14562 ( n6837, n7379, n6859 );
nor U14563 ( n7379, n927, n914 );
nor U14564 ( n8960, n8961, n8962 );
nand U14565 ( n8961, n8964, n11533 );
nand U14566 ( n8962, n74, n8963 );
buf U14567 ( n11388, n11389 );
nor U14568 ( n3987, n2652, n112 );
nor U14569 ( n4727, n948, n918 );
nor U14570 ( n7786, n924, n926 );
not U14571 ( n902, n6777 );
not U14572 ( n917, n6859 );
buf U14573 ( n11448, n11238 );
not U14574 ( n903, n5187 );
nor U14575 ( n4712, n5315, n4744 );
and U14576 ( n7359, n7379, n6859 );
not U14577 ( n941, n8253 );
not U14578 ( n346, n2658 );
not U14579 ( n1022, n8304 );
not U14580 ( n919, n6649 );
not U14581 ( n419, n3997 );
nand U14582 ( n1378, n1379, n391 );
not U14583 ( n118, n1866 );
nor U14584 ( n10236, n9694, n9693 );
nand U14585 ( n9690, n9691, n9692 );
nand U14586 ( n9692, n9693, n9694 );
nand U14587 ( n9691, n9695, n9696 );
nor U14588 ( n9696, n9697, n9698 );
nor U14589 ( n1170, n9447, n9448 );
nor U14590 ( n9447, n73, n11533 );
nand U14591 ( n9448, n9449, n9450 );
nand U14592 ( n9450, n9451, n353 );
nand U14593 ( n10240, n10251, n10252 );
nand U14594 ( n10251, n9574, n11263 );
nand U14595 ( n10252, n2665, n11259 );
and U14596 ( n10239, n10253, n10254 );
nand U14597 ( n10254, n9574, n11258 );
nand U14598 ( n10253, n2665, n11263 );
nor U14599 ( n9295, n45, n8749 );
nand U14600 ( n8722, n8723, n8724 );
nand U14601 ( n8723, n11508, n1962 );
nand U14602 ( n8724, n11506, n8725 );
nand U14603 ( n8725, n8726, n8727 );
nand U14604 ( n9064, n9283, n9284 );
nand U14605 ( n9283, n8790, n8793 );
nand U14606 ( n9284, n9285, n8792 );
or U14607 ( n9285, n8793, n8790 );
not U14608 ( n624, n4816 );
and U14609 ( n5197, n11232, n5196 );
or U14610 ( n11232, n619, n4884 );
not U14611 ( n46, n9291 );
nand U14612 ( n5191, n5199, n5200 );
nand U14613 ( n5200, n5201, n5202 );
nand U14614 ( n5199, n5204, n5205 );
nor U14615 ( n5201, n4878, n5203 );
nor U14616 ( n9580, n324, n118 );
nor U14617 ( n9575, n322, n9647 );
or U14618 ( n9647, n1898, n9580 );
nand U14619 ( n9578, n9579, n9574 );
nor U14620 ( n9579, n9580, n2665 );
nand U14621 ( n8622, n8623, n8624 );
nand U14622 ( n8623, n11508, n1984 );
nand U14623 ( n8624, n8625, n11506 );
xor U14624 ( n8625, n8626, n8627 );
nand U14625 ( n9656, n9664, n9665 );
nor U14626 ( n9665, n9666, n9667 );
nor U14627 ( n9664, n9668, n9669 );
nand U14628 ( n9667, n3959, n3879 );
and U14629 ( n4869, n4907, n4908 );
nand U14630 ( n4908, n11403, n4906 );
nand U14631 ( n4907, n624, n11391 );
nand U14632 ( n4870, n4904, n4905 );
nand U14633 ( n4904, n11392, n4906 );
nand U14634 ( n4905, n624, n11402 );
nand U14635 ( n9102, n9103, n9104 );
nand U14636 ( n9103, n11510, n2007 );
nand U14637 ( n9104, n9105, n9106 );
nor U14638 ( n9106, n9107, n9108 );
not U14639 ( n626, n4878 );
nand U14640 ( n10241, n10291, n10292 );
nand U14641 ( n10291, n11263, n1909 );
nand U14642 ( n10292, n1898, n11259 );
nand U14643 ( n10244, n10289, n10290 );
nand U14644 ( n10290, n1909, n11259 );
nand U14645 ( n10289, n1898, n11263 );
and U14646 ( n4839, n4875, n4876 );
nand U14647 ( n4876, n11403, n4877 );
nand U14648 ( n4875, n4878, n11391 );
nor U14649 ( n9552, n239, n1909 );
not U14650 ( n239, n1898 );
nand U14651 ( n1889, n2693, n2694 );
nor U14652 ( n2693, n2724, n2725 );
nor U14653 ( n2694, n2695, n2696 );
nand U14654 ( n2724, n2729, n2730 );
nand U14655 ( n2695, n2704, n2705 );
nand U14656 ( n2705, n2706, n2707 );
nor U14657 ( n2704, n2714, n2715 );
nor U14658 ( n2706, n2712, n2713 );
nand U14659 ( n8055, n8095, n8096 );
nand U14660 ( n8095, n601, n8098 );
nand U14661 ( n8096, n8097, n4691 );
or U14662 ( n8097, n8098, n601 );
nand U14663 ( n4840, n4880, n4881 );
nand U14664 ( n4880, n11392, n4877 );
nand U14665 ( n4881, n4878, n11402 );
nand U14666 ( n7381, n7431, n5273 );
nand U14667 ( n7431, n7432, n7433 );
nand U14668 ( n7433, n688, n4366 );
nor U14669 ( n7432, n7434, n7435 );
nand U14670 ( n6828, n6829, n6830 );
nor U14671 ( n6829, n6839, n6840 );
nor U14672 ( n6830, n6831, n6832 );
nor U14673 ( n6839, n6780, n6783 );
nor U14674 ( n2714, n2716, n2718 );
nand U14675 ( n2718, n2719, n232 );
not U14676 ( n242, n2665 );
nor U14677 ( n9454, n9477, n9478 );
nor U14678 ( n9478, n9479, n9480 );
nand U14679 ( n9479, n9556, n9557 );
nand U14680 ( n9480, n9481, n9482 );
nor U14681 ( n9481, n3007, n9457 );
nand U14682 ( n2110, n6140, n6141 );
nor U14683 ( n6141, n6142, n6143 );
nor U14684 ( n6140, n6147, n6148 );
nor U14685 ( n6142, n607, n11379 );
not U14686 ( n601, n5020 );
nand U14687 ( n8843, n8844, n8845 );
nand U14688 ( n8844, n11508, n2029 );
nand U14689 ( n8845, n11506, n8846 );
nand U14690 ( n8846, n8847, n8848 );
nand U14691 ( n5194, n5195, n5196 );
nor U14692 ( n5195, n1002, n4885 );
xnor U14693 ( n4815, n1004, n4816 );
nand U14694 ( n2725, n2726, n2727 );
nand U14695 ( n2726, n2728, n1939 );
nand U14696 ( n2727, n351, n2703 );
nor U14697 ( n9460, n1898, n322 );
xor U14698 ( n8790, n9303, n9149 );
nand U14699 ( n9303, n9304, n9305 );
nand U14700 ( n9304, n11500, n2537 );
nand U14701 ( n9305, n2512, n9152 );
nor U14702 ( n6688, n5306, n6689 );
nor U14703 ( n6689, n6690, n6691 );
nor U14704 ( n6690, n576, n6692 );
and U14705 ( n6126, n6670, n6671 );
nor U14706 ( n6670, n6705, n6706 );
nor U14707 ( n6671, n6672, n6673 );
nor U14708 ( n6705, n6692, n6713 );
nand U14709 ( n6673, n6674, n6675 );
nand U14710 ( n6675, n6676, n4897 );
nand U14711 ( n6674, n618, n6683 );
nand U14712 ( n6676, n6677, n6678 );
nand U14713 ( n6683, n6684, n6685 );
nand U14714 ( n6685, n6686, n617 );
nor U14715 ( n6684, n6687, n6688 );
nor U14716 ( n6687, n6693, n4897 );
not U14717 ( n629, n4640 );
nor U14718 ( n6775, n6776, n6764 );
nor U14719 ( n6693, n6694, n6686 );
nor U14720 ( n6694, n4199, n7685 );
nand U14721 ( n6686, n6772, n6773 );
nor U14722 ( n6772, n6778, n6779 );
nor U14723 ( n6773, n6774, n6775 );
nor U14724 ( n6778, n6780, n6764 );
xor U14725 ( n9063, n9278, n9149 );
nand U14726 ( n9278, n9279, n9280 );
nand U14727 ( n9279, n11500, n2516 );
nand U14728 ( n9280, n2501, n11286 );
nand U14729 ( n4862, n4895, n4896 );
nand U14730 ( n4896, n11403, n4897 );
nand U14731 ( n4895, n4199, n11391 );
nand U14732 ( n10250, n10307, n10308 );
nand U14733 ( n10308, n1939, n11315 );
nand U14734 ( n10307, n1923, n11263 );
and U14735 ( n10249, n10305, n10306 );
nand U14736 ( n10305, n11263, n1939 );
nand U14737 ( n10306, n1923, n11258 );
not U14738 ( n747, n4350 );
nor U14739 ( n7892, n4580, n747 );
and U14740 ( n4861, n4898, n4899 );
nand U14741 ( n4898, n11392, n4897 );
nand U14742 ( n4899, n4199, n11402 );
not U14743 ( n762, n5064 );
nor U14744 ( n8019, n4136, n762 );
not U14745 ( n227, n1934 );
nor U14746 ( n2794, n227, n1962 );
nor U14747 ( n9482, n9483, n9484 );
nand U14748 ( n9484, n9485, n9486 );
nand U14749 ( n9486, n9487, n9488 );
nand U14750 ( n9485, n323, n2665 );
nand U14751 ( n8919, n8920, n8921 );
nand U14752 ( n8920, n11509, n2046 );
nand U14753 ( n8921, n8922, n11505 );
xnor U14754 ( n8922, n8739, n8923 );
nand U14755 ( n9062, n9281, n9282 );
nand U14756 ( n9281, n11494, n2516 );
nand U14757 ( n9282, n11500, n2501 );
xnor U14758 ( n8702, n9308, n339 );
nand U14759 ( n9308, n9309, n9310 );
nand U14760 ( n9309, n11500, n2494 );
nand U14761 ( n9310, n2471, n11286 );
not U14762 ( n119, n9457 );
nand U14763 ( n6139, n6752, n6753 );
nand U14764 ( n6753, n932, n4182 );
nor U14765 ( n6752, n6754, n6755 );
nor U14766 ( n6755, n6756, n612 );
xnor U14767 ( n4807, n4885, n4884 );
nand U14768 ( n6712, n614, n6724 );
nand U14769 ( n6724, n4807, n6725 );
nand U14770 ( n6725, n617, n4897 );
nand U14771 ( n1924, n2757, n2758 );
nand U14772 ( n2758, n2728, n1962 );
nor U14773 ( n2757, n2759, n2760 );
nor U14774 ( n2759, n2779, n228 );
nor U14775 ( n2765, n2767, n2768 );
nor U14776 ( n2767, n2687, n344 );
nor U14777 ( n2768, n19, n2769 );
nand U14778 ( n2115, n6127, n6128 );
nor U14779 ( n6128, n6129, n6130 );
nor U14780 ( n6127, n6135, n6136 );
nor U14781 ( n6129, n617, n11379 );
nor U14782 ( n2771, n2772, n2773 );
nor U14783 ( n2772, n19, n2775 );
nor U14784 ( n2773, n19, n2774 );
nand U14785 ( n1919, n1921, n1922 );
nand U14786 ( n1922, n1923, n11518 );
nand U14787 ( n1921, n11514, n1924 );
nand U14788 ( n890, n1901, n1902 );
nor U14789 ( n1902, n1903, n1904 );
nor U14790 ( n1901, n1918, n1919 );
nand U14791 ( n1904, n1906, n1907 );
not U14792 ( n234, n1923 );
nor U14793 ( n2735, n234, n1939 );
not U14794 ( n972, n4580 );
nor U14795 ( n7912, n4350, n972 );
or U14796 ( n11233, n1008, n1007 );
nand U14797 ( n4865, n4886, n4887 );
nand U14798 ( n4886, n11392, n4884 );
nand U14799 ( n4887, n4885, n11402 );
nand U14800 ( n8792, n9286, n9287 );
nand U14801 ( n9286, n11494, n2537 );
nand U14802 ( n9287, n11500, n2512 );
not U14803 ( n607, n4063 );
nor U14804 ( n5305, n4182, n607 );
and U14805 ( n6742, n6790, n6791 );
nand U14806 ( n6790, n4182, n607 );
nand U14807 ( n6791, n5303, n606 );
not U14808 ( n606, n5305 );
nand U14809 ( n4863, n4882, n4883 );
nand U14810 ( n4883, n11403, n4884 );
nand U14811 ( n4882, n4885, n11391 );
nand U14812 ( n2796, n1962, n227 );
nand U14813 ( n6678, n4807, n6679 );
nand U14814 ( n6679, n6680, n6681 );
nand U14815 ( n6681, n4199, n6682 );
not U14816 ( n971, n4344 );
not U14817 ( n619, n4885 );
nor U14818 ( n2795, n247, n1984 );
not U14819 ( n247, n1968 );
not U14820 ( n973, n4038 );
nand U14821 ( n5259, n973, n4586 );
nor U14822 ( n8022, n5064, n968 );
nand U14823 ( n5255, n8020, n8021 );
nand U14824 ( n8020, n756, n4404 );
nand U14825 ( n8021, n8022, n5265 );
nand U14826 ( n5265, n969, n4141 );
nor U14827 ( n5206, n4906, n4816 );
not U14828 ( n636, n4311 );
nand U14829 ( n2687, n2801, n2802 );
nand U14830 ( n2801, n1934, n1962 );
nand U14831 ( n2802, n2803, n2804 );
nand U14832 ( n2804, n319, n227 );
nor U14833 ( n2782, n2784, n2785 );
nor U14834 ( n2785, n2739, n2769 );
nor U14835 ( n2784, n33, n344 );
nand U14836 ( n9276, n9306, n9307 );
nand U14837 ( n9306, n11494, n2494 );
nand U14838 ( n9307, n11500, n2471 );
not U14839 ( n756, n4141 );
nor U14840 ( n2786, n2799, n2800 );
nor U14841 ( n2799, n33, n2713 );
nor U14842 ( n2800, n33, n2778 );
nand U14843 ( n9364, n2545, n348 );
nand U14844 ( n9300, n11500, n3956 );
nand U14845 ( n2105, n6152, n6153 );
nor U14846 ( n6153, n6154, n6155 );
nor U14847 ( n6152, n6159, n6160 );
nor U14848 ( n6154, n629, n11379 );
xor U14849 ( n1863, n1866, n2659 );
nand U14850 ( n2659, n2668, n2669 );
nor U14851 ( n2668, n2665, n1898 );
nand U14852 ( n2555, n2655, n2656 );
nand U14853 ( n2656, n11417, n118 );
nor U14854 ( n2655, n281, n2657 );
nor U14855 ( n2657, n2658, n1863 );
not U14856 ( n617, n4199 );
nor U14857 ( n5306, n617, n4897 );
not U14858 ( n752, n4410 );
nand U14859 ( n6847, n4640, n4056 );
and U14860 ( n4850, n4902, n4903 );
nand U14861 ( n4903, n11403, n4182 );
nand U14862 ( n4902, n4063, n11391 );
nand U14863 ( n7894, n971, n4410 );
nor U14864 ( n2770, n2776, n2777 );
nor U14865 ( n2776, n2687, n2713 );
nor U14866 ( n2777, n2687, n2778 );
nand U14867 ( n8652, n8653, n8654 );
nand U14868 ( n8653, n11508, n2074 );
nand U14869 ( n8654, n8655, n11506 );
xnor U14870 ( n8655, n8656, n8657 );
nor U14871 ( n2789, n2739, n2774 );
nand U14872 ( n4852, n4900, n4901 );
nand U14873 ( n4900, n11392, n4182 );
nand U14874 ( n4901, n4063, n11402 );
nand U14875 ( n6854, n6855, n6856 );
nand U14876 ( n6855, n6860, n6803 );
nand U14877 ( n6856, n6857, n6803 );
nor U14878 ( n6860, n6858, n6692 );
nor U14879 ( n6897, n4604, n4311 );
not U14880 ( n741, n4586 );
nand U14881 ( n5253, n741, n4038 );
nand U14882 ( n6781, n4063, n4182 );
nand U14883 ( n1876, n2667, n2659 );
nand U14884 ( n2667, n2665, n2670 );
nand U14885 ( n2670, n2669, n239 );
nand U14886 ( n2559, n2663, n2664 );
nand U14887 ( n2664, n11417, n2665 );
nor U14888 ( n2663, n281, n2666 );
nor U14889 ( n2666, n2658, n1876 );
not U14890 ( n286, n3956 );
buf U14891 ( n11307, n11306 );
not U14892 ( n967, n4693 );
nor U14893 ( n6918, n6920, n6921 );
nor U14894 ( n6920, n4739, n6788 );
nor U14895 ( n6921, n6859, n6788 );
nand U14896 ( n3024, n3063, n3064 );
nand U14897 ( n3063, n2058, n2074 );
nand U14898 ( n3064, n3065, n3066 );
nand U14899 ( n3066, n313, n266 );
nand U14900 ( n3334, n3436, n3437 );
nand U14901 ( n3436, n2226, n2204 );
nand U14902 ( n3437, n3438, n3439 );
nand U14903 ( n3438, n304, n197 );
nand U14904 ( n2847, n3022, n3023 );
nand U14905 ( n3022, n2024, n2046 );
nand U14906 ( n3023, n3024, n3025 );
nand U14907 ( n3025, n314, n272 );
nand U14908 ( n3123, n3331, n3332 );
and U14909 ( n3331, n3336, n3337 );
nand U14910 ( n3332, n3333, n3334 );
nand U14911 ( n3336, n3339, n2159 );
nand U14912 ( n3065, n3120, n3121 );
and U14913 ( n3120, n3127, n3128 );
nand U14914 ( n3121, n3122, n3123 );
nand U14915 ( n3127, n2069, n2097 );
nor U14916 ( n3943, n45, n286 );
nor U14917 ( n3744, n3747, n3748 );
nor U14918 ( n3747, n2382, n2409 );
nand U14919 ( n3748, n3749, n154 );
and U14920 ( n3639, n3741, n3742 );
nand U14921 ( n3742, n3743, n2382 );
nor U14922 ( n3741, n3744, n3745 );
nor U14923 ( n3745, n294, n3746 );
nor U14924 ( n3816, n3818, n3819 );
nor U14925 ( n3818, n3820, n3822 );
nor U14926 ( n3819, n3820, n3821 );
nor U14927 ( n3820, n2471, n2494 );
nand U14928 ( n3749, n3807, n3808 );
nand U14929 ( n3808, n3809, n2426 );
nor U14930 ( n3807, n3810, n3811 );
nor U14931 ( n3811, n292, n3812 );
nor U14932 ( n3810, n3813, n3814 );
nor U14933 ( n3813, n2426, n2447 );
nand U14934 ( n3814, n3815, n166 );
nand U14935 ( n3815, n3816, n3817 );
nand U14936 ( n3439, n3484, n3485 );
nand U14937 ( n3484, n3487, n2238 );
nand U14938 ( n3485, n3486, n2253 );
nand U14939 ( n3486, n34, n193 );
not U14940 ( n253, n1979 );
nand U14941 ( n2914, n2007, n253 );
nor U14942 ( n2691, n1939, n1923 );
nor U14943 ( n8088, n539, n967 );
nand U14944 ( n7083, n7141, n7142 );
and U14945 ( n7141, n7148, n7149 );
nand U14946 ( n7142, n7143, n7144 );
nand U14947 ( n7148, n4268, n7151 );
nor U14948 ( n7837, n7840, n7841 );
nor U14949 ( n7840, n4046, n4211 );
nand U14950 ( n7841, n7842, n742 );
nand U14951 ( n7829, n7834, n7835 );
nand U14952 ( n7835, n7836, n4046 );
nor U14953 ( n7834, n7837, n7838 );
nor U14954 ( n7838, n974, n7839 );
nor U14955 ( n2798, n318, n1968 );
nor U14956 ( n3961, n3956, n45 );
nand U14957 ( n3910, n9627, n9628 );
nand U14958 ( n9627, n168, n2537 );
or U14959 ( n9628, n9537, n3961 );
nor U14960 ( n9394, n349, n356 );
not U14961 ( n349, n9376 );
not U14962 ( n168, n2512 );
nand U14963 ( n7069, n7070, n7071 );
nor U14964 ( n7070, n7079, n7080 );
nor U14965 ( n7071, n7072, n7073 );
nor U14966 ( n7079, n6780, n7023 );
not U14967 ( n736, n4046 );
nor U14968 ( n5198, n1001, n4199 );
buf U14969 ( n11300, n11299 );
and U14970 ( n10209, n10319, n10320 );
nand U14971 ( n10319, n11262, n1962 );
nand U14972 ( n10320, n1934, n11258 );
nand U14973 ( n10210, n10321, n10322 );
nand U14974 ( n10322, n1962, n11258 );
nand U14975 ( n10321, n1934, n11263 );
nand U14976 ( n2090, n6195, n6196 );
nor U14977 ( n6196, n6197, n6198 );
nor U14978 ( n6195, n6202, n6203 );
nor U14979 ( n6197, n646, n11379 );
not U14980 ( n272, n2024 );
nor U14981 ( n9476, n272, n2046 );
nor U14982 ( n9537, n2537, n168 );
nand U14983 ( n885, n1926, n1927 );
nor U14984 ( n1927, n1928, n1929 );
nor U14985 ( n1926, n1941, n1942 );
nand U14986 ( n1929, n1931, n1932 );
not U14987 ( n646, n4102 );
or U14988 ( n5275, n7032, n11234 );
and U14989 ( n11234, n646, n4094 );
nand U14990 ( n8802, n8803, n8804 );
nand U14991 ( n8803, n11508, n2118 );
nand U14992 ( n8804, n8805, n11506 );
nor U14993 ( n8805, n8806, n8807 );
buf U14994 ( n11313, n11310 );
nand U14995 ( n2545, n9391, n353 );
nor U14996 ( n9391, n356, n359 );
nand U14997 ( n2850, n1968, n1984 );
not U14998 ( n652, n4513 );
nor U14999 ( n8750, n8751, n8752 );
nor U15000 ( n8752, n321, n8753 );
nor U15001 ( n8751, n8749, n234 );
nor U15002 ( n6954, n6958, n6959 );
nor U15003 ( n6958, n4739, n6923 );
nor U15004 ( n6959, n6859, n6923 );
nand U15005 ( n6175, n6943, n6944 );
nand U15006 ( n6944, n932, n4305 );
nor U15007 ( n6943, n6945, n6946 );
nor U15008 ( n6945, n6960, n632 );
nor U15009 ( n6950, n6952, n6953 );
nor U15010 ( n6953, n521, n6780 );
nor U15011 ( n6952, n6692, n6923 );
nand U15012 ( n6665, n1008, n1007 );
nor U15013 ( n6963, n6965, n6966 );
nor U15014 ( n6966, n6780, n6894 );
and U15015 ( n6965, n6923, n927 );
nand U15016 ( n2100, n6164, n6165 );
nor U15017 ( n6165, n6166, n6167 );
nor U15018 ( n6164, n6171, n6172 );
nor U15019 ( n6166, n636, n11379 );
buf U15020 ( n11344, n11343 );
nor U15021 ( n6831, n6776, n6783 );
nand U15022 ( n9021, n9022, n9023 );
nand U15023 ( n9022, n11509, n2097 );
nand U15024 ( n9023, n9024, n11505 );
xnor U15025 ( n9024, n9025, n9026 );
nand U15026 ( n6518, n6110, n6648 );
nand U15027 ( n6648, n624, n6649 );
not U15028 ( n277, n2069 );
nand U15029 ( n2838, n2840, n2841 );
or U15030 ( n2841, n2803, n344 );
nor U15031 ( n2840, n2842, n2843 );
nor U15032 ( n2842, n2713, n2803 );
not U15033 ( n974, n4211 );
not U15034 ( n49, n2501 );
nor U15035 ( n9524, n2516, n49 );
and U15036 ( n4859, n4890, n4891 );
nand U15037 ( n4891, n11403, n4056 );
nand U15038 ( n4890, n4640, n11391 );
buf U15039 ( n11352, n11351 );
nand U15040 ( n1992, n2928, n2929 );
nand U15041 ( n2929, n2728, n2029 );
nor U15042 ( n2928, n2930, n2931 );
nor U15043 ( n2931, n249, n2932 );
nor U15044 ( n2948, n2950, n2951 );
nor U15045 ( n2951, n2769, n2916 );
nor U15046 ( n2950, n32, n344 );
nor U15047 ( n2952, n2960, n2961 );
nor U15048 ( n2960, n32, n2713 );
nor U15049 ( n2961, n32, n2778 );
not U15050 ( n266, n2058 );
nor U15051 ( n3014, n314, n2024 );
nand U15052 ( n8937, n9269, n9270 );
nand U15053 ( n9269, n11494, n2474 );
nand U15054 ( n9270, n11500, n2459 );
nand U15055 ( n4860, n4892, n4893 );
nand U15056 ( n4892, n11392, n4056 );
nand U15057 ( n4893, n4640, n11402 );
nand U15058 ( n875, n1971, n1972 );
nor U15059 ( n1972, n1973, n1974 );
nor U15060 ( n1971, n1986, n1987 );
nand U15061 ( n1974, n1976, n1977 );
xnor U15062 ( n8935, n9266, n339 );
nand U15063 ( n9266, n9267, n9268 );
nand U15064 ( n9267, n11499, n2474 );
nand U15065 ( n9268, n2459, n9152 );
not U15066 ( n638, n4393 );
buf U15067 ( n11305, n10472 );
nand U15068 ( n3941, n2537, n2512 );
buf U15069 ( n11484, n11481 );
and U15070 ( n10211, n10224, n10225 );
nand U15071 ( n10224, n11262, n1984 );
nand U15072 ( n10225, n1968, n11259 );
not U15073 ( n259, n2013 );
nand U15074 ( n2956, n2029, n259 );
nand U15075 ( n5298, n636, n4604 );
nor U15076 ( n1861, n1866, n1867 );
nand U15077 ( n2959, n316, n2013 );
nand U15078 ( n10212, n10226, n10227 );
nand U15079 ( n10227, n1984, n11258 );
nand U15080 ( n10226, n1968, n11263 );
and U15081 ( n2669, n2754, n2753 );
nor U15082 ( n2754, n1923, n1934 );
nand U15083 ( n6850, n4393, n4305 );
nand U15084 ( n2917, n1979, n317 );
nand U15085 ( n8971, n8972, n8973 );
nand U15086 ( n8972, n11509, n2136 );
nand U15087 ( n8973, n11507, n8974 );
nand U15088 ( n8974, n8975, n8976 );
nand U15089 ( n8086, n4691, n5020 );
nand U15090 ( n5302, n997, n4311 );
nand U15091 ( n5299, n638, n4305 );
nor U15092 ( n2903, n18, n2774 );
nand U15093 ( n9117, n9202, n9203 );
nand U15094 ( n9202, n11493, n1984 );
nand U15095 ( n9203, n1968, n11498 );
nand U15096 ( n1969, n2869, n2870 );
nor U15097 ( n2870, n2871, n2872 );
nor U15098 ( n2869, n2894, n2895 );
nor U15099 ( n2871, n2713, n2889 );
nand U15100 ( n2899, n2900, n2901 );
nor U15101 ( n2900, n2904, n2905 );
nor U15102 ( n2901, n2902, n2903 );
nor U15103 ( n2904, n18, n2769 );
nand U15104 ( n9822, n9847, n769 );
nand U15105 ( n5301, n996, n4393 );
xor U15106 ( n8891, n9311, n9149 );
nand U15107 ( n9311, n9312, n9313 );
nand U15108 ( n9312, n11500, n2447 );
nand U15109 ( n9313, n2426, n9152 );
not U15110 ( n968, n4136 );
buf U15111 ( n11455, n11452 );
not U15112 ( n669, n4468 );
nand U15113 ( n7149, n7150, n4507 );
or U15114 ( n7150, n7151, n4268 );
nand U15115 ( n1964, n1966, n1967 );
nand U15116 ( n1967, n1968, n11518 );
nand U15117 ( n1966, n11513, n1969 );
nand U15118 ( n880, n1948, n1949 );
nor U15119 ( n1949, n1951, n1952 );
nor U15120 ( n1948, n1963, n1964 );
nand U15121 ( n1951, n1958, n1959 );
nor U15122 ( n6900, n6780, n6902 );
nor U15123 ( n2939, n2943, n2944 );
nor U15124 ( n2943, n2713, n2882 );
nor U15125 ( n2944, n2778, n2882 );
buf U15126 ( n11457, n11452 );
nor U15127 ( n6903, n6776, n6902 );
nand U15128 ( n6194, n6992, n6993 );
nand U15129 ( n6993, n932, n4094 );
nor U15130 ( n6992, n6994, n6995 );
nor U15131 ( n6994, n7010, n4793 );
nor U15132 ( n7003, n7007, n7008 );
nor U15133 ( n7007, n6933, n4739 );
nor U15134 ( n7008, n6933, n6859 );
xor U15135 ( n1899, n1898, n2669 );
nor U15136 ( n6999, n7001, n7002 );
and U15137 ( n7002, n6844, n926 );
nor U15138 ( n7001, n6933, n6692 );
not U15139 ( n969, n4404 );
nor U15140 ( n2909, n2910, n2911 );
nor U15141 ( n2910, n2775, n2793 );
nor U15142 ( n2911, n2774, n2793 );
nor U15143 ( n3909, n2501, n288 );
nor U15144 ( n6955, n6956, n6957 );
nor U15145 ( n6956, n521, n6777 );
nor U15146 ( n6957, n521, n6776 );
and U15147 ( n7143, n7145, n666 );
nor U15148 ( n7145, n7146, n7147 );
nor U15149 ( n7147, n4268, n4507 );
nand U15150 ( n2095, n6183, n6184 );
nor U15151 ( n6184, n6185, n6186 );
nor U15152 ( n6183, n6190, n6191 );
nor U15153 ( n6185, n638, n11379 );
nor U15154 ( n2908, n2912, n2913 );
nor U15155 ( n2912, n2769, n2793 );
nor U15156 ( n2913, n2906, n2793 );
nand U15157 ( n6130, n6131, n6132 );
nand U15158 ( n6132, n11369, n4884 );
nand U15159 ( n6131, n584, n11370 );
not U15160 ( n584, n6134 );
nand U15161 ( n2835, n2719, n2803 );
not U15162 ( n723, n4118 );
nor U15163 ( n7642, n4111, n723 );
nand U15164 ( n5300, n994, n4102 );
nor U15165 ( n3100, n3074, n2774 );
nor U15166 ( n3101, n3074, n2769 );
nand U15167 ( n8709, n8710, n8711 );
nand U15168 ( n8710, n11508, n2163 );
nand U15169 ( n8711, n8712, n11506 );
xnor U15170 ( n8712, n98, n8713 );
nand U15171 ( n1285, n8706, n8707 );
nor U15172 ( n8706, n1857, n8716 );
nor U15173 ( n8707, n8708, n8709 );
nand U15174 ( n8716, n8717, n8718 );
nand U15175 ( n865, n2016, n2017 );
nor U15176 ( n2017, n2018, n2019 );
nor U15177 ( n2016, n2031, n2032 );
nand U15178 ( n2019, n2021, n2022 );
nand U15179 ( n4163, n4164, n4165 );
nand U15180 ( n4164, n11472, n4182 );
nand U15181 ( n4165, n11471, n4166 );
nand U15182 ( n4166, n4167, n4168 );
nand U15183 ( n3822, n2516, n2501 );
nor U15184 ( n7017, n7025, n7026 );
nor U15185 ( n7025, n4739, n7009 );
nor U15186 ( n7026, n7009, n6859 );
nor U15187 ( n7013, n7015, n7016 );
nor U15188 ( n7016, n6780, n6844 );
nor U15189 ( n7015, n7009, n6692 );
not U15190 ( n731, n4217 );
nand U15191 ( n5268, n731, n4209 );
nor U15192 ( n5248, n4209, n731 );
nand U15193 ( n8058, n5064, n4136 );
nand U15194 ( n6143, n6144, n6145 );
nand U15195 ( n6145, n11369, n4897 );
nand U15196 ( n6144, n11372, n6146 );
nor U15197 ( n1916, n2669, n2751 );
and U15198 ( n2751, n1923, n2752 );
nand U15199 ( n2752, n2753, n227 );
nand U15200 ( n6522, n6110, n6654 );
nand U15201 ( n6654, n4878, n6649 );
nand U15202 ( n1894, n1896, n1897 );
nand U15203 ( n1897, n1898, n11518 );
or U15204 ( n1896, n1899, n1864 );
nand U15205 ( n2085, n6207, n6208 );
nor U15206 ( n6208, n6209, n6210 );
nor U15207 ( n6207, n6214, n6215 );
nor U15208 ( n6209, n652, n11379 );
nor U15209 ( n5280, n4507, n657 );
not U15210 ( n657, n4268 );
not U15211 ( n702, n4290 );
nor U15212 ( n5231, n4490, n702 );
nor U15213 ( n7137, n7156, n7157 );
nor U15214 ( n7156, n4739, n7044 );
nor U15215 ( n7157, n6859, n7044 );
nor U15216 ( n7133, n7135, n7136 );
nor U15217 ( n7136, n518, n6780 );
nor U15218 ( n7135, n6692, n7044 );
nand U15219 ( n1928, n1936, n1937 );
nand U15220 ( n1936, n11441, n1939 );
nand U15221 ( n1937, n11443, n1938 );
not U15222 ( n164, n2459 );
nor U15223 ( n3812, n3809, n2426 );
xnor U15224 ( n4446, n539, n11296 );
nand U15225 ( n4543, n4688, n4689 );
nand U15226 ( n4688, n4239, n4691 );
nand U15227 ( n4689, n4234, n4690 );
or U15228 ( n4690, n4691, n4239 );
nand U15229 ( n4324, n4624, n4625 );
nand U15230 ( n4624, n4628, n4327 );
nand U15231 ( n4625, n4626, n4627 );
or U15232 ( n4627, n4327, n4628 );
nor U15233 ( n4684, n4687, n4134 );
nor U15234 ( n4687, n4135, n4404 );
nor U15235 ( n4620, n4623, n4364 );
nor U15236 ( n4623, n4365, n4558 );
nor U15237 ( n4676, n4677, n4678 );
and U15238 ( n4678, n4580, n4341 );
nor U15239 ( n4677, n4343, n4579 );
nor U15240 ( n4594, n4601, n4602 );
nor U15241 ( n4601, n4639, n631 );
nor U15242 ( n4602, n4603, n4599 );
nor U15243 ( n4639, n4598, n4056 );
and U15244 ( n4095, n4609, n4610 );
or U15245 ( n4609, n4505, n4506 );
nand U15246 ( n4610, n4611, n4096 );
nand U15247 ( n4611, n4506, n4505 );
nand U15248 ( n4234, n4238, n4692 );
nand U15249 ( n4692, n4236, n4693 );
nand U15250 ( n4590, n4591, n4592 );
nand U15251 ( n4591, n11474, n4604 );
nand U15252 ( n4592, n4593, n11469 );
nor U15253 ( n4593, n4594, n4595 );
nand U15254 ( n4187, n4606, n4607 );
or U15255 ( n4606, n4092, n4095 );
nand U15256 ( n4607, n4608, n4094 );
nand U15257 ( n4608, n4095, n4092 );
nand U15258 ( n4420, n4669, n4670 );
nand U15259 ( n4669, n4207, n4210 );
nand U15260 ( n4670, n4671, n4209 );
or U15261 ( n4671, n4210, n4207 );
nand U15262 ( n4077, n4666, n4667 );
nand U15263 ( n4666, n4418, n4420 );
nand U15264 ( n4667, n4668, n4112 );
or U15265 ( n4668, n4420, n4418 );
and U15266 ( n4343, n4679, n4680 );
nand U15267 ( n4679, n4401, n4403 );
nand U15268 ( n4680, n4681, n4344 );
or U15269 ( n4681, n4403, n4401 );
and U15270 ( n4152, n4615, n4616 );
nand U15271 ( n4615, n4555, n4557 );
nand U15272 ( n4616, n4617, n4153 );
or U15273 ( n4617, n4557, n4555 );
xnor U15274 ( n4598, n923, n4640 );
nor U15275 ( n4599, n4604, n4304 );
xor U15276 ( n9093, n9316, n9149 );
nand U15277 ( n9316, n9317, n9318 );
nand U15278 ( n9317, n11500, n2429 );
nand U15279 ( n9318, n2416, n11286 );
nor U15280 ( n5279, n4268, n992 );
xnor U15281 ( n4183, n4063, n11291 );
nand U15282 ( n4192, n4056, n634 );
nand U15283 ( n7216, n4468, n4262 );
not U15284 ( n279, n2103 );
nand U15285 ( n2853, n2013, n2029 );
nand U15286 ( n7942, n4141, n4404 );
nor U15287 ( n9542, n2471, n289 );
nor U15288 ( n3853, n2474, n2459 );
nor U15289 ( n2953, n2954, n2955 );
nor U15290 ( n2954, n2775, n2916 );
nor U15291 ( n2955, n2774, n2916 );
nand U15292 ( n3886, n289, n2471 );
nor U15293 ( n4171, n4182, n611 );
nand U15294 ( n7087, n7088, n7089 );
nand U15295 ( n7088, n7092, n7045 );
nand U15296 ( n7089, n7090, n7045 );
nor U15297 ( n7092, n7093, n6692 );
not U15298 ( n712, n4532 );
and U15299 ( n5241, n724, n7639 );
nand U15300 ( n7639, n712, n4284 );
nand U15301 ( n9172, n9180, n9181 );
nand U15302 ( n9180, n11493, n2097 );
nand U15303 ( n9181, n2069, n11498 );
nor U15304 ( n2986, n2988, n2989 );
nor U15305 ( n2989, n17, n2769 );
nor U15306 ( n2988, n344, n2847 );
nand U15307 ( n7021, n4102, n4094 );
not U15308 ( n977, n4112 );
nand U15309 ( n7643, n977, n4426 );
nand U15310 ( n2059, n3088, n3089 );
nand U15311 ( n3089, n2728, n2097 );
nor U15312 ( n3088, n3090, n3091 );
nor U15313 ( n3090, n3106, n262 );
nor U15314 ( n3177, n3179, n3180 );
nor U15315 ( n3180, n2769, n3006 );
and U15316 ( n3179, n3170, n338 );
nor U15317 ( n2990, n2994, n2995 );
nor U15318 ( n2994, n2713, n2847 );
nor U15319 ( n2995, n2778, n2847 );
nand U15320 ( n8894, n9261, n9262 );
nand U15321 ( n9261, n11494, n2447 );
nand U15322 ( n9262, n11499, n2426 );
nor U15323 ( n6970, n6776, n6894 );
nand U15324 ( n2009, n2011, n2012 );
nand U15325 ( n2012, n2013, n11518 );
nand U15326 ( n2011, n11513, n2014 );
nand U15327 ( n870, n1993, n1994 );
nor U15328 ( n1994, n1996, n1997 );
nor U15329 ( n1993, n2008, n2009 );
nand U15330 ( n1996, n2003, n2004 );
and U15331 ( n8628, n8763, n8764 );
nand U15332 ( n8763, n11493, n1962 );
nand U15333 ( n8764, n1934, n11498 );
nand U15334 ( n855, n2061, n2062 );
nor U15335 ( n2062, n2063, n2064 );
nor U15336 ( n2061, n2076, n2077 );
nand U15337 ( n2064, n2066, n2067 );
nand U15338 ( n2054, n2056, n2057 );
nand U15339 ( n2057, n2058, n11518 );
nand U15340 ( n2056, n11514, n2059 );
nand U15341 ( n860, n2038, n2039 );
nor U15342 ( n2039, n2041, n2042 );
nor U15343 ( n2038, n2053, n2054 );
nand U15344 ( n2042, n2043, n2044 );
and U15345 ( n4857, n5179, n5180 );
nand U15346 ( n5180, n11402, n4604 );
nand U15347 ( n5179, n4311, n11391 );
nand U15348 ( n4050, n4051, n4052 );
nand U15349 ( n4051, n11472, n4056 );
nand U15350 ( n4052, n4053, n11469 );
xnor U15351 ( n4053, n4054, n611 );
nand U15352 ( n7081, n4513, n4096 );
not U15353 ( n978, n4111 );
nor U15354 ( n7667, n4118, n978 );
buf U15355 ( n11486, n11481 );
buf U15356 ( n11385, n11243 );
nor U15357 ( n3786, n2416, n293 );
and U15358 ( n8851, n9207, n9208 );
nand U15359 ( n9207, n11493, n2007 );
nand U15360 ( n9208, n1979, n11498 );
nand U15361 ( n4858, n5177, n5178 );
nand U15362 ( n5177, n11395, n4604 );
nand U15363 ( n5178, n4311, n11402 );
not U15364 ( n674, n4159 );
nor U15365 ( n9555, n277, n2097 );
xor U15366 ( n8613, n9321, n9149 );
nand U15367 ( n9321, n9322, n9323 );
nand U15368 ( n9322, n11500, n2409 );
nand U15369 ( n9323, n2382, n9152 );
nand U15370 ( n3817, n2494, n2471 );
buf U15371 ( n11421, n11242 );
nor U15372 ( n3785, n2426, n292 );
nand U15373 ( n3778, n292, n2426 );
nand U15374 ( n9092, n9314, n9315 );
nand U15375 ( n9314, n11494, n2429 );
nand U15376 ( n9315, n11500, n2416 );
nor U15377 ( n7839, n7836, n4046 );
nand U15378 ( n6155, n6156, n6157 );
nand U15379 ( n6156, n11369, n4182 );
nand U15380 ( n6157, n11372, n6158 );
nand U15381 ( n7938, n4344, n4410 );
not U15382 ( n728, n4426 );
nand U15383 ( n5267, n728, n4112 );
nor U15384 ( n5235, n4284, n712 );
nand U15385 ( n5242, n702, n4490 );
xnor U15386 ( n10507, n766, n764 );
nand U15387 ( n9071, n9072, n9073 );
nand U15388 ( n9072, n11509, n2187 );
nand U15389 ( n9073, n9074, n11505 );
xnor U15390 ( n9074, n9075, n9076 );
nor U15391 ( n5204, n4063, n999 );
nand U15392 ( n3781, n293, n2416 );
nand U15393 ( n3861, n291, n2459 );
nand U15394 ( n4177, n4598, n4056 );
not U15395 ( n966, n4691 );
nand U15396 ( n4132, n4544, n4136 );
and U15397 ( n10180, n10193, n10194 );
nand U15398 ( n10193, n11262, n2029 );
nand U15399 ( n10194, n2013, n11258 );
nor U15400 ( n7209, n7211, n7212 );
nor U15401 ( n7211, n7213, n6780 );
nor U15402 ( n7212, n4739, n7029 );
nor U15403 ( n7213, n7197, n667 );
nand U15404 ( n3038, n3039, n3040 );
nand U15405 ( n3039, n3044, n3042 );
nand U15406 ( n3040, n3041, n3042 );
nor U15407 ( n3044, n3043, n2774 );
and U15408 ( n3165, n3272, n3273 );
nand U15409 ( n3272, n30, n2719 );
nand U15410 ( n3273, n30, n333 );
nor U15411 ( n3071, n3043, n2769 );
not U15412 ( n184, n2382 );
nand U15413 ( n10181, n10195, n10196 );
nand U15414 ( n10196, n2029, n11259 );
nand U15415 ( n10195, n2013, n11263 );
nand U15416 ( n4376, n4377, n4378 );
nand U15417 ( n4377, n11473, n4094 );
nand U15418 ( n4378, n11470, n4379 );
nand U15419 ( n4379, n4380, n4381 );
and U15420 ( n10202, n10217, n10218 );
nand U15421 ( n10218, n2007, n11258 );
nand U15422 ( n10217, n1979, n11263 );
nor U15423 ( n2991, n2992, n2993 );
nor U15424 ( n2992, n17, n2775 );
nor U15425 ( n2993, n17, n2774 );
and U15426 ( n2753, n2865, n2864 );
nor U15427 ( n2865, n1979, n1968 );
nand U15428 ( n2080, n6219, n6220 );
nor U15429 ( n6220, n6221, n6222 );
nor U15430 ( n6219, n6226, n6227 );
nor U15431 ( n6221, n657, n11379 );
nand U15432 ( n10203, n10215, n10216 );
nand U15433 ( n10215, n11262, n2007 );
nand U15434 ( n10216, n1979, n11259 );
nor U15435 ( n3015, n258, n3017 );
not U15436 ( n258, n2977 );
nor U15437 ( n3017, n3018, n3019 );
and U15438 ( n3018, n2847, n2719 );
not U15439 ( n706, n4084 );
nor U15440 ( n5238, n4661, n706 );
nor U15441 ( n9821, n708, n9822 );
nor U15442 ( n3109, n3112, n3113 );
nor U15443 ( n3112, n31, n344 );
nor U15444 ( n3113, n2769, n3103 );
nand U15445 ( n6198, n6199, n6200 );
nand U15446 ( n6200, n11368, n4305 );
nand U15447 ( n6199, n11372, n6201 );
nor U15448 ( n3115, n3116, n3117 );
nor U15449 ( n3116, n2775, n3103 );
nor U15450 ( n3117, n2774, n3103 );
nand U15451 ( n8612, n9319, n9320 );
nand U15452 ( n9319, n11494, n2409 );
nand U15453 ( n9320, n11500, n2382 );
nand U15454 ( n7217, n4151, n4159 );
or U15455 ( n4131, n4136, n4544 );
not U15456 ( n683, n4372 );
nor U15457 ( n5295, n4558, n683 );
nand U15458 ( n1973, n1981, n1982 );
nand U15459 ( n1981, n11441, n1984 );
nand U15460 ( n1982, n11443, n1983 );
nand U15461 ( n6167, n6168, n6169 );
nand U15462 ( n6169, n11369, n4056 );
nand U15463 ( n6168, n11372, n579 );
not U15464 ( n579, n6170 );
not U15465 ( n217, n2114 );
nor U15466 ( n7883, n4038, n4586 );
nand U15467 ( n4294, n4295, n4296 );
nand U15468 ( n4295, n11472, n4305 );
nand U15469 ( n4296, n11470, n4297 );
nand U15470 ( n4297, n4298, n4299 );
nand U15471 ( n3187, n2103, n2118 );
nor U15472 ( n7218, n7168, n7220 );
nor U15473 ( n7220, n7221, n7222 );
nand U15474 ( n7222, n7223, n7224 );
nor U15475 ( n7221, n567, n6692 );
nand U15476 ( n7934, n4350, n4580 );
and U15477 ( n4930, n5183, n5184 );
nand U15478 ( n5184, n11403, n4305 );
nand U15479 ( n5183, n4393, n11391 );
nor U15480 ( n5283, n4468, n991 );
nand U15481 ( n4931, n5181, n5182 );
nand U15482 ( n5181, n11392, n4305 );
nand U15483 ( n5182, n4393, n11402 );
nand U15484 ( n5271, n991, n4468 );
nor U15485 ( n7018, n7019, n7020 );
nor U15486 ( n7019, n6777, n6844 );
nor U15487 ( n7020, n6776, n6844 );
not U15488 ( n153, n2416 );
nor U15489 ( n3746, n3743, n2382 );
nand U15490 ( n4302, n4304, n4604 );
and U15491 ( n8979, n9185, n9186 );
nand U15492 ( n9185, n11493, n2118 );
nand U15493 ( n9186, n2103, n11498 );
buf U15494 ( n11485, n11481 );
nor U15495 ( n3769, n2429, n2416 );
not U15496 ( n133, n2327 );
nand U15497 ( n2099, n2101, n2102 );
nand U15498 ( n2102, n2103, n11518 );
nand U15499 ( n2101, n11514, n2104 );
nand U15500 ( n850, n2083, n2084 );
nor U15501 ( n2084, n2086, n2087 );
nor U15502 ( n2083, n2098, n2099 );
nand U15503 ( n2086, n2093, n2094 );
nor U15504 ( n3227, n2136, n2114 );
not U15505 ( n717, n4496 );
nand U15506 ( n5232, n717, n4078 );
nand U15507 ( n3216, n3222, n3223 );
nand U15508 ( n3222, n3220, n2719 );
nand U15509 ( n3223, n3220, n333 );
nor U15510 ( n3057, n2713, n3024 );
not U15511 ( n108, n8753 );
nand U15512 ( n8901, n8902, n8903 );
nand U15513 ( n8902, n11509, n2209 );
nand U15514 ( n8903, n8904, n11505 );
nor U15515 ( n8904, n8905, n8906 );
nand U15516 ( n1240, n8898, n8899 );
nor U15517 ( n8898, n1643, n8913 );
nor U15518 ( n8899, n8900, n8901 );
nand U15519 ( n8913, n8914, n8915 );
nor U15520 ( n3738, n2382, n294 );
not U15521 ( n287, n2537 );
nor U15522 ( n7190, n7193, n7194 );
and U15523 ( n7194, n7188, n7195 );
nor U15524 ( n7193, n4808, n7196 );
or U15525 ( n7196, n6780, n7197 );
xor U15526 ( n8776, n9324, n9149 );
nand U15527 ( n9324, n9325, n9326 );
nand U15528 ( n9325, n11501, n2386 );
nand U15529 ( n9326, n2372, n11286 );
xor U15530 ( n4387, n923, n4393 );
nor U15531 ( n9601, n2136, n217 );
nand U15532 ( n3188, n3263, n3264 );
nand U15533 ( n3263, n2719, n3146 );
nand U15534 ( n3264, n333, n3146 );
nor U15535 ( n3711, n2386, n179 );
not U15536 ( n179, n2372 );
nand U15537 ( n5229, n982, n4496 );
nand U15538 ( n6186, n6187, n6188 );
nand U15539 ( n6188, n11369, n4604 );
nand U15540 ( n6187, n578, n11370 );
not U15541 ( n578, n6189 );
nor U15542 ( n5294, n4159, n989 );
xnor U15543 ( n1946, n1934, n2753 );
nor U15544 ( n5296, n4564, n988 );
nand U15545 ( n845, n2106, n2107 );
nor U15546 ( n2107, n2108, n2109 );
nor U15547 ( n2106, n2121, n2122 );
nand U15548 ( n2108, n2116, n2117 );
xnor U15549 ( n4135, n4141, n923 );
nor U15550 ( n7436, n4327, n696 );
not U15551 ( n696, n4746 );
nor U15552 ( n3674, n2359, n2338 );
nand U15553 ( n5293, n988, n4564 );
nand U15554 ( n5292, n989, n4159 );
nor U15555 ( n3118, n31, n2713 );
nand U15556 ( n11286, n8753, n9360 );
nor U15557 ( n9549, n311, n2103 );
not U15558 ( n688, n4333 );
nor U15559 ( n3181, n3189, n3190 );
nor U15560 ( n3189, n2775, n3006 );
nor U15561 ( n3190, n2774, n3006 );
xor U15562 ( n4637, n4268, n923 );
nand U15563 ( n6210, n6211, n6212 );
nand U15564 ( n6212, n11368, n4094 );
nand U15565 ( n6211, n11371, n6213 );
nor U15566 ( n1961, n2753, n2862 );
and U15567 ( n2862, n1968, n2863 );
nand U15568 ( n2863, n2864, n253 );
nand U15569 ( n3193, n2103, n311 );
and U15570 ( n10165, n10173, n10174 );
nand U15571 ( n10173, n11262, n2046 );
nand U15572 ( n10174, n2024, n11258 );
xnor U15573 ( n8833, n9347, n9149 );
nand U15574 ( n9347, n9348, n9349 );
nand U15575 ( n9348, n11501, n2299 );
nand U15576 ( n9349, n2283, n11286 );
nor U15577 ( n7254, n7255, n6776 );
nand U15578 ( n10164, n10171, n10172 );
nand U15579 ( n10172, n2046, n11258 );
nand U15580 ( n10171, n2024, n11263 );
nand U15581 ( n2075, n6231, n6232 );
nor U15582 ( n6232, n6233, n6234 );
nor U15583 ( n6231, n6238, n6239 );
nor U15584 ( n6233, n669, n11379 );
nand U15585 ( n9360, n3969, n9302 );
nand U15586 ( n8738, n9121, n9122 );
nand U15587 ( n9121, n11493, n2029 );
nand U15588 ( n9122, n2013, n11498 );
nor U15589 ( n3252, n3248, n3261 );
nor U15590 ( n3261, n3262, n3188 );
nor U15591 ( n3262, n30, n2713 );
nand U15592 ( n7155, n4564, n4153 );
nor U15593 ( n7438, n4084, n983 );
nor U15594 ( n5289, n4372, n987 );
nand U15595 ( n3050, n2719, n3024 );
not U15596 ( n173, n2338 );
nor U15597 ( n3684, n2359, n173 );
xor U15598 ( n9014, n9337, n9149 );
nand U15599 ( n9337, n9338, n9339 );
nand U15600 ( n9338, n11501, n2277 );
nand U15601 ( n9339, n2249, n11286 );
nor U15602 ( n7303, n516, n6780 );
nand U15603 ( n6254, n7293, n7294 );
nand U15604 ( n7294, n932, n4153 );
nor U15605 ( n7293, n7295, n7296 );
nor U15606 ( n7295, n7310, n4799 );
nand U15607 ( n7299, n7300, n7301 );
nand U15608 ( n7301, n903, n7208 );
nor U15609 ( n7300, n7302, n7303 );
nor U15610 ( n7302, n6692, n7276 );
nor U15611 ( n9600, n2163, n204 );
not U15612 ( n204, n2148 );
nor U15613 ( n9529, n2372, n296 );
nor U15614 ( n7304, n7308, n7309 );
nor U15615 ( n7308, n4739, n7276 );
nor U15616 ( n7309, n6859, n7276 );
nand U15617 ( n2070, n6243, n6244 );
nor U15618 ( n6244, n6245, n6246 );
nor U15619 ( n6243, n6250, n6251 );
nor U15620 ( n6245, n674, n11379 );
nand U15621 ( n8659, n9126, n9127 );
nand U15622 ( n9126, n11493, n2046 );
nand U15623 ( n9127, n2024, n11498 );
and U15624 ( n4917, n4928, n4929 );
nand U15625 ( n4929, n11403, n4094 );
nand U15626 ( n4928, n4102, n11391 );
nand U15627 ( n3096, n31, n2719 );
not U15628 ( n188, n2249 );
nand U15629 ( n8862, n8863, n8864 );
nand U15630 ( n8863, n11509, n2226 );
nand U15631 ( n8864, n11506, n8865 );
nand U15632 ( n8865, n8866, n8867 );
nand U15633 ( n5273, n986, n4333 );
xnor U15634 ( n4093, n4094, n4095 );
nand U15635 ( n4088, n4089, n4090 );
nand U15636 ( n4089, n11472, n4096 );
nand U15637 ( n4090, n4091, n11469 );
xnor U15638 ( n4091, n4092, n4093 );
not U15639 ( n288, n2516 );
nor U15640 ( n7138, n7139, n7140 );
nor U15641 ( n7139, n518, n6777 );
nor U15642 ( n7140, n518, n6776 );
nand U15643 ( n4918, n4926, n4927 );
nand U15644 ( n4926, n11392, n4094 );
nand U15645 ( n4927, n4102, n11402 );
nand U15646 ( n9028, n9131, n9132 );
nand U15647 ( n9131, n11493, n2074 );
nand U15648 ( n9132, n2058, n11498 );
nor U15649 ( n7187, n7208, n6776 );
nor U15650 ( n7072, n6776, n7023 );
nand U15651 ( n2063, n2071, n2072 );
nand U15652 ( n2071, n11440, n2074 );
nand U15653 ( n2072, n2073, n11442 );
nand U15654 ( n1175, n9217, n9218 );
nor U15655 ( n9217, n1582, n9368 );
nor U15656 ( n9218, n9219, n9220 );
nand U15657 ( n9368, n9369, n9370 );
nand U15658 ( n9220, n9221, n9222 );
nand U15659 ( n9221, n11510, n2253 );
nand U15660 ( n9222, n9223, n11505 );
xor U15661 ( n9223, n9160, n9227 );
and U15662 ( n4938, n5171, n5172 );
nand U15663 ( n5171, n11395, n4507 );
nand U15664 ( n5172, n4268, n11402 );
and U15665 ( n8832, n9345, n9346 );
nand U15666 ( n9345, n11495, n2299 );
nand U15667 ( n9346, n11501, n2283 );
nor U15668 ( n9494, n2114, n309 );
nand U15669 ( n8779, n9254, n9255 );
nand U15670 ( n9254, n11494, n2386 );
nand U15671 ( n9255, n11499, n2372 );
and U15672 ( n2864, n2974, n2973 );
nor U15673 ( n2974, n2024, n2013 );
nand U15674 ( n4939, n5169, n5170 );
nand U15675 ( n5170, n11402, n4507 );
nand U15676 ( n5169, n4268, n11391 );
nor U15677 ( n7146, n4153, n4564 );
nor U15678 ( n7245, n7270, n4739 );
xnor U15679 ( n7270, n7226, n4809 );
not U15680 ( n982, n4078 );
nor U15681 ( n3562, n2299, n2283 );
not U15682 ( n137, n2283 );
nor U15683 ( n9545, n2299, n137 );
nand U15684 ( n3389, n124, n2209 );
not U15685 ( n124, n2193 );
nand U15686 ( n9013, n9340, n9341 );
nand U15687 ( n9340, n11495, n2277 );
nand U15688 ( n9341, n11501, n2249 );
nand U15689 ( n2149, n3297, n3298 );
nand U15690 ( n3298, n2728, n2187 );
nor U15691 ( n3297, n3299, n3300 );
nor U15692 ( n3299, n3314, n201 );
nor U15693 ( n3308, n3312, n3313 );
nor U15694 ( n3312, n2713, n3123 );
nor U15695 ( n3313, n2778, n3123 );
nand U15696 ( n6222, n6223, n6224 );
nand U15697 ( n6224, n11368, n4096 );
nand U15698 ( n6223, n11371, n6225 );
buf U15699 ( n11302, n11299 );
nor U15700 ( n3702, n2338, n297 );
nor U15701 ( n7434, n4746, n984 );
nor U15702 ( n9829, n9833, n9834 );
nand U15703 ( n9834, n9835, n9836 );
nor U15704 ( n9833, n9832, n9831 );
nand U15705 ( n9836, n2277, n11259 );
and U15706 ( n9970, n9981, n9982 );
nand U15707 ( n9981, n11260, n2516 );
nand U15708 ( n9982, n2501, n11315 );
nand U15709 ( n1931, n1934, n11518 );
nand U15710 ( n8631, n8632, n8633 );
nand U15711 ( n8633, n1933, n8634 );
nand U15712 ( n8632, n11524, n1934 );
nand U15713 ( n2144, n2146, n2147 );
nand U15714 ( n2147, n11518, n2148 );
nand U15715 ( n2146, n11514, n2149 );
nand U15716 ( n840, n2128, n2129 );
nor U15717 ( n2129, n2131, n2132 );
nor U15718 ( n2128, n2143, n2144 );
nand U15719 ( n2132, n2133, n2134 );
nand U15720 ( n3647, n2386, n2372 );
nand U15721 ( n4255, n664, n4507 );
nand U15722 ( n10003, n10019, n10020 );
nand U15723 ( n10019, n11261, n2494 );
nand U15724 ( n10020, n2471, n11315 );
nand U15725 ( n9971, n9983, n9984 );
nand U15726 ( n9984, n2516, n11315 );
nand U15727 ( n9983, n11260, n2501 );
nor U15728 ( n3271, n3274, n3275 );
nor U15729 ( n3274, n14, n2769 );
nor U15730 ( n3275, n14, n2906 );
xor U15731 ( n8984, n9182, n9149 );
nand U15732 ( n9182, n9183, n9184 );
nand U15733 ( n9183, n11499, n2136 );
nand U15734 ( n9184, n2114, n9152 );
and U15735 ( n10002, n10021, n10022 );
nand U15736 ( n10022, n2494, n11315 );
nand U15737 ( n10021, n11261, n2471 );
nand U15738 ( n10162, n10182, n10183 );
nand U15739 ( n10183, n2074, n11259 );
nand U15740 ( n10182, n2058, n11263 );
nand U15741 ( n9947, n9974, n9975 );
nand U15742 ( n9974, n11260, n2537 );
nand U15743 ( n9975, n2512, n11315 );
nor U15744 ( n3276, n3279, n3280 );
nor U15745 ( n3279, n14, n2775 );
nor U15746 ( n3280, n14, n2774 );
and U15747 ( n9946, n9972, n9973 );
nand U15748 ( n9973, n2537, n11315 );
nand U15749 ( n9972, n11260, n2512 );
xor U15750 ( n4092, n4102, n923 );
nand U15751 ( n4247, n4248, n4249 );
nand U15752 ( n4248, n11472, n4262 );
nand U15753 ( n4249, n4250, n11469 );
nor U15754 ( n4250, n4251, n4252 );
nor U15755 ( n9495, n2148, n308 );
nor U15756 ( n3317, n3319, n3320 );
nor U15757 ( n3320, n2769, n3282 );
and U15758 ( n3319, n3123, n2719 );
not U15759 ( n976, n4209 );
nor U15760 ( n7784, n4209, n4217 );
not U15761 ( n291, n2474 );
not U15762 ( n289, n2494 );
not U15763 ( n197, n2204 );
nand U15764 ( n9152, n8753, n9360 );
not U15765 ( n293, n2429 );
nand U15766 ( n9960, n10036, n10037 );
nand U15767 ( n10036, n11261, n2447 );
nand U15768 ( n10037, n2426, n11315 );
not U15769 ( n209, n2159 );
nand U15770 ( n3325, n209, n2187 );
nand U15771 ( n7376, n7377, n4558 );
nand U15772 ( n7377, n683, n7378 );
nor U15773 ( n10727, n827, n11302 );
not U15774 ( n827, n2431 );
nor U15775 ( n9944, n9948, n9949 );
nor U15776 ( n9948, n45, n9951 );
nor U15777 ( n9949, n9950, n11258 );
and U15778 ( n9950, n9951, n286 );
nand U15779 ( n8951, n9249, n9250 );
nand U15780 ( n9249, n11494, n2359 );
nand U15781 ( n9250, n11499, n2338 );
nand U15782 ( n10161, n10168, n10169 );
nand U15783 ( n10168, n11262, n2074 );
nand U15784 ( n10169, n2058, n11258 );
xnor U15785 ( n8949, n9246, n339 );
nand U15786 ( n9246, n9247, n9248 );
nand U15787 ( n9247, n11499, n2359 );
nand U15788 ( n9248, n2338, n11286 );
nor U15789 ( n9508, n2316, n144 );
not U15790 ( n144, n2294 );
nand U15791 ( n6266, n7346, n7347 );
nand U15792 ( n7347, n932, n4558 );
nor U15793 ( n7346, n7348, n7349 );
nor U15794 ( n7348, n7361, n4798 );
nor U15795 ( n3640, n2386, n2372 );
nand U15796 ( n4500, n4501, n4502 );
nand U15797 ( n4501, n11473, n4507 );
nand U15798 ( n4502, n4503, n11469 );
xor U15799 ( n4503, n4504, n4505 );
xnor U15800 ( n8912, n9163, n339 );
nand U15801 ( n9163, n9164, n9165 );
nand U15802 ( n9164, n11499, n2187 );
nand U15803 ( n9165, n2159, n9152 );
and U15804 ( n9959, n10038, n10039 );
nand U15805 ( n10039, n2447, n11315 );
nand U15806 ( n10038, n11261, n2426 );
nand U15807 ( n2065, n6255, n6256 );
nor U15808 ( n6256, n6257, n6258 );
nor U15809 ( n6255, n6262, n6263 );
nor U15810 ( n6257, n678, n11380 );
not U15811 ( n292, n2447 );
nand U15812 ( n2018, n2026, n2027 );
nand U15813 ( n2026, n11440, n2029 );
nand U15814 ( n2027, n11443, n2028 );
nand U15815 ( n3328, n307, n2159 );
nor U15816 ( n4579, n4580, n4341 );
nand U15817 ( n9962, n10006, n10007 );
nand U15818 ( n10006, n11261, n2474 );
nand U15819 ( n10007, n2459, n11315 );
nand U15820 ( n8993, n8994, n8995 );
nand U15821 ( n8994, n11509, n2299 );
nand U15822 ( n8995, n8996, n11505 );
nor U15823 ( n8996, n8997, n8998 );
nand U15824 ( n1210, n8990, n8991 );
nor U15825 ( n8990, n1544, n9015 );
nor U15826 ( n8991, n8992, n8993 );
nand U15827 ( n9015, n9016, n9017 );
and U15828 ( n4919, n4934, n4935 );
nand U15829 ( n4935, n11403, n4096 );
nand U15830 ( n4934, n4513, n11392 );
nand U15831 ( n2109, n2111, n2112 );
nand U15832 ( n2111, n11518, n2114 );
nand U15833 ( n2112, n11443, n2113 );
nor U15834 ( n3602, n2294, n299 );
nand U15835 ( n4920, n4936, n4937 );
nand U15836 ( n4936, n11392, n4096 );
nand U15837 ( n4937, n4513, n11402 );
or U15838 ( n4283, n4490, n4279 );
nand U15839 ( n8714, n9175, n9176 );
nand U15840 ( n9175, n11493, n2136 );
nand U15841 ( n9176, n11499, n2114 );
nand U15842 ( n3133, n2163, n2148 );
nand U15843 ( n835, n2151, n2152 );
nor U15844 ( n2152, n2153, n2154 );
nor U15845 ( n2151, n2166, n2167 );
nand U15846 ( n2153, n2161, n2162 );
nand U15847 ( n3357, n3363, n3364 );
nand U15848 ( n3363, n3369, n2719 );
nand U15849 ( n3364, n3361, n333 );
nor U15850 ( n3369, n3370, n3366 );
and U15851 ( n9961, n10004, n10005 );
nand U15852 ( n10005, n2474, n11315 );
nand U15853 ( n10004, n11260, n2459 );
nor U15854 ( n4675, n4211, n4037 );
nand U15855 ( n5140, n5167, n5168 );
nand U15856 ( n5167, n11395, n4262 );
nand U15857 ( n5168, n4468, n11402 );
buf U15858 ( n11312, n11310 );
nor U15859 ( n9509, n2283, n301 );
nand U15860 ( n6234, n6235, n6236 );
nand U15861 ( n6236, n11368, n4507 );
nand U15862 ( n6235, n11371, n6237 );
nand U15863 ( n3231, n3232, n3233 );
nand U15864 ( n3232, n2728, n2136 );
nand U15865 ( n3233, n3221, n352 );
nand U15866 ( n3421, n3422, n3423 );
nand U15867 ( n3423, n2719, n3334 );
nor U15868 ( n3422, n3424, n3425 );
nor U15869 ( n3424, n29, n2713 );
nand U15870 ( n8638, n8639, n8640 );
nand U15871 ( n8639, n11508, n2277 );
nand U15872 ( n8640, n8641, n11506 );
xnor U15873 ( n8641, n8642, n8643 );
xor U15874 ( n8870, n9148, n9149 );
nand U15875 ( n9148, n9150, n9151 );
nand U15876 ( n9150, n11498, n2209 );
nand U15877 ( n9151, n2193, n11286 );
xor U15878 ( n8679, n9327, n9149 );
nand U15879 ( n9327, n9328, n9329 );
nand U15880 ( n9328, n11501, n2342 );
nand U15881 ( n9329, n2327, n9152 );
xor U15882 ( n9011, n9342, n9149 );
nand U15883 ( n9342, n9343, n9344 );
nand U15884 ( n9343, n11501, n2316 );
nand U15885 ( n9344, n2294, n9152 );
nand U15886 ( n2189, n2191, n2192 );
nand U15887 ( n2192, n11519, n2193 );
nand U15888 ( n2191, n11514, n2194 );
nand U15889 ( n830, n2173, n2174 );
nor U15890 ( n2174, n2176, n2177 );
nor U15891 ( n2173, n2188, n2189 );
nand U15892 ( n2177, n2178, n2179 );
nor U15893 ( n9612, n2277, n188 );
xor U15894 ( n9075, n9166, n9149 );
nand U15895 ( n9166, n9167, n9168 );
nand U15896 ( n9167, n11499, n2163 );
nand U15897 ( n9168, n2148, n11286 );
nor U15898 ( n3446, n2204, n304 );
nand U15899 ( n3644, n2342, n2327 );
nor U15900 ( n3467, n3447, n2774 );
nand U15901 ( n3433, n3464, n3465 );
nor U15902 ( n3464, n3469, n3470 );
nor U15903 ( n3465, n3466, n3467 );
nor U15904 ( n3469, n3447, n2769 );
nor U15905 ( n3428, n3429, n3430 );
nor U15906 ( n3430, n2713, n3334 );
nor U15907 ( n3429, n3416, n3431 );
nor U15908 ( n3431, n3432, n3433 );
nand U15909 ( n5139, n5173, n5174 );
nand U15910 ( n5174, n11402, n4262 );
nand U15911 ( n5173, n4468, n11391 );
nor U15912 ( n3324, n2774, n3282 );
xnor U15913 ( n1991, n1979, n2864 );
nand U15914 ( n4455, n532, n4456 );
xnor U15915 ( n4456, n4262, n4457 );
nand U15916 ( n4450, n4451, n4452 );
nand U15917 ( n4451, n11473, n4151 );
nand U15918 ( n4452, n11470, n4453 );
nand U15919 ( n4453, n4454, n4455 );
and U15920 ( n9717, n10143, n10144 );
nand U15921 ( n10144, n2118, n11259 );
nand U15922 ( n10143, n2103, n11263 );
or U15923 ( n4699, n4078, n4489 );
nand U15924 ( n3337, n3338, n2187 );
nand U15925 ( n3338, n209, n122 );
and U15926 ( n9705, n10150, n10151 );
nand U15927 ( n10151, n2097, n11259 );
nand U15928 ( n10150, n2069, n11263 );
nand U15929 ( n3381, n306, n2193 );
nor U15930 ( n7410, n4366, n4333 );
and U15931 ( n9723, n9768, n9769 );
nand U15932 ( n9769, n2163, n11258 );
nand U15933 ( n9768, n11263, n2148 );
nand U15934 ( n9724, n9770, n9771 );
nand U15935 ( n9770, n11263, n2163 );
nand U15936 ( n9771, n2148, n11258 );
or U15937 ( n4035, n4038, n4575 );
nand U15938 ( n9146, n9161, n9162 );
nand U15939 ( n9161, n11493, n2187 );
nand U15940 ( n9162, n11498, n2159 );
nand U15941 ( n9718, n10141, n10142 );
nand U15942 ( n10141, n11262, n2118 );
nand U15943 ( n10142, n2103, n11259 );
nand U15944 ( n9706, n10152, n10153 );
nand U15945 ( n10152, n11262, n2097 );
nand U15946 ( n10153, n2069, n11259 );
xnor U15947 ( n4808, n4268, n4507 );
nand U15948 ( n2060, n6267, n6268 );
nor U15949 ( n6268, n6269, n6270 );
nor U15950 ( n6267, n6274, n6275 );
nor U15951 ( n6269, n683, n11380 );
nor U15952 ( n2006, n2864, n2971 );
and U15953 ( n2971, n2013, n2972 );
nand U15954 ( n2972, n2973, n272 );
nand U15955 ( n7378, n4366, n4333 );
not U15956 ( n983, n4661 );
not U15957 ( n87, n9302 );
nand U15958 ( n9012, n9335, n9336 );
nand U15959 ( n9335, n11495, n2316 );
nand U15960 ( n9336, n11501, n2294 );
nand U15961 ( n4459, n4149, n4151 );
nand U15962 ( n8869, n9153, n9154 );
nand U15963 ( n9153, n11493, n2209 );
nand U15964 ( n9154, n11499, n2193 );
nand U15965 ( n8825, n8826, n8827 );
nand U15966 ( n8826, n11508, n2316 );
nand U15967 ( n8827, n11506, n8828 );
nand U15968 ( n8828, n8829, n8830 );
xor U15969 ( n8642, n9350, n9149 );
nand U15970 ( n9350, n9351, n9352 );
nand U15971 ( n9351, n11501, n2253 );
nand U15972 ( n9352, n2238, n9152 );
xnor U15973 ( n4150, n4151, n4152 );
nand U15974 ( n6246, n6247, n6248 );
nand U15975 ( n6248, n11368, n4262 );
nand U15976 ( n6247, n11371, n6249 );
nand U15977 ( n4145, n4146, n4147 );
nand U15978 ( n4146, n11472, n4153 );
nand U15979 ( n4147, n11471, n4148 );
xor U15980 ( n4148, n4149, n4150 );
nand U15981 ( n3539, n2316, n2294 );
or U15982 ( n7365, n7144, n6780 );
or U15983 ( n7367, n7144, n6776 );
and U15984 ( n2973, n3086, n3085 );
nor U15985 ( n3086, n2058, n2069 );
nor U15986 ( n3388, n2238, n303 );
nand U15987 ( n4031, n4575, n4038 );
nand U15988 ( n4282, n4279, n4490 );
nor U15989 ( n10709, n807, n11302 );
not U15990 ( n807, n2387 );
nand U15991 ( n3482, n303, n2238 );
nand U15992 ( n10035, n10055, n10056 );
nand U15993 ( n10055, n11261, n2429 );
nand U15994 ( n10056, n2416, n11315 );
and U15995 ( n10034, n10057, n10058 );
nand U15996 ( n10058, n2429, n11315 );
nand U15997 ( n10057, n11261, n2416 );
not U15998 ( n294, n2409 );
nand U15999 ( n9036, n9037, n9038 );
nand U16000 ( n9037, n11509, n2342 );
nand U16001 ( n9038, n9039, n11505 );
xnor U16002 ( n9039, n9011, n9040 );
nand U16003 ( n1200, n9033, n9034 );
nor U16004 ( n9033, n1482, n9041 );
nor U16005 ( n9034, n9035, n9036 );
nand U16006 ( n9041, n9042, n9043 );
nand U16007 ( n7648, n4532, n4284 );
and U16008 ( n9713, n9725, n9726 );
nand U16009 ( n9725, n11261, n2136 );
nand U16010 ( n9726, n2114, n11259 );
nor U16011 ( n3368, n2209, n2193 );
nand U16012 ( n9866, n9921, n9922 );
nand U16013 ( n9921, n11260, n2359 );
nand U16014 ( n9922, n2338, n11258 );
nor U16015 ( n4461, n4151, n4149 );
nand U16016 ( n9877, n9899, n9900 );
nand U16017 ( n9899, n11260, n2386 );
nand U16018 ( n9900, n2372, n11259 );
nand U16019 ( n9880, n9901, n9902 );
nand U16020 ( n9902, n2386, n11315 );
nand U16021 ( n9901, n11260, n2372 );
not U16022 ( n772, n9913 );
nand U16023 ( n9714, n9728, n9729 );
nand U16024 ( n9729, n2136, n11258 );
nand U16025 ( n9728, n11263, n2114 );
nand U16026 ( n8682, n9241, n9242 );
nand U16027 ( n9241, n11494, n2342 );
nand U16028 ( n9242, n11499, n2327 );
nor U16029 ( n3527, n2249, n302 );
nor U16030 ( n3532, n2316, n2294 );
and U16031 ( n5131, n5164, n5165 );
nand U16032 ( n5165, n11402, n4153 );
nand U16033 ( n5164, n11395, n4564 );
xor U16034 ( n9160, n9353, n9149 );
nand U16035 ( n9353, n9358, n9359 );
nand U16036 ( n9358, n11498, n2226 );
nand U16037 ( n9359, n2204, n11286 );
nor U16038 ( n4664, n4661, n4071 );
nand U16039 ( n9078, n9139, n9140 );
nand U16040 ( n9139, n11493, n2163 );
nand U16041 ( n9140, n11498, n2148 );
nand U16042 ( n3536, n2277, n2249 );
nand U16043 ( n2217, n3458, n3459 );
nand U16044 ( n3459, n2728, n2253 );
nor U16045 ( n3458, n3460, n3461 );
nor U16046 ( n3461, n3456, n3462 );
and U16047 ( n9865, n9923, n9924 );
nand U16048 ( n9924, n2359, n11315 );
nand U16049 ( n9923, n11260, n2338 );
nand U16050 ( n5130, n5162, n5163 );
nand U16051 ( n5162, n11395, n4153 );
nand U16052 ( n5163, n11402, n4564 );
nand U16053 ( n825, n2196, n2197 );
nor U16054 ( n2197, n2198, n2199 );
nor U16055 ( n2196, n2211, n2212 );
nand U16056 ( n2198, n2206, n2207 );
not U16057 ( n298, n2342 );
nand U16058 ( n4325, n4322, n4366 );
xnor U16059 ( n4365, n4372, n923 );
not U16060 ( n984, n4327 );
not U16061 ( n193, n2238 );
nand U16062 ( n4944, n5143, n5144 );
nand U16063 ( n5144, n11404, n4151 );
nand U16064 ( n5143, n11395, n4159 );
nand U16065 ( n10073, n10091, n10092 );
nand U16066 ( n10092, n2299, n11315 );
nand U16067 ( n10091, n11261, n2283 );
not U16068 ( n678, n4564 );
not U16069 ( n979, n4284 );
nand U16070 ( n1976, n1979, n11518 );
nand U16071 ( n8856, n8857, n8858 );
nand U16072 ( n8858, n1978, n8634 );
nand U16073 ( n8857, n11524, n1979 );
and U16074 ( n10072, n10093, n10094 );
nand U16075 ( n10093, n11262, n2299 );
nand U16076 ( n10094, n2283, n11315 );
nand U16077 ( n4029, n4037, n4211 );
nand U16078 ( n4946, n5141, n5142 );
nand U16079 ( n5141, n11395, n4151 );
nand U16080 ( n5142, n11404, n4159 );
buf U16081 ( n11301, n11299 );
nand U16082 ( n9872, n9884, n9885 );
nand U16083 ( n9884, n11260, n2409 );
nand U16084 ( n9885, n2382, n11315 );
nand U16085 ( n4485, n4521, n4284 );
nand U16086 ( n7523, n4084, n4661 );
or U16087 ( n4326, n4366, n4322 );
nor U16088 ( n3444, n3418, n2769 );
nor U16089 ( n3417, n3418, n2774 );
nand U16090 ( n4551, n4552, n4553 );
nand U16091 ( n4552, n11473, n4558 );
nand U16092 ( n4553, n11470, n4554 );
xor U16093 ( n4554, n4555, n4556 );
nand U16094 ( n9748, n9757, n9758 );
nand U16095 ( n9757, n11263, n2187 );
nand U16096 ( n9758, n2159, n11258 );
nand U16097 ( n8645, n9233, n9234 );
nand U16098 ( n9233, n11494, n2253 );
nand U16099 ( n9234, n11499, n2238 );
nand U16100 ( n1864, n2536, n11513 );
nand U16101 ( n2539, n11410, n356 );
nand U16102 ( n1878, n81, n2547 );
nand U16103 ( n2547, n2548, n2539 );
nand U16104 ( n2548, n2549, n111 );
nor U16105 ( n2549, n2551, n2552 );
nand U16106 ( n2176, n2183, n2184 );
nand U16107 ( n2183, n11440, n2187 );
nand U16108 ( n2184, n2186, n11521 );
nand U16109 ( n2266, n2273, n2274 );
nand U16110 ( n2273, n11440, n2277 );
nand U16111 ( n2274, n2276, n11521 );
nand U16112 ( n2398, n2406, n2407 );
nand U16113 ( n2406, n11439, n2409 );
nand U16114 ( n2407, n2408, n11521 );
nand U16115 ( n2486, n2491, n2492 );
nand U16116 ( n2491, n11439, n2494 );
nand U16117 ( n2492, n2493, n11521 );
and U16118 ( n9873, n9886, n9887 );
nand U16119 ( n9887, n2409, n11259 );
nand U16120 ( n9886, n11260, n2382 );
not U16121 ( n296, n2386 );
nand U16122 ( n775, n2418, n2419 );
nor U16123 ( n2419, n2421, n2422 );
nor U16124 ( n2418, n2432, n2433 );
nand U16125 ( n2421, n2427, n2428 );
nand U16126 ( n815, n2241, n2242 );
nor U16127 ( n2242, n2243, n2244 );
nor U16128 ( n2241, n2256, n2257 );
nand U16129 ( n2243, n2251, n2252 );
nand U16130 ( n795, n2329, n2331 );
nor U16131 ( n2331, n2332, n2333 );
nor U16132 ( n2329, n2344, n2346 );
nand U16133 ( n2332, n2339, n2341 );
nand U16134 ( n805, n2286, n2287 );
nor U16135 ( n2287, n2288, n2289 );
nor U16136 ( n2286, n2301, n2302 );
nand U16137 ( n2288, n2296, n2297 );
nand U16138 ( n1867, n2534, n11513 );
nand U16139 ( n2021, n2024, n11518 );
nand U16140 ( n2066, n2069, n11518 );
nand U16141 ( n2154, n2156, n2157 );
nand U16142 ( n2156, n11519, n2159 );
nand U16143 ( n2157, n2158, n11442 );
nand U16144 ( n9159, n9228, n9229 );
nand U16145 ( n9228, n11494, n2226 );
nand U16146 ( n9229, n11499, n2204 );
nand U16147 ( n6258, n6259, n6260 );
nand U16148 ( n6260, n11368, n4151 );
nand U16149 ( n6259, n11371, n6261 );
nand U16150 ( n2422, n2423, n2424 );
nand U16151 ( n2424, n22, n11442 );
nand U16152 ( n2423, n11519, n2426 );
nand U16153 ( n2378, n2379, n2381 );
nand U16154 ( n2381, n23, n11442 );
nand U16155 ( n2379, n11519, n2382 );
nand U16156 ( n2323, n2324, n2326 );
nand U16157 ( n2324, n11514, n2328 );
nand U16158 ( n2326, n11519, n2327 );
nand U16159 ( n2412, n2413, n2414 );
nand U16160 ( n2413, n11514, n2417 );
nand U16161 ( n2414, n11519, n2416 );
nand U16162 ( n2368, n2369, n2371 );
nand U16163 ( n2369, n11514, n2373 );
nand U16164 ( n2371, n11519, n2372 );
nand U16165 ( n2333, n2334, n2336 );
nand U16166 ( n2336, n2337, n11442 );
nand U16167 ( n2334, n11519, n2338 );
nand U16168 ( n2234, n2236, n2237 );
nand U16169 ( n2236, n11514, n2239 );
nand U16170 ( n2237, n11519, n2238 );
nand U16171 ( n2279, n2281, n2282 );
nand U16172 ( n2281, n11514, n2284 );
nand U16173 ( n2282, n11519, n2283 );
nand U16174 ( n2289, n2291, n2292 );
nand U16175 ( n2292, n11434, n2293 );
nand U16176 ( n2291, n11519, n2294 );
nand U16177 ( n2244, n2246, n2247 );
nand U16178 ( n2247, n2248, n11442 );
nand U16179 ( n2246, n11519, n2249 );
nand U16180 ( n2199, n2201, n2202 );
nand U16181 ( n2202, n11435, n2203 );
nand U16182 ( n2201, n11519, n2204 );
nand U16183 ( n9745, n9755, n9756 );
nand U16184 ( n9756, n2187, n11258 );
nand U16185 ( n9755, n11263, n2159 );
nand U16186 ( n765, n2462, n2463 );
nor U16187 ( n2463, n2464, n2466 );
nor U16188 ( n2462, n2476, n2477 );
nand U16189 ( n2464, n2472, n2473 );
nand U16190 ( n4632, n4071, n4661 );
not U16191 ( n981, n4490 );
nand U16192 ( n2507, n2508, n2509 );
nand U16193 ( n2509, n11442, n2511 );
nand U16194 ( n2508, n11520, n2512 );
nand U16195 ( n2456, n2457, n2458 );
nand U16196 ( n2457, n11514, n2461 );
nand U16197 ( n2458, n11520, n2459 );
nand U16198 ( n2497, n2498, n2499 );
nand U16199 ( n2498, n11515, n2502 );
nand U16200 ( n2499, n11520, n2501 );
nand U16201 ( n2466, n2467, n2468 );
nand U16202 ( n2468, n11443, n2469 );
nand U16203 ( n2467, n11520, n2471 );
nand U16204 ( n2055, n6279, n6280 );
nor U16205 ( n6280, n6281, n6282 );
nor U16206 ( n6279, n6286, n6287 );
nor U16207 ( n6281, n688, n11380 );
nor U16208 ( n4488, n4284, n4521 );
nand U16209 ( n4480, n4489, n4078 );
nand U16210 ( n8675, n8676, n8677 );
nand U16211 ( n8676, n11508, n2359 );
nand U16212 ( n8677, n8678, n11506 );
xnor U16213 ( n8678, n8679, n8680 );
nand U16214 ( n3873, n3921, n45 );
nor U16215 ( n3921, n2512, n2501 );
nand U16216 ( n3294, n3400, n197 );
nor U16217 ( n3400, n3401, n2193 );
nand U16218 ( n3499, n3585, n137 );
nor U16219 ( n3585, n3586, n2294 );
nand U16220 ( n3723, n3797, n153 );
nor U16221 ( n3797, n3798, n2426 );
nand U16222 ( n3798, n3872, n164 );
nor U16223 ( n3872, n3873, n2471 );
nand U16224 ( n3662, n3722, n179 );
nor U16225 ( n3722, n3723, n2382 );
nand U16226 ( n3401, n3498, n193 );
nor U16227 ( n3498, n3499, n2249 );
nand U16228 ( n3205, n3293, n204 );
nor U16229 ( n3293, n3294, n2159 );
and U16230 ( n3085, n3204, n217 );
nor U16231 ( n3204, n2103, n3205 );
nand U16232 ( n3586, n3661, n173 );
nor U16233 ( n3661, n3662, n2327 );
nand U16234 ( n7480, n4746, n4327 );
nand U16235 ( n9868, n10113, n10114 );
nand U16236 ( n10114, n2342, n11259 );
nand U16237 ( n10113, n11262, n2327 );
nand U16238 ( n2050, n6291, n6292 );
nor U16239 ( n6292, n6293, n6294 );
nor U16240 ( n6291, n6298, n6299 );
nor U16241 ( n6293, n696, n11380 );
buf U16242 ( n11345, n11343 );
nand U16243 ( n9867, n10075, n10076 );
nand U16244 ( n10075, n11261, n2342 );
nand U16245 ( n10076, n2327, n11315 );
nand U16246 ( n9858, n10080, n10081 );
nand U16247 ( n10080, n11261, n2316 );
nand U16248 ( n10081, n2294, n11315 );
not U16249 ( n297, n2359 );
nor U16250 ( n10691, n809, n11302 );
not U16251 ( n809, n2343 );
not U16252 ( n986, n4366 );
nand U16253 ( n3375, n3376, n3377 );
nand U16254 ( n3376, n2728, n2209 );
nand U16255 ( n3377, n352, n3362 );
nand U16256 ( n2239, n3502, n3503 );
nand U16257 ( n3503, n2728, n2277 );
nor U16258 ( n3502, n3504, n3505 );
nor U16259 ( n3505, n191, n3506 );
buf U16260 ( n11304, n10472 );
nand U16261 ( n9855, n10078, n10079 );
nand U16262 ( n10079, n2316, n11315 );
nand U16263 ( n10078, n11261, n2294 );
buf U16264 ( n11353, n11351 );
xnor U16265 ( n2036, n2024, n2973 );
nand U16266 ( n6270, n6271, n6272 );
nand U16267 ( n6272, n11368, n4153 );
nand U16268 ( n6271, n562, n11370 );
not U16269 ( n562, n6273 );
and U16270 ( n5128, n5160, n5161 );
nand U16271 ( n5161, n11404, n4558 );
nand U16272 ( n5160, n11395, n4372 );
nand U16273 ( n5127, n5158, n5159 );
nand U16274 ( n5158, n11395, n4558 );
nand U16275 ( n5159, n11404, n4372 );
buf U16276 ( n11308, n11306 );
nand U16277 ( n4487, n4523, n4524 );
nand U16278 ( n4523, n4526, n4111 );
or U16279 ( n4524, n536, n4525 );
nand U16280 ( n4472, n4473, n4474 );
nand U16281 ( n4473, n11473, n4490 );
nand U16282 ( n4474, n4475, n11469 );
nor U16283 ( n4475, n4476, n4477 );
nor U16284 ( n2051, n2973, n3083 );
and U16285 ( n3083, n2058, n3084 );
nand U16286 ( n3084, n3085, n277 );
not U16287 ( n987, n4558 );
nand U16288 ( n4354, n4355, n4356 );
nand U16289 ( n4355, n11473, n4366 );
nand U16290 ( n4356, n4357, n11469 );
nor U16291 ( n4357, n4358, n4359 );
or U16292 ( n3520, n3385, n2769 );
nand U16293 ( n8945, n8946, n8947 );
nand U16294 ( n8946, n11509, n2386 );
nand U16295 ( n8947, n8948, n11505 );
xor U16296 ( n8948, n8949, n8950 );
nand U16297 ( n1225, n8942, n8943 );
nor U16298 ( n8942, n1413, n8953 );
nor U16299 ( n8943, n8944, n8945 );
nand U16300 ( n8953, n8954, n8955 );
not U16301 ( n302, n2277 );
nand U16302 ( n2045, n6311, n6312 );
nor U16303 ( n6312, n6313, n6314 );
nor U16304 ( n6311, n6318, n6319 );
nor U16305 ( n6313, n706, n11380 );
or U16306 ( n3522, n3385, n2774 );
not U16307 ( n299, n2316 );
nor U16308 ( n10655, n814, n11301 );
not U16309 ( n814, n2254 );
nand U16310 ( n9531, n9532, n9516 );
nor U16311 ( n9532, n9535, n9536 );
nor U16312 ( n9536, n287, n2512 );
nor U16313 ( n9535, n9537, n9538 );
nand U16314 ( n4703, n4704, n938 );
nor U16315 ( n4704, n951, n929 );
nand U16316 ( n4654, n4655, n4656 );
nand U16317 ( n4655, n11474, n4661 );
nand U16318 ( n4656, n11470, n4657 );
xor U16319 ( n4657, n4628, n4658 );
nor U16320 ( n10673, n812, n11301 );
not U16321 ( n812, n2293 );
nand U16322 ( n2284, n3592, n3593 );
nand U16323 ( n3593, n2728, n2316 );
nor U16324 ( n3592, n3594, n3595 );
nor U16325 ( n3595, n3596, n3597 );
and U16326 ( n9741, n10128, n10129 );
nand U16327 ( n10128, n11262, n2209 );
nand U16328 ( n10129, n2193, n11259 );
nor U16329 ( n4525, n4111, n4526 );
nand U16330 ( n9740, n10126, n10127 );
nand U16331 ( n10127, n2209, n11259 );
nand U16332 ( n10126, n11262, n2193 );
nand U16333 ( n4272, n4273, n4274 );
nand U16334 ( n4273, n11472, n4284 );
nand U16335 ( n4274, n11470, n4275 );
nand U16336 ( n4275, n4276, n4277 );
nor U16337 ( n5287, n5289, n5290 );
nor U16338 ( n5290, n986, n4333 );
nand U16339 ( n4315, n4316, n4317 );
nand U16340 ( n4316, n11473, n4327 );
nand U16341 ( n4317, n11470, n4318 );
nand U16342 ( n4318, n4319, n4320 );
nand U16343 ( n5036, n5057, n5058 );
nand U16344 ( n5057, n11393, n4038 );
nand U16345 ( n5058, n11403, n4586 );
nand U16346 ( n4968, n4998, n4999 );
nand U16347 ( n4998, n5017, n5015 );
nand U16348 ( n4999, n5000, n5001 );
nor U16349 ( n5017, n602, n5014 );
nand U16350 ( n4955, n4956, n4957 );
nor U16351 ( n4956, n5113, n5114 );
or U16352 ( n4957, n4952, n4951 );
and U16353 ( n5114, n4661, n11391 );
nand U16354 ( n6282, n6283, n6284 );
nand U16355 ( n6284, n11368, n4558 );
nand U16356 ( n6283, n11371, n6285 );
nand U16357 ( n8661, n8662, n8663 );
nand U16358 ( n8663, n2023, n8634 );
nand U16359 ( n8662, n11524, n2024 );
nand U16360 ( n5033, n5043, n5044 );
nand U16361 ( n5043, n11393, n4580 );
nand U16362 ( n5044, n11403, n4350 );
nand U16363 ( n2022, n11435, n2023 );
nand U16364 ( n1977, n11435, n1978 );
nand U16365 ( n2067, n11435, n2068 );
nand U16366 ( n2161, n11435, n2164 );
nand U16367 ( n2251, n11434, n2254 );
nand U16368 ( n2427, n11434, n2431 );
nand U16369 ( n2339, n11434, n2343 );
nand U16370 ( n2116, n11435, n2119 );
nand U16371 ( n2377, n2383, n2384 );
nand U16372 ( n2384, n11439, n2386 );
nand U16373 ( n2383, n11434, n2387 );
not U16374 ( n991, n4262 );
and U16375 ( n5037, n5059, n5060 );
nand U16376 ( n5059, n11393, n4586 );
nand U16377 ( n5060, n11403, n4038 );
and U16378 ( n5034, n5045, n5046 );
nand U16379 ( n5045, n11393, n4350 );
nand U16380 ( n5046, n11403, n4580 );
nand U16381 ( n1932, n11435, n1933 );
not U16382 ( n301, n2299 );
and U16383 ( n9803, n9807, n9808 );
nand U16384 ( n9807, n11263, n2253 );
nand U16385 ( n9808, n2238, n11259 );
xnor U16386 ( n4522, n4487, n4284 );
nand U16387 ( n4517, n4518, n4519 );
nand U16388 ( n4518, n11473, n4111 );
nand U16389 ( n4519, n11470, n4520 );
xnor U16390 ( n4520, n4521, n4522 );
not U16391 ( n989, n4151 );
not U16392 ( n988, n4153 );
nand U16393 ( n9831, n9837, n9838 );
nand U16394 ( n9837, n11263, n2277 );
nand U16395 ( n9838, n2249, n11259 );
nand U16396 ( n9804, n9809, n9810 );
nand U16397 ( n9810, n2253, n11259 );
nand U16398 ( n9809, n11263, n2238 );
and U16399 ( n5134, n5154, n5155 );
nand U16400 ( n5155, n11404, n4366 );
nand U16401 ( n5154, n11395, n4333 );
nand U16402 ( n6334, n7598, n7599 );
nand U16403 ( n7599, n932, n4490 );
nor U16404 ( n7598, n7600, n7601 );
nor U16405 ( n7601, n7359, n556 );
nand U16406 ( n8772, n8773, n8774 );
nand U16407 ( n8773, n11508, n2409 );
nand U16408 ( n8774, n8775, n11506 );
xnor U16409 ( n8775, n8776, n8777 );
nand U16410 ( n4981, n5055, n5056 );
nand U16411 ( n5056, n11403, n4217 );
nand U16412 ( n5055, n11393, n4209 );
nand U16413 ( n2040, n6323, n6324 );
nor U16414 ( n6324, n6325, n6326 );
nor U16415 ( n6323, n6330, n6331 );
nor U16416 ( n6325, n717, n11380 );
and U16417 ( n4980, n5053, n5054 );
nand U16418 ( n5053, n11393, n4217 );
nand U16419 ( n5054, n11403, n4209 );
nand U16420 ( n4067, n4068, n4069 );
nand U16421 ( n4068, n11472, n4078 );
nand U16422 ( n4069, n11469, n4070 );
xor U16423 ( n4070, n4071, n4072 );
and U16424 ( n9752, n9787, n9788 );
nand U16425 ( n9787, n11263, n2226 );
nand U16426 ( n9788, n2204, n11259 );
nor U16427 ( n3551, n2774, n3568 );
xnor U16428 ( n3568, n3526, n3560 );
nand U16429 ( n9753, n9789, n9790 );
nand U16430 ( n9790, n2226, n11259 );
nand U16431 ( n9789, n11263, n2204 );
and U16432 ( n4978, n5030, n5031 );
nand U16433 ( n5030, n11393, n4211 );
nand U16434 ( n5031, n11403, n4046 );
nand U16435 ( n5133, n5152, n5153 );
nand U16436 ( n5152, n11395, n4366 );
nand U16437 ( n5153, n11404, n4333 );
nand U16438 ( n6294, n6295, n6296 );
nand U16439 ( n6296, n11368, n4366 );
nand U16440 ( n6295, n11371, n6297 );
nand U16441 ( n9835, n11263, n2249 );
and U16442 ( n5051, n5079, n5080 );
nand U16443 ( n5080, n11404, n4426 );
nand U16444 ( n5079, n11394, n4112 );
nor U16445 ( n2096, n3085, n3202 );
and U16446 ( n3202, n2103, n3203 );
nand U16447 ( n3203, n217, n44 );
xnor U16448 ( n4110, n4111, n536 );
nand U16449 ( n6346, n7633, n7634 );
nand U16450 ( n7634, n932, n4284 );
nor U16451 ( n7633, n7635, n7636 );
nor U16452 ( n7636, n7359, n6341 );
nand U16453 ( n4106, n4107, n4108 );
nand U16454 ( n4107, n11472, n4112 );
nand U16455 ( n4108, n11471, n4109 );
xnor U16456 ( n4109, n722, n4110 );
xnor U16457 ( n2081, n2069, n3085 );
nand U16458 ( n4977, n5028, n5029 );
nand U16459 ( n5029, n11403, n4211 );
nand U16460 ( n5028, n11392, n4046 );
nand U16461 ( n2035, n6335, n6336 );
nor U16462 ( n6336, n6337, n6338 );
nor U16463 ( n6335, n6342, n6343 );
nor U16464 ( n6337, n702, n11380 );
nand U16465 ( n4996, n5039, n5040 );
nand U16466 ( n5039, n11393, n4410 );
nand U16467 ( n5040, n11403, n4344 );
not U16468 ( n304, n2226 );
nand U16469 ( n5052, n5081, n5082 );
nand U16470 ( n5081, n11394, n4426 );
nand U16471 ( n5082, n11404, n4112 );
nand U16472 ( n5093, n5101, n5102 );
nand U16473 ( n5101, n11394, n4490 );
nand U16474 ( n5102, n11404, n4290 );
nand U16475 ( n4997, n5047, n5048 );
nand U16476 ( n5048, n11403, n4410 );
nand U16477 ( n5047, n11393, n4344 );
nand U16478 ( n8597, n8598, n8599 );
nand U16479 ( n8598, n11508, n2429 );
nand U16480 ( n8599, n8600, n11505 );
nor U16481 ( n8600, n8601, n8602 );
nand U16482 ( n1315, n8594, n8595 );
nor U16483 ( n8594, n1383, n8615 );
nor U16484 ( n8595, n8596, n8597 );
nand U16485 ( n8615, n8616, n8617 );
and U16486 ( n5092, n5103, n5104 );
nand U16487 ( n5104, n11404, n4490 );
nand U16488 ( n5103, n11394, n4290 );
nor U16489 ( n10637, n787, n11301 );
not U16490 ( n787, n2203 );
and U16491 ( n4988, n5069, n5070 );
nand U16492 ( n5069, n11394, n4404 );
nand U16493 ( n5070, n11404, n4141 );
xnor U16494 ( n2126, n2114, n44 );
nor U16495 ( n2141, n44, n3291 );
and U16496 ( n3291, n2148, n3292 );
nand U16497 ( n3292, n209, n43 );
nor U16498 ( n5004, n4741, n598 );
not U16499 ( n598, n5008 );
nand U16500 ( n4990, n5065, n5066 );
nand U16501 ( n5066, n11404, n4136 );
nand U16502 ( n5065, n11393, n5064 );
nand U16503 ( n4993, n5062, n5063 );
nand U16504 ( n5062, n11393, n4136 );
nand U16505 ( n5063, n11403, n5064 );
nand U16506 ( n4989, n5067, n5068 );
nand U16507 ( n5068, n11404, n4404 );
nand U16508 ( n5067, n11393, n4141 );
nand U16509 ( n2030, n6347, n6348 );
nor U16510 ( n6348, n6349, n6350 );
nor U16511 ( n6347, n6354, n6355 );
nor U16512 ( n6349, n712, n11380 );
not U16513 ( n992, n4507 );
not U16514 ( n303, n2253 );
nand U16515 ( n6314, n6315, n6316 );
nand U16516 ( n6316, n11368, n4327 );
nand U16517 ( n6315, n11371, n6317 );
not U16518 ( n993, n4096 );
nand U16519 ( n5089, n5099, n5100 );
nand U16520 ( n5100, n11404, n4284 );
nand U16521 ( n5099, n11394, n4532 );
nand U16522 ( n9085, n9086, n9087 );
nand U16523 ( n9086, n11509, n2447 );
nand U16524 ( n9087, n11507, n9088 );
nand U16525 ( n9088, n9089, n9090 );
nand U16526 ( n5088, n5105, n5106 );
nand U16527 ( n5105, n11394, n4284 );
nand U16528 ( n5106, n11404, n4532 );
nand U16529 ( n8819, n8820, n8821 );
nand U16530 ( n8821, n2068, n8634 );
nand U16531 ( n8820, n11524, n2069 );
xnor U16532 ( n4419, n4420, n4112 );
nand U16533 ( n4414, n4415, n4416 );
nand U16534 ( n4415, n11473, n4209 );
nand U16535 ( n4416, n11470, n4417 );
xnor U16536 ( n4417, n4418, n4419 );
nor U16537 ( n2186, n43, n3398 );
and U16538 ( n3398, n2193, n3399 );
nand U16539 ( n3399, n197, n42 );
nand U16540 ( n4702, n929, n4705 );
buf U16541 ( n11456, n11452 );
nand U16542 ( n5588, n5926, n5927 );
nand U16543 ( n5927, n5928, n5929 );
nand U16544 ( n5926, n5936, n868 );
nand U16545 ( n5929, n5930, n5931 );
nand U16546 ( n5830, n5875, n5876 );
nand U16547 ( n5876, n5877, n5878 );
nand U16548 ( n5875, n5885, n891 );
nand U16549 ( n5878, n5879, n5880 );
not U16550 ( n857, n5461 );
nand U16551 ( n5714, n5899, n5900 );
nand U16552 ( n5900, n5901, n5902 );
nand U16553 ( n5899, n5909, n879 );
nand U16554 ( n5902, n5903, n5904 );
not U16555 ( n849, n5794 );
not U16556 ( n854, n5558 );
nand U16557 ( n5858, n5865, n5864 );
nand U16558 ( n5865, n5863, n5871 );
nand U16559 ( n5871, n897, n5861 );
not U16560 ( n964, n5869 );
nand U16561 ( n5016, n5071, n5072 );
nand U16562 ( n5071, n11394, n4691 );
nand U16563 ( n5072, n11404, n5020 );
not U16564 ( n306, n2209 );
and U16565 ( n5015, n5018, n5019 );
nand U16566 ( n5019, n11403, n4691 );
nand U16567 ( n5018, n11392, n5020 );
and U16568 ( n5096, n5109, n5110 );
nand U16569 ( n5110, n11404, n4078 );
nand U16570 ( n5109, n11394, n4496 );
nand U16571 ( n6326, n6327, n6328 );
nand U16572 ( n6327, n11368, n4661 );
nand U16573 ( n6328, n11371, n6329 );
nand U16574 ( n5097, n5107, n5108 );
nand U16575 ( n5107, n11394, n4078 );
nand U16576 ( n5108, n11404, n4496 );
nand U16577 ( n2025, n6359, n6360 );
nor U16578 ( n6360, n6361, n6362 );
nor U16579 ( n6359, n6366, n6367 );
nor U16580 ( n6361, n723, n11380 );
nand U16581 ( n8887, n8888, n8889 );
nand U16582 ( n8888, n11509, n2474 );
nand U16583 ( n8889, n8890, n11505 );
xnor U16584 ( n8890, n8891, n8892 );
nand U16585 ( n1245, n8884, n8885 );
nor U16586 ( n8884, n1323, n8895 );
nor U16587 ( n8885, n8886, n8887 );
nand U16588 ( n8895, n8896, n8897 );
and U16589 ( n5115, n5148, n5149 );
nand U16590 ( n5148, n11395, n4327 );
nand U16591 ( n5149, n11404, n4746 );
not U16592 ( n307, n2187 );
nand U16593 ( n5116, n5150, n5151 );
nand U16594 ( n5151, n11404, n4327 );
nand U16595 ( n5150, n11393, n4746 );
nand U16596 ( n6338, n6339, n6340 );
nand U16597 ( n6340, n11368, n4078 );
nand U16598 ( n6339, n554, n11370 );
not U16599 ( n554, n6341 );
or U16600 ( n11235, n939, n938 );
not U16601 ( n312, n2097 );
nor U16602 ( n2231, n42, n3496 );
and U16603 ( n3496, n2238, n3497 );
nand U16604 ( n3497, n188, n41 );
nand U16605 ( n6382, n7765, n7766 );
nand U16606 ( n7766, n932, n4209 );
nor U16607 ( n7765, n7767, n7768 );
nor U16608 ( n7768, n7359, n553 );
nand U16609 ( n5078, n5084, n5085 );
nand U16610 ( n5085, n11404, n4118 );
nand U16611 ( n5084, n11394, n4111 );
not U16612 ( n311, n2118 );
nor U16613 ( n10619, n789, n11301 );
not U16614 ( n789, n2164 );
and U16615 ( n5077, n5090, n5091 );
nand U16616 ( n5090, n11394, n4118 );
nand U16617 ( n5091, n11404, n4111 );
xnor U16618 ( n4208, n4209, n4210 );
nand U16619 ( n4203, n4204, n4205 );
nand U16620 ( n4204, n11472, n4211 );
nand U16621 ( n4205, n11470, n4206 );
xnor U16622 ( n4206, n4207, n4208 );
nand U16623 ( n2020, n6371, n6372 );
nor U16624 ( n6372, n6373, n6374 );
nor U16625 ( n6371, n6378, n6379 );
nor U16626 ( n6373, n728, n11380 );
not U16627 ( n309, n2136 );
nand U16628 ( n4952, n5111, n5112 );
nand U16629 ( n5112, n11404, n4661 );
nand U16630 ( n5111, n11394, n4084 );
nor U16631 ( n10572, n794, n11300 );
not U16632 ( n794, n2068 );
not U16633 ( n851, n5764 );
not U16634 ( n997, n4604 );
nand U16635 ( n2044, n11440, n2046 );
nand U16636 ( n2162, n11440, n2163 );
nand U16637 ( n2341, n11439, n2342 );
nand U16638 ( n2252, n11440, n2253 );
nand U16639 ( n2473, n11439, n2474 );
nand U16640 ( n2428, n11439, n2429 );
nand U16641 ( n2134, n11440, n2136 );
nand U16642 ( n2117, n11440, n2118 );
nand U16643 ( n2514, n11439, n2516 );
not U16644 ( n994, n4094 );
nand U16645 ( n2093, n11440, n2097 );
nand U16646 ( n2206, n11440, n2209 );
nand U16647 ( n2296, n11439, n2299 );
nand U16648 ( n1907, n11441, n1909 );
buf U16649 ( n11311, n11310 );
nand U16650 ( n2003, n11441, n2007 );
nand U16651 ( n1958, n11441, n1962 );
nand U16652 ( n8931, n8932, n8933 );
nand U16653 ( n8932, n11509, n2494 );
nand U16654 ( n8933, n8934, n11505 );
xor U16655 ( n8934, n8935, n8936 );
nand U16656 ( n6350, n6351, n6352 );
nand U16657 ( n6352, n11367, n4490 );
nand U16658 ( n6351, n11371, n6353 );
not U16659 ( n998, n4056 );
nor U16660 ( n10590, n792, n11301 );
not U16661 ( n792, n2119 );
not U16662 ( n308, n2163 );
nor U16663 ( n6513, n11402, n6515 );
nand U16664 ( n6111, n942, n6505 );
nand U16665 ( n6505, n6506, n4748 );
nand U16666 ( n6506, n6507, n952 );
not U16667 ( n952, n6508 );
buf U16668 ( n11370, n11373 );
nand U16669 ( n6442, n6443, n6444 );
nand U16670 ( n6443, n11367, n4580 );
nand U16671 ( n6444, n11370, n6445 );
buf U16672 ( n11371, n11373 );
nand U16673 ( n6490, n6491, n6492 );
nand U16674 ( n6491, n11367, n4691 );
nand U16675 ( n6492, n11371, n6493 );
nand U16676 ( n6466, n6467, n6468 );
nand U16677 ( n6467, n11367, n4404 );
nand U16678 ( n6468, n11370, n6469 );
nand U16679 ( n6398, n6399, n6400 );
nand U16680 ( n6399, n11367, n4209 );
nand U16681 ( n6400, n11371, n6401 );
nand U16682 ( n6478, n6479, n6480 );
nand U16683 ( n6480, n11367, n4136 );
nand U16684 ( n6479, n11370, n6481 );
nand U16685 ( n6454, n6455, n6456 );
nand U16686 ( n6456, n11367, n4344 );
nand U16687 ( n6455, n11370, n6457 );
nand U16688 ( n6374, n6375, n6376 );
nand U16689 ( n6376, n11367, n4111 );
nand U16690 ( n6375, n11370, n6377 );
nand U16691 ( n6422, n6423, n6424 );
nand U16692 ( n6424, n11367, n4038 );
nand U16693 ( n6423, n11370, n6425 );
nand U16694 ( n6386, n6387, n6388 );
nand U16695 ( n6388, n11367, n4112 );
nand U16696 ( n6387, n11370, n6389 );
nand U16697 ( n6410, n6411, n6412 );
nand U16698 ( n6412, n11367, n4211 );
nand U16699 ( n6411, n11370, n6413 );
nand U16700 ( n6362, n6363, n6364 );
nand U16701 ( n6364, n11367, n4284 );
nand U16702 ( n6363, n11371, n6365 );
buf U16703 ( n11372, n11373 );
nand U16704 ( n4036, n4577, n4578 );
nand U16705 ( n4577, n4341, n4580 );
or U16706 ( n4578, n4579, n4343 );
nand U16707 ( n4021, n4022, n4023 );
nand U16708 ( n4022, n11472, n4038 );
nand U16709 ( n4023, n4024, n11469 );
nor U16710 ( n4024, n4025, n4026 );
nand U16711 ( n8798, n81, n9396 );
nand U16712 ( n9396, n2539, n9397 );
nand U16713 ( n9397, n9225, n2534 );
nand U16714 ( n8896, n11525, n2426 );
nand U16715 ( n8616, n11524, n2382 );
nand U16716 ( n9042, n11525, n2294 );
nand U16717 ( n1290, n8686, n8687 );
nor U16718 ( n8687, n8688, n8689 );
nor U16719 ( n8686, n1232, n8703 );
nor U16720 ( n8688, n291, n11320 );
nand U16721 ( n8876, n11525, n2193 );
nand U16722 ( n8684, n11524, n2327 );
nand U16723 ( n8781, n11524, n2372 );
nand U16724 ( n9097, n11525, n2416 );
nand U16725 ( n8940, n11525, n2459 );
nand U16726 ( n8717, n11524, n2114 );
nand U16727 ( n9016, n11525, n2249 );
nand U16728 ( n8647, n11524, n2238 );
nand U16729 ( n8838, n11524, n2283 );
nand U16730 ( n8914, n11525, n2159 );
nand U16731 ( n9080, n11525, n2148 );
nand U16732 ( n8954, n11525, n2338 );
nor U16733 ( n2276, n41, n3583 );
and U16734 ( n3583, n2283, n3584 );
nand U16735 ( n3584, n144, n40 );
nand U16736 ( n7913, n7990, n7991 );
nand U16737 ( n7990, n752, n4344 );
nand U16738 ( n7991, n552, n7894 );
nand U16739 ( n9369, n11526, n2204 );
not U16740 ( n313, n2074 );
xnor U16741 ( n5829, n896, n5830 );
not U16742 ( n996, n4305 );
buf U16743 ( n11303, n10472 );
nand U16744 ( n6106, n11480, n4745 );
or U16745 ( n5787, n5763, n11236 );
and U16746 ( n11236, n5790, n5764 );
nor U16747 ( n6489, n539, n11379 );
nand U16748 ( n4156, n11465, n4159 );
nand U16749 ( n4568, n4569, n4570 );
nand U16750 ( n4569, n11473, n4580 );
nand U16751 ( n4570, n11469, n4571 );
nand U16752 ( n4571, n4572, n4573 );
nor U16753 ( n2321, n40, n3659 );
and U16754 ( n3659, n2327, n3660 );
nand U16755 ( n3660, n173, n39 );
nand U16756 ( n5762, n5763, n5764 );
nand U16757 ( n8689, n8690, n8691 );
nand U16758 ( n8690, n11508, n2516 );
nand U16759 ( n8691, n8692, n11506 );
nor U16760 ( n8692, n8693, n8694 );
not U16761 ( n314, n2046 );
nand U16762 ( n2461, n3875, n3876 );
nand U16763 ( n3876, n2728, n2494 );
nor U16764 ( n3875, n3877, n3878 );
and U16765 ( n3878, n331, n2453 );
nand U16766 ( n5934, n5928, n5554 );
nor U16767 ( n3972, n3961, n9540 );
buf U16768 ( n11333, n11334 );
nand U16769 ( n4337, n4338, n4339 );
nand U16770 ( n4338, n11473, n4344 );
nand U16771 ( n4339, n11470, n4340 );
xnor U16772 ( n4340, n4341, n4342 );
nor U16773 ( n10554, n797, n11301 );
not U16774 ( n797, n2023 );
nand U16775 ( n4561, n11465, n4564 );
nor U16776 ( n2364, n39, n3720 );
and U16777 ( n3720, n2372, n3721 );
nand U16778 ( n3721, n184, n38 );
nand U16779 ( n2482, n3896, n3897 );
nand U16780 ( n3897, n2728, n2516 );
nor U16781 ( n3896, n3898, n3899 );
and U16782 ( n3899, n331, n2469 );
not U16783 ( n999, n4182 );
nand U16784 ( n6450, n8013, n8014 );
nand U16785 ( n8014, n932, n4404 );
nor U16786 ( n8013, n8015, n8016 );
nor U16787 ( n8015, n7685, n8023 );
not U16788 ( n112, n9401 );
nand U16789 ( n9445, n113, n114 );
xor U16790 ( n8791, n8792, n8793 );
not U16791 ( n162, n2471 );
nand U16792 ( n2455, n4394, n4395 );
nor U16793 ( n4394, n4405, n4406 );
nor U16794 ( n4395, n4396, n4397 );
nand U16795 ( n4406, n4407, n4408 );
nand U16796 ( n4397, n4398, n4399 );
nand U16797 ( n4398, n11473, n4404 );
nand U16798 ( n4399, n11470, n4400 );
xor U16799 ( n4400, n4401, n4402 );
xor U16800 ( n1247, n8967, n46 );
xnor U16801 ( n8967, n339, n7 );
nor U16802 ( n2408, n38, n3795 );
and U16803 ( n3795, n2416, n3796 );
nand U16804 ( n3796, n158, n37 );
nor U16805 ( n3937, n2713, n3922 );
not U16806 ( n316, n2029 );
buf U16807 ( n11309, n11306 );
xnor U16808 ( n5733, n887, n5734 );
not U16809 ( n317, n2007 );
nand U16810 ( n4369, n11465, n4372 );
nor U16811 ( n10536, n799, n11300 );
not U16812 ( n799, n1978 );
nand U16813 ( n6462, n8047, n8048 );
nand U16814 ( n8048, n932, n4136 );
nor U16815 ( n8047, n8049, n8050 );
nor U16816 ( n8049, n7685, n8057 );
not U16817 ( n318, n1984 );
nand U16818 ( n4776, n4780, n504 );
not U16819 ( n504, n4781 );
nor U16820 ( n2452, n37, n3870 );
and U16821 ( n3870, n2459, n3871 );
nand U16822 ( n3871, n162, n36 );
buf U16823 ( n11346, n11343 );
nand U16824 ( n4122, n4123, n4124 );
nand U16825 ( n4123, n11472, n4136 );
nand U16826 ( n4124, n4125, n11469 );
nor U16827 ( n4125, n4126, n4127 );
nand U16828 ( n2515, n4119, n4120 );
nor U16829 ( n4119, n4137, n4138 );
nor U16830 ( n4120, n4121, n4122 );
nand U16831 ( n4138, n4139, n4140 );
nand U16832 ( n2523, n3954, n3955 );
nand U16833 ( n3955, n2728, n3956 );
nor U16834 ( n3954, n3957, n3958 );
nor U16835 ( n3957, n334, n3960 );
xnor U16836 ( n3960, n3961, n3962 );
xnor U16837 ( n3962, n168, n2537 );
buf U16838 ( n11397, n11390 );
nor U16839 ( n8966, n45, n8798 );
buf U16840 ( n11354, n11351 );
nor U16841 ( n9574, n323, n324 );
not U16842 ( n1001, n4897 );
nand U16843 ( n4330, n11465, n4333 );
or U16844 ( n5678, n5654, n11237 );
and U16845 ( n11237, n5681, n5655 );
nor U16846 ( n2493, n36, n3919 );
and U16847 ( n3919, n2501, n3920 );
nand U16848 ( n3920, n45, n168 );
nand U16849 ( n2652, n10809, n328 );
nor U16850 ( n10809, n11534, n87 );
nand U16851 ( n5653, n5654, n5655 );
nand U16852 ( n4039, n4714, n4712 );
nor U16853 ( n4714, n4715, n4716 );
nand U16854 ( n2445, n4436, n4437 );
nor U16855 ( n4436, n4441, n4442 );
nor U16856 ( n4437, n4438, n4439 );
nor U16857 ( n4442, n539, n4243 );
xor U16858 ( n6481, n4780, n8098 );
nand U16859 ( n6486, n8120, n8121 );
nand U16860 ( n8121, n932, n4693 );
nor U16861 ( n8120, n8122, n8123 );
nor U16862 ( n8122, n7685, n8124 );
not U16863 ( n158, n2426 );
nor U16864 ( n10518, n802, n11300 );
not U16865 ( n802, n1933 );
not U16866 ( n321, n1939 );
nand U16867 ( n5975, n6038, n6039 );
nand U16868 ( n6038, n6041, n6040 );
nand U16869 ( n6039, n942, n6040 );
nor U16870 ( n6041, n11282, n946 );
not U16871 ( n914, n4739 );
nand U16872 ( n6512, n5315, n6637 );
nand U16873 ( n6637, n914, n938 );
nand U16874 ( n5907, n5901, n5681 );
xnor U16875 ( n2522, n2512, n45 );
not U16876 ( n322, n1909 );
not U16877 ( n319, n1962 );
nor U16878 ( n6660, n1149, n11338 );
not U16879 ( n1004, n4906 );
not U16880 ( n937, n5439 );
nor U16881 ( n2672, n341, n356 );
nor U16882 ( n2551, n9376, n329 );
nand U16883 ( n4719, n11465, n4746 );
not U16884 ( n1003, n4877 );
nand U16885 ( n4081, n11464, n4084 );
and U16886 ( n11238, n9375, n11533 );
nor U16887 ( n3967, n45, n3968 );
nor U16888 ( n3968, n11491, n11417 );
nand U16889 ( n6632, n8133, n8134 );
nor U16890 ( n8134, n8135, n8136 );
nor U16891 ( n8133, n8139, n6504 );
nor U16892 ( n8136, n539, n11468 );
nand U16893 ( n6504, n8140, n8141 );
nand U16894 ( n8141, n6493, n6837 );
nand U16895 ( n8140, n4781, n6682 );
nor U16896 ( n5404, n859, n5419 );
nand U16897 ( n6493, n8098, n8143 );
nand U16898 ( n8143, n539, n4693 );
not U16899 ( n947, n4730 );
nand U16900 ( n4744, n8284, n946 );
nor U16901 ( n8284, n11282, n947 );
nand U16902 ( n4287, n11465, n4290 );
not U16903 ( n11429, n2556 );
nand U16904 ( n2556, n2650, n2651 );
nor U16905 ( n2650, n111, n2652 );
nand U16906 ( n5315, n6495, n6515 );
nand U16907 ( n5608, n5609, n877 );
not U16908 ( n877, n5610 );
nor U16909 ( n5609, n5589, n5611 );
nor U16910 ( n5611, n5590, n853 );
not U16911 ( n856, n5528 );
nand U16912 ( n4493, n11465, n4496 );
not U16913 ( n11389, n5318 );
nand U16914 ( n5318, n5976, n946 );
nor U16915 ( n5976, n11282, n4730 );
nand U16916 ( n5607, n5612, n5610 );
nor U16917 ( n5612, n5590, n5615 );
nor U16918 ( n5615, n5589, n5588 );
nor U16919 ( n6037, n11459, n1009 );
nor U16920 ( n1203, n9375, n1325 );
nand U16921 ( n1229, n284, n10808 );
nand U16922 ( n1325, n10815, n11533 );
nand U16923 ( n10815, n10816, n11420 );
nand U16924 ( n10816, n328, n10825 );
nand U16925 ( n10825, n329, n9302 );
nand U16926 ( n10801, n10810, n71 );
nor U16927 ( n10810, n11534, n328 );
nor U16928 ( n11285, n1253, n10800 );
not U16929 ( n933, n6040 );
buf U16930 ( n11413, n11244 );
nand U16931 ( n4529, n11464, n4532 );
nand U16932 ( n1194, n282, n10808 );
nand U16933 ( n4044, n4722, n4646 );
nor U16934 ( n4722, n4723, n4724 );
nor U16935 ( n4723, n4744, n4650 );
nor U16936 ( n4724, n11282, n4649 );
nand U16937 ( n4728, n4729, n4730 );
nand U16938 ( n4729, n11402, n4731 );
nand U16939 ( n4731, n929, n907 );
nor U16940 ( n1187, n1253, n10800 );
or U16941 ( n5551, n5527, n11239 );
and U16942 ( n11239, n5554, n5528 );
nand U16943 ( n4734, n8183, n6643 );
nor U16944 ( n8183, n953, n951 );
nand U16945 ( n5582, n5587, n5588 );
or U16946 ( n5587, n5589, n5590 );
nor U16947 ( n10794, n409, n1229 );
nor U16948 ( n1662, n359, n1229 );
nor U16949 ( n1647, n361, n1229 );
nor U16950 ( n1586, n366, n1229 );
nor U16951 ( n1548, n369, n1229 );
nor U16952 ( n1501, n378, n1229 );
nor U16953 ( n1486, n374, n1229 );
nor U16954 ( n1468, n387, n1229 );
nor U16955 ( n1417, n382, n1229 );
nor U16956 ( n1402, n388, n1229 );
nor U16957 ( n1387, n389, n1229 );
nor U16958 ( n1327, n393, n1229 );
nor U16959 ( n1207, n407, n1229 );
not U16960 ( n948, n4716 );
nor U16961 ( n9225, n2552, n111 );
nand U16962 ( n8795, n9365, n9366 );
nor U16963 ( n9365, n284, n109 );
nor U16964 ( n11284, n1253, n10800 );
not U16965 ( n1002, n4884 );
not U16966 ( n928, n6642 );
not U16967 ( n56, n1462 );
nand U16968 ( n1379, n1346, n1347 );
not U16969 ( n54, n1477 );
nand U16970 ( n1766, n51, n361 );
not U16971 ( n51, n1772 );
nand U16972 ( n4748, n6499, n929 );
nand U16973 ( n5526, n5527, n5528 );
not U16974 ( n11362, n6519 );
nand U16975 ( n6519, n6633, n6634 );
nor U16976 ( n6634, n6635, n6636 );
nor U16977 ( n6633, n4744, n6508 );
not U16978 ( n61, n1524 );
not U16979 ( n63, n1441 );
nand U16980 ( n1367, n1337, n1338 );
nand U16981 ( n1673, n58, n361 );
not U16982 ( n58, n1679 );
nor U16983 ( n6636, n953, n6512 );
nand U16984 ( n4042, n11464, n4046 );
nand U16985 ( n4139, n11465, n4141 );
nand U16986 ( n4115, n11465, n4118 );
nand U16987 ( n4583, n11464, n4586 );
nand U16988 ( n4347, n11465, n4350 );
nand U16989 ( n4407, n11465, n4410 );
nand U16990 ( n4214, n11465, n4217 );
nand U16991 ( n4423, n11465, n4426 );
buf U16992 ( n11321, n11318 );
nand U16993 ( n5883, n5877, n5790 );
nor U16994 ( n9386, n341, n359 );
nand U16995 ( n9113, n9224, n9225 );
nor U16996 ( n9224, n9226, n2652 );
nand U16997 ( n4061, n4646, n4647 );
nand U16998 ( n4647, n4648, n11527 );
nand U16999 ( n4648, n4649, n4650 );
nand U17000 ( n2538, n2672, n284 );
nand U17001 ( n4240, n4711, n4712 );
and U17002 ( n4711, n4713, n948 );
nand U17003 ( n3984, n341, n3985 );
nand U17004 ( n3985, n353, n356 );
not U17005 ( n337, n2774 );
nand U17006 ( n5482, n5483, n866 );
not U17007 ( n866, n5484 );
nor U17008 ( n5483, n5462, n5485 );
nor U17009 ( n5485, n5463, n857 );
nor U17010 ( n1631, n1632, n1633 );
nor U17011 ( n1632, n367, n1638 );
nor U17012 ( n1633, n1634, n1636 );
not U17013 ( n367, n1634 );
nand U17014 ( n1636, n1637, n1607 );
nand U17015 ( n1637, n52, n363 );
not U17016 ( n351, n2769 );
nor U17017 ( n9392, n356, n353 );
nor U17018 ( n9389, n352, n9390 );
nand U17019 ( n9390, n2769, n2545 );
and U17020 ( n9366, n9393, n9394 );
nor U17021 ( n9393, n341, n2652 );
nand U17022 ( n8618, n9371, n9372 );
and U17023 ( n9371, n8964, n8963 );
nand U17024 ( n9372, n9216, n11533 );
or U17025 ( n8794, n8618, n11534 );
nand U17026 ( n1638, n1639, n363 );
nor U17027 ( n1621, n1622, n1623 );
nand U17028 ( n1623, n1624, n1598 );
nand U17029 ( n1624, n59, n364 );
nand U17030 ( n8634, n8963, n9213 );
nand U17031 ( n9213, n9214, n11533 );
nand U17032 ( n9214, n74, n9215 );
nand U17033 ( n9215, n2534, n109 );
not U17034 ( n74, n9216 );
nor U17035 ( n4709, n4742, n929 );
or U17036 ( n4742, n4705, n939 );
nand U17037 ( n5481, n5486, n5484 );
nor U17038 ( n5486, n5463, n5489 );
nor U17039 ( n5489, n5462, n5461 );
nand U17040 ( n4243, n942, n4747 );
nand U17041 ( n4747, n4748, n4749 );
nand U17042 ( n4749, n949, n4745 );
and U17043 ( n1619, n1622, n11240 );
and U17044 ( n11240, n1627, n364 );
buf U17045 ( n11282, n11529 );
nand U17046 ( n8964, n9395, n2534 );
nor U17047 ( n9395, n9225, n2652 );
nand U17048 ( n8915, n2164, n8618 );
nand U17049 ( n9017, n2254, n8618 );
nand U17050 ( n9043, n2293, n8618 );
nand U17051 ( n8955, n2343, n8618 );
nand U17052 ( n8617, n2387, n8618 );
nand U17053 ( n8897, n2431, n8618 );
nand U17054 ( n8718, n2119, n8618 );
nand U17055 ( n9370, n2203, n8618 );
nand U17056 ( n4444, n942, n4706 );
nand U17057 ( n4706, n4707, n4708 );
nand U17058 ( n4708, n4709, n948 );
nand U17059 ( n4707, n949, n4710 );
not U17060 ( n11533, n10956 );
nand U17061 ( n5455, n5460, n5461 );
or U17062 ( n5460, n5462, n5463 );
not U17063 ( n924, n6776 );
nand U17064 ( n8184, n8185, n8186 );
nand U17065 ( n8186, n907, n938 );
xnor U17066 ( n8185, n939, n6642 );
nor U17067 ( n8146, n939, n907 );
not U17068 ( n926, n6780 );
nor U17069 ( n8144, n938, n929 );
not U17070 ( n338, n2713 );
not U17071 ( n927, n6692 );
nand U17072 ( n2550, n4007, n4008 );
nand U17073 ( n4008, n4009, n11384 );
nor U17074 ( n4009, n947, n11402 );
nand U17075 ( n1532, n53, n374 );
nor U17076 ( n5410, n858, n5413 );
nor U17077 ( n5413, n11459, n861 );
nand U17078 ( n2658, n353, n3969 );
nor U17079 ( n3471, n333, n3483 );
nand U17080 ( n3483, n344, n2713 );
nand U17081 ( n1512, n60, n374 );
xnor U17082 ( n5679, n961, n884 );
xnor U17083 ( n5552, n959, n872 );
nand U17084 ( n4650, n4745, n4734 );
xnor U17085 ( n5788, n963, n894 );
buf U17086 ( n11417, n11248 );
nor U17087 ( n2728, n329, n284 );
nor U17088 ( n8253, n4744, n954 );
not U17089 ( n381, n1724 );
not U17090 ( n379, n1816 );
nor U17091 ( n3556, n338, n2719 );
nor U17092 ( n8304, n11323, n11282 );
nand U17093 ( n1451, n55, n388 );
nand U17094 ( n4646, n4712, n4716 );
nand U17095 ( n1428, n62, n388 );
nand U17096 ( n6649, n921, n6497 );
not U17097 ( n921, n6499 );
nor U17098 ( n3997, n11408, n11534 );
nor U17099 ( n3596, n3603, n3604 );
nand U17100 ( n3603, n2774, n2769 );
nand U17101 ( n3604, n2906, n2775 );
not U17102 ( n373, n1708 );
not U17103 ( n372, n1799 );
nor U17104 ( n7473, n7484, n7485 );
nand U17105 ( n7484, n5187, n6780 );
nand U17106 ( n7485, n6776, n6777 );
buf U17107 ( n11342, n11339 );
nor U17108 ( n7430, n917, n7472 );
nand U17109 ( n7472, n4739, n6692 );
nand U17110 ( n1376, n1377, n1347 );
nand U17111 ( n1377, n57, n391 );
not U17112 ( n57, n1346 );
nor U17113 ( n1371, n1372, n1373 );
nor U17114 ( n1372, n396, n1378 );
nor U17115 ( n1373, n1374, n1376 );
not U17116 ( n396, n1374 );
nor U17117 ( n1361, n1362, n1363 );
nand U17118 ( n1363, n1364, n1338 );
nand U17119 ( n1364, n64, n392 );
not U17120 ( n64, n1337 );
and U17121 ( n1359, n1362, n11241 );
and U17122 ( n11241, n1367, n392 );
not U17123 ( n65, n1271 );
nand U17124 ( n1311, n1312, n1269 );
nand U17125 ( n1312, n65, n401 );
nor U17126 ( n1306, n1307, n1308 );
nor U17127 ( n1307, n398, n1313 );
nor U17128 ( n1308, n1309, n1311 );
not U17129 ( n398, n1309 );
not U17130 ( n357, n1763 );
nand U17131 ( n1332, n1336, n1337 );
nand U17132 ( n1336, n392, n1338 );
nor U17133 ( n1289, n1291, n1292 );
nand U17134 ( n1292, n1293, n1263 );
nand U17135 ( n1293, n67, n402 );
not U17136 ( n67, n1262 );
nand U17137 ( n1313, n1314, n401 );
nand U17138 ( n1314, n1271, n1269 );
nor U17139 ( n1288, n399, n1294 );
not U17140 ( n399, n1291 );
nand U17141 ( n1294, n1296, n402 );
nand U17142 ( n1296, n1262, n1263 );
not U17143 ( n404, n1321 );
not U17144 ( n364, n1628 );
not U17145 ( n363, n1641 );
not U17146 ( n406, n1303 );
not U17147 ( n402, n1297 );
not U17148 ( n401, n1316 );
not U17149 ( n392, n1368 );
not U17150 ( n391, n1381 );
and U17151 ( n1268, n1269, n401 );
not U17152 ( n376, n1529 );
nand U17153 ( n1261, n402, n1263 );
not U17154 ( n11527, n11528 );
buf U17155 ( n11283, n11529 );
not U17156 ( n411, n1254 );
nand U17157 ( n1866, n11421, n3999 );
not U17158 ( n708, n9848 );
nand U17159 ( n9686, n9648, n9387 );
nor U17160 ( n10269, n10270, n10271 );
nand U17161 ( n10271, n10272, n10258 );
nand U17162 ( n10272, n777, n1176 );
nand U17163 ( n10427, n766, n10509 );
nor U17164 ( n9564, n9650, n9651 );
nor U17165 ( n9651, n9356, n9652 );
nor U17166 ( n9650, n2769, n9686 );
xnor U17167 ( n9652, n359, n9653 );
nand U17168 ( n10047, n10051, n10417 );
nand U17169 ( n10417, n10049, n10014 );
and U17170 ( n9693, n10260, n10261 );
nand U17171 ( n10261, n9553, n11259 );
nand U17172 ( n10260, n118, n11263 );
nand U17173 ( n10390, n10392, n10393 );
nand U17174 ( n10393, n10394, n769 );
or U17175 ( n10392, n9822, n708 );
nand U17176 ( n10394, n9824, n9819 );
nand U17177 ( n9449, n9561, n9562 );
nand U17178 ( n9561, n9563, n9378 );
nand U17179 ( n9563, n9564, n9565 );
nor U17180 ( n9565, n9566, n9567 );
and U17181 ( n8309, n10266, n10267 );
nor U17182 ( n10266, n10281, n10282 );
nor U17183 ( n10267, n10268, n10269 );
nor U17184 ( n10282, n10270, n10275 );
nand U17185 ( n10425, n764, n10510 );
not U17186 ( n764, n10509 );
not U17187 ( n766, n10510 );
nand U17188 ( n9694, n10262, n10263 );
nand U17189 ( n10263, n11262, n9553 );
nand U17190 ( n10262, n118, n11258 );
nor U17191 ( n9566, n9648, n9649 );
nand U17192 ( n9649, n341, n9356 );
nor U17193 ( n10268, n10258, n10274 );
nand U17194 ( n10274, n10270, n10275 );
not U17195 ( n45, n2533 );
not U17196 ( n327, n4435 );
not U17197 ( n408, n9051 );
or U17198 ( n11242, n10803, n1249 );
not U17199 ( n7, n9292 );
nand U17200 ( n8793, n9288, n9289 );
nand U17201 ( n9288, n9291, n9292 );
nand U17202 ( n9289, n9290, n9149 );
nand U17203 ( n9290, n7, n46 );
nand U17204 ( n4816, n11385, n6650 );
nand U17205 ( n4758, n4761, n4762 );
nor U17206 ( n4762, n4763, n4764 );
nor U17207 ( n4761, n5185, n5186 );
nand U17208 ( n4764, n4765, n4760 );
nor U17209 ( n2395, n4756, n4757 );
and U17210 ( n4756, n4760, n946 );
nand U17211 ( n4757, n4758, n4759 );
nand U17212 ( n4759, n11530, n4760 );
nand U17213 ( n9301, n11286, n2533 );
xor U17214 ( n9291, n339, n9297 );
nor U17215 ( n9297, n9298, n9299 );
nor U17216 ( n9298, n9302, n10963 );
nand U17217 ( n9299, n9300, n9301 );
nand U17218 ( n9567, n9568, n3970 );
nand U17219 ( n9568, n9569, n9570 );
nor U17220 ( n9569, n9384, n329 );
nor U17221 ( n9570, n9477, n9571 );
nand U17222 ( n1310, n8619, n8620 );
nor U17223 ( n8619, n8630, n8631 );
nor U17224 ( n8620, n8621, n8622 );
nor U17225 ( n8630, P1_STATE_REG, n11121 );
nand U17226 ( n9668, n9670, n9671 );
xnor U17227 ( n9670, n2665, n2700 );
xnor U17228 ( n9671, n118, n9553 );
nor U17229 ( n4763, n4743, n4830 );
xor U17230 ( n4830, n4831, n4832 );
xnor U17231 ( n4832, n11402, n907 );
nand U17232 ( n4831, n4833, n4834 );
nor U17233 ( n4878, n6655, n11382 );
or U17234 ( n11243, n5314, n5869 );
nand U17235 ( n5869, n8157, n8158 );
nand U17236 ( n8098, n967, n5007 );
not U17237 ( n1013, n7955 );
not U17238 ( n1011, n8292 );
or U17239 ( n8158, n8159, n11455 );
nand U17240 ( n1884, n1886, n1887 );
or U17241 ( n1887, n11437, n1888 );
nand U17242 ( n1886, n11513, n1889 );
nand U17243 ( n895, n1881, n1882 );
nor U17244 ( n1881, n1893, n1894 );
nor U17245 ( n1882, n1883, n1884 );
nor U17246 ( n1893, n11511, n11143 );
nand U17247 ( n9457, n9550, n9551 );
nand U17248 ( n9550, n9553, n1866 );
nand U17249 ( n9551, n9552, n9463 );
nand U17250 ( n9463, n2700, n242 );
nor U17251 ( n9451, n73, n9452 );
xnor U17252 ( n9452, n9453, n9384 );
nand U17253 ( n9453, n9454, n9455 );
nand U17254 ( n9455, n9456, n119 );
nand U17255 ( n6148, n6149, n6150 );
nand U17256 ( n6150, n11375, n4062 );
nand U17257 ( n6149, n11480, n6151 );
nand U17258 ( n5020, n8125, n8126 );
nand U17259 ( n8126, n8127, n11384 );
nand U17260 ( n8125, n11383, n5437 );
nand U17261 ( n1255, n8840, n8841 );
nor U17262 ( n8840, n8855, n8856 );
nor U17263 ( n8841, n8842, n8843 );
nor U17264 ( n8855, P1_STATE_REG, n11108 );
nand U17265 ( n4765, n4766, n4767 );
nor U17266 ( n4766, n929, n4738 );
xnor U17267 ( n4767, n4768, n4769 );
nand U17268 ( n4768, n4770, n4771 );
nand U17269 ( n2696, n2697, n2698 );
nand U17270 ( n2698, n2699, n2700 );
nand U17271 ( n2697, n352, n2703 );
nand U17272 ( n2699, n2701, n2702 );
nand U17273 ( n2512, n9976, n9977 );
nand U17274 ( n9977, n9978, n11420 );
nand U17275 ( n9976, n11419, n1853 );
nand U17276 ( n2120, n6116, n6117 );
nor U17277 ( n6117, n6118, n6119 );
nor U17278 ( n6116, n6124, n6125 );
and U17279 ( n6118, n6113, n11375 );
nand U17280 ( n2501, n9985, n9986 );
nand U17281 ( n9986, n9048, n11420 );
nand U17282 ( n9985, n11419, n1192 );
nand U17283 ( n4350, n7992, n7993 );
nand U17284 ( n7993, n7994, n11384 );
nand U17285 ( n7992, n11383, n5533 );
nand U17286 ( n5064, n8099, n8100 );
nand U17287 ( n8100, n8101, n11385 );
nand U17288 ( n8099, n11383, n5459 );
nor U17289 ( n9456, n9458, n9459 );
nor U17290 ( n9459, n242, n2700 );
nor U17291 ( n9458, n9460, n9461 );
nand U17292 ( n9461, n9462, n9463 );
nand U17293 ( n2471, n10023, n10024 );
nand U17294 ( n10024, n8883, n11421 );
nand U17295 ( n10023, n11419, n1854 );
nor U17296 ( n4885, n6728, n11382 );
nand U17297 ( n6136, n6137, n6138 );
nand U17298 ( n6138, n11375, n4198 );
nand U17299 ( n6137, n11480, n6139 );
nand U17300 ( n4580, n8004, n8005 );
nor U17301 ( n8004, n8010, n8011 );
nor U17302 ( n8005, n8006, n8007 );
nor U17303 ( n8010, n11344, n10980 );
not U17304 ( n1008, n8169 );
and U17305 ( n8006, n4349, n11337 );
nor U17306 ( n9477, n1866, n9553 );
nand U17307 ( n4344, n8039, n8040 );
nor U17308 ( n8039, n8044, n8045 );
nor U17309 ( n8040, n8041, n8042 );
nor U17310 ( n8044, n11344, n10995 );
and U17311 ( n8041, n4409, n11337 );
nor U17312 ( n9913, n1177, n9894 );
nand U17313 ( n10436, n9913, n10434 );
and U17314 ( n10408, n9912, n10434 );
nand U17315 ( n9912, n9894, n1177 );
nand U17316 ( n4038, n7966, n7967 );
nor U17317 ( n7966, n7972, n7973 );
nor U17318 ( n7967, n7968, n7969 );
nor U17319 ( n7972, n11344, n11000 );
and U17320 ( n7968, n4585, n11337 );
nand U17321 ( n4141, n8062, n8063 );
nand U17322 ( n8063, n8064, n11385 );
nand U17323 ( n8062, n11383, n5488 );
nor U17324 ( n4311, n6975, n11382 );
not U17325 ( n116, n10844 );
nand U17326 ( n6160, n6161, n6162 );
nand U17327 ( n6162, n11375, n4645 );
nand U17328 ( n6161, n11480, n6163 );
nand U17329 ( n9302, n10837, n9446 );
nor U17330 ( n10837, n113, n9402 );
nand U17331 ( n4410, n8026, n8027 );
nand U17332 ( n8026, n8032, n11385 );
nand U17333 ( n8027, n11383, n5508 );
not U17334 ( n113, n9443 );
nand U17335 ( n6672, n6695, n6696 );
nand U17336 ( n6695, n6698, n11402 );
nand U17337 ( n6696, n6697, n4199 );
nor U17338 ( n6698, n1003, n6657 );
nand U17339 ( n1300, n8649, n8650 );
nor U17340 ( n8649, n8660, n8661 );
nor U17341 ( n8650, n8651, n8652 );
nor U17342 ( n8660, P1_STATE_REG, n11100 );
nand U17343 ( n4586, n7949, n7950 );
nand U17344 ( n7950, n7951, n11385 );
nand U17345 ( n7949, n11383, n5559 );
not U17346 ( n1007, n8172 );
nand U17347 ( n3956, n10765, n10766 );
nor U17348 ( n10766, n10767, n10768 );
nor U17349 ( n10765, n10771, n10772 );
nor U17350 ( n10767, n11305, n10964 );
nor U17351 ( n10771, n11307, n10963 );
not U17352 ( n326, n10770 );
nand U17353 ( n10471, n326, n10769 );
nand U17354 ( n4693, n8148, n8149 );
nor U17355 ( n8148, n8152, n8153 );
nor U17356 ( n8149, n8150, n8151 );
nor U17357 ( n8152, n11344, n10967 );
nor U17358 ( n8151, n11338, n10968 );
nand U17359 ( n905, n1858, n1859 );
nor U17360 ( n1858, n1868, n1869 );
nor U17361 ( n1859, n1861, n1862 );
nor U17362 ( n1869, n11513, n11131 );
not U17363 ( n539, n5007 );
nor U17364 ( n9376, n3970, n9384 );
not U17365 ( n354, n10828 );
nand U17366 ( n4046, n7895, n7896 );
nand U17367 ( n7895, n7900, n11385 );
nand U17368 ( n7896, n11383, n5586 );
nor U17369 ( n10768, n11300, n10965 );
nand U17370 ( n10485, n10769, n10770 );
nand U17371 ( n6203, n6204, n6205 );
nand U17372 ( n6205, n11375, n4101 );
nand U17373 ( n6204, n11480, n6206 );
not U17374 ( n356, n9356 );
nor U17375 ( n4102, n7094, n11382 );
nor U17376 ( n10468, n10770, n10769 );
nand U17377 ( n1265, n8799, n8800 );
nor U17378 ( n8799, n8818, n8819 );
nor U17379 ( n8800, n8801, n8802 );
nor U17380 ( n8818, P1_STATE_REG, n11077 );
nor U17381 ( n4513, n7159, n11382 );
nand U17382 ( n900, n1871, n1872 );
nor U17383 ( n1871, n1868, n1877 );
nor U17384 ( n1872, n1873, n1874 );
nor U17385 ( n1877, n11511, n11133 );
nand U17386 ( n6172, n6173, n6174 );
nand U17387 ( n6174, n11375, n4310 );
nand U17388 ( n6173, n11480, n6175 );
nand U17389 ( n6666, n1008, n8172 );
not U17390 ( n353, n3970 );
nand U17391 ( n4211, n7914, n7915 );
nor U17392 ( n7914, n7920, n7921 );
nor U17393 ( n7915, n7916, n7917 );
nor U17394 ( n7920, n11344, n11005 );
and U17395 ( n7916, n4045, n11337 );
nor U17396 ( n8150, n11352, n10966 );
nand U17397 ( n6662, n1007, n8169 );
nand U17398 ( n2459, n10008, n10009 );
nand U17399 ( n10009, n8668, n11421 );
nand U17400 ( n10008, n11419, n1273 );
nor U17401 ( n4393, n7033, n11382 );
nand U17402 ( n8547, n10044, n10045 );
nand U17403 ( n10045, n10046, n10047 );
nand U17404 ( n10044, n773, n10048 );
not U17405 ( n773, n10046 );
nand U17406 ( n10048, n10049, n10050 );
nand U17407 ( n10050, n751, n10051 );
not U17408 ( n751, n10014 );
not U17409 ( n359, n9384 );
nand U17410 ( n2130, n6102, n6103 );
nor U17411 ( n6102, n6104, n6105 );
nor U17412 ( n6105, n11478, n11151 );
nor U17413 ( n6104, n4816, n11380 );
nand U17414 ( n4691, n8165, n8166 );
nor U17415 ( n8165, n8170, n8171 );
nor U17416 ( n8166, n8167, n8168 );
nor U17417 ( n8170, n11344, n10986 );
nor U17418 ( n8168, n11338, n10987 );
nor U17419 ( n9847, n10397, n10107 );
nand U17420 ( n10041, n8570, n11421 );
nand U17421 ( n10040, n11419, n1304 );
nor U17422 ( n8116, n11338, n10992 );
nand U17423 ( n4136, n8113, n8114 );
nor U17424 ( n8113, n8117, n8118 );
nor U17425 ( n8114, n8115, n8116 );
nor U17426 ( n8117, n11344, n10991 );
xnor U17427 ( n8529, n9892, n9893 );
xnor U17428 ( n9893, n1177, n9894 );
nand U17429 ( n2537, n10757, n10758 );
nor U17430 ( n10758, n10759, n10760 );
nor U17431 ( n10757, n10761, n10762 );
nor U17432 ( n10759, n11305, n10974 );
nor U17433 ( n10761, n11307, n10973 );
not U17434 ( n769, n9823 );
nand U17435 ( n2125, n6107, n6103 );
nor U17436 ( n6107, n6114, n6115 );
nor U17437 ( n6115, n11477, n11154 );
nor U17438 ( n6114, n626, n11379 );
nand U17439 ( n4404, n8074, n8075 );
nor U17440 ( n8074, n8078, n8079 );
nor U17441 ( n8075, n8076, n8077 );
nor U17442 ( n8078, n11344, n10985 );
nand U17443 ( n6191, n6192, n6193 );
nand U17444 ( n6193, n11375, n4392 );
nand U17445 ( n6192, n11480, n6194 );
buf U17446 ( n11487, n11482 );
buf U17447 ( n11482, n11483 );
nand U17448 ( n4118, n7743, n7744 );
nand U17449 ( n7744, n7745, n11385 );
nand U17450 ( n7743, n11383, n5660 );
nand U17451 ( n2516, n10749, n10750 );
nor U17452 ( n10750, n10751, n10752 );
nor U17453 ( n10749, n10753, n10754 );
nor U17454 ( n10751, n11305, n10975 );
nor U17455 ( n10760, n11300, n10972 );
nand U17456 ( n4217, n7847, n7848 );
nand U17457 ( n7848, n7849, n11385 );
nand U17458 ( n7847, n11383, n5614 );
nand U17459 ( n6215, n6216, n6217 );
nand U17460 ( n6217, n11375, n4512 );
nand U17461 ( n6216, n11480, n6218 );
nor U17462 ( n10752, n11300, n10976 );
nand U17463 ( n8484, n10099, n10100 );
nand U17464 ( n10100, n10101, n10102 );
nand U17465 ( n10099, n767, n10105 );
nand U17466 ( n10102, n10103, n10104 );
nand U17467 ( n10105, n768, n10106 );
nand U17468 ( n10106, n708, n10103 );
nand U17469 ( n4290, n7649, n7650 );
nand U17470 ( n7649, n11383, n5701 );
nand U17471 ( n7650, n7651, n11384 );
nand U17472 ( n8577, n9989, n9990 );
nand U17473 ( n9990, n774, n9991 );
nor U17474 ( n9989, n9993, n9994 );
not U17475 ( n774, n9992 );
nand U17476 ( n2416, n10059, n10060 );
nand U17477 ( n10060, n8475, n11421 );
nand U17478 ( n10059, n11419, n1829 );
nand U17479 ( n2494, n10741, n10742 );
nor U17480 ( n10742, n10743, n10744 );
nor U17481 ( n10741, n10745, n10746 );
nor U17482 ( n10743, n11305, n10981 );
nor U17483 ( n10745, n11307, n10982 );
nand U17484 ( n4209, n7861, n7862 );
nor U17485 ( n7861, n7867, n7868 );
nor U17486 ( n7862, n7863, n7864 );
nor U17487 ( n7867, n11344, n11017 );
and U17488 ( n7863, n4216, n11337 );
nor U17489 ( n8167, n11352, n10984 );
nand U17490 ( n4111, n7756, n7757 );
nor U17491 ( n7756, n7762, n7763 );
nor U17492 ( n7757, n7758, n7759 );
nor U17493 ( n7762, n11344, n11015 );
and U17494 ( n7758, n4117, n11337 );
nand U17495 ( n8519, n9907, n9908 );
nand U17496 ( n9908, n9909, n9910 );
nand U17497 ( n9907, n771, n9914 );
nand U17498 ( n9910, n772, n9911 );
nand U17499 ( n9914, n9912, n9915 );
or U17500 ( n9915, n9892, n9913 );
nand U17501 ( n4532, n7702, n7703 );
nand U17502 ( n7703, n11383, n5685 );
nand U17503 ( n7702, n7707, n11384 );
nand U17504 ( n4112, n7813, n7814 );
nor U17505 ( n7813, n7819, n7820 );
nor U17506 ( n7814, n7815, n7816 );
nor U17507 ( n7819, n11344, n11018 );
and U17508 ( n7815, n4425, n11337 );
nor U17509 ( n8314, P2_STATE_REG, n6655 );
nor U17510 ( n8007, n11352, n10979 );
nor U17511 ( n8115, n11352, n10989 );
nor U17512 ( n4003, n11533, n4006 );
nor U17513 ( n8076, n11352, n10983 );
nand U17514 ( n9911, n9892, n9912 );
nand U17515 ( n4159, n7322, n7323 );
nand U17516 ( n7323, n11383, n4769 );
nand U17517 ( n7322, n7324, n11384 );
nand U17518 ( n10104, n9848, n768 );
nand U17519 ( n2382, n9888, n9889 );
nand U17520 ( n9889, n8383, n11420 );
nand U17521 ( n9888, n11419, n1369 );
nor U17522 ( n8042, n11352, n10988 );
nand U17523 ( n4426, n7787, n7788 );
nand U17524 ( n7787, n7792, n11385 );
nand U17525 ( n7788, n11383, n5635 );
nor U17526 ( n7969, n11352, n10998 );
nand U17527 ( n1190, n9068, n9069 );
nor U17528 ( n9068, n1658, n9079 );
nor U17529 ( n9069, n9070, n9071 );
nand U17530 ( n9079, n9080, n9081 );
nand U17531 ( n1952, n1953, n1954 );
nand U17532 ( n1954, n11435, n1956 );
nand U17533 ( n1953, n1957, n11442 );
nand U17534 ( n6227, n6228, n6229 );
nand U17535 ( n6229, n11375, n4267 );
nand U17536 ( n6228, n11480, n6230 );
nand U17537 ( n4084, n7576, n7577 );
nand U17538 ( n7577, n11383, n5744 );
nand U17539 ( n7576, n7582, n11384 );
nand U17540 ( n4372, n7440, n7441 );
nand U17541 ( n7441, n11383, n5817 );
nand U17542 ( n7440, n7445, n11384 );
nand U17543 ( n2114, n9730, n9731 );
nand U17544 ( n9730, n11419, n9384 );
nand U17545 ( n9731, n6307, n11420 );
nand U17546 ( n2327, n10115, n10116 );
nand U17547 ( n10116, n8258, n11421 );
nand U17548 ( n10115, n11419, n1443 );
nand U17549 ( n4496, n7612, n7613 );
nand U17550 ( n7612, n11383, n5721 );
nand U17551 ( n7613, n7614, n11384 );
nor U17552 ( n8321, P2_STATE_REG, n6728 );
nand U17553 ( n8753, n9361, n9302 );
nand U17554 ( n9361, n9362, n353 );
nor U17555 ( n9362, n9357, n9363 );
nor U17556 ( n9363, n359, n9356 );
nor U17557 ( n4014, P1_STATE_REG, n4015 );
nand U17558 ( n2372, n9903, n9904 );
nand U17559 ( n9904, n8274, n11420 );
nand U17560 ( n9903, n11419, n1442 );
nand U17561 ( n8766, n8767, n8768 );
nand U17562 ( n8768, n1912, n8634 );
nand U17563 ( n8767, n11524, n1923 );
nand U17564 ( n4284, n7717, n7718 );
nor U17565 ( n7717, n7723, n7724 );
nor U17566 ( n7718, n7719, n7720 );
nor U17567 ( n7723, n11344, n11028 );
and U17568 ( n7719, n4531, n11337 );
nand U17569 ( n4564, n7382, n7383 );
nand U17570 ( n7383, n11383, n5837 );
nand U17571 ( n7382, n7388, n11384 );
nand U17572 ( n4746, n7530, n7531 );
nand U17573 ( n7531, n11383, n5769 );
nand U17574 ( n7530, n7535, n11384 );
nand U17575 ( n4195, n4196, n4197 );
nand U17576 ( n4197, n4061, n4198 );
nand U17577 ( n4196, n4199, n11464 );
nand U17578 ( n2338, n9925, n9926 );
nand U17579 ( n9926, n8266, n11420 );
nand U17580 ( n9925, n11419, n1436 );
nand U17581 ( n4333, n7489, n7490 );
nand U17582 ( n7490, n11383, n5795 );
nand U17583 ( n7489, n7496, n11384 );
nand U17584 ( n2283, n10095, n10096 );
nand U17585 ( n10095, n11419, n1519 );
nand U17586 ( n10096, n7797, n11421 );
not U17587 ( n341, n9387 );
nor U17588 ( n9357, n9384, n341 );
nand U17589 ( n6239, n6240, n6241 );
nand U17590 ( n6241, n11375, n4467 );
nand U17591 ( n6240, n11480, n6242 );
nand U17592 ( n2249, n9839, n9840 );
nand U17593 ( n9839, n11419, n1704 );
nand U17594 ( n9840, n7330, n11420 );
nand U17595 ( n2148, n9772, n9773 );
nand U17596 ( n9772, n11419, n1681 );
nand U17597 ( n9773, n6435, n11420 );
nor U17598 ( n7917, n11352, n11004 );
nand U17599 ( n6251, n6252, n6253 );
nand U17600 ( n6253, n11375, n4158 );
nand U17601 ( n6252, n11480, n6254 );
nand U17602 ( n1250, n8859, n8860 );
nor U17603 ( n8859, n1609, n8875 );
nor U17604 ( n8860, n8861, n8862 );
nand U17605 ( n8875, n8876, n8877 );
nor U17606 ( n8329, P2_STATE_REG, n6792 );
nand U17607 ( n1997, n1998, n1999 );
nand U17608 ( n1999, n11435, n2001 );
nand U17609 ( n1998, n11443, n2002 );
nand U17610 ( n2474, n10733, n10734 );
nor U17611 ( n10734, n10735, n10736 );
nor U17612 ( n10733, n10737, n10738 );
nor U17613 ( n10736, n11305, n11007 );
nor U17614 ( n10737, n11307, n11009 );
nand U17615 ( n4490, n7669, n7670 );
nor U17616 ( n7669, n7675, n7676 );
nor U17617 ( n7670, n7671, n7672 );
nor U17618 ( n7675, n11345, n11033 );
and U17619 ( n7671, n4289, n11337 );
nor U17620 ( n4220, n11533, n4223 );
nand U17621 ( n9354, n3970, n9356 );
or U17622 ( n9355, n9356, n9357 );
nand U17623 ( n4078, n7624, n7625 );
nor U17624 ( n7624, n7630, n7631 );
nor U17625 ( n7625, n7626, n7627 );
nor U17626 ( n7630, n11345, n11039 );
and U17627 ( n7626, n4495, n11337 );
nand U17628 ( n2193, n10130, n10131 );
nand U17629 ( n10130, n11419, n1781 );
nand U17630 ( n10131, n6572, n11421 );
nor U17631 ( n10735, n828, n11302 );
not U17632 ( n828, n2448 );
nand U17633 ( n2447, n10725, n10726 );
nor U17634 ( n10726, n10727, n10728 );
nor U17635 ( n10725, n10729, n10730 );
nor U17636 ( n10728, n11305, n11011 );
nor U17637 ( n10729, n11307, n11012 );
nand U17638 ( n4058, n4059, n4060 );
nand U17639 ( n4060, n4061, n4062 );
nand U17640 ( n4059, n4063, n11464 );
nand U17641 ( n2204, n9791, n9792 );
nand U17642 ( n9791, n11419, n1576 );
nand U17643 ( n9792, n6611, n11420 );
nand U17644 ( n2429, n10716, n10717 );
nor U17645 ( n10717, n10718, n10719 );
nor U17646 ( n10716, n10721, n10722 );
nor U17647 ( n10719, n11305, n11020 );
nor U17648 ( n10721, n11307, n11023 );
nand U17649 ( n2159, n9759, n9760 );
nand U17650 ( n9759, n11419, n1629 );
nand U17651 ( n9760, n6537, n11420 );
nand U17652 ( n9951, n286, n9952 );
nand U17653 ( n9952, n11260, n2533 );
nand U17654 ( n2294, n10082, n10083 );
nand U17655 ( n10082, n11419, n1479 );
nand U17656 ( n10083, n8252, n11421 );
nand U17657 ( n6263, n6264, n6265 );
nand U17658 ( n6265, n11375, n4563 );
nand U17659 ( n6264, n11480, n6266 );
nand U17660 ( n2087, n2088, n2089 );
nand U17661 ( n2089, n11435, n2091 );
nand U17662 ( n2088, n2092, n11442 );
nor U17663 ( n10718, n817, n11302 );
not U17664 ( n817, n2403 );
nor U17665 ( n7864, n11352, n11014 );
nand U17666 ( n1305, n8635, n8636 );
nor U17667 ( n8635, n1563, n8646 );
nor U17668 ( n8636, n8637, n8638 );
nand U17669 ( n8646, n8647, n8648 );
nor U17670 ( n7759, n11352, n11013 );
nor U17671 ( n8339, n11527, n6861 );
nor U17672 ( n7816, n11352, n11016 );
nor U17673 ( n4431, n11533, n4432 );
nand U17674 ( n245, n4427, n4428 );
nand U17675 ( n4428, n3997, n4429 );
nor U17676 ( n4427, n4430, n4431 );
nor U17677 ( n4430, n4433, n10961 );
nand U17678 ( n9210, n9211, n9212 );
nand U17679 ( n9212, n1956, n8634 );
nand U17680 ( n9211, n11526, n1968 );
nor U17681 ( n3969, n9387, n9356 );
nand U17682 ( n4642, n4643, n4644 );
nand U17683 ( n4644, n4061, n4645 );
nand U17684 ( n4643, n4640, n11464 );
nand U17685 ( n2409, n10707, n10708 );
nor U17686 ( n10708, n10709, n10710 );
nor U17687 ( n10707, n10712, n10713 );
nor U17688 ( n10710, n11305, n11024 );
nor U17689 ( n10712, n11307, n11025 );
nand U17690 ( n6275, n6276, n6277 );
nand U17691 ( n6277, n11376, n4371 );
nand U17692 ( n6276, n11480, n6278 );
nand U17693 ( n4661, n7589, n7590 );
nor U17694 ( n7589, n7595, n7596 );
nor U17695 ( n7590, n7591, n7592 );
nor U17696 ( n7595, n11345, n11050 );
and U17697 ( n7591, n4083, n11337 );
nand U17698 ( n1260, n8822, n8823 );
nor U17699 ( n8822, n1497, n8837 );
nor U17700 ( n8823, n8824, n8825 );
nand U17701 ( n8837, n8838, n8839 );
nand U17702 ( n2238, n9811, n9812 );
nand U17703 ( n9811, n11419, n1561 );
nand U17704 ( n9812, n6733, n11420 );
nand U17705 ( n2510, n4142, n4143 );
nor U17706 ( n4142, n4154, n4155 );
nor U17707 ( n4143, n4144, n4145 );
nand U17708 ( n4155, n4156, n4157 );
nor U17709 ( n8346, P2_STATE_REG, n6924 );
nor U17710 ( n4752, P1_STATE_REG, n4755 );
nand U17711 ( n2342, n10680, n10681 );
nor U17712 ( n10681, n10682, n10683 );
nor U17713 ( n10680, n10685, n10686 );
nor U17714 ( n10683, n11304, n11041 );
nor U17715 ( n10685, n11307, n11043 );
not U17716 ( n771, n9909 );
nand U17717 ( n4327, n7546, n7547 );
nor U17718 ( n7546, n7552, n7553 );
nor U17719 ( n7547, n7548, n7549 );
nor U17720 ( n7552, n11345, n11057 );
and U17721 ( n7548, n4721, n11337 );
nand U17722 ( n2386, n10698, n10699 );
nor U17723 ( n10699, n10700, n10701 );
nor U17724 ( n10698, n10703, n10704 );
nor U17725 ( n10701, n11304, n11032 );
nor U17726 ( n10682, n811, n11301 );
not U17727 ( n811, n2317 );
nor U17728 ( n7720, n11352, n11027 );
nand U17729 ( n2415, n4548, n4549 );
nor U17730 ( n4548, n4559, n4560 );
nor U17731 ( n4549, n4550, n4551 );
nand U17732 ( n4560, n4561, n4562 );
or U17733 ( n11244, n11258, n3970 );
nor U17734 ( n9727, n9387, n359 );
nand U17735 ( n790, n2352, n2353 );
nor U17736 ( n2352, n2367, n2368 );
nor U17737 ( n2353, n2354, n2356 );
nor U17738 ( n2367, n11512, n11032 );
nand U17739 ( n800, n2308, n2309 );
nor U17740 ( n2308, n2322, n2323 );
nor U17741 ( n2309, n2311, n2312 );
nor U17742 ( n2322, n11512, n11041 );
nand U17743 ( n820, n2218, n2219 );
nor U17744 ( n2218, n2233, n2234 );
nor U17745 ( n2219, n2221, n2222 );
nor U17746 ( n2233, n11513, n11071 );
nand U17747 ( n810, n2263, n2264 );
nor U17748 ( n2263, n2278, n2279 );
nor U17749 ( n2264, n2266, n2267 );
nor U17750 ( n2278, n11512, n11049 );
nand U17751 ( n770, n2439, n2441 );
nor U17752 ( n2439, n2454, n2456 );
nor U17753 ( n2441, n2442, n2443 );
nor U17754 ( n2454, n11511, n11007 );
nand U17755 ( n780, n2396, n2397 );
nor U17756 ( n2396, n2411, n2412 );
nor U17757 ( n2397, n2398, n2399 );
nor U17758 ( n2411, n11512, n11020 );
nand U17759 ( n760, n2483, n2484 );
nor U17760 ( n2483, n2496, n2497 );
nor U17761 ( n2484, n2486, n2487 );
nor U17762 ( n2496, n11511, n10975 );
nand U17763 ( n4307, n4308, n4309 );
nand U17764 ( n4309, n4310, n4061 );
nand U17765 ( n4308, n4311, n11464 );
nand U17766 ( n785, n2374, n2376 );
nor U17767 ( n2374, n2388, n2389 );
nor U17768 ( n2376, n2377, n2378 );
nor U17769 ( n2388, n11511, n11024 );
nand U17770 ( n755, n2503, n2504 );
nor U17771 ( n2504, n2506, n2507 );
nor U17772 ( n2503, n2517, n2518 );
nand U17773 ( n2506, n2513, n2514 );
nand U17774 ( n2359, n10689, n10690 );
nor U17775 ( n10690, n10691, n10692 );
nor U17776 ( n10689, n10694, n10695 );
nor U17777 ( n10692, n11304, n11044 );
nor U17778 ( n10694, n11307, n11045 );
nand U17779 ( n6287, n6288, n6289 );
nand U17780 ( n6289, n11376, n4332 );
nand U17781 ( n6288, n11480, n6290 );
nor U17782 ( n10700, n808, n11302 );
not U17783 ( n808, n2361 );
nand U17784 ( n1295, n8672, n8673 );
nor U17785 ( n8672, n1464, n8683 );
nor U17786 ( n8673, n8674, n8675 );
nand U17787 ( n8683, n8684, n8685 );
nand U17788 ( n6299, n6300, n6301 );
nand U17789 ( n6301, n11376, n4721 );
nand U17790 ( n6300, n11479, n6302 );
nand U17791 ( n4366, n7506, n7507 );
nor U17792 ( n7506, n7512, n7513 );
nor U17793 ( n7507, n7508, n7509 );
nor U17794 ( n7512, n11345, n11061 );
and U17795 ( n7508, n4332, n11337 );
nor U17796 ( n8357, P2_STATE_REG, n6975 );
nor U17797 ( n7672, n11353, n11031 );
nor U17798 ( n5337, P1_STATE_REG, n5340 );
nand U17799 ( n8925, n8926, n8927 );
nand U17800 ( n8927, n2001, n8634 );
nand U17801 ( n8926, n11525, n2013 );
nand U17802 ( n4389, n4390, n4391 );
nand U17803 ( n4391, n4392, n4061 );
nand U17804 ( n4390, n4393, n11464 );
nand U17805 ( n2277, n10653, n10654 );
nor U17806 ( n10654, n10655, n10656 );
nor U17807 ( n10653, n10658, n10659 );
nor U17808 ( n10656, n11304, n11046 );
nor U17809 ( n10658, n11308, n11047 );
nor U17810 ( n7627, n11353, n11036 );
nand U17811 ( n2435, n4469, n4470 );
nor U17812 ( n4469, n4491, n4492 );
nor U17813 ( n4470, n4471, n4472 );
nand U17814 ( n4492, n4493, n4494 );
nand U17815 ( n2299, n10662, n10663 );
nor U17816 ( n10663, n10664, n10665 );
nor U17817 ( n10662, n10667, n10668 );
nor U17818 ( n10665, n11304, n11049 );
nor U17819 ( n10667, n11308, n11051 );
nand U17820 ( n4558, n7457, n7458 );
nor U17821 ( n7457, n7463, n7464 );
nor U17822 ( n7458, n7459, n7460 );
nor U17823 ( n7463, n11345, n11064 );
nand U17824 ( n2465, n4351, n4352 );
nor U17825 ( n4351, n4367, n4368 );
nor U17826 ( n4352, n4353, n4354 );
nand U17827 ( n4368, n4369, n4370 );
and U17828 ( n7459, n4371, n11337 );
nand U17829 ( n6319, n6320, n6321 );
nand U17830 ( n6321, n11376, n4083 );
nand U17831 ( n6320, n11479, n6322 );
nand U17832 ( n2316, n10671, n10672 );
nor U17833 ( n10672, n10673, n10674 );
nor U17834 ( n10671, n10676, n10677 );
nor U17835 ( n10674, n11304, n11052 );
nor U17836 ( n9538, n9539, n9540 );
nor U17837 ( n9539, n3961, n9356 );
not U17838 ( n954, n8243 );
not U17839 ( n957, n8352 );
not U17840 ( n951, n6645 );
nor U17841 ( n10664, n813, n11301 );
not U17842 ( n813, n2271 );
nand U17843 ( n2400, n4651, n4652 );
nor U17844 ( n4651, n4717, n4718 );
nor U17845 ( n4652, n4653, n4654 );
nand U17846 ( n4718, n4719, n4720 );
not U17847 ( n768, n10107 );
nor U17848 ( n8364, P2_STATE_REG, n7033 );
nor U17849 ( n5364, P1_STATE_REG, n5365 );
not U17850 ( n767, n10101 );
nand U17851 ( n2485, n4269, n4270 );
nor U17852 ( n4269, n4285, n4286 );
nor U17853 ( n4270, n4271, n4272 );
nand U17854 ( n4286, n4287, n4288 );
nand U17855 ( n8246, n956, n8280 );
not U17856 ( n956, n8281 );
nand U17857 ( n2475, n4312, n4313 );
nor U17858 ( n4312, n4328, n4329 );
nor U17859 ( n4313, n4314, n4315 );
nand U17860 ( n4329, n4330, n4331 );
nor U17861 ( n9820, n9823, n9824 );
nand U17862 ( n2267, n2268, n2269 );
nand U17863 ( n2268, n11443, n2272 );
nand U17864 ( n2269, n11434, n2271 );
nand U17865 ( n2399, n2401, n2402 );
nand U17866 ( n2401, n11442, n2404 );
nand U17867 ( n2402, n11434, n2403 );
nand U17868 ( n2179, n11435, n2181 );
nand U17869 ( n2312, n2313, n2314 );
nand U17870 ( n2314, n11439, n2316 );
nand U17871 ( n2313, n11434, n2317 );
nand U17872 ( n2356, n2357, n2358 );
nand U17873 ( n2358, n11439, n2359 );
nand U17874 ( n2357, n11434, n2361 );
nand U17875 ( n2443, n2444, n2446 );
nand U17876 ( n2446, n11439, n2447 );
nand U17877 ( n2444, n11434, n2448 );
nand U17878 ( n2133, n11435, n2137 );
nand U17879 ( n2043, n11435, n2047 );
nand U17880 ( n2222, n2223, n2224 );
nand U17881 ( n2224, n11440, n2226 );
nand U17882 ( n2223, n11435, n2227 );
nand U17883 ( n2472, n11434, n11002 );
nand U17884 ( n750, n2524, n2526 );
nor U17885 ( n2526, n2527, n2528 );
nor U17886 ( n2524, n2541, n2542 );
nor U17887 ( n2527, n10965, n11437 );
nand U17888 ( n4262, n7284, n7285 );
nor U17889 ( n7284, n7290, n7291 );
nor U17890 ( n7285, n7286, n7287 );
nor U17891 ( n7290, n11345, n11082 );
and U17892 ( n7286, n4467, n11337 );
nand U17893 ( n1906, n11434, n1912 );
nand U17894 ( n2425, n4514, n4515 );
nor U17895 ( n4514, n4527, n4528 );
nor U17896 ( n4515, n4516, n4517 );
nand U17897 ( n4528, n4529, n4530 );
nand U17898 ( n4151, n7337, n7338 );
nor U17899 ( n7337, n7343, n7344 );
nor U17900 ( n7338, n7339, n7340 );
nor U17901 ( n7343, n11345, n11078 );
and U17902 ( n7339, n4158, n11337 );
nand U17903 ( n4153, n7395, n7396 );
nor U17904 ( n7395, n7401, n7402 );
nor U17905 ( n7396, n7397, n7398 );
nor U17906 ( n7401, n11345, n11070 );
and U17907 ( n7397, n4563, n11337 );
nand U17908 ( n4098, n4099, n4100 );
nand U17909 ( n4100, n4101, n4061 );
nand U17910 ( n4099, n4102, n11464 );
nor U17911 ( n7592, n11353, n11048 );
nor U17912 ( n9540, n286, n2533 );
nand U17913 ( n1275, n8769, n8770 );
nor U17914 ( n8769, n1398, n8780 );
nor U17915 ( n8770, n8771, n8772 );
nand U17916 ( n8780, n8781, n8782 );
nand U17917 ( n6331, n6332, n6333 );
nand U17918 ( n6333, n11376, n4495 );
nand U17919 ( n6332, n11480, n6334 );
nand U17920 ( n2530, n4064, n4065 );
nor U17921 ( n4064, n4079, n4080 );
nor U17922 ( n4065, n4066, n4067 );
nand U17923 ( n4080, n4081, n4082 );
nand U17924 ( n2520, n4103, n4104 );
nor U17925 ( n4103, n4113, n4114 );
nor U17926 ( n4104, n4105, n4106 );
nand U17927 ( n4114, n4115, n4116 );
nor U17928 ( n8374, P2_STATE_REG, n7094 );
nor U17929 ( n5391, n11533, n5392 );
nand U17930 ( n6343, n6344, n6345 );
nand U17931 ( n6345, n11376, n4289 );
nand U17932 ( n6344, n11479, n6346 );
nand U17933 ( n2226, n10635, n10636 );
nor U17934 ( n10636, n10637, n10638 );
nor U17935 ( n10635, n10640, n10641 );
nor U17936 ( n10638, n11304, n11067 );
nand U17937 ( n9030, n9031, n9032 );
nand U17938 ( n9032, n2047, n8634 );
nand U17939 ( n9031, n11525, n2058 );
nand U17940 ( n4509, n4510, n4511 );
nand U17941 ( n4511, n4512, n4061 );
nand U17942 ( n4510, n4513, n11464 );
nor U17943 ( n7549, n11353, n11056 );
nand U17944 ( n2528, n2529, n2531 );
nand U17945 ( n2529, n11439, n2537 );
nand U17946 ( n2531, n2532, n2533 );
nand U17947 ( n2532, n1864, n1867 );
nand U17948 ( n5008, n5011, n5012 );
nand U17949 ( n5011, n11392, n4693 );
nand U17950 ( n5012, n11403, n5007 );
nor U17951 ( n5001, n5002, n5003 );
nor U17952 ( n5002, n5008, n5010 );
nor U17953 ( n5003, n5004, n5005 );
nand U17954 ( n5010, n939, n4738 );
nand U17955 ( n6355, n6356, n6357 );
nand U17956 ( n6357, n11376, n4531 );
nand U17957 ( n6356, n11479, n6358 );
nand U17958 ( n4507, n7234, n7235 );
nor U17959 ( n7234, n7240, n7241 );
nor U17960 ( n7235, n7236, n7237 );
nor U17961 ( n7240, n11345, n11096 );
and U17962 ( n7236, n4267, n11337 );
nand U17963 ( n2253, n10644, n10645 );
nor U17964 ( n10645, n10646, n10647 );
nor U17965 ( n10644, n10649, n10650 );
nor U17966 ( n10647, n11304, n11071 );
nand U17967 ( n4096, n7169, n7170 );
nor U17968 ( n7169, n7175, n7176 );
nor U17969 ( n7170, n7171, n7172 );
nor U17970 ( n7175, n11345, n11099 );
and U17971 ( n7171, n4512, n11337 );
nor U17972 ( n8387, P2_STATE_REG, n7159 );
nor U17973 ( n5571, n11533, n5574 );
nor U17974 ( n10646, n816, n11301 );
not U17975 ( n816, n2227 );
nand U17976 ( n1185, n9082, n9083 );
nor U17977 ( n9082, n1349, n9096 );
nor U17978 ( n9083, n9084, n9085 );
nand U17979 ( n9096, n9097, n9098 );
nand U17980 ( n2209, n10626, n10627 );
nor U17981 ( n10627, n10628, n10629 );
nor U17982 ( n10626, n10631, n10632 );
nor U17983 ( n10629, n11304, n11075 );
nor U17984 ( n10631, n11308, n11076 );
nor U17985 ( n2166, n11513, n11084 );
nor U17986 ( n2143, n11513, n11092 );
nor U17987 ( n2121, n11513, n11086 );
nor U17988 ( n2211, n11513, n11067 );
nor U17989 ( n2098, n11513, n11090 );
nor U17990 ( n2053, n11513, n11104 );
nor U17991 ( n7509, n11353, n11060 );
nand U17992 ( n2450, n4411, n4412 );
nor U17993 ( n4411, n4421, n4422 );
nor U17994 ( n4412, n4413, n4414 );
nand U17995 ( n4422, n4423, n4424 );
nand U17996 ( n4264, n4265, n4266 );
nand U17997 ( n4266, n4267, n4061 );
nand U17998 ( n4265, n4268, n11464 );
not U17999 ( n938, n4738 );
nand U18000 ( n4705, n938, n4769 );
nor U18001 ( n2541, n11511, n10964 );
nor U18002 ( n2432, n11511, n11011 );
nor U18003 ( n2188, n11512, n11075 );
nor U18004 ( n2256, n11512, n11046 );
nor U18005 ( n2476, n11511, n10981 );
nor U18006 ( n2344, n11512, n11044 );
nor U18007 ( n2301, n11511, n11052 );
nor U18008 ( n2517, n11511, n10974 );
nor U18009 ( n10628, n788, n11301 );
not U18010 ( n788, n2181 );
nor U18011 ( n1918, n11512, n11138 );
nor U18012 ( n2031, n11512, n11107 );
nor U18013 ( n2008, n11512, n11122 );
nor U18014 ( n1986, n11511, n11123 );
nor U18015 ( n1963, n11512, n11126 );
nor U18016 ( n2076, n11512, n11088 );
nor U18017 ( n1941, n11511, n11136 );
nand U18018 ( n5632, n5917, n5918 );
nand U18019 ( n5918, n5589, n5613 );
nor U18020 ( n5917, n5919, n5920 );
nor U18021 ( n5920, n5921, n5614 );
nand U18022 ( n5734, n5896, n5897 );
nand U18023 ( n5896, n5712, n5714 );
nand U18024 ( n5897, n886, n5898 );
or U18025 ( n5898, n5712, n5714 );
nand U18026 ( n5850, n5872, n5873 );
nand U18027 ( n5872, n5828, n5830 );
nand U18028 ( n5873, n896, n5874 );
or U18029 ( n5874, n5828, n5830 );
nand U18030 ( n5558, n5944, n5945 );
nand U18031 ( n5945, n5462, n5487 );
nor U18032 ( n5944, n5946, n5947 );
nor U18033 ( n5947, n5948, n5488 );
nand U18034 ( n5794, n5893, n5894 );
nand U18035 ( n5893, n5732, n5734 );
nand U18036 ( n5894, n887, n5895 );
or U18037 ( n5895, n5732, n5734 );
nor U18038 ( n5946, n5949, n5950 );
nor U18039 ( n5949, n864, n5487 );
or U18040 ( n5950, n857, n5463 );
nor U18041 ( n5919, n5922, n5923 );
nor U18042 ( n5922, n876, n5613 );
or U18043 ( n5923, n853, n5590 );
nand U18044 ( n5854, n5855, n5856 );
nand U18045 ( n5855, n5439, n4769 );
nand U18046 ( n5856, n5408, n5857 );
nand U18047 ( n5857, n5858, n5859 );
nor U18048 ( n5885, n849, n5890 );
nor U18049 ( n5890, n888, n5743 );
nor U18050 ( n5936, n854, n5941 );
nor U18051 ( n5941, n867, n5507 );
and U18052 ( n5909, n5632, n11245 );
or U18053 ( n11245, n878, n5634 );
nand U18054 ( n5461, n5953, n5954 );
nand U18055 ( n5953, n5444, n5445 );
nand U18056 ( n5954, n863, n5955 );
or U18057 ( n5955, n5444, n5445 );
or U18058 ( n5861, n5848, n5850 );
nand U18059 ( n2135, n5851, n5852 );
nor U18060 ( n5851, n4154, n6033 );
nor U18061 ( n5852, n5853, n5854 );
nand U18062 ( n6033, n6034, n6035 );
not U18063 ( n929, n4743 );
nor U18064 ( n5005, n5006, n5007 );
nor U18065 ( n5006, n967, n11406 );
nand U18066 ( n5863, n5848, n5850 );
nand U18067 ( n5859, n904, n5860 );
not U18068 ( n904, n5864 );
nand U18069 ( n5860, n5861, n5862 );
nand U18070 ( n5862, n5863, n5837 );
nor U18071 ( n7460, n11353, n11063 );
nand U18072 ( n6367, n6368, n6369 );
nand U18073 ( n6369, n11376, n4117 );
nand U18074 ( n6368, n11479, n6370 );
xnor U18075 ( n5849, n5850, n5837 );
nand U18076 ( n2140, n5831, n5832 );
nor U18077 ( n5832, n5833, n5834 );
nor U18078 ( n5831, n4559, n5844 );
nor U18079 ( n5833, n5418, n5841 );
nand U18080 ( n2187, n10617, n10618 );
nor U18081 ( n10618, n10619, n10620 );
nor U18082 ( n10617, n10622, n10623 );
nor U18083 ( n10620, n11304, n11084 );
nor U18084 ( n10622, n11308, n11085 );
nand U18085 ( n4094, n7104, n7105 );
nor U18086 ( n7104, n7110, n7111 );
nor U18087 ( n7105, n7106, n7107 );
nor U18088 ( n7110, n11345, n11103 );
and U18089 ( n7106, n4101, n11337 );
not U18090 ( n939, n5009 );
nand U18091 ( n2097, n10570, n10571 );
nor U18092 ( n10571, n10572, n10573 );
nor U18093 ( n10570, n10575, n10576 );
nor U18094 ( n10573, n11303, n11088 );
nor U18095 ( n8397, P2_STATE_REG, n7227 );
buf U18096 ( n11458, n11453 );
buf U18097 ( n11453, n11454 );
nor U18098 ( n5807, P1_STATE_REG, n5810 );
nand U18099 ( n2118, n10579, n10580 );
nor U18100 ( n10580, n10581, n10582 );
nor U18101 ( n10579, n10584, n10585 );
nor U18102 ( n10582, n11303, n11090 );
nand U18103 ( n8987, n8988, n8989 );
nand U18104 ( n8989, n2091, n8634 );
nand U18105 ( n8988, n11525, n2103 );
nand U18106 ( n6379, n6380, n6381 );
nand U18107 ( n6381, n11376, n4425 );
nand U18108 ( n6380, n11479, n6382 );
nand U18109 ( n2500, n4200, n4201 );
nor U18110 ( n4200, n4212, n4213 );
nor U18111 ( n4201, n4202, n4203 );
nand U18112 ( n4213, n4214, n4215 );
nand U18113 ( n2136, n10588, n10589 );
nor U18114 ( n10589, n10590, n10591 );
nor U18115 ( n10588, n10593, n10594 );
nor U18116 ( n10591, n11304, n11086 );
nor U18117 ( n10593, n11308, n11087 );
xnor U18118 ( n5767, n5768, n851 );
nand U18119 ( n5764, n5791, n5792 );
nand U18120 ( n5791, n5794, n5743 );
nand U18121 ( n5792, n888, n5793 );
or U18122 ( n5793, n5794, n5743 );
nand U18123 ( n5757, n5758, n5759 );
nand U18124 ( n5758, n5439, n5769 );
nand U18125 ( n5759, n5408, n5760 );
nand U18126 ( n5760, n5761, n5762 );
nor U18127 ( n5761, n5765, n5766 );
nor U18128 ( n5765, n5769, n5770 );
nor U18129 ( n5766, n893, n5767 );
nand U18130 ( n5770, n5768, n851 );
nand U18131 ( n2155, n5754, n5755 );
nor U18132 ( n5754, n4717, n5774 );
nor U18133 ( n5755, n5756, n5757 );
nand U18134 ( n5774, n5775, n5776 );
nand U18135 ( n4464, n4465, n4466 );
nand U18136 ( n4466, n4467, n4061 );
nand U18137 ( n4465, n4468, n11464 );
nand U18138 ( n4604, n6983, n6984 );
nor U18139 ( n6983, n6989, n6990 );
nor U18140 ( n6984, n6985, n6986 );
nor U18141 ( n6989, n11346, n11114 );
and U18142 ( n6985, n4310, n11337 );
nor U18143 ( n10581, n793, n11301 );
not U18144 ( n793, n2091 );
nand U18145 ( n1230, n8928, n8929 );
nor U18146 ( n8928, n1274, n8939 );
nor U18147 ( n8929, n8930, n8931 );
nand U18148 ( n8939, n8940, n8941 );
xnor U18149 ( n8189, n8410, n10996 );
nand U18150 ( n4056, n6934, n6935 );
nor U18151 ( n6934, n6940, n6941 );
nor U18152 ( n6935, n6936, n6937 );
nor U18153 ( n6940, n11346, n11117 );
and U18154 ( n6936, n4645, n11337 );
nand U18155 ( n2163, n10597, n10598 );
nor U18156 ( n10598, n10599, n10600 );
nor U18157 ( n10597, n10602, n10603 );
nor U18158 ( n10600, n11304, n11092 );
nor U18159 ( n10602, n11308, n11093 );
nor U18160 ( n6507, n6509, n6510 );
nor U18161 ( n6510, n6511, n6512 );
nor U18162 ( n6509, n6513, n6514 );
nand U18163 ( n6514, n928, n6511 );
and U18164 ( n6122, n6494, n11479 );
and U18165 ( n6494, n4769, n6495 );
nand U18166 ( n1995, n6439, n6440 );
nor U18167 ( n6439, n6446, n6447 );
nor U18168 ( n6440, n6441, n6442 );
nor U18169 ( n6446, n11479, n10988 );
nand U18170 ( n1975, n6487, n6488 );
nor U18171 ( n6487, n6500, n6501 );
nor U18172 ( n6488, n6489, n6490 );
nand U18173 ( n6501, n6502, n6503 );
nand U18174 ( n1985, n6463, n6464 );
nor U18175 ( n6463, n6470, n6471 );
nor U18176 ( n6464, n6465, n6466 );
nand U18177 ( n6471, n6472, n6473 );
nand U18178 ( n2010, n6395, n6396 );
nor U18179 ( n6395, n6402, n6403 );
nor U18180 ( n6396, n6397, n6398 );
nor U18181 ( n6402, n11479, n11004 );
nand U18182 ( n1980, n6475, n6476 );
nor U18183 ( n6475, n6482, n6483 );
nor U18184 ( n6476, n6477, n6478 );
nand U18185 ( n6483, n6484, n6485 );
nand U18186 ( n2000, n6419, n6420 );
nor U18187 ( n6419, n6426, n6427 );
nor U18188 ( n6420, n6421, n6422 );
nor U18189 ( n6426, n11479, n10979 );
nand U18190 ( n2005, n6407, n6408 );
nor U18191 ( n6407, n6414, n6415 );
nor U18192 ( n6408, n6409, n6410 );
nor U18193 ( n6414, n11479, n10998 );
nand U18194 ( n2015, n6383, n6384 );
nor U18195 ( n6383, n6390, n6391 );
nor U18196 ( n6384, n6385, n6386 );
nor U18197 ( n6390, n11479, n11014 );
nand U18198 ( n1990, n6451, n6452 );
nor U18199 ( n6451, n6458, n6459 );
nor U18200 ( n6452, n6453, n6454 );
nor U18201 ( n6458, n11479, n10983 );
nand U18202 ( n2540, n4018, n4019 );
nor U18203 ( n4018, n4040, n4041 );
nor U18204 ( n4019, n4020, n4021 );
nand U18205 ( n4041, n4042, n4043 );
nor U18206 ( n7398, n11353, n11069 );
not U18207 ( n873, n8539 );
nand U18208 ( n8703, n8704, n8705 );
nand U18209 ( n8705, n8618, n11002 );
nand U18210 ( n8704, n11524, n2471 );
nor U18211 ( n10599, n791, n11301 );
not U18212 ( n791, n2137 );
nand U18213 ( n2074, n10561, n10562 );
nor U18214 ( n10562, n10563, n10564 );
nor U18215 ( n10561, n10566, n10567 );
nor U18216 ( n10564, n11303, n11104 );
nand U18217 ( n6391, n6392, n6393 );
nand U18218 ( n6393, n11376, n4216 );
nand U18219 ( n6392, n11479, n6394 );
nand U18220 ( n6415, n6416, n6417 );
nand U18221 ( n6417, n11376, n4585 );
nand U18222 ( n6416, n11480, n6418 );
nor U18223 ( n7287, n11353, n11080 );
nor U18224 ( n8404, n11527, n7277 );
nor U18225 ( n6179, P1_STATE_REG, n6180 );
nor U18226 ( n7340, n11353, n11079 );
nand U18227 ( n2145, n5811, n5812 );
nor U18228 ( n5812, n5813, n5814 );
nor U18229 ( n5811, n4367, n5824 );
nor U18230 ( n5813, n5418, n5821 );
nand U18231 ( n4305, n7047, n7048 );
nor U18232 ( n7047, n7053, n7054 );
nor U18233 ( n7048, n7049, n7050 );
nor U18234 ( n7053, n11346, n11120 );
and U18235 ( n7049, n4392, n11337 );
nand U18236 ( n5783, n5784, n5785 );
nand U18237 ( n5784, n5439, n5795 );
nand U18238 ( n5785, n5408, n5786 );
xor U18239 ( n5786, n5787, n5788 );
nand U18240 ( n2150, n5780, n5781 );
nor U18241 ( n5780, n4328, n5799 );
nor U18242 ( n5781, n5782, n5783 );
nand U18243 ( n5799, n5800, n5801 );
nor U18244 ( n5463, n5458, n862 );
and U18245 ( n5462, n862, n5458 );
nor U18246 ( n5948, n5462, n5487 );
nor U18247 ( n10563, n796, n11300 );
not U18248 ( n796, n2047 );
nand U18249 ( n2410, n4565, n4566 );
nor U18250 ( n4565, n4581, n4582 );
nor U18251 ( n4566, n4567, n4568 );
nand U18252 ( n4582, n4583, n4584 );
nand U18253 ( n6403, n6404, n6405 );
nand U18254 ( n6405, n11376, n4045 );
nand U18255 ( n6404, n11480, n6406 );
nand U18256 ( n2046, n10552, n10553 );
nor U18257 ( n10553, n10554, n10555 );
nor U18258 ( n10552, n10557, n10558 );
nor U18259 ( n10555, n11303, n11107 );
nor U18260 ( n7237, n11353, n11094 );
nand U18261 ( n5928, n959, n5559 );
nor U18262 ( n5930, n5527, n5933 );
nor U18263 ( n5933, n5934, n5935 );
nand U18264 ( n5935, n867, n5507 );
not U18265 ( n959, n5932 );
nand U18266 ( n2470, n4334, n4335 );
nor U18267 ( n4334, n4345, n4346 );
nor U18268 ( n4335, n4336, n4337 );
nand U18269 ( n4346, n4347, n4348 );
nand U18270 ( n5554, n5532, n5533 );
xnor U18271 ( n7899, n1013, n10978 );
nor U18272 ( n7172, n11353, n11097 );
nand U18273 ( n6427, n6428, n6429 );
nand U18274 ( n6429, n11377, n4349 );
nand U18275 ( n6428, n11480, n6430 );
and U18276 ( n8415, n11283, n7324 );
and U18277 ( n6306, n11534, n6307 );
nand U18278 ( n4182, n6868, n6869 );
nor U18279 ( n6868, n6874, n6875 );
nor U18280 ( n6869, n6870, n6871 );
nor U18281 ( n6874, n11346, n11141 );
and U18282 ( n6870, n4062, n11337 );
nand U18283 ( n1195, n9052, n9053 );
nor U18284 ( n9052, n9066, n9067 );
nor U18285 ( n9053, n9054, n9055 );
nor U18286 ( n9066, n289, n11319 );
nand U18287 ( n5738, n5739, n5740 );
nand U18288 ( n5739, n5439, n5744 );
nand U18289 ( n5740, n5408, n5741 );
xnor U18290 ( n5741, n849, n5742 );
nand U18291 ( n2160, n5735, n5736 );
nor U18292 ( n5735, n4079, n5748 );
nor U18293 ( n5736, n5737, n5738 );
nand U18294 ( n5748, n5749, n5750 );
nand U18295 ( n10897, n783, n11106 );
not U18296 ( n783, n10903 );
nor U18297 ( ADD_1068_U4, n10894, n10895 );
nor U18298 ( n10895, n781, n10896 );
nor U18299 ( n10894, n10900, n10901 );
not U18300 ( n781, n10900 );
nor U18301 ( n5527, n5533, n5532 );
nand U18302 ( n6447, n6448, n6449 );
nand U18303 ( n6449, n11377, n4409 );
nand U18304 ( n6448, n11480, n6450 );
not U18305 ( n883, n8487 );
nand U18306 ( n8009, n10970, n10958 );
nand U18307 ( n3981, n9405, n9406 );
nor U18308 ( n9405, n9424, n9425 );
nor U18309 ( n9406, n9407, n9408 );
nand U18310 ( n9424, n9434, n9435 );
nand U18311 ( n9408, n9409, n9410 );
nand U18312 ( n9409, n112, n9414 );
nand U18313 ( n9410, n112, n9411 );
nand U18314 ( n9414, n9415, n9416 );
not U18315 ( n114, n9446 );
nand U18316 ( n9401, n9441, n9442 );
nand U18317 ( n9442, n9443, n11111 );
nor U18318 ( n9441, n9402, n9444 );
nor U18319 ( n9444, n11111, n9445 );
or U18320 ( n2552, n3981, n3979 );
nand U18321 ( n9425, n9426, n9427 );
nand U18322 ( n9426, n112, n9431 );
nand U18323 ( n9427, n112, n9428 );
nand U18324 ( n9431, n9432, n9433 );
buf U18325 ( n11390, n4879 );
nand U18326 ( n4879, n4738, n5009 );
nand U18327 ( n10896, n10897, n10898 );
nand U18328 ( n10898, n10899, n11110 );
nand U18329 ( n9407, n9417, n9418 );
nand U18330 ( n9417, n112, n9422 );
nand U18331 ( n9418, n112, n9419 );
nand U18332 ( n9422, n9423, n11128 );
not U18333 ( n863, n5437 );
nand U18334 ( n5517, n6088, n6089 );
nand U18335 ( n6088, n5497, n5488 );
nand U18336 ( n6089, n6090, n10983 );
or U18337 ( n6090, n5497, n5488 );
nand U18338 ( n5473, n6094, n6095 );
nand U18339 ( n6094, n861, n5437 );
nand U18340 ( n6095, n6096, n10984 );
nand U18341 ( n6096, n863, n5424 );
nand U18342 ( n5693, n6067, n6068 );
nand U18343 ( n6067, n5670, n5660 );
nand U18344 ( n6068, n6069, n11013 );
or U18345 ( n6069, n5670, n5660 );
nand U18346 ( n5726, n6061, n6062 );
nand U18347 ( n6061, n5706, n5701 );
nand U18348 ( n6062, n6063, n11031 );
or U18349 ( n6063, n5706, n5701 );
nand U18350 ( n5778, n6055, n6056 );
nand U18351 ( n6055, n5753, n5744 );
nand U18352 ( n6056, n6057, n11048 );
or U18353 ( n6057, n5753, n5744 );
nand U18354 ( n5822, n6049, n6050 );
nand U18355 ( n6049, n5804, n5795 );
nand U18356 ( n6050, n6051, n11060 );
or U18357 ( n6051, n5804, n5795 );
nand U18358 ( n5842, n6046, n6047 );
nand U18359 ( n6046, n5822, n5817 );
nand U18360 ( n6047, n6048, n11063 );
or U18361 ( n6048, n5822, n5817 );
nand U18362 ( n5643, n6073, n6074 );
nand U18363 ( n6073, n5624, n5614 );
nand U18364 ( n6074, n6075, n11014 );
or U18365 ( n6075, n5624, n5614 );
nand U18366 ( n5598, n6079, n6080 );
nand U18367 ( n6079, n5568, n5559 );
nand U18368 ( n6080, n6081, n10998 );
or U18369 ( n6081, n5568, n5559 );
nand U18370 ( n5542, n6085, n6086 );
nand U18371 ( n6085, n5517, n5508 );
nand U18372 ( n6086, n6087, n10988 );
or U18373 ( n6087, n5517, n5508 );
nand U18374 ( n5497, n6091, n6092 );
nand U18375 ( n6091, n5473, n5459 );
nand U18376 ( n6092, n6093, n10989 );
or U18377 ( n6093, n5473, n5459 );
nand U18378 ( n5706, n6064, n6065 );
nand U18379 ( n6064, n5693, n5685 );
nand U18380 ( n6065, n6066, n11027 );
or U18381 ( n6066, n5693, n5685 );
nand U18382 ( n6035, n6036, n934 );
xnor U18383 ( n6036, n6042, n5868 );
nand U18384 ( n6042, n6043, n6044 );
nand U18385 ( n6043, n5842, n5837 );
nand U18386 ( n6044, n6045, n11069 );
or U18387 ( n6045, n5842, n5837 );
nand U18388 ( n5670, n6070, n6071 );
nand U18389 ( n6070, n5643, n5635 );
nand U18390 ( n6071, n6072, n11016 );
or U18391 ( n6072, n5643, n5635 );
nand U18392 ( n5753, n6058, n6059 );
nand U18393 ( n6058, n5726, n5721 );
nand U18394 ( n6059, n6060, n11036 );
or U18395 ( n6060, n5726, n5721 );
nand U18396 ( n5804, n6052, n6053 );
nand U18397 ( n6052, n5778, n5769 );
nand U18398 ( n6053, n6054, n11056 );
or U18399 ( n6054, n5778, n5769 );
nand U18400 ( n5568, n6082, n6083 );
nand U18401 ( n6082, n5542, n5533 );
nand U18402 ( n6083, n6084, n10979 );
or U18403 ( n6084, n5542, n5533 );
nand U18404 ( n5624, n6076, n6077 );
nand U18405 ( n6076, n5598, n5586 );
nand U18406 ( n6077, n6078, n11004 );
or U18407 ( n6078, n5598, n5586 );
nand U18408 ( n1270, n8783, n8784 );
nor U18409 ( n8783, n8796, n8797 );
nor U18410 ( n8784, n8785, n8786 );
nor U18411 ( n8796, n288, n11320 );
xnor U18412 ( n8882, n408, n10971 );
nand U18413 ( n4897, n6805, n6806 );
nor U18414 ( n6805, n6812, n6813 );
nor U18415 ( n6806, n6807, n6808 );
nor U18416 ( n6812, n11346, n11146 );
nor U18417 ( n5853, n5419, n5977 );
xor U18418 ( n5977, n5978, n5870 );
nand U18419 ( n5978, n5979, n5980 );
nand U18420 ( n5979, n5840, n5837 );
nand U18421 ( n5704, n6000, n6001 );
nand U18422 ( n6000, n5687, n5685 );
nand U18423 ( n6001, n6002, n11028 );
or U18424 ( n6002, n5687, n5685 );
nand U18425 ( n5491, n6027, n6028 );
nand U18426 ( n6027, n5465, n5459 );
nand U18427 ( n6028, n6029, n10991 );
or U18428 ( n6029, n5465, n5459 );
nand U18429 ( n5617, n6012, n6013 );
nand U18430 ( n6012, n5592, n5586 );
nand U18431 ( n6013, n6014, n11005 );
or U18432 ( n6014, n5592, n5586 );
nand U18433 ( n5637, n6009, n6010 );
nand U18434 ( n6009, n5617, n5614 );
nand U18435 ( n6010, n6011, n11017 );
or U18436 ( n6011, n5617, n5614 );
nand U18437 ( n5819, n5985, n5986 );
nand U18438 ( n5985, n5797, n5795 );
nand U18439 ( n5986, n5987, n11061 );
or U18440 ( n5987, n5797, n5795 );
nand U18441 ( n5723, n5997, n5998 );
nand U18442 ( n5997, n5704, n5701 );
nand U18443 ( n5998, n5999, n11033 );
or U18444 ( n5999, n5704, n5701 );
nand U18445 ( n5465, n6030, n6031 );
nand U18446 ( n6030, n859, n5437 );
nand U18447 ( n6031, n6032, n10986 );
nand U18448 ( n6032, n863, n5412 );
nand U18449 ( n5510, n6024, n6025 );
nand U18450 ( n6024, n5491, n5488 );
nand U18451 ( n6025, n6026, n10985 );
or U18452 ( n6026, n5491, n5488 );
nand U18453 ( n5663, n6006, n6007 );
nand U18454 ( n6006, n5637, n5635 );
nand U18455 ( n6007, n6008, n11018 );
or U18456 ( n6008, n5637, n5635 );
nand U18457 ( n5797, n5988, n5989 );
nand U18458 ( n5988, n5772, n5769 );
nand U18459 ( n5989, n5990, n11057 );
or U18460 ( n5990, n5772, n5769 );
nand U18461 ( n5536, n6021, n6022 );
nand U18462 ( n6021, n5510, n5508 );
nand U18463 ( n6022, n6023, n10995 );
or U18464 ( n6023, n5510, n5508 );
nand U18465 ( n5980, n5981, n11070 );
or U18466 ( n5981, n5840, n5837 );
nand U18467 ( n5746, n5994, n5995 );
nand U18468 ( n5994, n5723, n5721 );
nand U18469 ( n5995, n5996, n11039 );
or U18470 ( n5996, n5723, n5721 );
nand U18471 ( n5772, n5991, n5992 );
nand U18472 ( n5991, n5746, n5744 );
nand U18473 ( n5992, n5993, n11050 );
or U18474 ( n5993, n5746, n5744 );
nand U18475 ( n5840, n5982, n5983 );
nand U18476 ( n5982, n5819, n5817 );
nand U18477 ( n5983, n5984, n11064 );
or U18478 ( n5984, n5819, n5817 );
nand U18479 ( n5592, n6015, n6016 );
nand U18480 ( n6015, n5561, n5559 );
nand U18481 ( n6016, n6017, n11000 );
or U18482 ( n6017, n5561, n5559 );
nand U18483 ( n5561, n6018, n6019 );
nand U18484 ( n6018, n5536, n5533 );
nand U18485 ( n6019, n6020, n10980 );
or U18486 ( n6020, n5536, n5533 );
nand U18487 ( n5687, n6003, n6004 );
nand U18488 ( n6003, n5663, n5660 );
nand U18489 ( n6004, n6005, n11015 );
or U18490 ( n6005, n5663, n5660 );
and U18491 ( n6807, n4198, n11337 );
nor U18492 ( n1242, n1247, n1248 );
nand U18493 ( n1248, n282, n1249 );
nand U18494 ( n1186, n1239, n1241 );
nor U18495 ( n1239, n1251, n11445 );
nor U18496 ( n1241, n1242, n1243 );
nor U18497 ( n1251, n1253, n411 );
nand U18498 ( n1237, n1238, n1186 );
nand U18499 ( n1238, n1187, n1256 );
nand U18500 ( n1256, n1257, n1258 );
nand U18501 ( n1257, n1261, n1262 );
nand U18502 ( n985, n1233, n1234 );
nor U18503 ( n1233, n1274, n1276 );
nor U18504 ( n1234, n1236, n1237 );
nand U18505 ( n1276, n1277, n1278 );
nand U18506 ( n995, n1179, n1181 );
nor U18507 ( n1179, n1198, n1199 );
nor U18508 ( n1181, n1182, n1183 );
nor U18509 ( n1198, P1_STATE_REG, n10976 );
nand U18510 ( n11287, n8157, n8158 );
and U18511 ( n8422, n11283, n7388 );
and U18512 ( n6434, n11534, n6435 );
nand U18513 ( n2029, n10543, n10544 );
nor U18514 ( n10544, n10545, n10546 );
nor U18515 ( n10543, n10548, n10549 );
nor U18516 ( n10546, n11303, n11122 );
nand U18517 ( n2165, n5715, n5716 );
nor U18518 ( n5716, n5717, n5718 );
nor U18519 ( n5715, n4491, n5728 );
nor U18520 ( n5717, n5418, n5725 );
nand U18521 ( n2007, n10534, n10535 );
nor U18522 ( n10535, n10536, n10537 );
nor U18523 ( n10534, n10539, n10540 );
nor U18524 ( n10537, n11303, n11123 );
nor U18525 ( n7107, n11353, n11101 );
nand U18526 ( n5931, n872, n5932 );
nor U18527 ( n10545, n798, n11300 );
not U18528 ( n798, n2001 );
nand U18529 ( n6459, n6460, n6461 );
nand U18530 ( n6461, n11377, n10958 );
nand U18531 ( n6460, n11480, n6462 );
nand U18532 ( n1984, n10525, n10526 );
nor U18533 ( n10526, n10527, n10528 );
nor U18534 ( n10525, n10530, n10531 );
nor U18535 ( n10528, n11303, n11126 );
nand U18536 ( n5834, n5835, n5836 );
nand U18537 ( n5836, n5439, n5837 );
nand U18538 ( n5835, n5838, n936 );
xnor U18539 ( n5838, n5839, n5840 );
nor U18540 ( n4781, n8088, n8147 );
nor U18541 ( n8147, n4693, n5007 );
xnor U18542 ( n5658, n5655, n5659 );
nand U18543 ( n5655, n5682, n5683 );
nand U18544 ( n5682, n5632, n5634 );
nand U18545 ( n5683, n878, n5684 );
or U18546 ( n5684, n5632, n5634 );
nand U18547 ( n5648, n5649, n5650 );
nand U18548 ( n5649, n5439, n5660 );
nand U18549 ( n5650, n5408, n5651 );
nand U18550 ( n5651, n5652, n5653 );
nor U18551 ( n5652, n5656, n5657 );
nor U18552 ( n5656, n5660, n5661 );
nor U18553 ( n5657, n882, n5658 );
or U18554 ( n5661, n5659, n5655 );
nand U18555 ( n2180, n5645, n5646 );
nor U18556 ( n5645, n4113, n5665 );
nor U18557 ( n5646, n5647, n5648 );
nand U18558 ( n5665, n5666, n5667 );
not U18559 ( n111, n3986 );
nor U18560 ( n10527, n801, n11300 );
not U18561 ( n801, n1956 );
nor U18562 ( n1868, n1878, n1879 );
nand U18563 ( n1220, n8956, n8957 );
nor U18564 ( n8957, n8958, n8959 );
nor U18565 ( n8956, n8965, n8966 );
nor U18566 ( n8958, n8960, n10965 );
nor U18567 ( n6482, n11479, n10984 );
nor U18568 ( n6470, n11479, n10989 );
nor U18569 ( n6125, n11477, n11148 );
nor U18570 ( n6500, n11477, n10966 );
nor U18571 ( n6286, n11478, n11060 );
nor U18572 ( n6354, n11478, n11027 );
nor U18573 ( n6318, n11478, n11048 );
nor U18574 ( n6298, n11478, n11056 );
nor U18575 ( n6366, n11478, n11013 );
nor U18576 ( n6342, n11478, n11031 );
nor U18577 ( n6262, n11478, n11069 );
nor U18578 ( n6274, n11478, n11063 );
nor U18579 ( n6330, n11478, n11036 );
nor U18580 ( n6378, n11478, n11016 );
nor U18581 ( n6250, n11478, n11079 );
nor U18582 ( n6214, n11477, n11097 );
nor U18583 ( n6202, n11477, n11101 );
nor U18584 ( n6190, n11477, n11118 );
nor U18585 ( n6171, n11477, n11112 );
nor U18586 ( n6159, n11477, n11115 );
nor U18587 ( n6147, n11477, n11139 );
nor U18588 ( n6238, n11477, n11080 );
nor U18589 ( n6226, n11477, n11094 );
nor U18590 ( n6135, n11477, n11144 );
nor U18591 ( n6986, n11354, n11112 );
not U18592 ( n324, n9553 );
nor U18593 ( n5590, n5585, n874 );
xnor U18594 ( n7706, n8487, n11010 );
xnor U18595 ( n5713, n5714, n5701 );
nand U18596 ( n2170, n5695, n5696 );
nor U18597 ( n5696, n5697, n5698 );
nor U18598 ( n5695, n4285, n5708 );
nor U18599 ( n5697, n5418, n5705 );
and U18600 ( n5589, n874, n5585 );
nor U18601 ( n5921, n5589, n5613 );
nand U18602 ( n5674, n5675, n5676 );
nand U18603 ( n5675, n5439, n5685 );
nand U18604 ( n5676, n5408, n5677 );
xor U18605 ( n5677, n5678, n5679 );
nand U18606 ( n2175, n5671, n5672 );
nor U18607 ( n5671, n4527, n5689 );
nor U18608 ( n5672, n5673, n5674 );
nand U18609 ( n5689, n5690, n5691 );
nor U18610 ( n6937, n11354, n11115 );
not U18611 ( n323, n2700 );
nor U18612 ( n7050, n11354, n11118 );
and U18613 ( n8432, n11283, n7445 );
and U18614 ( n6534, n11534, n6537 );
nand U18615 ( n5814, n5815, n5816 );
nand U18616 ( n5816, n5439, n5817 );
nand U18617 ( n5815, n5818, n936 );
xor U18618 ( n5818, n5819, n5820 );
nand U18619 ( n1962, n10516, n10517 );
nor U18620 ( n10517, n10518, n10519 );
nor U18621 ( n10516, n10521, n10522 );
nor U18622 ( n10519, n11303, n11136 );
nand U18623 ( n2420, n4533, n4534 );
nor U18624 ( n4533, n4546, n4547 );
nor U18625 ( n4534, n4535, n4536 );
nor U18626 ( n4547, n762, n4243 );
nand U18627 ( n3990, n9402, n114 );
nand U18628 ( n1939, n10491, n10492 );
nor U18629 ( n10492, n10493, n10494 );
nor U18630 ( n10491, n10496, n10497 );
nor U18631 ( n10494, n11303, n11138 );
nand U18632 ( n6040, n6097, n4007 );
nor U18633 ( n6097, n6099, n6100 );
nor U18634 ( n6100, n4730, n4733 );
nor U18635 ( n6099, n11402, n11382 );
nor U18636 ( n6515, n4769, n939 );
nand U18637 ( n2230, n5402, n5403 );
nor U18638 ( n5402, n5420, n5421 );
nor U18639 ( n5403, n5404, n5405 );
nor U18640 ( n5420, n11527, n10968 );
nand U18641 ( n2495, n4224, n4225 );
nor U18642 ( n4225, n4226, n4227 );
nor U18643 ( n4224, n4241, n4242 );
nor U18644 ( n4226, n967, n4240 );
nand U18645 ( n5428, n5429, n5430 );
nand U18646 ( n5430, n863, n5431 );
nand U18647 ( n5429, n5436, n5437 );
nand U18648 ( n5431, n5432, n5433 );
nand U18649 ( n5436, n5438, n937 );
nor U18650 ( n5438, n5440, n5441 );
nor U18651 ( n5441, n5418, n5435 );
nor U18652 ( n5440, n5419, n5434 );
nand U18653 ( n2225, n5425, n5426 );
nor U18654 ( n5425, n5446, n5447 );
nor U18655 ( n5426, n5427, n5428 );
nor U18656 ( n5447, n11527, n10987 );
nand U18657 ( n5681, n962, n5660 );
not U18658 ( n962, n5659 );
nor U18659 ( n5903, n5654, n5906 );
nor U18660 ( n5906, n5907, n5908 );
nand U18661 ( n5908, n878, n5634 );
not U18662 ( n953, n6511 );
nand U18663 ( n6508, n6643, n6644 );
xnor U18664 ( n6644, n953, n6645 );
nand U18665 ( n5433, n936, n5434 );
nand U18666 ( n5901, n961, n5685 );
not U18667 ( n961, n5905 );
nand U18668 ( n5432, n934, n5435 );
nand U18669 ( n1909, n10481, n10482 );
nor U18670 ( n10482, n10483, n10484 );
nor U18671 ( n10481, n10487, n10488 );
nor U18672 ( n10484, n11303, n11143 );
nor U18673 ( n10493, n803, n11300 );
not U18674 ( n803, n1912 );
xnor U18675 ( n8382, n9897, n11008 );
not U18676 ( n394, n9897 );
and U18677 ( n8439, n11283, n7496 );
nand U18678 ( n8207, n8208, n8209 );
nand U18679 ( n8208, n954, n8213 );
nand U18680 ( n8209, n954, n8210 );
nand U18681 ( n8213, n8214, n8215 );
and U18682 ( n6643, n8204, n8205 );
nor U18683 ( n8204, n8223, n8224 );
nor U18684 ( n8205, n8206, n8207 );
nand U18685 ( n8223, n8233, n8234 );
and U18686 ( n6571, n11534, n6572 );
nand U18687 ( n8224, n8225, n8226 );
nand U18688 ( n8225, n954, n8230 );
nand U18689 ( n8226, n954, n8227 );
nand U18690 ( n8230, n8231, n8232 );
not U18691 ( n889, n8445 );
nand U18692 ( n8206, n8216, n8217 );
nand U18693 ( n8216, n954, n8221 );
nand U18694 ( n8217, n954, n8218 );
nand U18695 ( n8221, n8222, n11134 );
nor U18696 ( n5654, n5660, n962 );
nand U18697 ( n4906, n6658, n6659 );
nor U18698 ( n6658, n6663, n6664 );
nor U18699 ( n6659, n6660, n6661 );
nor U18700 ( n6663, n11346, n11153 );
nand U18701 ( n5439, n5973, n5974 );
nand U18702 ( n5973, n11388, n5314 );
nand U18703 ( n5974, n1009, n5975 );
not U18704 ( n386, n10090 );
nor U18705 ( n10483, n11300, n1888 );
nand U18706 ( n8242, n956, n8269 );
nor U18707 ( n6103, n11246, n11247 );
and U18708 ( n11246, n11376, n6113 );
nor U18709 ( n11247, n6110, n6111 );
nand U18710 ( n5718, n5719, n5720 );
nand U18711 ( n5720, n5439, n5721 );
nand U18712 ( n5719, n5722, n936 );
xor U18713 ( n5722, n5723, n5724 );
nand U18714 ( n5698, n5699, n5700 );
nand U18715 ( n5700, n5439, n5701 );
nand U18716 ( n5699, n5702, n936 );
xnor U18717 ( n5702, n5703, n5704 );
nand U18718 ( n2185, n5625, n5626 );
nor U18719 ( n5626, n5627, n5628 );
nor U18720 ( n5625, n4421, n5639 );
nor U18721 ( n5627, n5419, n5636 );
nand U18722 ( n2190, n5600, n5601 );
nor U18723 ( n5601, n5602, n5603 );
nor U18724 ( n5600, n4212, n5619 );
nor U18725 ( n5602, n5419, n5616 );
nand U18726 ( n2195, n5575, n5576 );
nor U18727 ( n5576, n5577, n5578 );
nor U18728 ( n5575, n4040, n5594 );
nor U18729 ( n5577, n5419, n5591 );
nand U18730 ( n2200, n5544, n5545 );
nor U18731 ( n5545, n5546, n5547 );
nor U18732 ( n5544, n4581, n5563 );
nor U18733 ( n5546, n5419, n5560 );
nand U18734 ( n2205, n5518, n5519 );
nor U18735 ( n5519, n5520, n5521 );
nor U18736 ( n5518, n4345, n5538 );
nor U18737 ( n5520, n5419, n5535 );
nand U18738 ( n2210, n5499, n5500 );
nor U18739 ( n5500, n5501, n5502 );
nor U18740 ( n5499, n4405, n5512 );
nor U18741 ( n5501, n5419, n5509 );
nand U18742 ( n2215, n5474, n5475 );
nor U18743 ( n5475, n5476, n5477 );
nor U18744 ( n5474, n4137, n5493 );
nor U18745 ( n5476, n5419, n5490 );
nand U18746 ( n2220, n5448, n5449 );
nor U18747 ( n5449, n5450, n5451 );
nor U18748 ( n5448, n5467, n5468 );
nor U18749 ( n5450, n5419, n5464 );
nand U18750 ( n4877, n6700, n6701 );
nor U18751 ( n6700, n6703, n6704 );
nor U18752 ( n6701, n6660, n6702 );
nor U18753 ( n6703, n11346, n11156 );
nand U18754 ( n3993, n9402, n113 );
nor U18755 ( n9375, n9302, n9378 );
nand U18756 ( n5628, n5629, n5630 );
nand U18757 ( n5629, n5439, n5635 );
nand U18758 ( n5630, n5408, n5631 );
xnor U18759 ( n5631, n5632, n5633 );
nand U18760 ( n5603, n5604, n5605 );
nand U18761 ( n5605, n5408, n5606 );
nand U18762 ( n5604, n5439, n5614 );
nand U18763 ( n5606, n5607, n5608 );
nand U18764 ( n5578, n5579, n5580 );
nand U18765 ( n5580, n5408, n5581 );
nand U18766 ( n5579, n5439, n5586 );
nand U18767 ( n5581, n5582, n5583 );
nand U18768 ( n5547, n5548, n5549 );
nand U18769 ( n5549, n5408, n5550 );
nand U18770 ( n5548, n5439, n5559 );
xor U18771 ( n5550, n5551, n5552 );
nand U18772 ( n5521, n5522, n5523 );
nand U18773 ( n5523, n5408, n5524 );
nand U18774 ( n5522, n5439, n5533 );
nand U18775 ( n5524, n5525, n5526 );
nand U18776 ( n5502, n5503, n5504 );
nand U18777 ( n5504, n5408, n5505 );
nand U18778 ( n5503, n5439, n5508 );
xnor U18779 ( n5505, n854, n5506 );
nand U18780 ( n5477, n5478, n5479 );
nand U18781 ( n5479, n5408, n5480 );
nand U18782 ( n5478, n5439, n5488 );
nand U18783 ( n5480, n5481, n5482 );
nand U18784 ( n5451, n5452, n5453 );
nand U18785 ( n5453, n5408, n5454 );
nand U18786 ( n5452, n5439, n5459 );
nand U18787 ( n5454, n5455, n5456 );
nor U18788 ( n6871, n11354, n11139 );
xnor U18789 ( n7534, n8445, n11038 );
nand U18790 ( n4884, n6746, n6747 );
nor U18791 ( n6746, n6749, n6750 );
nor U18792 ( n6747, n6660, n6748 );
nor U18793 ( n6749, n11346, n11150 );
nor U18794 ( n5647, n5419, n5662 );
xnor U18795 ( n5662, n5663, n5664 );
xnor U18796 ( n5664, n11015, n882 );
nor U18797 ( n5737, n5419, n5745 );
xnor U18798 ( n5745, n5746, n5747 );
xnor U18799 ( n5747, n11050, n888 );
nor U18800 ( n6808, n11354, n11144 );
nand U18801 ( n4730, n8288, n8281 );
nor U18802 ( n8288, n8280, n8269 );
not U18803 ( n11425, n2660 );
nand U18804 ( n2660, n3977, n2651 );
nor U18805 ( n3977, n2652, n3986 );
and U18806 ( n2651, n3978, n3979 );
nor U18807 ( n3978, n3980, n3981 );
nor U18808 ( n3980, n3982, n3983 );
nand U18809 ( n3983, n3984, n349 );
nor U18810 ( n10711, n10720, n11003 );
not U18811 ( n281, n1879 );
nand U18812 ( n5904, n884, n5905 );
and U18813 ( n8450, n11283, n7535 );
xnor U18814 ( n5531, n5532, n856 );
nand U18815 ( n5528, n5555, n5556 );
nand U18816 ( n5555, n5558, n5507 );
nand U18817 ( n5556, n867, n5557 );
or U18818 ( n5557, n5558, n5507 );
nor U18819 ( n5525, n5529, n5530 );
nor U18820 ( n5529, n5533, n5534 );
nor U18821 ( n5530, n871, n5531 );
nand U18822 ( n5534, n5532, n856 );
xor U18823 ( n2431, n10720, n11003 );
and U18824 ( n8457, n11283, n7582 );
and U18825 ( n6608, n11534, n6611 );
and U18826 ( n6732, n11534, n6733 );
nor U18827 ( n5427, n5442, n944 );
xnor U18828 ( n5442, n5443, n5444 );
not U18829 ( n944, n5408 );
xnor U18830 ( n5443, n863, n858 );
xor U18831 ( n2254, n10648, n11042 );
nor U18832 ( n10693, n10702, n10955 );
nor U18833 ( n10675, n10684, n11026 );
nor U18834 ( n10657, n10666, n11030 );
xnor U18835 ( n8251, n10090, n11037 );
nor U18836 ( n6495, n4743, n938 );
nor U18837 ( n6661, n11354, n11151 );
xor U18838 ( n2387, n10702, n10955 );
nand U18839 ( n1005, n10779, n10780 );
nor U18840 ( n10779, n10790, n10791 );
nor U18841 ( n10780, n10781, n10782 );
nor U18842 ( n10791, n11533, n10965 );
nand U18843 ( n10786, n11285, n10964 );
not U18844 ( n328, n9378 );
nor U18845 ( n6702, n11354, n11154 );
xnor U18846 ( n6610, n9800, n11055 );
nand U18847 ( n1278, n69, n1273 );
nand U18848 ( n1663, n1664, n1666 );
nand U18849 ( n1666, n1667, n1187 );
nand U18850 ( n1664, n1759, n70 );
nor U18851 ( n1667, n1668, n1669 );
nand U18852 ( n1502, n1503, n1504 );
nand U18853 ( n1504, n1506, n11285 );
nand U18854 ( n1503, n1526, n70 );
nor U18855 ( n1506, n1507, n1508 );
nand U18856 ( n1418, n1419, n1421 );
nand U18857 ( n1421, n1422, n1187 );
nand U18858 ( n1419, n1444, n70 );
nor U18859 ( n1422, n1423, n1424 );
nand U18860 ( n910, n1659, n1661 );
nor U18861 ( n1659, n1856, n1857 );
nor U18862 ( n1661, n1662, n1663 );
nor U18863 ( n1856, n10959, n71 );
and U18864 ( n4649, n4725, n4726 );
nor U18865 ( n4725, n4732, n4733 );
nor U18866 ( n4726, n4727, n4728 );
and U18867 ( n4732, n4734, n4710 );
and U18868 ( n8481, n11283, n7651 );
and U18869 ( n7796, n11534, n7797 );
nand U18870 ( n10795, n10796, n10797 );
nand U18871 ( n10797, n11284, n10798 );
nand U18872 ( n10796, n70, n10804 );
xnor U18873 ( n10798, n1254, n10799 );
nand U18874 ( n1648, n1649, n1651 );
nand U18875 ( n1651, n1187, n1652 );
nand U18876 ( n1649, n70, n1654 );
xnor U18877 ( n1652, n58, n1653 );
nand U18878 ( n1587, n1588, n1589 );
nand U18879 ( n1589, n11284, n1591 );
nand U18880 ( n1588, n70, n1599 );
nand U18881 ( n1591, n1592, n1593 );
nand U18882 ( n1568, n1569, n1571 );
nand U18883 ( n1571, n11285, n1572 );
nand U18884 ( n1569, n70, n1577 );
xor U18885 ( n1572, n1573, n1574 );
nand U18886 ( n1549, n1551, n1552 );
nand U18887 ( n1552, n1187, n1553 );
nand U18888 ( n1551, n70, n1557 );
xor U18889 ( n1553, n1554, n1556 );
nand U18890 ( n1487, n1488, n1489 );
nand U18891 ( n1489, n11284, n1491 );
nand U18892 ( n1488, n70, n1493 );
xnor U18893 ( n1491, n60, n1492 );
nand U18894 ( n1469, n1471, n1472 );
nand U18895 ( n1472, n11285, n1473 );
nand U18896 ( n1471, n70, n1476 );
xnor U18897 ( n1473, n61, n1474 );
nand U18898 ( n1403, n1404, n1406 );
nand U18899 ( n1406, n1187, n1407 );
nand U18900 ( n1404, n70, n1409 );
xnor U18901 ( n1407, n62, n1408 );
nand U18902 ( n1388, n1389, n1391 );
nand U18903 ( n1391, n11284, n1392 );
nand U18904 ( n1389, n70, n1394 );
xnor U18905 ( n1392, n63, n1393 );
nand U18906 ( n1328, n1329, n1330 );
nand U18907 ( n1330, n11285, n1331 );
nand U18908 ( n1329, n70, n1339 );
nand U18909 ( n1331, n1332, n1333 );
nand U18910 ( n1208, n1209, n1211 );
nand U18911 ( n1211, n11284, n1212 );
nand U18912 ( n1209, n70, n1221 );
nand U18913 ( n1212, n1213, n1214 );
nand U18914 ( n1000, n10792, n10793 );
nor U18915 ( n10792, n10813, n10814 );
nor U18916 ( n10793, n10794, n10795 );
nor U18917 ( n10814, n11533, n10972 );
nand U18918 ( n915, n1644, n1646 );
nor U18919 ( n1644, n1657, n1658 );
nor U18920 ( n1646, n1647, n1648 );
nor U18921 ( n1657, n71, n11106 );
nand U18922 ( n5583, n5584, n853 );
xnor U18923 ( n5584, n5585, n5586 );
and U18924 ( n1567, n1576, n69 );
and U18925 ( n1613, n1629, n69 );
and U18926 ( n1353, n1369, n69 );
and U18927 ( n1282, n1304, n69 );
xor U18928 ( n2068, n10565, n11077 );
nor U18929 ( n10574, n10583, n11072 );
nor U18930 ( n10639, n10648, n11042 );
nor U18931 ( n10621, n10630, n11059 );
nor U18932 ( n10592, n10601, n11066 );
xor U18933 ( n2343, n10684, n11026 );
nor U18934 ( n6748, n11354, n11148 );
and U18935 ( n8466, n11283, n7614 );
and U18936 ( n7327, n11534, n7330 );
nor U18937 ( n4438, n4440, n10968 );
nand U18938 ( n4716, n8203, n6643 );
nor U18939 ( n8203, n6645, n6511 );
nor U18940 ( n10556, n11077, n10565 );
xor U18941 ( n2293, n10666, n11030 );
not U18942 ( n1149, n6113 );
xor U18943 ( n2203, n10630, n11059 );
nor U18944 ( n6642, n4743, n4738 );
nand U18945 ( n1558, n1789, n1791 );
nand U18946 ( n1791, n1792, n1793 );
nand U18947 ( n1789, n1802, n372 );
nand U18948 ( n1793, n1794, n1796 );
nand U18949 ( n1477, n1806, n1807 );
nand U18950 ( n1807, n1808, n1809 );
nand U18951 ( n1806, n1818, n379 );
nand U18952 ( n1809, n1811, n1812 );
nand U18953 ( n1639, n1606, n1607 );
nand U18954 ( n1346, n1831, n1832 );
nand U18955 ( n1832, n1316, n1304 );
nor U18956 ( n1831, n1833, n1834 );
nor U18957 ( n1834, n1836, n11012 );
nand U18958 ( n1772, n1773, n1774 );
nand U18959 ( n1774, n1641, n1629 );
nor U18960 ( n1773, n1776, n1777 );
nor U18961 ( n1777, n1778, n11085 );
nand U18962 ( n1462, n1822, n1823 );
nand U18963 ( n1823, n1381, n1369 );
nor U18964 ( n1822, n1824, n1826 );
nor U18965 ( n1826, n1827, n11025 );
nor U18966 ( n1759, n1761, n1762 );
nor U18967 ( n1762, n1763, n1764 );
nor U18968 ( n1761, n357, n1769 );
nand U18969 ( n1764, n1766, n1767 );
nor U18970 ( n6499, n5009, n4705 );
and U18971 ( n8492, n11283, n7707 );
nand U18972 ( n4424, n4425, n4044 );
nand U18973 ( n4116, n4117, n4044 );
nand U18974 ( n4530, n4531, n4044 );
nand U18975 ( n4288, n4289, n4044 );
nand U18976 ( n4494, n4495, n4044 );
nand U18977 ( n4082, n4083, n4044 );
nand U18978 ( n4157, n4158, n4044 );
nand U18979 ( n4562, n4563, n4044 );
nand U18980 ( n4370, n4371, n4044 );
nand U18981 ( n4331, n4332, n4044 );
nand U18982 ( n4720, n4721, n4044 );
nand U18983 ( n1189, n1756, n1757 );
nand U18984 ( n1757, n1254, n1758 );
not U18985 ( n409, n1853 );
nand U18986 ( n1554, n1697, n1698 );
nand U18987 ( n1698, n1699, n1701 );
nand U18988 ( n1697, n1711, n373 );
nand U18989 ( n1701, n1702, n1703 );
nand U18990 ( n1627, n1597, n1598 );
nand U18991 ( n1337, n1738, n1739 );
nand U18992 ( n1739, n1297, n1304 );
nor U18993 ( n1738, n1741, n1742 );
nor U18994 ( n1742, n1743, n11011 );
nand U18995 ( n1758, n409, n10974 );
nand U18996 ( n1679, n1682, n1683 );
nand U18997 ( n1683, n1628, n1629 );
nor U18998 ( n1682, n1684, n1686 );
nor U18999 ( n1686, n1687, n11084 );
nand U19000 ( n1441, n1731, n1732 );
nand U19001 ( n1732, n1368, n1369 );
nor U19002 ( n1731, n1733, n1734 );
nor U19003 ( n1734, n1736, n11024 );
nand U19004 ( n1524, n1714, n1716 );
nand U19005 ( n1716, n1717, n1718 );
nand U19006 ( n1714, n1727, n381 );
nand U19007 ( n1718, n1719, n1721 );
nand U19008 ( n1768, n1681, n1772 );
nand U19009 ( n1767, n1768, n11093 );
not U19010 ( n861, n5424 );
nand U19011 ( n4043, n4044, n4045 );
nand U19012 ( n4215, n4044, n4216 );
nand U19013 ( n4584, n4044, n4585 );
nand U19014 ( n4348, n4044, n4349 );
nand U19015 ( n4408, n4044, n4409 );
nand U19016 ( n4140, n4044, n10958 );
not U19017 ( n859, n5412 );
and U19018 ( n8249, n11534, n8252 );
not U19019 ( n407, n1854 );
nand U19020 ( n1219, n407, n10981 );
nor U19021 ( n1236, n1264, n1194 );
nor U19022 ( n1264, n1266, n1267 );
nor U19023 ( n1266, n1271, n1272 );
nor U19024 ( n1267, n65, n1268 );
nand U19025 ( n1228, n407, n10982 );
not U19026 ( n862, n5459 );
nand U19027 ( n8614, n9367, n9366 );
nor U19028 ( n9367, n1249, n109 );
nor U19029 ( n1669, n1671, n1672 );
nand U19030 ( n1672, n1673, n1674 );
nand U19031 ( n1674, n1676, n11092 );
nand U19032 ( n1676, n1681, n1679 );
nor U19033 ( n10281, n10273, n10283 );
nand U19034 ( n10283, n10270, n1176 );
not U19035 ( n371, n9800 );
not U19036 ( n777, n10273 );
not U19037 ( n946, n4733 );
nand U19038 ( n5877, n963, n5795 );
not U19039 ( n963, n5881 );
nor U19040 ( n5879, n5763, n5882 );
nor U19041 ( n5882, n5883, n5884 );
nand U19042 ( n5884, n888, n5743 );
xor U19043 ( n2023, n10547, n11100 );
not U19044 ( n898, n8410 );
nand U19045 ( n5790, n5768, n5769 );
xor U19046 ( n2119, n10583, n11072 );
nor U19047 ( n9381, n9382, n9356 );
nor U19048 ( n9382, n336, n9383 );
nand U19049 ( n9383, n2774, n2713 );
and U19050 ( n9226, n9379, n9380 );
nor U19051 ( n9379, n9388, n332 );
nor U19052 ( n9380, n2536, n9381 );
nor U19053 ( n9388, n9389, n9387 );
nor U19054 ( n6635, n6511, n6638 );
nand U19055 ( n6638, n6639, n4742 );
nand U19056 ( n6639, n6640, n6641 );
nand U19057 ( n6641, n6642, n4769 );
and U19058 ( n4007, n6098, n11527 );
nand U19059 ( n6098, n11385, n4733 );
not U19060 ( n284, n1249 );
not U19061 ( n864, n5488 );
nor U19062 ( n1303, n10981, n407 );
nor U19063 ( n1321, n10982, n407 );
nor U19064 ( n5763, n5769, n5768 );
xor U19065 ( n2164, n10601, n11066 );
nor U19066 ( n3982, n341, n9356 );
xor U19067 ( n1978, n10529, n11108 );
nor U19068 ( n10538, n11100, n10547 );
nor U19069 ( n10520, n11108, n10529 );
xnor U19070 ( n4713, n11459, n5314 );
nor U19071 ( n4741, n938, n5009 );
and U19072 ( n8499, n11283, n7745 );
and U19073 ( n8257, n11534, n8258 );
nor U19074 ( n10486, n10495, n11121 );
nor U19075 ( n9385, n341, n353 );
not U19076 ( n403, n1273 );
nor U19077 ( n1297, n11007, n403 );
nor U19078 ( n1743, n1297, n1304 );
nor U19079 ( n1316, n11009, n403 );
nor U19080 ( n1836, n1316, n1304 );
xor U19081 ( n1933, n10495, n11121 );
nor U19082 ( n10813, n71, n10962 );
nand U19083 ( n6110, n6656, n11402 );
nor U19084 ( n6656, n1004, n6657 );
nand U19085 ( n1263, n403, n11007 );
nand U19086 ( n1269, n403, n11009 );
not U19087 ( n867, n5508 );
not U19088 ( n52, n1606 );
nand U19089 ( n9216, n9373, n9374 );
nor U19090 ( n9374, n9375, n2551 );
nor U19091 ( n9373, n9377, n9378 );
nor U19092 ( n9377, n9226, n9225 );
nand U19093 ( n5880, n894, n5881 );
and U19094 ( n8516, n11283, n7849 );
and U19095 ( n8509, n11283, n7792 );
and U19096 ( n8273, n11534, n8274 );
not U19097 ( n59, n1597 );
and U19098 ( n8263, n11534, n8266 );
buf U19099 ( n11529, n11531 );
and U19100 ( n11248, n3969, n3970 );
nand U19101 ( n9081, n2137, n8618 );
nand U19102 ( n8877, n2181, n8618 );
nand U19103 ( n8648, n2227, n8618 );
nand U19104 ( n8839, n2271, n8618 );
nand U19105 ( n8685, n2317, n8618 );
nand U19106 ( n8782, n2361, n8618 );
nand U19107 ( n9098, n2403, n8618 );
nand U19108 ( n8941, n2448, n8618 );
not U19109 ( n1009, n5314 );
and U19110 ( n8526, n11283, n7900 );
nand U19111 ( n1599, n1601, n1602 );
nand U19112 ( n1601, n1604, n1606 );
nand U19113 ( n1602, n1603, n52 );
nand U19114 ( n1604, n363, n1607 );
not U19115 ( n872, n5559 );
nand U19116 ( n5456, n5457, n857 );
xnor U19117 ( n5457, n5458, n5459 );
and U19118 ( n8380, n11534, n8383 );
nand U19119 ( n6640, n928, n5009 );
not U19120 ( n393, n1829 );
nor U19121 ( n1368, n11020, n393 );
nor U19122 ( n1736, n1368, n1369 );
nor U19123 ( n1381, n11023, n393 );
nor U19124 ( n1827, n1381, n1369 );
nor U19125 ( n8145, n939, n929 );
nand U19126 ( n1592, n1596, n1597 );
nand U19127 ( n1596, n364, n1598 );
nand U19128 ( n4710, n4735, n4736 );
nor U19129 ( n4735, n4740, n4741 );
nor U19130 ( n4736, n917, n4737 );
nor U19131 ( n4740, n4742, n4743 );
nand U19132 ( n1338, n393, n11020 );
nand U19133 ( n1347, n393, n11023 );
not U19134 ( n874, n5586 );
nor U19135 ( n4737, n4738, n4739 );
nor U19136 ( n8142, n4769, n5009 );
not U19137 ( n858, n5445 );
not U19138 ( n53, n1538 );
nor U19139 ( n1526, n1527, n1528 );
nor U19140 ( n1528, n1529, n1531 );
nor U19141 ( n1527, n376, n1536 );
nand U19142 ( n1531, n1532, n1533 );
and U19143 ( n8533, n11283, n7951 );
and U19144 ( n8474, n11535, n8475 );
xor U19145 ( n5484, n5487, n5488 );
xor U19146 ( n5610, n5613, n5614 );
nor U19147 ( n2536, n2658, n9384 );
nand U19148 ( n1534, n1519, n1538 );
nand U19149 ( n1533, n1534, n11051 );
not U19150 ( n60, n1518 );
not U19151 ( n388, n1436 );
nand U19152 ( n1724, n1728, n1717 );
nand U19153 ( n1728, n388, n11044 );
nand U19154 ( n1816, n1819, n1808 );
nand U19155 ( n1819, n388, n11045 );
not U19156 ( n907, n4769 );
nor U19157 ( n1508, n1509, n1511 );
nand U19158 ( n1511, n1512, n1513 );
nand U19159 ( n1513, n1514, n11049 );
nand U19160 ( n1514, n1519, n1518 );
not U19161 ( n382, n1443 );
nand U19162 ( n1717, n382, n11041 );
nand U19163 ( n1808, n382, n11043 );
not U19164 ( n876, n5614 );
xnor U19165 ( n5633, n878, n5634 );
xnor U19166 ( n5506, n5507, n5508 );
nand U19167 ( n5313, n11460, n5314 );
and U19168 ( n8543, n11530, n7994 );
and U19169 ( n8567, n11535, n8570 );
xnor U19170 ( n5742, n5743, n5744 );
and U19171 ( n8551, n11530, n8032 );
and U19172 ( n8667, n11535, n8668 );
not U19173 ( n878, n5635 );
and U19174 ( n2534, n9398, n341 );
nor U19175 ( n9398, n353, n9356 );
nand U19176 ( n4745, n6497, n6498 );
nand U19177 ( n6498, n6499, n4743 );
nand U19178 ( n5864, n5866, n5867 );
nand U19179 ( n5867, n5868, n11287 );
nand U19180 ( n5866, n5870, n11460 );
nor U19181 ( n8561, n8067, n11450 );
buf U19182 ( n11323, n11322 );
not U19183 ( n55, n1457 );
nor U19184 ( n1444, n1446, n1447 );
nor U19185 ( n1447, n1448, n1449 );
nor U19186 ( n1446, n383, n1454 );
nand U19187 ( n1449, n1451, n1452 );
nor U19188 ( n8573, n11449, n8578 );
nand U19189 ( n8578, n8106, n8105 );
and U19190 ( n9047, n11535, n9048 );
nand U19191 ( n1453, n1436, n1457 );
nand U19192 ( n1452, n1453, n11045 );
not U19193 ( n62, n1434 );
not U19194 ( n374, n1519 );
nand U19195 ( n1708, n1699, n1712 );
nand U19196 ( n1712, n374, n11049 );
nand U19197 ( n1799, n1792, n1803 );
nand U19198 ( n1803, n374, n11051 );
nor U19199 ( n1254, n10964, n10957 );
nor U19200 ( n1424, n1426, n1427 );
nand U19201 ( n1427, n1428, n1429 );
nand U19202 ( n1429, n1431, n11044 );
nand U19203 ( n1431, n1436, n1434 );
not U19204 ( n378, n1704 );
nand U19205 ( n1699, n378, n11046 );
nand U19206 ( n1792, n378, n11047 );
nand U19207 ( n6497, n8137, n939 );
nor U19208 ( n8137, n4738, n4769 );
nor U19209 ( n4433, n4434, n11408 );
nor U19210 ( n4434, n4435, n11490 );
buf U19211 ( n11408, n11407 );
not U19212 ( n73, n9562 );
and U19213 ( n8880, n11535, n8883 );
nand U19214 ( n5411, n5412, n11460 );
not U19215 ( n884, n5685 );
nand U19216 ( n1253, n1249, n10803 );
nand U19217 ( n10455, n10456, n10457 );
nor U19218 ( n10457, n341, n9378 );
nor U19219 ( n10456, n1253, n348 );
and U19220 ( n8583, n11530, n8127 );
and U19221 ( n10500, n11535, n9978 );
nand U19222 ( n6718, n8138, n939 );
nor U19223 ( n8138, n907, n4743 );
nor U19224 ( n305, n3987, n11128 );
nor U19225 ( n380, n3987, n11129 );
not U19226 ( n282, n10803 );
not U19227 ( n886, n5701 );
nand U19228 ( n10454, n341, n9378 );
xnor U19229 ( n5560, n5561, n5562 );
xnor U19230 ( n5562, n11000, n872 );
nor U19231 ( n1530, n8253, n11134 );
nor U19232 ( n1605, n8253, n11135 );
not U19233 ( n888, n5744 );
not U19234 ( n887, n5721 );
not U19235 ( n366, n1781 );
nor U19236 ( n1628, n11075, n366 );
nor U19237 ( n1687, n1628, n1629 );
nor U19238 ( n1641, n11076, n366 );
nor U19239 ( n1778, n1641, n1629 );
nand U19240 ( n1339, n1341, n1342 );
nand U19241 ( n1341, n1344, n1346 );
nand U19242 ( n1342, n1343, n57 );
nand U19243 ( n1344, n391, n1347 );
nand U19244 ( n1598, n366, n11075 );
nand U19245 ( n1607, n366, n11076 );
not U19246 ( n894, n5795 );
nand U19247 ( n1271, n404, n1317 );
nand U19248 ( n1317, n1228, n1226 );
nand U19249 ( n5312, n4733, n11527 );
xnor U19250 ( n1671, n359, n11086 );
xnor U19251 ( n1763, n359, n11087 );
nand U19252 ( n4016, n4017, n3998 );
nand U19253 ( n1262, n406, n1298 );
nand U19254 ( n1298, n1219, n1217 );
nor U19255 ( n1383, P1_STATE_REG, n10955 );
buf U19256 ( n11324, n11322 );
not U19257 ( n387, n1479 );
not U19258 ( n389, n1442 );
not U19259 ( n361, n1681 );
xnor U19260 ( n5868, n4769, n11079 );
nand U19261 ( n8325, n8175, n8305 );
not U19262 ( n896, n5817 );
nand U19263 ( n1221, n1222, n1223 );
nand U19264 ( n1222, n1227, n1226 );
nand U19265 ( n1223, n1224, n66 );
nand U19266 ( n1227, n1228, n404 );
not U19267 ( n66, n1226 );
nand U19268 ( n5366, n5367, n116 );
xor U19269 ( n1622, n1629, n11084 );
xor U19270 ( n1634, n1629, n11085 );
nand U19271 ( n8333, n8164, n8163 );
nand U19272 ( n8350, n8293, n8292 );
nand U19273 ( n1213, n1218, n1217 );
nand U19274 ( n1218, n1219, n406 );
not U19275 ( n897, n5837 );
buf U19276 ( n11409, n11407 );
xor U19277 ( n1362, n1369, n11024 );
xor U19278 ( n1291, n1304, n11011 );
xor U19279 ( n1374, n1369, n11025 );
xor U19280 ( n1309, n1304, n11012 );
nand U19281 ( n5393, n5394, n5395 );
xnor U19282 ( n1509, n378, n11046 );
xnor U19283 ( n1529, n378, n11047 );
nand U19284 ( n8368, n8300, n957 );
nor U19285 ( n1643, n11533, n11066 );
nor U19286 ( n1544, n11533, n11042 );
nor U19287 ( n1482, n11533, n11030 );
nor U19288 ( n1413, n11533, n11026 );
nor U19289 ( n1323, n11533, n11003 );
nor U19290 ( n1232, n11533, n11002 );
nor U19291 ( n1857, n11533, n11072 );
nor U19292 ( n1582, P1_STATE_REG, n11059 );
nor U19293 ( n4137, n11527, n10958 );
nor U19294 ( n4405, n11527, n10970 );
nor U19295 ( n5467, n11527, n10992 );
not U19296 ( n369, n1561 );
not U19297 ( n893, n5769 );
not U19298 ( n871, n5533 );
xnor U19299 ( n1574, n1576, n11067 );
not U19300 ( n882, n5660 );
not U19301 ( n383, n1448 );
nand U19302 ( n6181, n6182, n354 );
nand U19303 ( n10799, n1756, n1758 );
nand U19304 ( n8391, n8202, n8201 );
nand U19305 ( n6308, n6309, n6310 );
nand U19306 ( n8408, n8197, n8196 );
nand U19307 ( n6436, n6437, n6438 );
nand U19308 ( n8426, n7387, n898 );
nand U19309 ( n6573, n6574, n6575 );
nand U19310 ( n6734, n6735, n371 );
nand U19311 ( n8443, n7495, n7494 );
buf U19312 ( n11535, n11536 );
buf U19313 ( n11530, n11531 );
nand U19314 ( n8461, n7581, n889 );
nand U19315 ( n7798, n7799, n7800 );
nand U19316 ( n8259, n8260, n386 );
nand U19317 ( n8485, n7656, n7655 );
nand U19318 ( n8503, n7749, n883 );
nand U19319 ( n8275, n8276, n8277 );
nand U19320 ( n8476, n8477, n394 );
nand U19321 ( n8520, n7854, n7853 );
nand U19322 ( n8537, n7956, n7955 );
nand U19323 ( n8669, n8670, n8671 );
nand U19324 ( n8555, n8031, n873 );
nand U19325 ( n9049, n9050, n9051 );
nand U19326 ( n9991, n10425, n10426 );
nand U19327 ( n10426, SI_1_, n10427 );
nand U19328 ( n9892, n10409, n10410 );
nand U19329 ( n10409, n10063, n10065 );
nand U19330 ( n10410, SI_6_, n10411 );
or U19331 ( n10411, n10065, n10063 );
nand U19332 ( n9848, n10398, n10399 );
nand U19333 ( n10398, n10119, n10121 );
nand U19334 ( n10399, SI_10_, n10400 );
or U19335 ( n10400, n10121, n10119 );
nand U19336 ( n10014, n10418, n10419 );
nand U19337 ( n10418, SI_3_, n10029 );
nand U19338 ( n10419, n10027, n10420 );
or U19339 ( n10420, n10029, SI_3_ );
nand U19340 ( n10135, n10383, n10384 );
nand U19341 ( n10383, n9795, n9797 );
nand U19342 ( n10384, SI_15_, n10385 );
or U19343 ( n10385, n9797, n9795 );
nand U19344 ( n9777, n10373, n10374 );
nand U19345 ( n10373, n9763, n9765 );
nand U19346 ( n10374, SI_17_, n10375 );
or U19347 ( n10375, n9765, n9763 );
nand U19348 ( n10148, n10363, n10364 );
nand U19349 ( n10363, n9734, n9736 );
nand U19350 ( n10364, SI_19_, n10365 );
or U19351 ( n10365, n9736, n9734 );
nand U19352 ( n10187, n10353, n10354 );
nand U19353 ( n10353, n10156, n10158 );
nand U19354 ( n10354, SI_21_, n10355 );
or U19355 ( n10355, n10158, n10156 );
nand U19356 ( n10200, n10343, n10344 );
nand U19357 ( n10343, n10177, n10179 );
nand U19358 ( n10344, SI_23_, n10345 );
or U19359 ( n10345, n10179, n10177 );
nand U19360 ( n10231, n10333, n10334 );
nand U19361 ( n10333, n10221, n10223 );
nand U19362 ( n10334, SI_25_, n10335 );
or U19363 ( n10335, n10223, n10221 );
nand U19364 ( n10302, n10312, n10313 );
nand U19365 ( n10312, n10316, n10315 );
nand U19366 ( n10313, SI_27_, n10314 );
or U19367 ( n10314, n10315, n10316 );
nand U19368 ( n9795, n10388, n10389 );
nand U19369 ( n10388, SI_14_, n9817 );
nand U19370 ( n10389, n10390, n10391 );
or U19371 ( n10391, n9817, SI_14_ );
nand U19372 ( n10063, n10414, n10415 );
nand U19373 ( n10414, SI_5_, n10052 );
nand U19374 ( n10415, n10047, n10416 );
or U19375 ( n10416, n10052, SI_5_ );
nand U19376 ( n10119, n10403, n10404 );
nand U19377 ( n10403, SI_9_, n9931 );
nand U19378 ( n10404, n9929, n10405 );
or U19379 ( n10405, n9931, SI_9_ );
nand U19380 ( n9763, n10378, n10379 );
nand U19381 ( n10378, n10135, n10136 );
nand U19382 ( n10379, SI_16_, n10380 );
or U19383 ( n10380, n10136, n10135 );
nand U19384 ( n9734, n10368, n10369 );
nand U19385 ( n10368, n9777, n9778 );
nand U19386 ( n10369, SI_18_, n10370 );
or U19387 ( n10370, n9778, n9777 );
nand U19388 ( n10156, n10358, n10359 );
nand U19389 ( n10358, n10148, n10149 );
nand U19390 ( n10359, SI_20_, n10360 );
or U19391 ( n10360, n10149, n10148 );
nand U19392 ( n10177, n10348, n10349 );
nand U19393 ( n10348, n10187, n10188 );
nand U19394 ( n10349, SI_22_, n10350 );
or U19395 ( n10350, n10188, n10187 );
nand U19396 ( n10221, n10338, n10339 );
nand U19397 ( n10338, n10200, n10201 );
nand U19398 ( n10339, SI_24_, n10340 );
or U19399 ( n10340, n10201, n10200 );
nand U19400 ( n10316, n10328, n10329 );
nand U19401 ( n10328, n10231, n10232 );
nand U19402 ( n10329, SI_26_, n10330 );
or U19403 ( n10330, n10232, n10231 );
nand U19404 ( n10280, n10298, n10299 );
nand U19405 ( n10298, n10302, n10301 );
nand U19406 ( n10299, SI_28_, n10300 );
or U19407 ( n10300, n10301, n10302 );
nand U19408 ( n10513, n10609, n10610 );
nand U19409 ( n10610, P1_DATAO_REG_0_, n11330 );
nand U19410 ( n10609, P2_DATAO_REG_0_, n11325 );
nand U19411 ( n10027, n10421, n9992 );
nand U19412 ( n10421, n9991, n10422 );
or U19413 ( n10422, n9996, SI_2_ );
nand U19414 ( n9929, n10406, n10407 );
and U19415 ( n10406, n10435, n10436 );
nand U19416 ( n10407, n10408, n9892 );
nand U19417 ( n10435, SI_8_, n9916 );
not U19418 ( n11336, n8308 );
nand U19419 ( n8308, n10611, n10612 );
nand U19420 ( n10612, n10613, n10959 );
nand U19421 ( n10611, n10614, P2_ADDR_REG_19_ );
nand U19422 ( n10509, SI_0_, n10513 );
nand U19423 ( n3999, n10264, n10265 );
nand U19424 ( n10265, P2_DATAO_REG_31_, n11265 );
nand U19425 ( n10264, n8309, n8308 );
nor U19426 ( n10614, P2_RD_REG, n10959 );
nand U19427 ( n10258, n10276, n10277 );
nand U19428 ( n10276, n10280, n10279 );
nand U19429 ( n10277, SI_29_, n10278 );
or U19430 ( n10278, n10279, n10280 );
nand U19431 ( n10510, n10511, n10512 );
nand U19432 ( n10512, P1_DATAO_REG_1_, n11330 );
nand U19433 ( n10511, P2_DATAO_REG_1_, n11325 );
nor U19434 ( n10613, P2_ADDR_REG_19_, P1_RD_REG );
nand U19435 ( n9996, n10423, n10424 );
nand U19436 ( n10424, P1_DATAO_REG_2_, n11330 );
nand U19437 ( n10423, P2_DATAO_REG_2_, n11326 );
xor U19438 ( n8317, n10257, n10258 );
xnor U19439 ( n10257, SI_30_, n777 );
and U19440 ( n4006, n10255, n10256 );
nand U19441 ( n10255, P2_DATAO_REG_30_, n11265 );
nand U19442 ( n10256, n8317, n8308 );
nand U19443 ( n7800, n10853, n10090 );
nor U19444 ( n10853, P1_IR_REG_12_, P1_IR_REG_11_ );
nand U19445 ( n8277, n10855, n9897 );
nor U19446 ( n10855, P1_IR_REG_8_, P1_IR_REG_7_ );
nand U19447 ( n8671, n10857, n408 );
nor U19448 ( n10857, P1_IR_REG_4_, P1_IR_REG_3_ );
nand U19449 ( n6575, n10851, n9800 );
nor U19450 ( n10851, P1_IR_REG_16_, P1_IR_REG_15_ );
nand U19451 ( n4435, n10843, n10844 );
nor U19452 ( n10843, P1_IR_REG_26_, P1_IR_REG_25_ );
nor U19453 ( n10090, n10854, n8277 );
or U19454 ( n10854, P1_IR_REG_9_, P1_IR_REG_10_ );
nor U19455 ( n9800, n10852, n7800 );
or U19456 ( n10852, P1_IR_REG_14_, P1_IR_REG_13_ );
nor U19457 ( n9897, n10856, n8671 );
or U19458 ( n10856, P1_IR_REG_6_, P1_IR_REG_5_ );
or U19459 ( n6438, n11249, n6575 );
or U19460 ( n11249, P1_IR_REG_18_, P1_IR_REG_17_ );
nor U19461 ( n10828, n6310, P1_IR_REG_20_ );
nand U19462 ( n2533, n9953, n9954 );
nand U19463 ( n9954, n9955, n11420 );
nand U19464 ( n9953, P1_IR_REG_0_, n11419 );
nand U19465 ( n9051, n10858, n10957 );
nor U19466 ( n10858, P1_IR_REG_2_, P1_IR_REG_1_ );
nand U19467 ( n10832, n10849, n10828 );
nor U19468 ( n10849, P1_IR_REG_22_, P1_IR_REG_21_ );
nand U19469 ( n4222, n10819, n10776 );
nand U19470 ( n10819, P1_IR_REG_28_, n10821 );
nand U19471 ( n10821, n327, n10961 );
nor U19472 ( n10844, n5395, P1_IR_REG_24_ );
nand U19473 ( n9292, n9293, n9294 );
nand U19474 ( n9294, P1_IR_REG_0_, n87 );
nor U19475 ( n9293, n9295, n9296 );
nor U19476 ( n9296, n286, n8753 );
or U19477 ( n6310, n6438, P1_IR_REG_19_ );
or U19478 ( n5395, n10832, P1_IR_REG_23_ );
nand U19479 ( n1249, n10817, n10818 );
nand U19480 ( n10817, P1_IR_REG_28_, n11487 );
or U19481 ( n10818, n4222, n11484 );
nand U19482 ( n1280, n8719, n8720 );
nor U19483 ( n8719, n8765, n8766 );
nor U19484 ( n8720, n8721, n8722 );
and U19485 ( n8765, n11535, P1_REG3_REG_28_ );
nand U19486 ( n9992, SI_2_, n9996 );
nand U19487 ( n6650, n8306, n8307 );
nand U19488 ( n8307, P1_DATAO_REG_31_, n8308 );
nand U19489 ( n8306, n8309, n11267 );
nand U19490 ( n10029, n10428, n10429 );
nand U19491 ( n10429, P1_DATAO_REG_3_, n11330 );
nand U19492 ( n10428, P2_DATAO_REG_3_, n11326 );
nand U19493 ( n10776, n10820, n327 );
nor U19494 ( n10820, P1_IR_REG_28_, P1_IR_REG_27_ );
nand U19495 ( n1180, n9099, n9100 );
nor U19496 ( n9099, n9209, n9210 );
nor U19497 ( n9100, n9101, n9102 );
and U19498 ( n9209, n11535, P1_REG3_REG_26_ );
nand U19499 ( n10012, n10430, n10431 );
nand U19500 ( n10431, P1_DATAO_REG_4_, n11330 );
nand U19501 ( n10430, P2_DATAO_REG_4_, n11326 );
or U19502 ( n10049, n10012, SI_4_ );
nand U19503 ( n10803, n10822, n10823 );
nand U19504 ( n10823, P1_IR_REG_27_, n10824 );
nand U19505 ( n10822, n4429, P1_IR_REG_31_ );
nand U19506 ( n10824, P1_IR_REG_31_, n4435 );
nor U19507 ( n4429, P1_IR_REG_27_, n327 );
and U19508 ( n6655, n8315, n8316 );
nand U19509 ( n8315, P1_DATAO_REG_30_, n11327 );
nand U19510 ( n8316, n11333, n8317 );
xnor U19511 ( n8324, n10280, n10295 );
xnor U19512 ( n10295, SI_29_, n10279 );
and U19513 ( n4015, n10293, n10294 );
nand U19514 ( n10293, P2_DATAO_REG_29_, n11266 );
nand U19515 ( n10294, n8324, n11328 );
nand U19516 ( n10051, SI_4_, n10012 );
nand U19517 ( n735, n2560, n2561 );
nand U19518 ( n2560, P1_REG1_REG_29_, n11426 );
nand U19519 ( n2561, n11279, n2562 );
nand U19520 ( n575, n2676, n2677 );
nand U19521 ( n2676, P1_REG0_REG_29_, n11422 );
nand U19522 ( n2677, n11276, n2562 );
xor U19523 ( n8159, n1011, P2_IR_REG_27_ );
nand U19524 ( n7494, n8444, n8445 );
nor U19525 ( n8444, P2_IR_REG_16_, P2_IR_REG_15_ );
nand U19526 ( n7655, n8486, n8487 );
nor U19527 ( n8486, P2_IR_REG_12_, P2_IR_REG_11_ );
nand U19528 ( n7853, n8521, n1013 );
nor U19529 ( n8521, P2_IR_REG_8_, P2_IR_REG_7_ );
nand U19530 ( n8105, n8579, n10960 );
nor U19531 ( n8579, P2_IR_REG_2_, P2_IR_REG_1_ );
or U19532 ( n8201, n11250, n8196 );
or U19533 ( n11250, P2_IR_REG_22_, P2_IR_REG_21_ );
nand U19534 ( n8196, n8409, n8410 );
nor U19535 ( n8409, P2_IR_REG_20_, P2_IR_REG_19_ );
nor U19536 ( n8445, n8462, n7655 );
or U19537 ( n8462, P2_IR_REG_14_, P2_IR_REG_13_ );
nor U19538 ( n8410, n8427, n7494 );
or U19539 ( n8427, P2_IR_REG_18_, P2_IR_REG_17_ );
nor U19540 ( n8487, n8504, n7853 );
or U19541 ( n8504, P2_IR_REG_9_, P2_IR_REG_10_ );
nand U19542 ( n8292, n8351, n8352 );
nor U19543 ( n8351, P2_IR_REG_26_, P2_IR_REG_25_ );
nand U19544 ( n5007, n8154, n8155 );
nand U19545 ( n8155, n8156, n11384 );
nand U19546 ( n8154, P2_IR_REG_0_, n11383 );
nand U19547 ( n7955, n8538, n8539 );
nor U19548 ( n8538, P2_IR_REG_6_, P2_IR_REG_5_ );
nor U19549 ( n8539, n8556, n8105 );
or U19550 ( n8556, P2_IR_REG_4_, P2_IR_REG_3_ );
nor U19551 ( n8352, n8369, n8201 );
or U19552 ( n8369, P2_IR_REG_24_, P2_IR_REG_23_ );
nand U19553 ( n1950, n6529, n6530 );
nand U19554 ( n6529, P2_REG1_REG_27_, n11359 );
nand U19555 ( n6530, n11273, n6531 );
nand U19556 ( n1790, n6793, n6794 );
nand U19557 ( n6793, P2_REG0_REG_27_, n11355 );
nand U19558 ( n6794, n11270, n6531 );
nand U19559 ( n10052, n10432, n10433 );
nand U19560 ( n10433, P1_DATAO_REG_5_, n11264 );
nand U19561 ( n10432, P2_DATAO_REG_5_, n11325 );
nand U19562 ( n5314, n8160, n8161 );
nand U19563 ( n8160, P2_IR_REG_28_, n11457 );
nand U19564 ( n8161, n8162, P2_IR_REG_31_ );
and U19565 ( n8162, n8163, n8164 );
nand U19566 ( n8163, n8334, n1011 );
nor U19567 ( n8334, P2_IR_REG_28_, P2_IR_REG_27_ );
xor U19568 ( n8349, n10230, n10231 );
xor U19569 ( n10230, SI_26_, n10232 );
and U19570 ( n6924, n8347, n8348 );
nand U19571 ( n8347, P1_DATAO_REG_26_, n11326 );
nand U19572 ( n8348, n11333, n8349 );
nand U19573 ( n1960, n6523, n6524 );
nand U19574 ( n6523, P2_REG1_REG_29_, n11359 );
nand U19575 ( n6524, n11273, n6525 );
nand U19576 ( n1800, n6667, n6668 );
nand U19577 ( n6667, P2_REG0_REG_29_, n11355 );
nand U19578 ( n6668, n11270, n6525 );
nand U19579 ( n8164, P2_IR_REG_28_, n8335 );
or U19580 ( n8335, n8292, P2_IR_REG_27_ );
xor U19581 ( n8332, n10311, n10302 );
xor U19582 ( n10311, SI_28_, n10301 );
and U19583 ( n6792, n8330, n8331 );
nand U19584 ( n8330, P1_DATAO_REG_28_, n8308 );
nand U19585 ( n8331, n11333, n8332 );
and U19586 ( n4223, n10309, n10310 );
nand U19587 ( n10309, P2_DATAO_REG_28_, n11266 );
nand U19588 ( n10310, n8332, n11327 );
xnor U19589 ( n8342, n10316, n10325 );
xnor U19590 ( n10325, SI_27_, n10315 );
and U19591 ( n4432, n10323, n10324 );
nand U19592 ( n10323, P2_DATAO_REG_27_, n11330 );
nand U19593 ( n10324, n8342, n11328 );
nand U19594 ( n1235, n8916, n8917 );
nor U19595 ( n8916, n8924, n8925 );
nor U19596 ( n8917, n8918, n8919 );
and U19597 ( n8924, n11535, P1_REG3_REG_24_ );
nand U19598 ( n1795, n6736, n6737 );
nand U19599 ( n6736, P2_REG0_REG_28_, n11355 );
nand U19600 ( n6737, n11270, n6528 );
nand U19601 ( n1955, n6526, n6527 );
nand U19602 ( n6526, P2_REG1_REG_28_, n6519 );
nand U19603 ( n6527, n11273, n6528 );
and U19604 ( n6728, n8322, n8323 );
nand U19605 ( n8322, P1_DATAO_REG_29_, n11328 );
nand U19606 ( n8323, n11333, n8324 );
nand U19607 ( n730, n2563, n2564 );
nand U19608 ( n2563, P1_REG1_REG_28_, n11426 );
nand U19609 ( n2564, n11279, n2565 );
nand U19610 ( n570, n2743, n2744 );
nand U19611 ( n2743, P1_REG0_REG_28_, n11422 );
nand U19612 ( n2744, n11276, n2565 );
nand U19613 ( n10065, n10412, n10413 );
nand U19614 ( n10413, P1_DATAO_REG_6_, n11330 );
nand U19615 ( n10412, P2_DATAO_REG_6_, n11326 );
xnor U19616 ( n8178, n8305, P2_IR_REG_30_ );
nand U19617 ( n8169, n8176, n8177 );
nand U19618 ( n8176, P2_IR_REG_30_, n11457 );
or U19619 ( n8177, n8178, n11455 );
or U19620 ( n8305, n8163, P2_IR_REG_29_ );
and U19621 ( n6861, n8340, n8341 );
nand U19622 ( n8340, P1_DATAO_REG_27_, n11327 );
nand U19623 ( n8341, n11333, n8342 );
and U19624 ( n9894, n10437, n10438 );
nand U19625 ( n10438, P1_DATAO_REG_7_, n11264 );
nand U19626 ( n10437, P2_DATAO_REG_7_, n11325 );
nand U19627 ( n9916, n10439, n10440 );
nand U19628 ( n10440, P1_DATAO_REG_8_, n11264 );
nand U19629 ( n10439, P2_DATAO_REG_8_, n11325 );
or U19630 ( n10434, n9916, SI_8_ );
and U19631 ( n4755, n10228, n10229 );
nand U19632 ( n10228, P2_DATAO_REG_26_, n11265 );
nand U19633 ( n10229, n8349, n8308 );
xnor U19634 ( n8360, n10221, n10222 );
xnor U19635 ( n10222, SI_25_, n10223 );
and U19636 ( n6975, n8358, n8359 );
nand U19637 ( n8358, P1_DATAO_REG_25_, n11325 );
nand U19638 ( n8359, n11333, n8360 );
nand U19639 ( n1945, n6538, n6539 );
nand U19640 ( n6538, P2_REG1_REG_26_, n11359 );
nand U19641 ( n6539, n11273, n6540 );
nand U19642 ( n1785, n6862, n6863 );
nand U19643 ( n6862, P2_REG0_REG_26_, n11355 );
nand U19644 ( n6863, n11270, n6540 );
nand U19645 ( n4754, n10842, n4435 );
nand U19646 ( n10842, P1_IR_REG_26_, n10845 );
or U19647 ( n10845, n116, P1_IR_REG_25_ );
nor U19648 ( n9402, n11251, n11252 );
and U19649 ( n11251, P1_IR_REG_26_, n11487 );
nor U19650 ( n11252, n4754, n11484 );
nand U19651 ( n745, n2553, n2554 );
nand U19652 ( n2553, P1_REG1_REG_31_, n2556 );
nand U19653 ( n2554, n11279, n2555 );
nand U19654 ( n585, n2653, n2654 );
nand U19655 ( n2653, P1_REG0_REG_31_, n2660 );
nand U19656 ( n2654, n11276, n2555 );
nand U19657 ( n9443, n10846, n10847 );
nand U19658 ( n10846, P1_IR_REG_24_, n11485 );
nand U19659 ( n10847, n10848, P1_IR_REG_31_ );
and U19660 ( n10848, n116, n5367 );
nand U19661 ( n8172, n8173, n8174 );
nand U19662 ( n8173, P2_IR_REG_29_, n11457 );
nand U19663 ( n8174, P2_IR_REG_31_, n8175 );
nand U19664 ( n8175, P2_IR_REG_29_, n8163 );
xnor U19665 ( n5339, P1_IR_REG_25_, n116 );
nand U19666 ( n9446, n10838, n10839 );
nand U19667 ( n10838, P1_IR_REG_25_, n11487 );
or U19668 ( n10839, n5339, n11484 );
nand U19669 ( n740, n2557, n2558 );
nand U19670 ( n2557, P1_REG1_REG_30_, n11426 );
nand U19671 ( n2558, n11279, n2559 );
nand U19672 ( n580, n2661, n2662 );
nand U19673 ( n2661, P1_REG0_REG_30_, n11422 );
nand U19674 ( n2662, n11276, n2559 );
xnor U19675 ( n4005, n3998, P1_IR_REG_30_ );
nand U19676 ( n10770, n10777, n10778 );
nand U19677 ( n10777, P1_IR_REG_30_, n11486 );
or U19678 ( n10778, n4005, n11484 );
or U19679 ( n3998, n10776, P1_IR_REG_29_ );
and U19680 ( n5340, n10219, n10220 );
nand U19681 ( n10219, P2_DATAO_REG_25_, n11265 );
nand U19682 ( n10220, n8360, n8308 );
nand U19683 ( n9931, n10441, n10442 );
nand U19684 ( n10442, P1_DATAO_REG_9_, n11264 );
nand U19685 ( n10441, P2_DATAO_REG_9_, n11325 );
nand U19686 ( n3970, n10461, n10462 );
nand U19687 ( n10461, P1_IR_REG_20_, n11486 );
nand U19688 ( n10462, n10463, P1_IR_REG_31_ );
and U19689 ( n10463, n354, n6182 );
nand U19690 ( n1930, n6547, n6548 );
nand U19691 ( n6547, P2_REG1_REG_23_, n11359 );
nand U19692 ( n6548, n11273, n6549 );
nand U19693 ( n1770, n7034, n7035 );
nand U19694 ( n7034, P2_REG0_REG_23_, n11355 );
nand U19695 ( n7035, n11270, n6549 );
xnor U19696 ( n8377, n10177, n10178 );
xnor U19697 ( n10178, SI_23_, n10179 );
and U19698 ( n5392, n10175, n10176 );
nand U19699 ( n10175, P2_DATAO_REG_23_, n11267 );
nand U19700 ( n10176, n8377, n11327 );
nand U19701 ( n565, n2805, n2806 );
nand U19702 ( n2805, P1_REG0_REG_27_, n2660 );
nand U19703 ( n2806, n11276, n2568 );
nand U19704 ( n725, n2566, n2567 );
nand U19705 ( n2566, P1_REG1_REG_27_, n2556 );
nand U19706 ( n2567, n11279, n2568 );
nand U19707 ( n10826, P1_IR_REG_21_, n11487 );
or U19708 ( n10827, n5809, n11484 );
xor U19709 ( n5809, n10828, P1_IR_REG_21_ );
and U19710 ( n7094, n8375, n8376 );
nand U19711 ( n8375, P1_DATAO_REG_23_, n11328 );
nand U19712 ( n8376, n11333, n8377 );
nand U19713 ( n5367, P1_IR_REG_24_, n5395 );
nand U19714 ( n10769, n10773, n10774 );
nand U19715 ( n10773, P1_IR_REG_29_, n11486 );
nand U19716 ( n10774, n10775, P1_IR_REG_31_ );
and U19717 ( n10775, n3998, n4017 );
and U19718 ( n10772, n11313, P1_REG0_REG_0_ );
xor U19719 ( n8390, n10186, n10187 );
xor U19720 ( n10186, SI_22_, n10188 );
and U19721 ( n7159, n8388, n8389 );
nand U19722 ( n8388, P1_DATAO_REG_22_, n11327 );
nand U19723 ( n8389, n11268, n8390 );
nand U19724 ( n1940, n6541, n6542 );
nand U19725 ( n6541, P2_REG1_REG_25_, n6519 );
nand U19726 ( n6542, n11273, n6543 );
nand U19727 ( n1780, n6925, n6926 );
nand U19728 ( n6925, P2_REG0_REG_25_, n11355 );
nand U19729 ( n6926, n11270, n6543 );
nor U19730 ( n8153, n11348, n10969 );
nand U19731 ( n1205, n9018, n9019 );
nor U19732 ( n9018, n9029, n9030 );
nor U19733 ( n9019, n9020, n9021 );
and U19734 ( n9029, n11535, P1_REG3_REG_22_ );
nand U19735 ( n1970, n6516, n6517 );
nand U19736 ( n6516, P2_REG1_REG_31_, n11359 );
nand U19737 ( n6517, n11273, n6518 );
nand U19738 ( n1810, n6646, n6647 );
nand U19739 ( n6646, P2_REG0_REG_31_, n6651 );
nand U19740 ( n6647, n11270, n6518 );
xnor U19741 ( n8400, n10156, n10157 );
xnor U19742 ( n10157, SI_21_, n10158 );
and U19743 ( n5810, n10154, n10155 );
nand U19744 ( n10154, P2_DATAO_REG_21_, n11267 );
nand U19745 ( n10155, n8400, n11327 );
nand U19746 ( n9384, n10458, n10459 );
nand U19747 ( n10458, P1_IR_REG_19_, n11486 );
nand U19748 ( n10459, n10460, P1_IR_REG_31_ );
and U19749 ( n10460, n6310, n6309 );
nand U19750 ( n6182, P1_IR_REG_20_, n6310 );
nand U19751 ( n715, n2572, n2573 );
nand U19752 ( n2572, P1_REG1_REG_25_, n2556 );
nand U19753 ( n2573, n11279, n2574 );
nand U19754 ( n555, n2918, n2919 );
nand U19755 ( n2918, P1_REG0_REG_25_, n2660 );
nand U19756 ( n2919, n11276, n2574 );
and U19757 ( n5574, n10184, n10185 );
nand U19758 ( n10184, P2_DATAO_REG_22_, n11267 );
nand U19759 ( n10185, n8390, n11327 );
nand U19760 ( n4017, P1_IR_REG_29_, n10776 );
xor U19761 ( n8367, n10199, n10200 );
xor U19762 ( n10199, SI_24_, n10201 );
and U19763 ( n7033, n8365, n8366 );
nand U19764 ( n8365, P1_DATAO_REG_24_, n8308 );
nand U19765 ( n8366, n11333, n8367 );
buf U19766 ( n11483, n421 );
not U19767 ( n421, P1_IR_REG_31_ );
nand U19768 ( n10108, n10447, n10448 );
nand U19769 ( n10448, P1_DATAO_REG_12_, n11330 );
nand U19770 ( n10447, P2_DATAO_REG_12_, n11325 );
nor U19771 ( n10397, n10108, SI_12_ );
nor U19772 ( n9824, n11253, n11254 );
and U19773 ( n11253, SI_12_, n10108 );
nor U19774 ( n11254, n10103, n10397 );
nand U19775 ( n6309, P1_IR_REG_19_, n6438 );
nand U19776 ( n10121, n10401, n10402 );
nand U19777 ( n10402, P1_DATAO_REG_10_, n11330 );
nand U19778 ( n10401, P2_DATAO_REG_10_, n11326 );
nand U19779 ( n7994, n8545, n8546 );
nand U19780 ( n8545, P1_DATAO_REG_5_, n11328 );
nand U19781 ( n8546, n11268, n8547 );
and U19782 ( n5365, n10197, n10198 );
nand U19783 ( n10197, P2_DATAO_REG_24_, n11265 );
nand U19784 ( n10198, n8367, n8308 );
nand U19785 ( n1215, n8968, n8969 );
nor U19786 ( n8968, n8986, n8987 );
nor U19787 ( n8969, n8970, n8971 );
and U19788 ( n8986, n11535, P1_REG3_REG_20_ );
nand U19789 ( n10087, n10445, n10446 );
nand U19790 ( n10446, P1_DATAO_REG_11_, n11264 );
nand U19791 ( n10445, P2_DATAO_REG_11_, n11325 );
nand U19792 ( n10103, SI_11_, n10087 );
nand U19793 ( n720, n2569, n2570 );
nand U19794 ( n2569, P1_REG1_REG_26_, n2556 );
nand U19795 ( n2570, n11279, n2571 );
nand U19796 ( n560, n2854, n2855 );
nand U19797 ( n2854, P1_REG0_REG_26_, n2660 );
nand U19798 ( n2855, n11276, n2571 );
nor U19799 ( n10107, n10087, SI_11_ );
buf U19800 ( n11454, n1021 );
not U19801 ( n1021, P2_IR_REG_31_ );
xor U19802 ( n8407, n10147, n10148 );
xor U19803 ( n10147, SI_20_, n10149 );
and U19804 ( n7277, n8405, n8406 );
nand U19805 ( n8405, P1_DATAO_REG_20_, n11328 );
nand U19806 ( n8406, n11269, n8407 );
nand U19807 ( n7900, n8527, n8528 );
nand U19808 ( n8527, P1_DATAO_REG_7_, n11328 );
nand U19809 ( n8528, n11268, n8529 );
nand U19810 ( n8157, P2_IR_REG_27_, n11457 );
nand U19811 ( n9845, n10443, n10444 );
nand U19812 ( n10444, P1_DATAO_REG_13_, n11264 );
nand U19813 ( n10443, P2_DATAO_REG_13_, n11325 );
nor U19814 ( n9823, n9845, SI_13_ );
nand U19815 ( n1935, n6544, n6545 );
nand U19816 ( n6544, P2_REG1_REG_24_, n6519 );
nand U19817 ( n6545, n11273, n6546 );
nand U19818 ( n1775, n6976, n6977 );
nand U19819 ( n6976, P2_REG0_REG_24_, n11355 );
nand U19820 ( n6977, n11270, n6546 );
nor U19821 ( n8077, P2_REG3_REG_3_, n11338 );
and U19822 ( n7227, n8398, n8399 );
nand U19823 ( n8398, P1_DATAO_REG_21_, n11328 );
nand U19824 ( n8399, n11269, n8400 );
nand U19825 ( n705, n2578, n2579 );
nand U19826 ( n2578, P1_REG1_REG_23_, n11426 );
nand U19827 ( n2579, n11279, n2580 );
nand U19828 ( n545, n3026, n3027 );
nand U19829 ( n3026, P1_REG0_REG_23_, n11422 );
nand U19830 ( n3027, n11276, n2580 );
nor U19831 ( n10753, n11307, n10977 );
xnor U19832 ( n8502, n10119, n10120 );
xnor U19833 ( n10120, SI_10_, n10121 );
nand U19834 ( n7745, n8500, n8501 );
nand U19835 ( n8500, P1_DATAO_REG_10_, n11328 );
nand U19836 ( n8501, n11269, n8502 );
nand U19837 ( n2505, n4160, n4161 );
nor U19838 ( n4160, n4194, n4195 );
nor U19839 ( n4161, n4162, n4163 );
and U19840 ( n4194, n11282, P2_REG3_REG_28_ );
nand U19841 ( n1925, n6550, n6551 );
nand U19842 ( n6550, P2_REG1_REG_22_, n11359 );
nand U19843 ( n6551, n11273, n6552 );
nand U19844 ( n1765, n7095, n7096 );
nand U19845 ( n7095, P2_REG0_REG_22_, n11355 );
nand U19846 ( n7096, n11270, n6552 );
nand U19847 ( n1805, n6652, n6653 );
nand U19848 ( n6652, P2_REG0_REG_30_, n6651 );
nand U19849 ( n6653, n11270, n6522 );
nand U19850 ( n1965, n6520, n6521 );
nand U19851 ( n6520, P2_REG1_REG_30_, n6519 );
nand U19852 ( n6521, n11273, n6522 );
nor U19853 ( n8171, n11348, n10994 );
nand U19854 ( n7651, n8482, n8483 );
nand U19855 ( n8482, P1_DATAO_REG_12_, n11326 );
nand U19856 ( n8483, n11269, n8484 );
nor U19857 ( n9994, SI_2_, n9995 );
xnor U19858 ( n9995, n9991, n9996 );
nand U19859 ( n8101, n8575, n8576 );
nand U19860 ( n8575, P1_DATAO_REG_2_, n11328 );
nand U19861 ( n8576, n11268, n8577 );
nand U19862 ( n2405, n4587, n4588 );
nor U19863 ( n4587, n4641, n4642 );
nor U19864 ( n4588, n4589, n4590 );
and U19865 ( n4641, n11283, P2_REG3_REG_26_ );
nor U19866 ( n8118, n11348, n10997 );
nand U19867 ( n9819, SI_13_, n9845 );
nor U19868 ( n8011, n11348, n10990 );
and U19869 ( n10762, n11313, P1_REG0_REG_1_ );
nor U19870 ( n8079, n11348, n10993 );
xnor U19871 ( n8536, n10063, n10064 );
xnor U19872 ( n10064, SI_6_, n10065 );
nand U19873 ( n7951, n8534, n8535 );
nand U19874 ( n8534, P1_DATAO_REG_6_, n11328 );
nand U19875 ( n8535, n11268, n8536 );
and U19876 ( n6180, n10145, n10146 );
nand U19877 ( n10145, P2_DATAO_REG_20_, n11267 );
nand U19878 ( n10146, n8407, n11328 );
nor U19879 ( n8045, n11348, n10999 );
and U19880 ( n10754, n11313, P1_REG0_REG_2_ );
xnor U19881 ( n8495, n9848, n10086 );
xnor U19882 ( n10086, SI_11_, n10087 );
nand U19883 ( n7707, n8493, n8494 );
nand U19884 ( n8493, P1_DATAO_REG_11_, n11326 );
nand U19885 ( n8494, n11333, n8495 );
nand U19886 ( n7849, n8517, n8518 );
nand U19887 ( n8517, P1_DATAO_REG_8_, n11328 );
nand U19888 ( n8518, n11268, n8519 );
nand U19889 ( n265, n3994, n3995 );
nand U19890 ( n3995, n3996, n3997 );
nand U19891 ( n3994, n3999, n11534 );
nor U19892 ( n3996, P1_IR_REG_30_, n3998 );
nand U19893 ( n1490, n8301, n8302 );
nand U19894 ( n8302, n8303, n8304 );
nand U19895 ( n8301, n6650, n11282 );
nor U19896 ( n8303, P2_IR_REG_30_, n8305 );
nand U19897 ( n710, n2575, n2576 );
nand U19898 ( n2575, P1_REG1_REG_24_, n2556 );
nand U19899 ( n2576, n11279, n2577 );
nand U19900 ( n550, n2963, n2964 );
nand U19901 ( n2963, P1_REG0_REG_24_, n2660 );
nand U19902 ( n2964, n11276, n2577 );
nand U19903 ( n695, n2584, n2585 );
nand U19904 ( n2584, P1_REG1_REG_21_, n11426 );
nand U19905 ( n2585, n11279, n2586 );
nand U19906 ( n700, n2581, n2582 );
nand U19907 ( n2581, P1_REG1_REG_22_, n11426 );
nand U19908 ( n2582, n11279, n2583 );
nand U19909 ( n540, n3075, n3076 );
nand U19910 ( n3075, P1_REG0_REG_22_, n11422 );
nand U19911 ( n3076, n11276, n2583 );
nand U19912 ( n535, n3134, n3135 );
nand U19913 ( n3134, P1_REG0_REG_21_, n11422 );
nand U19914 ( n3135, n11276, n2586 );
nand U19915 ( n1485, n8310, n8311 );
nand U19916 ( n8311, n11324, P2_IR_REG_30_ );
nor U19917 ( n8310, n8313, n8314 );
nor U19918 ( n8313, n8178, n11450 );
nand U19919 ( n2535, n4047, n4048 );
nor U19920 ( n4047, n4057, n4058 );
nor U19921 ( n4048, n4049, n4050 );
and U19922 ( n4057, n11283, P2_REG3_REG_27_ );
nor U19923 ( n7973, n11348, n11001 );
nand U19924 ( n260, n4000, n4001 );
nand U19925 ( n4001, n11408, P1_IR_REG_30_ );
nor U19926 ( n4000, n4003, n4004 );
nor U19927 ( n4004, n4005, n11490 );
nor U19928 ( n10744, P1_REG3_REG_3_, n11300 );
nor U19929 ( n9993, n9991, n9997 );
nand U19930 ( n9997, n776, SI_2_ );
not U19931 ( n776, n9996 );
xnor U19932 ( n8418, n9734, n9735 );
xnor U19933 ( n9735, SI_19_, n9736 );
nand U19934 ( n7324, n8416, n8417 );
nand U19935 ( n8416, P1_DATAO_REG_19_, n11326 );
nand U19936 ( n8417, n11269, n8418 );
xnor U19937 ( n8554, n10012, n10013 );
xnor U19938 ( n10013, SI_4_, n10014 );
nand U19939 ( n8032, n8552, n8553 );
nand U19940 ( n8552, P1_DATAO_REG_4_, n11328 );
nand U19941 ( n8553, n11268, n8554 );
nand U19942 ( n8127, n8585, n8586 );
nand U19943 ( n8585, P1_DATAO_REG_1_, n11328 );
nand U19944 ( n8586, n11268, n8587 );
nand U19945 ( n8587, n10505, n10506 );
nand U19946 ( n10505, SI_1_, n10508 );
nand U19947 ( n10506, n10507, n1178 );
nand U19948 ( n10508, n10425, n10427 );
nand U19949 ( n9817, n10449, n10450 );
nand U19950 ( n10450, P1_DATAO_REG_14_, n11330 );
nand U19951 ( n10449, P2_DATAO_REG_14_, n11325 );
and U19952 ( n10746, n11313, P1_REG0_REG_3_ );
nand U19953 ( n1920, n6553, n6554 );
nand U19954 ( n6553, P2_REG1_REG_21_, n11359 );
nand U19955 ( n6554, n11273, n6555 );
nand U19956 ( n1760, n7160, n7161 );
nand U19957 ( n7160, P2_REG0_REG_21_, n11355 );
nand U19958 ( n7161, n11270, n6555 );
nand U19959 ( n9048, n9987, n9988 );
nand U19960 ( n9987, P2_DATAO_REG_2_, n11330 );
nand U19961 ( n9988, n8577, n11327 );
nand U19962 ( n2460, n4373, n4374 );
nor U19963 ( n4373, n4388, n4389 );
nor U19964 ( n4374, n4375, n4376 );
and U19965 ( n4388, n11282, P2_REG3_REG_24_ );
nand U19966 ( n7582, n8458, n8459 );
nand U19967 ( n8458, P1_DATAO_REG_14_, n11326 );
nand U19968 ( n8459, n11269, n8460 );
xnor U19969 ( n8460, n9815, n9816 );
xnor U19970 ( n9816, SI_14_, n9817 );
nand U19971 ( n9815, n9818, n9819 );
nor U19972 ( n9818, n9820, n9821 );
xnor U19973 ( n8435, n9763, n9764 );
xnor U19974 ( n9764, SI_17_, n9765 );
nand U19975 ( n7445, n8433, n8434 );
nand U19976 ( n8433, P1_DATAO_REG_17_, n11326 );
nand U19977 ( n8434, n11269, n8435 );
nand U19978 ( n6307, n9732, n9733 );
nand U19979 ( n9732, P2_DATAO_REG_19_, n11267 );
nand U19980 ( n9733, n8418, n11328 );
nand U19981 ( n2480, n4291, n4292 );
nor U19982 ( n4291, n4306, n4307 );
nor U19983 ( n4292, n4293, n4294 );
and U19984 ( n4306, n11282, P2_REG3_REG_25_ );
xor U19985 ( n8593, SI_0_, n10513 );
nand U19986 ( n9955, n10607, n10608 );
nand U19987 ( n10607, P2_DATAO_REG_0_, n11266 );
nand U19988 ( n10608, n8593, n11325 );
xnor U19989 ( n8512, n9929, n9930 );
xnor U19990 ( n9930, SI_9_, n9931 );
nand U19991 ( n7792, n8510, n8511 );
nand U19992 ( n8510, P1_DATAO_REG_9_, n11328 );
nand U19993 ( n8511, n11269, n8512 );
xnor U19994 ( n8564, n10027, n10028 );
xnor U19995 ( n10028, SI_3_, n10029 );
nand U19996 ( n8064, n8562, n8563 );
nand U19997 ( n8562, P1_DATAO_REG_3_, n11328 );
nand U19998 ( n8563, n11269, n8564 );
nand U19999 ( n690, n2587, n2588 );
nand U20000 ( n2587, P1_REG1_REG_20_, n11426 );
nand U20001 ( n2588, n11279, n2589 );
nand U20002 ( n530, n3194, n3195 );
nand U20003 ( n3194, P1_REG0_REG_20_, n11422 );
nand U20004 ( n3195, n11276, n2589 );
xnor U20005 ( n10046, SI_5_, n10052 );
nand U20006 ( n7614, n8468, n8469 );
nand U20007 ( n8468, P1_DATAO_REG_13_, n11326 );
nand U20008 ( n8469, n11269, n8470 );
xnor U20009 ( n8470, n9843, n9844 );
xnor U20010 ( n9844, SI_13_, n9845 );
nand U20011 ( n9843, n9824, n9846 );
nand U20012 ( n9846, n9847, n9848 );
nand U20013 ( n1480, n8318, n8319 );
nand U20014 ( n8319, n11324, P2_IR_REG_29_ );
nor U20015 ( n8318, n8320, n8321 );
nor U20016 ( n8320, n11449, n8325 );
nand U20017 ( n255, n4011, n4012 );
nand U20018 ( n4012, n11408, P1_IR_REG_29_ );
nor U20019 ( n4011, n4013, n4014 );
nor U20020 ( n4013, n11488, n4016 );
nand U20021 ( n8156, n8591, n8592 );
nand U20022 ( n8591, P1_DATAO_REG_0_, n11328 );
nand U20023 ( n8592, n8593, n11267 );
nand U20024 ( n525, n3238, n3239 );
nand U20025 ( n3238, P1_REG0_REG_19_, n11422 );
nand U20026 ( n3239, n11277, n2592 );
nand U20027 ( n685, n2590, n2591 );
nand U20028 ( n2590, P1_REG1_REG_19_, n11426 );
nand U20029 ( n2591, n11280, n2592 );
nand U20030 ( n9797, n10386, n10387 );
nand U20031 ( n10387, P1_DATAO_REG_15_, n11330 );
nand U20032 ( n10386, P2_DATAO_REG_15_, n11326 );
xor U20033 ( n8425, n9776, n9777 );
xor U20034 ( n9776, SI_18_, n9778 );
nand U20035 ( n7388, n8423, n8424 );
nand U20036 ( n8423, P1_DATAO_REG_18_, n11326 );
nand U20037 ( n8424, n11269, n8425 );
xnor U20038 ( n8453, n9795, n9796 );
xnor U20039 ( n9796, SI_15_, n9797 );
nand U20040 ( n7535, n8451, n8452 );
nand U20041 ( n8451, P1_DATAO_REG_15_, n11326 );
nand U20042 ( n8452, n11269, n8453 );
xor U20043 ( n8442, n10134, n10135 );
xor U20044 ( n10134, SI_16_, n10136 );
nand U20045 ( n7496, n8440, n8441 );
nand U20046 ( n8440, P1_DATAO_REG_16_, n11326 );
nand U20047 ( n8441, n11269, n8442 );
not U20048 ( n1177, SI_7_ );
nand U20049 ( n9978, n10503, n10504 );
nand U20050 ( n10503, P2_DATAO_REG_1_, n11330 );
nand U20051 ( n10504, n8587, n11325 );
nand U20052 ( n8883, n10025, n10026 );
nand U20053 ( n10025, P2_DATAO_REG_3_, n11266 );
nand U20054 ( n10026, n8564, n11327 );
nand U20055 ( n7797, n10097, n10098 );
nand U20056 ( n10097, P2_DATAO_REG_12_, n11265 );
nand U20057 ( n10098, n8484, n11327 );
nor U20058 ( n7921, n11348, n11006 );
nand U20059 ( n1915, n6556, n6557 );
nand U20060 ( n6556, P2_REG1_REG_20_, n11359 );
nand U20061 ( n6557, n11273, n6558 );
nand U20062 ( n1755, n7228, n7229 );
nand U20063 ( n7228, P2_REG0_REG_20_, n11355 );
nand U20064 ( n7229, n11270, n6558 );
nand U20065 ( n9387, n10829, n10830 );
nand U20066 ( n10829, P1_IR_REG_22_, n11487 );
or U20067 ( n10830, n5573, n11484 );
nand U20068 ( n5573, n10831, n10832 );
nand U20069 ( n10831, P1_IR_REG_22_, n10833 );
or U20070 ( n10833, n354, P1_IR_REG_21_ );
nand U20071 ( n7330, n9841, n9842 );
nand U20072 ( n9841, P2_DATAO_REG_13_, n11267 );
nand U20073 ( n9842, n8470, n11327 );
nand U20074 ( n1910, n6559, n6560 );
nand U20075 ( n6559, P2_REG1_REG_19_, n11359 );
nand U20076 ( n6560, n11274, n6561 );
nand U20077 ( n1750, n7278, n7279 );
nand U20078 ( n7278, P2_REG0_REG_19_, n11355 );
nand U20079 ( n7279, n11271, n6561 );
nand U20080 ( n6435, n9774, n9775 );
nand U20081 ( n9774, P2_DATAO_REG_18_, n11267 );
nand U20082 ( n9775, n8425, n11328 );
nand U20083 ( n2525, n4085, n4086 );
nor U20084 ( n4085, n4097, n4098 );
nor U20085 ( n4086, n4087, n4088 );
and U20086 ( n4097, n11282, P2_REG3_REG_23_ );
nand U20087 ( n1475, n8326, n8327 );
nand U20088 ( n8327, n11324, P2_IR_REG_28_ );
nor U20089 ( n8326, n8328, n8329 );
nor U20090 ( n8328, n11449, n8333 );
nand U20091 ( n250, n4218, n4219 );
nand U20092 ( n4219, n11408, P1_IR_REG_28_ );
nor U20093 ( n4218, n4220, n4221 );
nor U20094 ( n4221, n4222, n11490 );
nand U20095 ( n8258, n10117, n10118 );
nand U20096 ( n10117, P2_DATAO_REG_10_, n11267 );
nand U20097 ( n10118, n8502, n11326 );
nand U20098 ( n6572, n10132, n10133 );
nand U20099 ( n10132, P2_DATAO_REG_16_, n11267 );
nand U20100 ( n10133, n8442, n11327 );
nand U20101 ( n680, n2593, n2594 );
nand U20102 ( n2593, P1_REG1_REG_18_, n11426 );
nand U20103 ( n2594, n11280, n2595 );
nand U20104 ( n520, n3283, n3284 );
nand U20105 ( n3283, P1_REG0_REG_18_, n11422 );
nand U20106 ( n3284, n11277, n2595 );
nand U20107 ( n10136, n10381, n10382 );
nand U20108 ( n10382, P1_DATAO_REG_16_, n11265 );
nand U20109 ( n10381, P2_DATAO_REG_16_, n11326 );
nand U20110 ( n8383, n9890, n9891 );
nand U20111 ( n9890, P2_DATAO_REG_7_, n11268 );
nand U20112 ( n9891, n8529, n11327 );
and U20113 ( n10738, n11313, P1_REG0_REG_4_ );
nand U20114 ( n2490, n4244, n4245 );
nor U20115 ( n4244, n4263, n4264 );
nor U20116 ( n4245, n4246, n4247 );
and U20117 ( n4263, n11282, P2_REG3_REG_21_ );
nand U20118 ( n8668, n10010, n10011 );
nand U20119 ( n10010, P2_DATAO_REG_4_, n11266 );
nand U20120 ( n10011, n8554, n11327 );
nand U20121 ( n6611, n9793, n9794 );
nand U20122 ( n9793, P2_DATAO_REG_15_, n11268 );
nand U20123 ( n9794, n8453, n11328 );
nand U20124 ( n8274, n9905, n9906 );
nand U20125 ( n9905, P2_DATAO_REG_8_, n11268 );
nand U20126 ( n9906, n8519, n11327 );
nand U20127 ( n6537, n9761, n9762 );
nand U20128 ( n9761, P2_DATAO_REG_17_, n11267 );
nand U20129 ( n9762, n8435, n11328 );
nand U20130 ( n8252, n10084, n10085 );
nand U20131 ( n10084, P2_DATAO_REG_11_, n11266 );
nand U20132 ( n10085, n8495, n11327 );
nand U20133 ( n1905, n6562, n6563 );
nand U20134 ( n6562, P2_REG1_REG_18_, n11359 );
nand U20135 ( n6563, n11274, n6564 );
nand U20136 ( n1745, n7331, n7332 );
nand U20137 ( n7331, P2_REG0_REG_18_, n11355 );
nand U20138 ( n7332, n11271, n6564 );
nand U20139 ( n2430, n4497, n4498 );
nor U20140 ( n4497, n4508, n4509 );
nor U20141 ( n4498, n4499, n4500 );
and U20142 ( n4508, n11282, P2_REG3_REG_22_ );
nand U20143 ( n8570, n10042, n10043 );
nand U20144 ( n10042, P2_DATAO_REG_5_, n11266 );
nand U20145 ( n10043, n8547, n11327 );
nor U20146 ( n7868, n11348, n11021 );
nor U20147 ( n7763, n11348, n11019 );
nor U20148 ( n7820, n11348, n11022 );
and U20149 ( n10730, n11313, P1_REG0_REG_5_ );
nand U20150 ( n675, n2596, n2597 );
nand U20151 ( n2596, P1_REG1_REG_17_, n11426 );
nand U20152 ( n2597, n11280, n2598 );
nand U20153 ( n515, n3340, n3341 );
nand U20154 ( n3340, P1_REG0_REG_17_, n11422 );
nand U20155 ( n3341, n11277, n2598 );
nand U20156 ( n8475, n10061, n10062 );
nand U20157 ( n10061, P2_DATAO_REG_6_, n11266 );
nand U20158 ( n10062, n8536, n11327 );
and U20159 ( n10722, n11312, P1_REG0_REG_6_ );
nand U20160 ( n8266, n9927, n9928 );
nand U20161 ( n9927, P2_DATAO_REG_9_, n11268 );
nand U20162 ( n9928, n8512, n11327 );
nand U20163 ( n670, n2599, n2600 );
nand U20164 ( n2599, P1_REG1_REG_16_, n11426 );
nand U20165 ( n2600, n11280, n2601 );
nand U20166 ( n510, n3390, n3391 );
nand U20167 ( n3390, P1_REG0_REG_16_, n11422 );
nand U20168 ( n3391, n11277, n2601 );
nand U20169 ( n1470, n8336, n8337 );
nand U20170 ( n8337, n11324, P2_IR_REG_27_ );
nor U20171 ( n8336, n8338, n8339 );
nor U20172 ( n8338, n8159, n11450 );
nand U20173 ( n9765, n10376, n10377 );
nand U20174 ( n10377, P1_DATAO_REG_17_, n11265 );
nand U20175 ( n10376, P2_DATAO_REG_17_, n11326 );
nand U20176 ( n2440, n4447, n4448 );
nor U20177 ( n4447, n4463, n4464 );
nor U20178 ( n4448, n4449, n4450 );
and U20179 ( n4463, n11282, P2_REG3_REG_20_ );
nand U20180 ( n1900, n6565, n6566 );
nand U20181 ( n6565, P2_REG1_REG_17_, n11359 );
nand U20182 ( n6566, n11274, n6567 );
nand U20183 ( n1740, n7389, n7390 );
nand U20184 ( n7389, P2_REG0_REG_17_, n11355 );
nand U20185 ( n7390, n11271, n6567 );
nand U20186 ( n6733, n9813, n9814 );
nand U20187 ( n9813, P2_DATAO_REG_14_, n11268 );
nand U20188 ( n9814, n8460, n11327 );
and U20189 ( n10713, n11312, P1_REG0_REG_7_ );
nand U20190 ( n1465, n8343, n8344 );
nand U20191 ( n8344, n11324, P2_IR_REG_26_ );
nor U20192 ( n8343, n8345, n8346 );
nor U20193 ( n8345, n11449, n8350 );
nand U20194 ( n240, n4750, n4751 );
nand U20195 ( n4751, n11408, P1_IR_REG_26_ );
nor U20196 ( n4750, n4752, n4753 );
nor U20197 ( n4753, n4754, n11490 );
nand U20198 ( n505, n3448, n3449 );
nand U20199 ( n3448, P1_REG0_REG_15_, n11422 );
nand U20200 ( n3449, n11277, n2604 );
nand U20201 ( n665, n2602, n2603 );
nand U20202 ( n2602, P1_REG1_REG_15_, n11426 );
nand U20203 ( n2603, n11280, n2604 );
nor U20204 ( n7724, n11348, n11029 );
xnor U20205 ( n9909, SI_8_, n9916 );
nand U20206 ( n9778, n10371, n10372 );
nand U20207 ( n10372, P1_DATAO_REG_18_, n11265 );
nand U20208 ( n10371, P2_DATAO_REG_18_, n11326 );
nor U20209 ( n10703, n11307, n11034 );
nand U20210 ( n1895, n6576, n6577 );
nand U20211 ( n6576, P2_REG1_REG_16_, n11359 );
nand U20212 ( n6577, n11274, n6578 );
nand U20213 ( n1735, n7446, n7447 );
nand U20214 ( n7446, P2_REG0_REG_16_, n11355 );
nand U20215 ( n7447, n11271, n6578 );
and U20216 ( n10686, n11312, P1_REG0_REG_10_ );
and U20217 ( n10704, n11312, P1_REG0_REG_8_ );
nand U20218 ( n1890, n6579, n6580 );
nand U20219 ( n6579, P2_REG1_REG_15_, n11359 );
nand U20220 ( n6580, n11274, n6581 );
nand U20221 ( n1730, n7497, n7498 );
nand U20222 ( n7497, P2_REG0_REG_15_, n11355 );
nand U20223 ( n7498, n11271, n6581 );
nor U20224 ( n7676, n11349, n11035 );
nand U20225 ( n500, n3488, n3489 );
nand U20226 ( n3488, P1_REG0_REG_14_, n11422 );
nand U20227 ( n3489, n11277, n2607 );
nand U20228 ( n660, n2605, n2606 );
nand U20229 ( n2605, P1_REG1_REG_14_, n11426 );
nand U20230 ( n2606, n11280, n2607 );
nand U20231 ( n495, n3540, n3541 );
nand U20232 ( n3540, P1_REG0_REG_13_, n11422 );
nand U20233 ( n3541, n11277, n2610 );
nand U20234 ( n655, n2608, n2609 );
nand U20235 ( n2608, P1_REG1_REG_13_, n11426 );
nand U20236 ( n2609, n11280, n2610 );
nand U20237 ( n1460, n8354, n8355 );
nand U20238 ( n8355, n11324, P2_IR_REG_25_ );
nor U20239 ( n8354, n8356, n8357 );
nor U20240 ( n8356, n8296, n11450 );
nor U20241 ( n7631, n11349, n11040 );
and U20242 ( n10695, n11312, P1_REG0_REG_9_ );
nand U20243 ( n235, n5335, n5336 );
nand U20244 ( n5336, n11408, P1_IR_REG_25_ );
nor U20245 ( n5335, n5337, n5338 );
nor U20246 ( n5338, n5339, n11489 );
nand U20247 ( n9736, n10366, n10367 );
nand U20248 ( n10367, P1_DATAO_REG_19_, n11265 );
nand U20249 ( n10366, P2_DATAO_REG_19_, n11326 );
nand U20250 ( n1885, n6582, n6583 );
nand U20251 ( n6582, P2_REG1_REG_14_, n11359 );
nand U20252 ( n6583, n11274, n6584 );
nand U20253 ( n1725, n7536, n7537 );
nand U20254 ( n7536, P2_REG0_REG_14_, n11355 );
nand U20255 ( n7537, n11271, n6584 );
nor U20256 ( n10676, n11307, n11053 );
not U20257 ( n1178, SI_1_ );
nand U20258 ( n8243, n8281, n8282 );
nand U20259 ( n8282, n8283, n8269 );
xnor U20260 ( n8283, n8280, P2_B_REG );
nand U20261 ( n8281, n8289, n8290 );
nand U20262 ( n8289, P2_IR_REG_26_, n11458 );
nand U20263 ( n8290, n8291, P2_IR_REG_31_ );
and U20264 ( n8291, n8292, n8293 );
nand U20265 ( n8293, P2_IR_REG_26_, n8353 );
or U20266 ( n8353, n957, P2_IR_REG_25_ );
nand U20267 ( n6645, n8244, n8245 );
nand U20268 ( n8245, n8246, n8243 );
nand U20269 ( n8244, P2_D_REG_0_, n954 );
and U20270 ( n8280, n8297, n8298 );
nand U20271 ( n8297, P2_IR_REG_24_, n11456 );
nand U20272 ( n8298, n8299, P2_IR_REG_31_ );
and U20273 ( n8299, n957, n8300 );
xnor U20274 ( n8296, P2_IR_REG_25_, n957 );
nor U20275 ( n8269, n11255, n11256 );
and U20276 ( n11255, P2_IR_REG_25_, n11458 );
nor U20277 ( n11256, n8296, n11455 );
and U20278 ( n10668, n11312, P1_REG0_REG_12_ );
and U20279 ( n10659, n11312, P1_REG0_REG_13_ );
nand U20280 ( n8300, P2_IR_REG_24_, n8370 );
or U20281 ( n8370, n8201, P2_IR_REG_23_ );
nand U20282 ( n650, n2611, n2612 );
nand U20283 ( n2611, P1_REG1_REG_12_, n11426 );
nand U20284 ( n2612, n11280, n2613 );
nand U20285 ( n490, n3575, n3576 );
nand U20286 ( n3575, P1_REG0_REG_12_, n11422 );
nand U20287 ( n3576, n11277, n2613 );
nand U20288 ( n1455, n8361, n8362 );
nand U20289 ( n8362, n11324, P2_IR_REG_24_ );
nor U20290 ( n8361, n8363, n8364 );
nor U20291 ( n8363, n11449, n8368 );
nand U20292 ( n230, n5361, n5362 );
nand U20293 ( n5362, n11408, P1_IR_REG_24_ );
nor U20294 ( n5361, n5363, n5364 );
nor U20295 ( n5363, n11488, n5366 );
and U20296 ( n10677, n11312, P1_REG0_REG_11_ );
xnor U20297 ( n10101, SI_12_, n10108 );
nand U20298 ( n10149, n10361, n10362 );
nand U20299 ( n10362, P1_DATAO_REG_20_, n11265 );
nand U20300 ( n10361, P2_DATAO_REG_20_, n11326 );
nand U20301 ( n2513, P1_REG3_REG_1_, n11434 );
nand U20302 ( n2487, n2488, n2489 );
nand U20303 ( n2488, n20, n11442 );
nand U20304 ( n2489, n11434, P1_REG3_REG_2_ );
nor U20305 ( n7596, n11349, n11054 );
nand U20306 ( n480, n3651, n3652 );
nand U20307 ( n3651, P1_REG0_REG_10_, n2660 );
nand U20308 ( n3652, n11277, n2619 );
nand U20309 ( n640, n2617, n2618 );
nand U20310 ( n2617, P1_REG1_REG_10_, n2556 );
nand U20311 ( n2618, n11280, n2619 );
nand U20312 ( n1720, n7583, n7584 );
nand U20313 ( n7583, P2_REG0_REG_13_, n11355 );
nand U20314 ( n7584, n11271, n6587 );
nand U20315 ( n1880, n6585, n6586 );
nand U20316 ( n6585, P2_REG1_REG_13_, n11359 );
nand U20317 ( n6586, n11274, n6587 );
nand U20318 ( n5437, n8128, n8129 );
nand U20319 ( n8129, P2_IR_REG_31_, n8130 );
nand U20320 ( n8128, P2_IR_REG_1_, n11457 );
nand U20321 ( n1875, n6588, n6589 );
nand U20322 ( n6588, P2_REG1_REG_12_, n11359 );
nand U20323 ( n6589, n11274, n6590 );
nand U20324 ( n1715, n7618, n7619 );
nand U20325 ( n7618, P2_REG0_REG_12_, n11355 );
nand U20326 ( n7619, n11271, n6590 );
nand U20327 ( n1450, n8371, n8372 );
nand U20328 ( n8372, n11324, P2_IR_REG_23_ );
nor U20329 ( n8371, n8373, n8374 );
nor U20330 ( n8373, n8287, n11450 );
nand U20331 ( n225, n5388, n5389 );
nand U20332 ( n5389, n11408, P1_IR_REG_23_ );
nor U20333 ( n5388, n5390, n5391 );
nor U20334 ( n5390, n11488, n5393 );
nor U20335 ( n7553, n11349, n11058 );
nand U20336 ( n645, n2614, n2615 );
nand U20337 ( n2614, P1_REG1_REG_11_, n2556 );
nand U20338 ( n2615, n11280, n2616 );
nand U20339 ( n485, n3609, n3610 );
nand U20340 ( n3609, P1_REG0_REG_11_, n2660 );
nand U20341 ( n3610, n11277, n2616 );
nand U20342 ( n635, n2620, n2621 );
nand U20343 ( n2620, P1_REG1_REG_9_, n2556 );
nand U20344 ( n2621, n11280, n2622 );
nor U20345 ( n10640, n11308, n11068 );
nand U20346 ( n475, n3685, n3686 );
nand U20347 ( n3685, P1_REG0_REG_9_, n2660 );
nand U20348 ( n3686, n11277, n2622 );
nand U20349 ( n5533, n7995, n7996 );
nand U20350 ( n7995, P2_IR_REG_5_, n11457 );
or U20351 ( n7996, n7997, n11455 );
nand U20352 ( n10158, n10356, n10357 );
nand U20353 ( n10357, P1_DATAO_REG_21_, n11265 );
nand U20354 ( n10356, P2_DATAO_REG_21_, n11326 );
nand U20355 ( n5459, n8102, n8103 );
nand U20356 ( n8103, n8104, P2_IR_REG_31_ );
nand U20357 ( n8102, P2_IR_REG_2_, n11457 );
and U20358 ( n8104, n8105, n8106 );
nand U20359 ( n1870, n6591, n6592 );
nand U20360 ( n6591, P2_REG1_REG_11_, n6519 );
nand U20361 ( n6592, n11274, n6593 );
nand U20362 ( n1710, n7657, n7658 );
nand U20363 ( n7657, P2_REG0_REG_11_, n6651 );
nand U20364 ( n7658, n11271, n6593 );
and U20365 ( n10641, n11312, P1_REG0_REG_15_ );
nor U20366 ( n10649, n11308, n11074 );
nand U20367 ( n1445, n8384, n8385 );
nand U20368 ( n8385, n11324, P2_IR_REG_22_ );
nor U20369 ( n8384, n8386, n8387 );
nor U20370 ( n8386, n11450, n8391 );
nor U20371 ( n7513, n11349, n11062 );
nand U20372 ( n220, n5569, n5570 );
nand U20373 ( n5570, n11408, P1_IR_REG_22_ );
nor U20374 ( n5569, n5571, n5572 );
nor U20375 ( n5572, n5573, n11489 );
and U20376 ( n10650, n11312, P1_REG0_REG_14_ );
nand U20377 ( n5488, n8065, n8066 );
nand U20378 ( n8065, P2_IR_REG_3_, n11457 );
or U20379 ( n8066, n8067, n11455 );
nand U20380 ( n1192, n9998, n9999 );
nand U20381 ( n9999, n10000, P1_IR_REG_31_ );
nand U20382 ( n9998, P1_IR_REG_2_, n11485 );
and U20383 ( n10000, n9051, n9050 );
xnor U20384 ( n8192, P2_IR_REG_21_, n8196 );
nand U20385 ( n4738, n8190, n8191 );
nand U20386 ( n8190, P2_IR_REG_21_, n11458 );
or U20387 ( n8191, n8192, n11455 );
nand U20388 ( n470, n3712, n3713 );
nand U20389 ( n3712, P1_REG0_REG_8_, n2660 );
nand U20390 ( n3713, n11277, n2625 );
nand U20391 ( n630, n2623, n2624 );
nand U20392 ( n2623, P1_REG1_REG_8_, n2556 );
nand U20393 ( n2624, n11280, n2625 );
nor U20394 ( n7464, n11349, n11065 );
nand U20395 ( n5508, n8028, n8029 );
nand U20396 ( n8029, n8030, P2_IR_REG_31_ );
nand U20397 ( n8028, P2_IR_REG_4_, n11457 );
and U20398 ( n8030, n873, n8031 );
nand U20399 ( n1853, n10811, n10812 );
nand U20400 ( n10812, P1_IR_REG_31_, n10502 );
nand U20401 ( n10811, P1_IR_REG_1_, n11487 );
nand U20402 ( n5445, n5956, P2_IR_REG_0_ );
nor U20403 ( n5956, n5957, n5958 );
nor U20404 ( n5957, n11287, n10967 );
nor U20405 ( n5958, n11459, n10966 );
nand U20406 ( n4743, n8193, n8194 );
nand U20407 ( n8193, P2_IR_REG_20_, n11458 );
nand U20408 ( n8194, n8195, P2_IR_REG_31_ );
and U20409 ( n8195, n8196, n8197 );
nand U20410 ( n8197, P2_IR_REG_20_, n8411 );
nand U20411 ( n8411, n8410, n10996 );
nand U20412 ( n465, n3750, n3751 );
nand U20413 ( n3750, P1_REG0_REG_7_, n2660 );
nand U20414 ( n3751, n11278, n2628 );
nand U20415 ( n625, n2626, n2627 );
nand U20416 ( n2626, P1_REG1_REG_7_, n2556 );
nand U20417 ( n2627, n11281, n2628 );
nand U20418 ( n5559, n7952, n7953 );
nand U20419 ( n7953, n7954, P2_IR_REG_31_ );
nand U20420 ( n7952, P2_IR_REG_6_, n11457 );
and U20421 ( n7954, n7955, n7956 );
and U20422 ( n10632, n11312, P1_REG0_REG_16_ );
nand U20423 ( n1865, n6594, n6595 );
nand U20424 ( n6594, P2_REG1_REG_10_, n6519 );
nand U20425 ( n6595, n11274, n6596 );
nand U20426 ( n1705, n7708, n7709 );
nand U20427 ( n7708, P2_REG0_REG_10_, n6651 );
nand U20428 ( n7709, n11271, n6596 );
nand U20429 ( n5844, n5845, n5846 );
nand U20430 ( n5845, P2_ADDR_REG_18_, n933 );
nand U20431 ( n5846, n5408, n5847 );
xor U20432 ( n5847, n5848, n5849 );
nand U20433 ( n5586, n7897, n7898 );
nand U20434 ( n7897, P2_IR_REG_7_, n11456 );
or U20435 ( n7898, n7899, n11456 );
nand U20436 ( n1854, n10030, n10031 );
nand U20437 ( n10030, P1_IR_REG_3_, n11485 );
or U20438 ( n10031, n8882, n11485 );
nand U20439 ( n5009, n8198, n8199 );
nand U20440 ( n8198, P2_IR_REG_22_, n11458 );
nand U20441 ( n8199, n8200, P2_IR_REG_31_ );
and U20442 ( n8200, n8201, n8202 );
nand U20443 ( n8202, P2_IR_REG_22_, n8393 );
or U20444 ( n8393, n8196, P2_IR_REG_21_ );
nor U20445 ( n10575, n11308, n11089 );
nand U20446 ( n1440, n8394, n8395 );
nand U20447 ( n8395, n11324, P2_IR_REG_21_ );
nor U20448 ( n8394, n8396, n8397 );
nor U20449 ( n8396, n8192, n11450 );
nand U20450 ( n1860, n6597, n6598 );
nand U20451 ( n6597, P2_REG1_REG_9_, n6519 );
nand U20452 ( n6598, n11274, n6599 );
nand U20453 ( n1700, n7750, n7751 );
nand U20454 ( n7750, P2_REG0_REG_9_, n6651 );
nand U20455 ( n7751, n11271, n6599 );
nand U20456 ( n215, n5805, n5806 );
nand U20457 ( n5806, n11408, P1_IR_REG_21_ );
nor U20458 ( n5805, n5807, n5808 );
nor U20459 ( n5808, n5809, n11489 );
nor U20460 ( n10584, n11308, n11091 );
nand U20461 ( n10188, n10351, n10352 );
nand U20462 ( n10352, P1_DATAO_REG_22_, n11264 );
nand U20463 ( n10351, P2_DATAO_REG_22_, n11326 );
nor U20464 ( n7402, n11349, n11073 );
and U20465 ( n10576, n11311, P1_REG0_REG_21_ );
nand U20466 ( n5444, n5959, n5960 );
nand U20467 ( n5959, P2_REG2_REG_1_, n11287 );
nand U20468 ( n5960, P2_REG1_REG_1_, n11459 );
and U20469 ( n10623, n11312, P1_REG0_REG_17_ );
nand U20470 ( n8187, P2_IR_REG_19_, n11458 );
or U20471 ( n8188, n8189, n11455 );
nand U20472 ( n460, n3787, n3788 );
nand U20473 ( n3787, P1_REG0_REG_6_, n2660 );
nand U20474 ( n3788, n11278, n2631 );
nand U20475 ( n620, n2629, n2630 );
nand U20476 ( n2629, P1_REG1_REG_6_, n2556 );
nand U20477 ( n2630, n11281, n2631 );
nor U20478 ( n7291, n11349, n11081 );
and U20479 ( n10585, n11311, P1_REG0_REG_20_ );
nor U20480 ( n7344, n11349, n11083 );
xnor U20481 ( n7997, P2_IR_REG_5_, n873 );
and U20482 ( n10594, n11311, P1_REG0_REG_19_ );
nand U20483 ( n1855, n6600, n6601 );
nand U20484 ( n6600, P2_REG1_REG_8_, n6519 );
nand U20485 ( n6601, n11274, n6602 );
nand U20486 ( n1695, n7801, n7802 );
nand U20487 ( n7801, P2_REG0_REG_8_, n6651 );
nand U20488 ( n7802, n11271, n6602 );
nand U20489 ( n1845, n6612, n6613 );
nand U20490 ( n6612, P2_REG1_REG_6_, n6519 );
nand U20491 ( n6613, n11275, n6614 );
nand U20492 ( n1685, n7901, n7902 );
nand U20493 ( n7901, P2_REG0_REG_6_, n6651 );
nand U20494 ( n7902, n11272, n6614 );
nor U20495 ( n10566, n11308, n11105 );
nand U20496 ( n1435, n8401, n8402 );
nand U20497 ( n8402, n11323, P2_IR_REG_20_ );
nor U20498 ( n8401, n8403, n8404 );
nor U20499 ( n8403, n11450, n8408 );
nand U20500 ( n210, n6176, n6177 );
nand U20501 ( n6177, n11408, P1_IR_REG_20_ );
nor U20502 ( n6176, n6178, n6179 );
nor U20503 ( n6178, n11488, n6181 );
nand U20504 ( n5824, n5825, n5826 );
nand U20505 ( n5825, P2_ADDR_REG_17_, n933 );
nand U20506 ( n5826, n5408, n5827 );
xnor U20507 ( n5827, n5828, n5829 );
and U20508 ( n10603, n11312, P1_REG0_REG_18_ );
nand U20509 ( n5458, n5951, n5952 );
nand U20510 ( n5951, P2_REG2_REG_2_, n5869 );
nand U20511 ( n5952, P2_REG1_REG_2_, n11459 );
and U20512 ( n10567, n11311, P1_REG0_REG_22_ );
nand U20513 ( n455, n3834, n3835 );
nand U20514 ( n3834, P1_REG0_REG_5_, n2660 );
nand U20515 ( n3835, n11278, n2634 );
nand U20516 ( n615, n2632, n2633 );
nand U20517 ( n2632, P1_REG1_REG_5_, n2556 );
nand U20518 ( n2633, n11281, n2634 );
nand U20519 ( n10179, n10346, n10347 );
nand U20520 ( n10347, P1_DATAO_REG_23_, n11264 );
nand U20521 ( n10346, P2_DATAO_REG_23_, n11327 );
nand U20522 ( n5660, n7746, n7747 );
nand U20523 ( n7747, n7748, P2_IR_REG_31_ );
nand U20524 ( n7746, P2_IR_REG_10_, n11456 );
and U20525 ( n7748, n883, n7749 );
nand U20526 ( n5614, n7850, n7851 );
nand U20527 ( n7851, n7852, P2_IR_REG_31_ );
nand U20528 ( n7850, P2_IR_REG_8_, n11456 );
and U20529 ( n7852, n7853, n7854 );
nand U20530 ( n1850, n6603, n6604 );
nand U20531 ( n6603, P2_REG1_REG_7_, n6519 );
nand U20532 ( n6604, n11275, n6605 );
nand U20533 ( n1690, n7855, n7856 );
nand U20534 ( n7855, P2_REG0_REG_7_, n6651 );
nand U20535 ( n7856, n11272, n6605 );
nand U20536 ( n5487, n5961, n5962 );
nand U20537 ( n5961, P2_REG2_REG_3_, n5869 );
nand U20538 ( n5962, P2_REG1_REG_3_, n11459 );
xnor U20539 ( n8130, P2_IR_REG_1_, n10960 );
nor U20540 ( n7241, n11349, n11095 );
nand U20541 ( n7956, P2_IR_REG_6_, n8540 );
or U20542 ( n8540, n873, P2_IR_REG_5_ );
nor U20543 ( n10557, n11308, n11109 );
nor U20544 ( n7176, n11349, n11098 );
nand U20545 ( n450, n3862, n3863 );
nand U20546 ( n3862, P1_REG0_REG_4_, n2660 );
nand U20547 ( n3863, n11278, n2637 );
nand U20548 ( n610, n2635, n2636 );
nand U20549 ( n2635, P1_REG1_REG_4_, n2556 );
nand U20550 ( n2636, n11281, n2637 );
nand U20551 ( n5932, n5939, n5940 );
nand U20552 ( n5939, P2_REG2_REG_6_, n5869 );
nand U20553 ( n5940, P2_REG1_REG_6_, n11459 );
nand U20554 ( n1304, n10053, n10054 );
nand U20555 ( n10053, P1_IR_REG_5_, n11486 );
or U20556 ( n10054, n8569, n11484 );
and U20557 ( n5532, n5937, n5938 );
nand U20558 ( n5937, P2_REG2_REG_5_, n11287 );
nand U20559 ( n5938, P2_REG1_REG_5_, n11459 );
nand U20560 ( n8106, P2_IR_REG_2_, n8580 );
or U20561 ( n8580, P2_IR_REG_0_, P2_IR_REG_1_ );
nand U20562 ( n1840, n6615, n6616 );
nand U20563 ( n6615, P2_REG1_REG_5_, n6519 );
nand U20564 ( n6616, n11275, n6617 );
nand U20565 ( n1680, n7957, n7958 );
nand U20566 ( n7957, P2_REG0_REG_5_, n6651 );
nand U20567 ( n7958, n11272, n6617 );
nand U20568 ( n1273, n10015, n10016 );
nand U20569 ( n10016, n10017, P1_IR_REG_31_ );
nand U20570 ( n10015, P1_IR_REG_4_, n11486 );
and U20571 ( n10017, n8671, n8670 );
nand U20572 ( n5635, n7789, n7790 );
nand U20573 ( n7789, P2_IR_REG_9_, n11456 );
or U20574 ( n7790, n7791, n11455 );
nand U20575 ( n1430, n8412, n8413 );
nand U20576 ( n8413, n11323, P2_IR_REG_19_ );
nor U20577 ( n8412, n8414, n8415 );
nor U20578 ( n8414, n8189, n11450 );
nand U20579 ( n5507, n5942, n5943 );
nand U20580 ( n5942, P2_REG2_REG_4_, n11287 );
nand U20581 ( n5943, P2_REG1_REG_4_, n11459 );
nand U20582 ( n205, n6303, n6304 );
nand U20583 ( n6304, n11408, P1_IR_REG_19_ );
nor U20584 ( n6303, n6305, n6306 );
nor U20585 ( n6305, n11488, n6308 );
nand U20586 ( n605, n2638, n2639 );
nand U20587 ( n2638, P1_REG1_REG_3_, n2556 );
nand U20588 ( n2639, n11281, n2640 );
nand U20589 ( n445, n3887, n3888 );
nand U20590 ( n3887, P1_REG0_REG_3_, n2660 );
nand U20591 ( n3888, n11278, n2640 );
and U20592 ( n10558, n11311, P1_REG0_REG_23_ );
nand U20593 ( n9055, n9056, n9057 );
nand U20594 ( n9056, P1_REG3_REG_2_, n8794 );
nand U20595 ( n9057, n11507, n9058 );
nand U20596 ( n9058, n9059, n9060 );
nand U20597 ( n10201, n10341, n10342 );
nand U20598 ( n10342, P1_DATAO_REG_24_, n11264 );
nand U20599 ( n10341, P2_DATAO_REG_24_, n11327 );
nand U20600 ( n8031, P2_IR_REG_4_, n8557 );
or U20601 ( n8557, n8105, P2_IR_REG_3_ );
nand U20602 ( n10879, n10949, n10950 );
nand U20603 ( n10949, P1_ADDR_REG_2_, n10876 );
nand U20604 ( n10950, P2_ADDR_REG_2_, n10951 );
or U20605 ( n10951, n10876, P1_ADDR_REG_2_ );
nand U20606 ( n10883, n10943, n10944 );
nand U20607 ( n10943, P1_ADDR_REG_4_, n10880 );
nand U20608 ( n10944, P2_ADDR_REG_4_, n10945 );
or U20609 ( n10945, n10880, P1_ADDR_REG_4_ );
nand U20610 ( n10889, n10937, n10938 );
nand U20611 ( n10937, P1_ADDR_REG_6_, n10884 );
nand U20612 ( n10938, P2_ADDR_REG_6_, n10939 );
or U20613 ( n10939, n10884, P1_ADDR_REG_6_ );
nand U20614 ( n10893, n10931, n10932 );
nand U20615 ( n10931, P1_ADDR_REG_8_, n10890 );
nand U20616 ( n10932, P2_ADDR_REG_8_, n10933 );
or U20617 ( n10933, n10890, P1_ADDR_REG_8_ );
nand U20618 ( n10862, n10925, n10926 );
nand U20619 ( n10925, P1_ADDR_REG_10_, n10859 );
nand U20620 ( n10926, P2_ADDR_REG_10_, n10927 );
or U20621 ( n10927, n10859, P1_ADDR_REG_10_ );
nand U20622 ( n10866, n10919, n10920 );
nand U20623 ( n10919, P1_ADDR_REG_12_, n10863 );
nand U20624 ( n10920, P2_ADDR_REG_12_, n10921 );
or U20625 ( n10921, n10863, P1_ADDR_REG_12_ );
nand U20626 ( n10870, n10913, n10914 );
nand U20627 ( n10913, P1_ADDR_REG_14_, n10867 );
nand U20628 ( n10914, P2_ADDR_REG_14_, n10915 );
or U20629 ( n10915, n10867, P1_ADDR_REG_14_ );
nand U20630 ( n10874, n10907, n10908 );
nand U20631 ( n10907, P1_ADDR_REG_16_, n10871 );
nand U20632 ( n10908, P2_ADDR_REG_16_, n10909 );
or U20633 ( n10909, n10871, P1_ADDR_REG_16_ );
nand U20634 ( n10876, n10952, n10953 );
or U20635 ( n10952, n10886, n10962 );
nand U20636 ( n10953, P2_ADDR_REG_1_, n10954 );
nand U20637 ( n10954, n10962, n10886 );
nand U20638 ( n10880, n10946, n10947 );
nand U20639 ( n10946, P1_ADDR_REG_3_, n10879 );
nand U20640 ( n10947, P2_ADDR_REG_3_, n10948 );
or U20641 ( n10948, n10879, P1_ADDR_REG_3_ );
nand U20642 ( n10884, n10940, n10941 );
nand U20643 ( n10940, P1_ADDR_REG_5_, n10883 );
nand U20644 ( n10941, P2_ADDR_REG_5_, n10942 );
or U20645 ( n10942, n10883, P1_ADDR_REG_5_ );
nand U20646 ( n10890, n10934, n10935 );
nand U20647 ( n10934, P1_ADDR_REG_7_, n10889 );
nand U20648 ( n10935, P2_ADDR_REG_7_, n10936 );
or U20649 ( n10936, n10889, P1_ADDR_REG_7_ );
nand U20650 ( n10859, n10928, n10929 );
nand U20651 ( n10928, P1_ADDR_REG_9_, n10893 );
nand U20652 ( n10929, P2_ADDR_REG_9_, n10930 );
or U20653 ( n10930, n10893, P1_ADDR_REG_9_ );
nand U20654 ( n10863, n10922, n10923 );
nand U20655 ( n10922, P1_ADDR_REG_11_, n10862 );
nand U20656 ( n10923, P2_ADDR_REG_11_, n10924 );
or U20657 ( n10924, n10862, P1_ADDR_REG_11_ );
nand U20658 ( n10867, n10916, n10917 );
nand U20659 ( n10916, P1_ADDR_REG_13_, n10866 );
nand U20660 ( n10917, P2_ADDR_REG_13_, n10918 );
or U20661 ( n10918, n10866, P1_ADDR_REG_13_ );
nand U20662 ( n10871, n10910, n10911 );
nand U20663 ( n10910, P1_ADDR_REG_15_, n10870 );
nand U20664 ( n10911, P2_ADDR_REG_15_, n10912 );
or U20665 ( n10912, n10870, P1_ADDR_REG_15_ );
nand U20666 ( n10886, P1_ADDR_REG_0_, P2_ADDR_REG_0_ );
nand U20667 ( n10903, n10904, n10905 );
nand U20668 ( n10904, P1_ADDR_REG_17_, n10874 );
nand U20669 ( n10905, P2_ADDR_REG_17_, n10906 );
or U20670 ( n10906, n10874, P1_ADDR_REG_17_ );
nand U20671 ( n10901, n10899, n10902 );
nand U20672 ( n10902, P2_ADDR_REG_18_, n10897 );
xnor U20673 ( n8067, n8105, P2_IR_REG_3_ );
nand U20674 ( n1835, n6618, n6619 );
nand U20675 ( n6618, P2_REG1_REG_4_, n6519 );
nand U20676 ( n6619, n11275, n6620 );
nand U20677 ( n1675, n7998, n7999 );
nand U20678 ( n7998, P2_REG0_REG_4_, n6651 );
nand U20679 ( n7999, n11272, n6620 );
nand U20680 ( n4585, n7919, n7970 );
nand U20681 ( n7970, P2_REG3_REG_6_, n7971 );
or U20682 ( n7971, n8009, P2_REG3_REG_5_ );
or U20683 ( n7919, n7971, P2_REG3_REG_6_ );
nand U20684 ( n4349, n7971, n8008 );
nand U20685 ( n8008, P2_REG3_REG_5_, n8009 );
xnor U20686 ( n10502, P1_IR_REG_1_, n10957 );
nand U20687 ( n9050, P1_IR_REG_2_, n10001 );
or U20688 ( n10001, P1_IR_REG_0_, P1_IR_REG_1_ );
nand U20689 ( n7749, P2_IR_REG_10_, n8505 );
or U20690 ( n8505, n7853, P2_IR_REG_9_ );
nand U20691 ( n10899, P1_ADDR_REG_18_, n10903 );
nand U20692 ( n9435, n112, n9436 );
nand U20693 ( n9436, n9437, n11129 );
nor U20694 ( n9437, P1_D_REG_24_, P1_D_REG_23_ );
nand U20695 ( n8786, n8787, n8788 );
nand U20696 ( n8787, P1_REG3_REG_1_, n8794 );
nand U20697 ( n8788, n8789, n11506 );
xor U20698 ( n8789, n8790, n8791 );
nand U20699 ( n9434, n112, n9438 );
nand U20700 ( n9438, n9439, n9440 );
nor U20701 ( n9439, P1_D_REG_19_, P1_D_REG_18_ );
nor U20702 ( n9440, P1_D_REG_21_, P1_D_REG_20_ );
nand U20703 ( n5685, n7704, n7705 );
nand U20704 ( n7704, P2_IR_REG_11_, n11456 );
or U20705 ( n7705, n7706, n11455 );
nor U20706 ( n7111, n11349, n11102 );
nand U20707 ( n1183, n1184, n1186 );
nand U20708 ( n1184, n11285, n1188 );
xnor U20709 ( n1188, n1189, n1191 );
xnor U20710 ( n1191, P1_REG2_REG_2_, n1192 );
nand U20711 ( n600, n2641, n2642 );
nand U20712 ( n2641, P1_REG1_REG_2_, n2556 );
nand U20713 ( n2642, n11281, n2643 );
nand U20714 ( n440, n3911, n3912 );
nand U20715 ( n3911, P1_REG0_REG_2_, n2660 );
nand U20716 ( n3912, n11278, n2643 );
nand U20717 ( n4409, n8009, n8043 );
nand U20718 ( n8043, P2_REG3_REG_4_, P2_REG3_REG_3_ );
nand U20719 ( n1425, n8419, n8420 );
nand U20720 ( n8420, n11323, P2_IR_REG_18_ );
nor U20721 ( n8419, n8421, n8422 );
nor U20722 ( n8421, n11450, n8426 );
and U20723 ( n3979, n9403, n9404 );
nand U20724 ( n9404, n3990, n9401 );
nand U20725 ( n9403, P1_D_REG_1_, n112 );
nand U20726 ( n200, n6431, n6432 );
nand U20727 ( n6432, n11408, P1_IR_REG_18_ );
nor U20728 ( n6431, n6433, n6434 );
nor U20729 ( n6433, n11488, n6436 );
nor U20730 ( n10548, n11309, n11124 );
nand U20731 ( n1829, n10066, n10067 );
nand U20732 ( n10067, n10068, P1_IR_REG_31_ );
nand U20733 ( n10066, P1_IR_REG_6_, n11486 );
and U20734 ( n10068, n394, n8477 );
nand U20735 ( n5728, n5729, n5730 );
nand U20736 ( n5729, P2_ADDR_REG_13_, n933 );
nand U20737 ( n5730, n5408, n5731 );
xnor U20738 ( n5731, n5732, n5733 );
nand U20739 ( n1369, n9895, n9896 );
nand U20740 ( n9895, P1_IR_REG_7_, n11485 );
or U20741 ( n9896, n8382, n11484 );
nor U20742 ( n10539, n11309, n11125 );
nand U20743 ( n10223, n10336, n10337 );
nand U20744 ( n10337, P1_DATAO_REG_25_, n11264 );
nand U20745 ( n10336, P2_DATAO_REG_25_, n11328 );
nand U20746 ( n7854, P2_IR_REG_8_, n8522 );
nand U20747 ( n8522, n1013, n10978 );
nand U20748 ( n1830, n6621, n6622 );
nand U20749 ( n6621, P2_REG1_REG_3_, n6519 );
nand U20750 ( n6622, n11275, n6623 );
nand U20751 ( n1670, n8033, n8034 );
nand U20752 ( n8033, P2_REG0_REG_3_, n6651 );
nand U20753 ( n8034, n11272, n6623 );
nand U20754 ( n5701, n7652, n7653 );
nand U20755 ( n7653, n7654, P2_IR_REG_31_ );
nand U20756 ( n7652, P2_IR_REG_12_, n11456 );
and U20757 ( n7654, n7655, n7656 );
nor U20758 ( n10530, n11309, n11127 );
xor U20759 ( n5841, n5842, n5843 );
xnor U20760 ( n5843, P2_REG2_REG_18_, n897 );
xnor U20761 ( ADD_1068_U55, n783, n10875 );
xnor U20762 ( n10875, n11110, P1_ADDR_REG_18_ );
nor U20763 ( n6990, n11350, n11113 );
nand U20764 ( n4045, n7866, n7918 );
nand U20765 ( n7918, P2_REG3_REG_7_, n7919 );
or U20766 ( n7866, n7919, P2_REG3_REG_7_ );
and U20767 ( n10549, n11311, P1_REG0_REG_24_ );
nand U20768 ( n4117, n7722, n7760 );
nand U20769 ( n7760, P2_REG3_REG_10_, n7761 );
or U20770 ( n7818, n7866, P2_REG3_REG_8_ );
or U20771 ( n7761, n7818, P2_REG3_REG_9_ );
and U20772 ( n10540, n11311, P1_REG0_REG_25_ );
nand U20773 ( n3986, n9399, n9400 );
nand U20774 ( n9400, n3993, n9401 );
nand U20775 ( n9399, P1_D_REG_0_, n112 );
nor U20776 ( n6941, n11350, n11116 );
or U20777 ( n7722, n7761, P2_REG3_REG_10_ );
nand U20778 ( n595, n2644, n2645 );
nand U20779 ( n2644, P1_REG1_REG_1_, n2556 );
nand U20780 ( n2645, n11281, n2646 );
nand U20781 ( n435, n3945, n3946 );
nand U20782 ( n3945, P1_REG0_REG_1_, n2660 );
nand U20783 ( n3946, n11278, n2646 );
nor U20784 ( n7054, n11350, n11119 );
xnor U20785 ( n7791, P2_IR_REG_9_, n7853 );
nand U20786 ( n9553, n10466, n10467 );
nand U20787 ( n10467, P1_REG0_REG_31_, n11311 );
nor U20788 ( n10466, n10469, n10470 );
nor U20789 ( n10469, n11303, n11131 );
nor U20790 ( n10470, n11309, n11130 );
nand U20791 ( n5585, n5924, n5925 );
nand U20792 ( n5924, P2_REG2_REG_7_, n5869 );
nand U20793 ( n5925, P2_REG1_REG_7_, n11459 );
nand U20794 ( n5708, n5709, n5710 );
nand U20795 ( n5709, P2_ADDR_REG_12_, n933 );
nand U20796 ( n5710, n5408, n5711 );
xor U20797 ( n5711, n5712, n5713 );
and U20798 ( n10531, n11311, P1_REG0_REG_26_ );
nand U20799 ( n4425, n7761, n7817 );
nand U20800 ( n7817, P2_REG3_REG_9_, n7818 );
nand U20801 ( n1442, n9917, n9918 );
nand U20802 ( n9918, n9919, P1_IR_REG_31_ );
nand U20803 ( n9917, P1_IR_REG_8_, n11486 );
and U20804 ( n9919, n8277, n8276 );
nand U20805 ( n1825, n6624, n6625 );
nand U20806 ( n6624, P2_REG1_REG_2_, n6519 );
nand U20807 ( n6625, n11275, n6626 );
nand U20808 ( n1665, n8068, n8069 );
nand U20809 ( n8068, P2_REG0_REG_2_, n6651 );
nand U20810 ( n8069, n11272, n6626 );
nand U20811 ( n2700, n10475, n10476 );
nand U20812 ( n10476, P1_REG0_REG_30_, n11311 );
nor U20813 ( n10475, n10477, n10478 );
nor U20814 ( n10477, n11303, n11133 );
nor U20815 ( n10478, n11309, n11132 );
nand U20816 ( n1420, n8429, n8430 );
nand U20817 ( n8430, n11323, P2_IR_REG_17_ );
nor U20818 ( n8429, n8431, n8432 );
nor U20819 ( n8431, n7444, n11450 );
xnor U20820 ( n8569, P1_IR_REG_5_, n8671 );
nand U20821 ( n195, n6532, n6533 );
nand U20822 ( n6533, n11408, P1_IR_REG_17_ );
nor U20823 ( n6532, n6534, n6535 );
nor U20824 ( n6535, n6536, n11489 );
nand U20825 ( n7656, P2_IR_REG_12_, n8488 );
nand U20826 ( n8488, n8487, n11010 );
nand U20827 ( n590, n2647, n2648 );
nand U20828 ( n2647, P1_REG1_REG_0_, n2556 );
nand U20829 ( n2648, n11281, n2649 );
nand U20830 ( n430, n3963, n3964 );
nand U20831 ( n3963, P1_REG0_REG_0_, n2660 );
nand U20832 ( n3964, n11278, n2649 );
nand U20833 ( n10232, n10331, n10332 );
nand U20834 ( n10332, P1_DATAO_REG_26_, n11264 );
nand U20835 ( n10331, P2_DATAO_REG_26_, n11327 );
nor U20836 ( n10521, n11309, n11137 );
nand U20837 ( n1443, n10122, n10123 );
nand U20838 ( n10123, n10124, P1_IR_REG_31_ );
nand U20839 ( n10122, P1_IR_REG_10_, n11486 );
and U20840 ( n10124, n386, n8260 );
xor U20841 ( n5821, n5822, n5823 );
xnor U20842 ( n5823, n896, P2_REG2_REG_17_ );
nand U20843 ( n5613, n5963, n5964 );
nand U20844 ( n5963, P2_REG2_REG_8_, n11287 );
nand U20845 ( n5964, P2_REG1_REG_8_, n11459 );
nand U20846 ( n4216, n7818, n7865 );
nand U20847 ( n7865, P2_REG3_REG_8_, n7866 );
nand U20848 ( n4536, n4537, n4538 );
nand U20849 ( n4537, P2_REG3_REG_2_, n906 );
nand U20850 ( n4538, n11469, n4539 );
nand U20851 ( n4539, n4540, n4541 );
nand U20852 ( n8670, P1_IR_REG_4_, n10018 );
nand U20853 ( n10018, n408, n10971 );
nand U20854 ( n5721, n7615, n7616 );
nand U20855 ( n7615, P2_IR_REG_13_, n11456 );
or U20856 ( n7616, n7617, n11455 );
nand U20857 ( n1436, n9932, n9933 );
nand U20858 ( n9932, P1_IR_REG_9_, n11485 );
or U20859 ( n9933, n8265, n11484 );
nand U20860 ( n4531, n7674, n7721 );
nand U20861 ( n7721, P2_REG3_REG_11_, n7722 );
xnor U20862 ( ADD_1068_U56, n10873, n10874 );
xnor U20863 ( n10873, P2_ADDR_REG_17_, P1_ADDR_REG_17_ );
nand U20864 ( n1820, n6627, n6628 );
nand U20865 ( n6627, P2_REG1_REG_1_, n6519 );
nand U20866 ( n6628, n11275, n6629 );
nand U20867 ( n1660, n8107, n8108 );
nand U20868 ( n8107, P2_REG0_REG_1_, n6651 );
nand U20869 ( n8108, n11272, n6629 );
nand U20870 ( n5405, n5406, n5407 );
nand U20871 ( n5407, n5408, n5409 );
nand U20872 ( n5406, P2_IR_REG_0_, n5414 );
nand U20873 ( n5409, n5410, n5411 );
nor U20874 ( n10496, n11309, n11142 );
nand U20875 ( n5414, n5415, n937 );
nor U20876 ( n5415, n5416, n5417 );
nor U20877 ( n5417, P2_REG2_REG_0_, n5418 );
nor U20878 ( n5416, P2_REG1_REG_0_, n5419 );
or U20879 ( n7674, n7722, P2_REG3_REG_11_ );
nand U20880 ( n4495, n7594, n7628 );
nand U20881 ( n7628, P2_REG3_REG_13_, n7629 );
or U20882 ( n7629, n7674, P2_REG3_REG_12_ );
and U20883 ( n10522, n11311, P1_REG0_REG_27_ );
nand U20884 ( n5659, n5910, n5911 );
nand U20885 ( n5910, P2_REG2_REG_10_, n11287 );
nand U20886 ( n5911, P2_REG1_REG_10_, n11459 );
nand U20887 ( n6511, n8240, n8241 );
nand U20888 ( n8241, n8242, n8243 );
nand U20889 ( n8240, P2_D_REG_1_, n954 );
nand U20890 ( n5905, n5912, n5913 );
nand U20891 ( n5912, P2_REG2_REG_11_, n5869 );
nand U20892 ( n5913, P2_REG1_REG_11_, n11459 );
nand U20893 ( n4289, n7629, n7673 );
nand U20894 ( n7673, P2_REG3_REG_12_, n7674 );
and U20895 ( n10497, n11311, P1_REG0_REG_28_ );
nand U20896 ( n5744, n7578, n7579 );
nand U20897 ( n7579, n7580, P2_IR_REG_31_ );
nand U20898 ( n7578, P2_IR_REG_14_, n11456 );
and U20899 ( n7580, n889, n7581 );
or U20900 ( n7594, n7629, P2_REG3_REG_13_ );
nor U20901 ( n10487, n11309, n11147 );
nand U20902 ( n8477, P1_IR_REG_6_, n10069 );
or U20903 ( n10069, n8671, P1_IR_REG_5_ );
nand U20904 ( n6503, n11375, P2_REG3_REG_0_ );
nand U20905 ( n1415, n8436, n8437 );
nand U20906 ( n8437, n11323, P2_IR_REG_16_ );
nor U20907 ( n8436, n8438, n8439 );
nor U20908 ( n8438, n11449, n8443 );
nand U20909 ( n190, n6568, n6569 );
nand U20910 ( n6569, n11408, P1_IR_REG_16_ );
nor U20911 ( n6568, n6570, n6571 );
nor U20912 ( n6570, n11488, n6573 );
nand U20913 ( n6485, n11377, P2_REG3_REG_1_ );
nand U20914 ( n6473, n11377, P2_REG3_REG_2_ );
nand U20915 ( n5634, n5915, n5916 );
nand U20916 ( n5915, P2_REG2_REG_9_, n11287 );
nand U20917 ( n5916, P2_REG1_REG_9_, n11459 );
nand U20918 ( n8234, n954, n8235 );
nand U20919 ( n8235, n8236, n11135 );
nor U20920 ( n8236, P2_D_REG_24_, P2_D_REG_23_ );
nand U20921 ( n7581, P2_IR_REG_14_, n8463 );
or U20922 ( n8463, n7655, P2_IR_REG_13_ );
nand U20923 ( n8233, n954, n8237 );
nand U20924 ( n8237, n8238, n8239 );
nor U20925 ( n8238, P2_D_REG_19_, P2_D_REG_18_ );
nor U20926 ( n8239, P2_D_REG_21_, P2_D_REG_20_ );
xnor U20927 ( n7617, P2_IR_REG_13_, n7655 );
and U20928 ( n10488, n11311, P1_REG0_REG_29_ );
nand U20929 ( n4227, n4228, n4229 );
nand U20930 ( n4228, P2_REG3_REG_1_, n906 );
nand U20931 ( n4229, n11470, n4230 );
nand U20932 ( n4230, n4231, n4232 );
nand U20933 ( n5801, n5802, n934 );
xnor U20934 ( n5802, n5803, n5804 );
xnor U20935 ( n5803, n894, P2_REG2_REG_16_ );
nand U20936 ( n10315, n10326, n10327 );
nand U20937 ( n10327, P1_DATAO_REG_27_, n11264 );
nand U20938 ( n10326, P2_DATAO_REG_27_, n11327 );
nand U20939 ( n5691, n5692, n934 );
xor U20940 ( n5692, n5693, n5694 );
xnor U20941 ( n5694, P2_REG2_REG_11_, n5685 );
nand U20942 ( n5667, n5668, n934 );
xnor U20943 ( n5668, n5669, n5670 );
xnor U20944 ( n5669, P2_REG2_REG_10_, n882 );
nand U20945 ( n5776, n5777, n934 );
xor U20946 ( n5777, n5778, n5779 );
xnor U20947 ( n5779, P2_REG2_REG_15_, n5769 );
nand U20948 ( n5750, n5751, n934 );
xnor U20949 ( n5751, n5752, n5753 );
xnor U20950 ( n5752, P2_REG2_REG_14_, n888 );
nand U20951 ( n5639, n5640, n5641 );
nand U20952 ( n5640, P2_ADDR_REG_9_, n933 );
nand U20953 ( n5641, n5642, n934 );
xor U20954 ( n5642, n5643, n5644 );
nand U20955 ( n5619, n5620, n5621 );
nand U20956 ( n5620, P2_ADDR_REG_8_, n933 );
nand U20957 ( n5621, n5622, n934 );
xnor U20958 ( n5622, n5623, n5624 );
nand U20959 ( n5594, n5595, n5596 );
nand U20960 ( n5595, P2_ADDR_REG_7_, n933 );
nand U20961 ( n5596, n5597, n934 );
xor U20962 ( n5597, n5598, n5599 );
nand U20963 ( n5563, n5564, n5565 );
nand U20964 ( n5564, P2_ADDR_REG_6_, n933 );
nand U20965 ( n5565, n5566, n934 );
xnor U20966 ( n5566, n5567, n5568 );
nand U20967 ( n5538, n5539, n5540 );
nand U20968 ( n5539, P2_ADDR_REG_5_, n933 );
nand U20969 ( n5540, n5541, n934 );
xor U20970 ( n5541, n5542, n5543 );
nand U20971 ( n5512, n5513, n5514 );
nand U20972 ( n5513, P2_ADDR_REG_4_, n933 );
nand U20973 ( n5514, n5515, n934 );
xnor U20974 ( n5515, n5516, n5517 );
nand U20975 ( n5493, n5494, n5495 );
nand U20976 ( n5494, P2_ADDR_REG_3_, n933 );
nand U20977 ( n5495, n5496, n934 );
xor U20978 ( n5496, n5497, n5498 );
nand U20979 ( n5468, n5469, n5470 );
nand U20980 ( n5469, P2_ADDR_REG_2_, n933 );
nand U20981 ( n5470, n5471, n934 );
xnor U20982 ( n5471, n5472, n5473 );
nand U20983 ( n8260, P1_IR_REG_10_, n10125 );
or U20984 ( n10125, n8277, P1_IR_REG_9_ );
nand U20985 ( n5421, n5422, n5423 );
nand U20986 ( n5422, P2_ADDR_REG_0_, n933 );
nand U20987 ( n5423, n934, n5424 );
nand U20988 ( n1704, n9849, n9850 );
nand U20989 ( n9849, P1_IR_REG_13_, n11485 );
or U20990 ( n9850, n7329, n11484 );
nor U20991 ( n6875, n11350, n11140 );
nor U20992 ( n5782, n5419, n5796 );
xnor U20993 ( n5796, n5797, n5798 );
xnor U20994 ( n5798, P2_REG1_REG_16_, n5795 );
xor U20995 ( ADD_1068_U57, n10871, n10872 );
xor U20996 ( n10872, P2_ADDR_REG_16_, P1_ADDR_REG_16_ );
nand U20997 ( n4083, n7551, n7593 );
nand U20998 ( n7593, P2_REG3_REG_14_, n7594 );
nand U20999 ( n1479, n10088, n10089 );
nand U21000 ( n10088, P1_IR_REG_11_, n11486 );
or U21001 ( n10089, n8251, n11485 );
nand U21002 ( n1519, n10109, n10110 );
nand U21003 ( n10110, n10111, P1_IR_REG_31_ );
nand U21004 ( n10109, P1_IR_REG_12_, n11486 );
and U21005 ( n10111, n7800, n7799 );
nand U21006 ( n1815, n6630, n6631 );
nand U21007 ( n6630, P2_REG1_REG_0_, n6519 );
nand U21008 ( n6631, n11275, n6632 );
nand U21009 ( n1655, n8131, n8132 );
nand U21010 ( n8131, P2_REG0_REG_0_, n6651 );
nand U21011 ( n8132, n11272, n6632 );
nand U21012 ( n5769, n7532, n7533 );
nand U21013 ( n7532, P2_IR_REG_15_, n11456 );
or U21014 ( n7533, n7534, n11455 );
or U21015 ( n7551, n7594, P2_REG3_REG_14_ );
nor U21016 ( n6813, n11350, n11145 );
xnor U21017 ( n7329, P1_IR_REG_13_, n7800 );
nand U21018 ( n8276, P1_IR_REG_8_, n9920 );
nand U21019 ( n9920, n9897, n11008 );
nor U21020 ( n5673, n5419, n5686 );
xor U21021 ( n5686, n5687, n5688 );
xnor U21022 ( n5688, n884, P2_REG1_REG_11_ );
nor U21023 ( n5756, n5419, n5771 );
xor U21024 ( n5771, n5772, n5773 );
xnor U21025 ( n5773, n893, P2_REG1_REG_15_ );
xnor U21026 ( n8265, P1_IR_REG_9_, n8277 );
nand U21027 ( n4467, n7239, n7288 );
nand U21028 ( n7288, P2_REG3_REG_20_, n7289 );
or U21029 ( n7239, n7289, P2_REG3_REG_20_ );
or U21030 ( n7462, n7511, P2_REG3_REG_16_ );
or U21031 ( n7400, n7462, P2_REG3_REG_17_ );
or U21032 ( n7511, n7551, P2_REG3_REG_15_ );
or U21033 ( n7342, n7400, P2_REG3_REG_18_ );
or U21034 ( n7289, n7342, P2_REG3_REG_19_ );
nand U21035 ( n4721, n7511, n7550 );
nand U21036 ( n7550, P2_REG3_REG_15_, n7551 );
xnor U21037 ( n2448, P1_REG3_REG_4_, n11002 );
nand U21038 ( n7799, P1_IR_REG_12_, n10112 );
nand U21039 ( n10112, n10090, n11037 );
xor U21040 ( n2403, P1_REG3_REG_6_, n10711 );
nand U21041 ( n10720, P1_REG3_REG_4_, P1_REG3_REG_3_ );
nand U21042 ( n1879, n2671, n2672 );
nor U21043 ( n2671, n324, n2673 );
nor U21044 ( n2673, n11418, n2675 );
nor U21045 ( n2675, P1_B_REG, n1249 );
nand U21046 ( n1410, n8447, n8448 );
nand U21047 ( n8448, n11323, P2_IR_REG_15_ );
nor U21048 ( n8447, n8449, n8450 );
nor U21049 ( n8449, n7534, n11450 );
nand U21050 ( n4332, n7462, n7510 );
nand U21051 ( n7510, P2_REG3_REG_16_, n7511 );
nand U21052 ( n1405, n8454, n8455 );
nand U21053 ( n8455, n11323, P2_IR_REG_14_ );
nor U21054 ( n8454, n8456, n8457 );
nor U21055 ( n8456, n11449, n8461 );
nor U21056 ( n6664, n11350, n11152 );
nand U21057 ( n185, n6606, n6607 );
nand U21058 ( n6607, n11408, P1_IR_REG_15_ );
nor U21059 ( n6606, n6608, n6609 );
nor U21060 ( n6609, n6610, n11489 );
nand U21061 ( n180, n6729, n6730 );
nand U21062 ( n6730, n11408, P1_IR_REG_14_ );
nor U21063 ( n6729, n6731, n6732 );
nor U21064 ( n6731, n11488, n6734 );
nand U21065 ( n4371, n7400, n7461 );
nand U21066 ( n7461, P2_REG3_REG_17_, n7462 );
nand U21067 ( n10301, n10317, n10318 );
nand U21068 ( n10318, P1_DATAO_REG_28_, n11266 );
nand U21069 ( n10317, P2_DATAO_REG_28_, n11328 );
nand U21070 ( n10702, n10711, P1_REG3_REG_6_ );
nand U21071 ( n10684, n10693, P1_REG3_REG_8_ );
nand U21072 ( n10666, n10675, P1_REG3_REG_10_ );
nand U21073 ( n10648, n10657, P1_REG3_REG_12_ );
nand U21074 ( n4158, n7289, n7341 );
nand U21075 ( n7341, P2_REG3_REG_19_, n7342 );
xor U21076 ( n2317, P1_REG3_REG_10_, n10675 );
nand U21077 ( n4645, n6873, n6938 );
nand U21078 ( n6938, P2_REG3_REG_26_, n6939 );
or U21079 ( n6939, n6988, P2_REG3_REG_25_ );
or U21080 ( n7109, n7174, P2_REG3_REG_22_ );
or U21081 ( n6873, n6939, P2_REG3_REG_26_ );
or U21082 ( n7052, n7109, P2_REG3_REG_23_ );
or U21083 ( n7174, n7239, P2_REG3_REG_21_ );
or U21084 ( n6988, n7052, P2_REG3_REG_24_ );
nor U21085 ( n6704, n11350, n11155 );
nand U21086 ( n4512, n7109, n7173 );
nand U21087 ( n7173, P2_REG3_REG_22_, n7174 );
xnor U21088 ( ADD_1068_U58, n10869, n10870 );
xnor U21089 ( n10869, P2_ADDR_REG_15_, P1_ADDR_REG_15_ );
nand U21090 ( n5817, n7442, n7443 );
nand U21091 ( n7442, P2_IR_REG_17_, n11456 );
or U21092 ( n7443, n7444, n11455 );
xnor U21093 ( n7444, P2_IR_REG_17_, n7494 );
nor U21094 ( n10782, n10783, n10957 );
nor U21095 ( n10783, n10784, n10785 );
nor U21096 ( n10784, P1_REG1_REG_0_, n1194 );
nand U21097 ( n10785, n10786, n1229 );
nand U21098 ( n5795, n7491, n7492 );
nand U21099 ( n7491, P2_IR_REG_16_, n11457 );
nand U21100 ( n7492, n7493, P2_IR_REG_31_ );
and U21101 ( n7493, n7494, n7495 );
nand U21102 ( n7495, P2_IR_REG_16_, n8446 );
nand U21103 ( n8446, n8445, n11038 );
nand U21104 ( n1095, n10615, n10616 );
nand U21105 ( n10616, n11447, n2187 );
nand U21106 ( n10615, P1_DATAO_REG_17_, n11445 );
nand U21107 ( n1085, n10633, n10634 );
nand U21108 ( n10634, n11448, n2226 );
nand U21109 ( n10633, P1_DATAO_REG_15_, n11445 );
nand U21110 ( n1100, n10595, n10596 );
nand U21111 ( n10596, n11447, n2163 );
nand U21112 ( n10595, P1_DATAO_REG_18_, n11445 );
nand U21113 ( n1115, n10568, n10569 );
nand U21114 ( n10569, n11447, n2097 );
nand U21115 ( n10568, P1_DATAO_REG_21_, n11445 );
nand U21116 ( n1080, n10642, n10643 );
nand U21117 ( n10643, n11448, n2253 );
nand U21118 ( n10642, P1_DATAO_REG_14_, n11445 );
nand U21119 ( n1140, n10523, n10524 );
nand U21120 ( n10524, n11447, n1984 );
nand U21121 ( n10523, P1_DATAO_REG_26_, n11445 );
nand U21122 ( n1130, n10541, n10542 );
nand U21123 ( n10542, n11447, n2029 );
nand U21124 ( n10541, P1_DATAO_REG_24_, n11445 );
nand U21125 ( n1125, n10550, n10551 );
nand U21126 ( n10551, n11447, n2046 );
nand U21127 ( n10550, P1_DATAO_REG_23_, n11445 );
nand U21128 ( n1120, n10559, n10560 );
nand U21129 ( n10560, n11447, n2074 );
nand U21130 ( n10559, P1_DATAO_REG_22_, n11445 );
nand U21131 ( n1150, n10489, n10490 );
nand U21132 ( n10490, n11447, n1939 );
nand U21133 ( n10489, P1_DATAO_REG_28_, n11445 );
nand U21134 ( n1110, n10577, n10578 );
nand U21135 ( n10578, n11447, n2118 );
nand U21136 ( n10577, P1_DATAO_REG_20_, n11445 );
nand U21137 ( n1165, n10464, n10465 );
nand U21138 ( n10465, n11448, n9553 );
nand U21139 ( n10464, P1_DATAO_REG_31_, n11445 );
nand U21140 ( n1135, n10532, n10533 );
nand U21141 ( n10533, n11447, n2007 );
nand U21142 ( n10532, P1_DATAO_REG_25_, n11445 );
nand U21143 ( n1160, n10473, n10474 );
nand U21144 ( n10474, n11447, n2700 );
nand U21145 ( n10473, P1_DATAO_REG_30_, n11445 );
nand U21146 ( n1155, n10479, n10480 );
nand U21147 ( n10480, n11447, n1909 );
nand U21148 ( n10479, P1_DATAO_REG_29_, n11445 );
nand U21149 ( n1105, n10586, n10587 );
nand U21150 ( n10587, n11447, n2136 );
nand U21151 ( n10586, P1_DATAO_REG_19_, n11445 );
nand U21152 ( n1090, n10624, n10625 );
nand U21153 ( n10625, n11448, n2209 );
nand U21154 ( n10624, P1_DATAO_REG_16_, n11445 );
nand U21155 ( n1075, n10651, n10652 );
nand U21156 ( n10652, n11448, n2277 );
nand U21157 ( n10651, P1_DATAO_REG_13_, n11445 );
nand U21158 ( n1145, n10514, n10515 );
nand U21159 ( n10515, n11447, n1962 );
nand U21160 ( n10514, P1_DATAO_REG_27_, n11445 );
nand U21161 ( n5690, P2_ADDR_REG_11_, n933 );
nand U21162 ( n5666, P2_ADDR_REG_10_, n933 );
nand U21163 ( n5800, P2_ADDR_REG_16_, n933 );
nand U21164 ( n5775, P2_ADDR_REG_15_, n933 );
nand U21165 ( n5749, P2_ADDR_REG_14_, n933 );
nand U21166 ( n9378, n10834, n10835 );
nand U21167 ( n10834, P1_IR_REG_23_, n11487 );
nand U21168 ( n10835, n10836, P1_IR_REG_31_ );
and U21169 ( n10836, n5395, n5394 );
nand U21170 ( n4310, n6939, n6987 );
nand U21171 ( n6987, P2_REG3_REG_25_, n6988 );
nand U21172 ( n6034, n933, P2_ADDR_REG_19_ );
nand U21173 ( n1060, n10678, n10679 );
nand U21174 ( n10679, n11448, n2342 );
nand U21175 ( n10678, P1_DATAO_REG_10_, n11446 );
nand U21176 ( n1040, n10714, n10715 );
nand U21177 ( n10715, n11448, n2429 );
nand U21178 ( n10714, P1_DATAO_REG_6_, n11446 );
nand U21179 ( n1035, n10723, n10724 );
nand U21180 ( n10724, n11448, n2447 );
nand U21181 ( n10723, P1_DATAO_REG_5_, n11446 );
nand U21182 ( n1030, n10731, n10732 );
nand U21183 ( n10732, n11448, n2474 );
nand U21184 ( n10731, P1_DATAO_REG_4_, n11446 );
nand U21185 ( n1065, n10669, n10670 );
nand U21186 ( n10670, n11448, n2316 );
nand U21187 ( n10669, P1_DATAO_REG_11_, n11446 );
nand U21188 ( n1050, n10696, n10697 );
nand U21189 ( n10697, n11448, n2386 );
nand U21190 ( n10696, P1_DATAO_REG_8_, n11446 );
nand U21191 ( n1015, n10755, n10756 );
nand U21192 ( n10756, n11448, n2537 );
nand U21193 ( n10755, P1_DATAO_REG_1_, n11446 );
nand U21194 ( n1025, n10739, n10740 );
nand U21195 ( n10740, n11448, n2494 );
nand U21196 ( n10739, P1_DATAO_REG_3_, n11446 );
nand U21197 ( n1055, n10687, n10688 );
nand U21198 ( n10688, n11448, n2359 );
nand U21199 ( n10687, P1_DATAO_REG_9_, n11446 );
nand U21200 ( n1045, n10705, n10706 );
nand U21201 ( n10706, n11448, n2409 );
nand U21202 ( n10705, P1_DATAO_REG_7_, n11446 );
nand U21203 ( n1020, n10747, n10748 );
nand U21204 ( n10748, n11448, n2516 );
nand U21205 ( n10747, P1_DATAO_REG_2_, n11446 );
nand U21206 ( n1070, n10660, n10661 );
nand U21207 ( n10661, n11448, n2299 );
nand U21208 ( n10660, P1_DATAO_REG_12_, n11446 );
nand U21209 ( n1010, n10763, n10764 );
nand U21210 ( n10764, n11448, n3956 );
nand U21211 ( n10763, P1_DATAO_REG_0_, n11446 );
xor U21212 ( n2271, P1_REG3_REG_12_, n10657 );
nand U21213 ( n4267, n7174, n7238 );
nand U21214 ( n7238, P2_REG3_REG_21_, n7239 );
nand U21215 ( n1576, n9798, n9799 );
nand U21216 ( n9798, P1_IR_REG_15_, n11485 );
or U21217 ( n9799, n6610, n11484 );
nand U21218 ( n1199, n1201, n1202 );
nand U21219 ( n1201, P1_ADDR_REG_2_, n1203 );
nand U21220 ( n1202, n69, n1192 );
nor U21221 ( n6750, n11350, n11149 );
nand U21222 ( n920, n1611, n1612 );
nor U21223 ( n1611, n1642, n1643 );
nor U21224 ( n1612, n1613, n1614 );
and U21225 ( n1642, n1203, P1_ADDR_REG_17_ );
nand U21226 ( n970, n1351, n1352 );
nor U21227 ( n1351, n1382, n1383 );
nor U21228 ( n1352, n1353, n1354 );
and U21229 ( n1382, n1203, P1_ADDR_REG_7_ );
nand U21230 ( n980, n1279, n1281 );
nor U21231 ( n1279, n1322, n1323 );
nor U21232 ( n1281, n1282, n1283 );
and U21233 ( n1322, n1203, P1_ADDR_REG_5_ );
and U21234 ( n5446, n933, P2_ADDR_REG_1_ );
nand U21235 ( n940, n1498, n1499 );
nor U21236 ( n1498, n1543, n1544 );
nor U21237 ( n1499, n1501, n1502 );
and U21238 ( n1543, n1203, P1_ADDR_REG_13_ );
nand U21239 ( n955, n1414, n1416 );
nor U21240 ( n1414, n1463, n1464 );
nor U21241 ( n1416, n1417, n1418 );
and U21242 ( n1463, n1203, P1_ADDR_REG_10_ );
nand U21243 ( n1395, n8478, n8479 );
nand U21244 ( n8479, n11323, P2_IR_REG_12_ );
nor U21245 ( n8478, n8480, n8481 );
nor U21246 ( n8480, n11449, n8485 );
nand U21247 ( n4563, n7342, n7399 );
nand U21248 ( n7399, P2_REG3_REG_18_, n7400 );
nand U21249 ( n170, n7793, n7794 );
nand U21250 ( n7794, n11409, P1_IR_REG_12_ );
nor U21251 ( n7793, n7795, n7796 );
nor U21252 ( n7795, n11488, n7798 );
nand U21253 ( n950, n1466, n1467 );
nor U21254 ( n1466, n1481, n1482 );
nor U21255 ( n1467, n1468, n1469 );
and U21256 ( n1481, n1203, P1_ADDR_REG_11_ );
nand U21257 ( n960, n1399, n1401 );
nor U21258 ( n1399, n1412, n1413 );
nor U21259 ( n1401, n1402, n1403 );
and U21260 ( n1412, n1203, P1_ADDR_REG_9_ );
nand U21261 ( n990, n1204, n1206 );
nor U21262 ( n1204, n1231, n1232 );
nor U21263 ( n1206, n1207, n1208 );
and U21264 ( n1231, n1203, P1_ADDR_REG_3_ );
nand U21265 ( n930, n1564, n1566 );
nor U21266 ( n1564, n1581, n1582 );
nor U21267 ( n1566, n1567, n1568 );
and U21268 ( n1581, n1203, P1_ADDR_REG_15_ );
nor U21269 ( n10781, P1_IR_REG_0_, n10787 );
nor U21270 ( n10787, n10788, n10789 );
and U21271 ( n10788, P1_REG2_REG_0_, n1187 );
nor U21272 ( n10789, n10963, n1194 );
nand U21273 ( n925, n1583, n1584 );
nor U21274 ( n1583, n1608, n1609 );
nor U21275 ( n1584, n1586, n1587 );
and U21276 ( n1608, n1203, P1_ADDR_REG_16_ );
nand U21277 ( n935, n1546, n1547 );
nor U21278 ( n1546, n1562, n1563 );
nor U21279 ( n1547, n1548, n1549 );
and U21280 ( n1562, n1203, P1_ADDR_REG_14_ );
nand U21281 ( n945, n1483, n1484 );
nor U21282 ( n1483, n1496, n1497 );
nor U21283 ( n1484, n1486, n1487 );
and U21284 ( n1496, n1203, P1_ADDR_REG_12_ );
nand U21285 ( n965, n1384, n1386 );
nor U21286 ( n1384, n1397, n1398 );
nor U21287 ( n1386, n1387, n1388 );
and U21288 ( n1397, n1203, P1_ADDR_REG_8_ );
nand U21289 ( n975, n1324, n1326 );
nor U21290 ( n1324, n1348, n1349 );
nor U21291 ( n1326, n1327, n1328 );
and U21292 ( n1348, n1203, P1_ADDR_REG_6_ );
nand U21293 ( n10630, n10639, P1_REG3_REG_14_ );
nand U21294 ( n10601, n10621, P1_REG3_REG_16_ );
nand U21295 ( n10583, n10592, P1_REG3_REG_18_ );
nand U21296 ( n10565, P1_REG3_REG_20_, n10574 );
nand U21297 ( n5394, P1_IR_REG_23_, n10832 );
nand U21298 ( n5712, n5965, n5966 );
nand U21299 ( n5965, P2_REG2_REG_12_, n5869 );
nand U21300 ( n5966, P2_REG1_REG_12_, n11459 );
nand U21301 ( n1400, n8464, n8465 );
nand U21302 ( n8465, n11323, P2_IR_REG_13_ );
nor U21303 ( n8464, n8466, n8467 );
nor U21304 ( n8467, n7617, n11451 );
nand U21305 ( n4101, n7052, n7108 );
nand U21306 ( n7108, P2_REG3_REG_23_, n7109 );
nand U21307 ( n175, n7325, n7326 );
nand U21308 ( n7326, n11408, P1_IR_REG_13_ );
nor U21309 ( n7325, n7327, n7328 );
nor U21310 ( n7328, n7329, n11489 );
xor U21311 ( n2361, P1_REG3_REG_8_, n10693 );
nand U21312 ( n10279, n10296, n10297 );
nand U21313 ( n10297, P1_DATAO_REG_29_, n11266 );
nand U21314 ( n10296, P2_DATAO_REG_29_, n11328 );
xor U21315 ( n2047, P1_REG3_REG_22_, n10556 );
nor U21316 ( n6113, n6811, P2_REG3_REG_28_ );
nand U21317 ( n4198, n1149, n6810 );
nand U21318 ( n6810, P2_REG3_REG_28_, n6811 );
or U21319 ( n6811, n6873, P2_REG3_REG_27_ );
xor U21320 ( ADD_1068_U59, n10867, n10868 );
xor U21321 ( n10868, P2_ADDR_REG_14_, P1_ADDR_REG_14_ );
nand U21322 ( n6574, P1_IR_REG_16_, n10140 );
nand U21323 ( n10140, n9800, n11055 );
nand U21324 ( n1781, n10137, n10138 );
nand U21325 ( n10137, P1_IR_REG_16_, n11486 );
nand U21326 ( n10138, n10139, P1_IR_REG_31_ );
and U21327 ( n10139, n6575, n6574 );
nand U21328 ( n1196, n1848, n1849 );
nand U21329 ( n1849, n1851, P1_REG1_REG_0_ );
nor U21330 ( n1851, n1852, n10957 );
nor U21331 ( n1852, P1_REG1_REG_1_, n1853 );
nand U21332 ( n1606, n1782, n1783 );
nand U21333 ( n1782, n1578, n1576 );
nand U21334 ( n1783, P1_REG1_REG_15_, n1784 );
or U21335 ( n1784, n1578, n1576 );
nor U21336 ( n1824, n1828, n1379 );
nor U21337 ( n1828, P1_REG1_REG_7_, n1369 );
nor U21338 ( n1776, n1779, n1639 );
nor U21339 ( n1779, P1_REG1_REG_17_, n1629 );
nor U21340 ( n1833, n1837, n1838 );
nor U21341 ( n1837, P1_REG1_REG_5_, n1304 );
nand U21342 ( n1838, n1839, n1269 );
nand U21343 ( n1839, n1841, n1842 );
nand U21344 ( n1769, n1768, n1771 );
nand U21345 ( n1771, P1_REG1_REG_18_, n1766 );
nand U21346 ( n1578, n1786, n1787 );
nand U21347 ( n1786, n1558, n1561 );
nand U21348 ( n1787, P1_REG1_REG_14_, n1788 );
or U21349 ( n1788, n1558, n1561 );
nor U21350 ( n1841, n1321, n1844 );
nor U21351 ( n1844, n1846, n1847 );
nor U21352 ( n1846, P1_REG1_REG_2_, n1192 );
nand U21353 ( n1847, n1228, n1196 );
nor U21354 ( n1818, n56, n1821 );
nor U21355 ( n1821, P1_REG1_REG_8_, n1442 );
nor U21356 ( n1802, n54, n1804 );
nor U21357 ( n1804, P1_REG1_REG_11_, n1479 );
xor U21358 ( n2091, P1_REG3_REG_20_, n10574 );
nand U21359 ( n1390, n8489, n8490 );
nand U21360 ( n8490, n11323, P2_IR_REG_11_ );
nor U21361 ( n8489, n8491, n8492 );
nor U21362 ( n8491, n7706, n11451 );
nand U21363 ( n1573, n1693, n1694 );
nand U21364 ( n1693, n1554, n1561 );
nand U21365 ( n1694, P1_REG2_REG_14_, n1696 );
or U21366 ( n1696, n1554, n1561 );
nor U21367 ( n1668, n358, n1677 );
not U21368 ( n358, n1671 );
nand U21369 ( n1677, n1676, n1678 );
nand U21370 ( n1678, P1_REG2_REG_18_, n1673 );
nor U21371 ( n1741, n1744, n1746 );
nor U21372 ( n1744, P1_REG2_REG_5_, n1304 );
nand U21373 ( n1746, n1747, n1263 );
nand U21374 ( n1747, n1748, n1749 );
nor U21375 ( n1733, n1737, n1367 );
nor U21376 ( n1737, P1_REG2_REG_7_, n1369 );
nor U21377 ( n1684, n1688, n1627 );
nor U21378 ( n1688, P1_REG2_REG_17_, n1629 );
nor U21379 ( n1748, n1303, n1752 );
nor U21380 ( n1752, n1753, n1754 );
nor U21381 ( n1753, P1_REG2_REG_2_, n1192 );
nand U21382 ( n1754, n1219, n1189 );
nor U21383 ( n1727, n63, n1729 );
nor U21384 ( n1729, P1_REG2_REG_8_, n1442 );
nor U21385 ( n1711, n61, n1713 );
nor U21386 ( n1713, P1_REG2_REG_11_, n1479 );
nand U21387 ( n1597, n1689, n1691 );
nand U21388 ( n1689, n1573, n1576 );
nand U21389 ( n1691, P1_REG2_REG_15_, n1692 );
or U21390 ( n1692, n1573, n1576 );
nor U21391 ( n5424, n10966, P2_IR_REG_0_ );
nor U21392 ( n5412, n10967, P2_IR_REG_0_ );
nand U21393 ( n165, n8247, n8248 );
nand U21394 ( n8248, n11409, P1_IR_REG_11_ );
nor U21395 ( n8247, n8249, n8250 );
nor U21396 ( n8250, n8251, n11489 );
nor U21397 ( n1182, n1193, n1194 );
xor U21398 ( n1193, n1196, n1197 );
xnor U21399 ( n1197, P1_REG1_REG_2_, n1192 );
xnor U21400 ( n10270, n10284, SI_31_ );
nand U21401 ( n10284, n10285, n10286 );
nand U21402 ( n10286, P1_DATAO_REG_31_, n11266 );
nand U21403 ( n10285, P2_DATAO_REG_31_, n11326 );
nand U21404 ( n4062, n6811, n6872 );
nand U21405 ( n6872, P2_REG3_REG_27_, n6873 );
nand U21406 ( n4392, n6988, n7051 );
nand U21407 ( n7051, P2_REG3_REG_24_, n7052 );
nand U21408 ( n1561, n9825, n9826 );
nand U21409 ( n9825, P1_IR_REG_14_, n11485 );
nand U21410 ( n9826, n9827, P1_IR_REG_31_ );
and U21411 ( n9827, n371, n6735 );
nand U21412 ( n10273, n10287, n10288 );
nand U21413 ( n10288, P1_DATAO_REG_30_, n11266 );
nand U21414 ( n10287, P2_DATAO_REG_30_, n11327 );
nand U21415 ( n5837, n7384, n7385 );
nand U21416 ( n7384, P2_IR_REG_18_, n11457 );
nand U21417 ( n7385, n7386, P2_IR_REG_31_ );
and U21418 ( n7386, n898, n7387 );
nand U21419 ( n7387, P2_IR_REG_18_, n8428 );
or U21420 ( n8428, n7494, P2_IR_REG_17_ );
xnor U21421 ( n8287, n8201, P2_IR_REG_23_ );
nand U21422 ( n4733, n8285, n8286 );
nand U21423 ( n8285, P2_IR_REG_23_, n11458 );
or U21424 ( n8286, n11458, n8287 );
nand U21425 ( n5881, n5888, n5889 );
nand U21426 ( n5888, P2_REG2_REG_16_, n11287 );
nand U21427 ( n5889, P2_REG1_REG_16_, n11460 );
nand U21428 ( n10547, P1_REG3_REG_22_, n10556 );
and U21429 ( n5768, n5886, n5887 );
nand U21430 ( n5886, P2_REG2_REG_15_, n5869 );
nand U21431 ( n5887, P2_REG1_REG_15_, n11460 );
nand U21432 ( n6735, P1_IR_REG_14_, n9828 );
or U21433 ( n9828, n7800, P1_IR_REG_13_ );
nand U21434 ( n10275, SI_30_, n10273 );
nand U21435 ( n5732, n5967, n5968 );
nand U21436 ( n5967, P2_REG2_REG_13_, n11287 );
nand U21437 ( n5968, P2_REG1_REG_13_, n11459 );
xor U21438 ( n2181, P1_REG3_REG_16_, n10621 );
xor U21439 ( n5725, n5726, n5727 );
xnor U21440 ( n5727, n887, P2_REG2_REG_13_ );
nand U21441 ( n1749, n1751, P1_REG2_REG_2_ );
and U21442 ( n1751, n1192, n1219 );
nand U21443 ( n1842, n1843, P1_REG1_REG_2_ );
and U21444 ( n1843, n1192, n1228 );
xnor U21445 ( n6536, P1_IR_REG_17_, n6575 );
nand U21446 ( n1629, n9766, n9767 );
nand U21447 ( n9766, P1_IR_REG_17_, n11485 );
or U21448 ( n9767, n6536, n11484 );
nand U21449 ( n1756, P1_REG2_REG_1_, n1853 );
nand U21450 ( n5743, n5891, n5892 );
nand U21451 ( n5891, P2_REG2_REG_14_, n5869 );
nand U21452 ( n5892, P2_REG1_REG_14_, n11460 );
nand U21453 ( n1848, P1_REG1_REG_1_, n1853 );
nand U21454 ( n2290, n5370, n5371 );
nand U21455 ( n5370, P2_DATAO_REG_11_, n11386 );
nand U21456 ( n5371, n11388, n4284 );
nand U21457 ( n1681, n9779, n9780 );
nand U21458 ( n9779, P1_IR_REG_18_, n11485 );
nand U21459 ( n9780, n9781, P1_IR_REG_31_ );
and U21460 ( n9781, n6438, n6437 );
nand U21461 ( n6437, P1_IR_REG_18_, n9782 );
or U21462 ( n9782, n6575, P1_IR_REG_17_ );
nand U21463 ( n2280, n5374, n5375 );
nand U21464 ( n5375, n11388, n4112 );
nand U21465 ( n5374, P2_DATAO_REG_9_, n11386 );
nand U21466 ( n2300, n5359, n5360 );
nand U21467 ( n5360, n11388, n4078 );
nand U21468 ( n5359, P2_DATAO_REG_13_, n11386 );
nand U21469 ( n2240, n5398, n5399 );
nand U21470 ( n5399, n11388, n4691 );
nand U21471 ( n5398, P2_DATAO_REG_1_, n11386 );
nand U21472 ( n2255, n5384, n5385 );
nand U21473 ( n5385, n11388, n4344 );
nand U21474 ( n5384, P2_DATAO_REG_4_, n11386 );
nand U21475 ( n2235, n5400, n5401 );
nand U21476 ( n5401, n11388, n4693 );
nand U21477 ( n5400, P2_DATAO_REG_0_, n11386 );
nand U21478 ( n2275, n5376, n5377 );
nand U21479 ( n5377, n11388, n4209 );
nand U21480 ( n5376, P2_DATAO_REG_8_, n11386 );
nand U21481 ( n2260, n5382, n5383 );
nand U21482 ( n5383, n11388, n4580 );
nand U21483 ( n5382, P2_DATAO_REG_5_, n11386 );
nand U21484 ( n2270, n5378, n5379 );
nand U21485 ( n5379, n11388, n4211 );
nand U21486 ( n5378, P2_DATAO_REG_7_, n11386 );
nand U21487 ( n2245, n5396, n5397 );
nand U21488 ( n5397, n11388, n4136 );
nand U21489 ( n5396, P2_DATAO_REG_2_, n11386 );
nand U21490 ( n2285, n5372, n5373 );
nand U21491 ( n5373, n11388, n4111 );
nand U21492 ( n5372, P2_DATAO_REG_10_, n11386 );
nand U21493 ( n2295, n5368, n5369 );
nand U21494 ( n5369, n11388, n4490 );
nand U21495 ( n5368, P2_DATAO_REG_12_, n11386 );
nand U21496 ( n2305, n5357, n5358 );
nand U21497 ( n5358, n11388, n4661 );
nand U21498 ( n5357, P2_DATAO_REG_14_, n11386 );
nand U21499 ( n2315, n5353, n5354 );
nand U21500 ( n5354, n11388, n4366 );
nand U21501 ( n5353, P2_DATAO_REG_16_, n11386 );
nand U21502 ( n2320, n5351, n5352 );
nand U21503 ( n5352, n11387, n4558 );
nand U21504 ( n5351, P2_DATAO_REG_17_, n11386 );
nand U21505 ( n2265, n5380, n5381 );
nand U21506 ( n5381, n11388, n4038 );
nand U21507 ( n5380, P2_DATAO_REG_6_, n11386 );
nand U21508 ( n2310, n5355, n5356 );
nand U21509 ( n5356, n11388, n4327 );
nand U21510 ( n5355, P2_DATAO_REG_15_, n11386 );
nand U21511 ( n2325, n5349, n5350 );
nand U21512 ( n5350, n11387, n4153 );
nand U21513 ( n5349, P2_DATAO_REG_18_, n11386 );
nand U21514 ( n2250, n5386, n5387 );
nand U21515 ( n5387, n11388, n4404 );
nand U21516 ( n5386, P2_DATAO_REG_3_, n11386 );
xor U21517 ( n2227, P1_REG3_REG_14_, n10639 );
nand U21518 ( n2345, n5341, n5342 );
nand U21519 ( n5341, P2_DATAO_REG_22_, n11386 );
nand U21520 ( n5342, n11387, n4096 );
nand U21521 ( n2355, n5331, n5332 );
nand U21522 ( n5331, P2_DATAO_REG_24_, n11386 );
nand U21523 ( n5332, n11387, n4305 );
nand U21524 ( n2340, n5343, n5344 );
nand U21525 ( n5343, P2_DATAO_REG_21_, n11386 );
nand U21526 ( n5344, n11387, n4507 );
nand U21527 ( n2335, n5345, n5346 );
nand U21528 ( n5345, P2_DATAO_REG_20_, n5318 );
nand U21529 ( n5346, n11387, n4262 );
nand U21530 ( n2365, n5327, n5328 );
nand U21531 ( n5327, P2_DATAO_REG_26_, n5318 );
nand U21532 ( n5328, n11387, n4056 );
nand U21533 ( n2370, n5325, n5326 );
nand U21534 ( n5325, P2_DATAO_REG_27_, n5318 );
nand U21535 ( n5326, n11387, n4182 );
nand U21536 ( n2360, n5329, n5330 );
nand U21537 ( n5329, P2_DATAO_REG_25_, n5318 );
nand U21538 ( n5330, n11387, n4604 );
nand U21539 ( n2375, n5323, n5324 );
nand U21540 ( n5324, n11387, n4897 );
nand U21541 ( n5323, P2_DATAO_REG_28_, n5318 );
nand U21542 ( n2330, n5347, n5348 );
nand U21543 ( n5347, P2_DATAO_REG_19_, n5318 );
nand U21544 ( n5348, n11387, n4151 );
nand U21545 ( n2380, n5321, n5322 );
nand U21546 ( n5322, n11387, n4884 );
nand U21547 ( n5321, P2_DATAO_REG_29_, n5318 );
nand U21548 ( n2390, n5316, n5317 );
nand U21549 ( n5317, n11388, n4906 );
nand U21550 ( n5316, P2_DATAO_REG_31_, n5318 );
nand U21551 ( n2350, n5333, n5334 );
nand U21552 ( n5334, n11387, n4094 );
nand U21553 ( n5333, P2_DATAO_REG_23_, n5318 );
nand U21554 ( n2385, n5319, n5320 );
nand U21555 ( n5320, n11387, n4877 );
nand U21556 ( n5319, P2_DATAO_REG_30_, n5318 );
xnor U21557 ( ADD_1068_U60, n10865, n10866 );
xnor U21558 ( n10865, P2_ADDR_REG_13_, P1_ADDR_REG_13_ );
nand U21559 ( n10529, P1_REG3_REG_24_, n10538 );
xnor U21560 ( n1654, n51, n1656 );
xnor U21561 ( n1656, n361, P1_REG1_REG_18_ );
xor U21562 ( n1956, P1_REG3_REG_26_, n10520 );
nand U21563 ( n1385, n8496, n8497 );
nand U21564 ( n8497, n11323, P2_IR_REG_10_ );
nor U21565 ( n8496, n8498, n8499 );
nor U21566 ( n8498, n11449, n8503 );
nand U21567 ( n160, n8254, n8255 );
nand U21568 ( n8255, n11409, P1_IR_REG_10_ );
nor U21569 ( n8254, n8256, n8257 );
nor U21570 ( n8256, n11488, n8259 );
xor U21571 ( n1912, P1_REG3_REG_28_, n10486 );
nand U21572 ( n10495, P1_REG3_REG_26_, n10520 );
xor U21573 ( n2137, P1_REG3_REG_18_, n10592 );
xor U21574 ( n2001, P1_REG3_REG_24_, n10538 );
xnor U21575 ( n5705, n5706, n5707 );
xnor U21576 ( n5707, P2_REG2_REG_12_, n5701 );
nand U21577 ( n1375, n8513, n8514 );
nand U21578 ( n8514, n11323, P2_IR_REG_8_ );
nor U21579 ( n8513, n8515, n8516 );
nor U21580 ( n8515, n11449, n8520 );
nand U21581 ( n1380, n8506, n8507 );
nand U21582 ( n8507, n11323, P2_IR_REG_9_ );
nor U21583 ( n8506, n8508, n8509 );
nor U21584 ( n8508, n7791, n11451 );
nand U21585 ( n150, n8270, n8271 );
nand U21586 ( n8271, n11409, P1_IR_REG_8_ );
nor U21587 ( n8270, n8272, n8273 );
nor U21588 ( n8272, n11488, n8275 );
xor U21589 ( ADD_1068_U61, n10863, n10864 );
xor U21590 ( n10864, P2_ADDR_REG_12_, P1_ADDR_REG_12_ );
nand U21591 ( n155, n8261, n8262 );
nand U21592 ( n8262, n11409, P1_IR_REG_9_ );
nor U21593 ( n8261, n8263, n8264 );
nor U21594 ( n8264, n8265, n11489 );
nand U21595 ( n1277, P1_ADDR_REG_4_, n1203 );
not U21596 ( n11532, P2_STATE_REG );
nand U21597 ( n1888, n10486, P1_REG3_REG_28_ );
and U21598 ( n10790, n1203, P1_ADDR_REG_0_ );
or U21599 ( n2702, n11433, P1_B_REG );
not U21600 ( n11537, P1_STATE_REG );
nand U21601 ( n1370, n8523, n8524 );
nand U21602 ( n8524, n11323, P2_IR_REG_7_ );
nor U21603 ( n8523, n8525, n8526 );
nor U21604 ( n8525, n7899, n11451 );
nand U21605 ( n145, n8378, n8379 );
nand U21606 ( n8379, n11409, P1_IR_REG_7_ );
nor U21607 ( n8378, n8380, n8381 );
nor U21608 ( n8381, n8382, n11489 );
nand U21609 ( n1593, n1594, n59 );
xnor U21610 ( n1594, n366, P1_REG2_REG_16_ );
nand U21611 ( n270, n3991, n3992 );
nand U21612 ( n3992, n3987, n3993 );
nand U21613 ( n3991, P1_D_REG_0_, n11502 );
nand U21614 ( n275, n3988, n3989 );
nand U21615 ( n3989, n3987, n3990 );
nand U21616 ( n3988, P1_D_REG_1_, n11502 );
nand U21617 ( n5828, n5969, n5970 );
nand U21618 ( n5969, P2_REG2_REG_17_, n5869 );
nand U21619 ( n5970, P2_REG1_REG_17_, n11459 );
and U21620 ( n280, n11502, P1_D_REG_2_ );
and U21621 ( n290, n11502, P1_D_REG_4_ );
and U21622 ( n300, n11502, P1_D_REG_6_ );
and U21623 ( n315, n11502, P1_D_REG_9_ );
and U21624 ( n325, n11502, P1_D_REG_11_ );
and U21625 ( n335, n11502, P1_D_REG_13_ );
and U21626 ( n345, n11503, P1_D_REG_15_ );
and U21627 ( n355, n11503, P1_D_REG_17_ );
and U21628 ( n365, n11503, P1_D_REG_19_ );
and U21629 ( n375, n11503, P1_D_REG_21_ );
and U21630 ( n390, n11503, P1_D_REG_24_ );
and U21631 ( n400, n11503, P1_D_REG_26_ );
and U21632 ( n285, n11502, P1_D_REG_3_ );
and U21633 ( n295, n11502, P1_D_REG_5_ );
and U21634 ( n310, n11502, P1_D_REG_8_ );
and U21635 ( n320, n11502, P1_D_REG_10_ );
and U21636 ( n330, n11502, P1_D_REG_12_ );
and U21637 ( n6657, n11385, n6699 );
nand U21638 ( n6699, n6037, n11157 );
and U21639 ( n340, n11503, P1_D_REG_14_ );
and U21640 ( n350, n11503, P1_D_REG_16_ );
and U21641 ( n360, n11503, P1_D_REG_18_ );
and U21642 ( n370, n11503, P1_D_REG_20_ );
and U21643 ( n385, n11503, P1_D_REG_23_ );
and U21644 ( n395, n11503, P1_D_REG_25_ );
and U21645 ( n405, n11503, P1_D_REG_27_ );
and U21646 ( n410, n11504, P1_D_REG_28_ );
and U21647 ( n425, n11504, P1_D_REG_31_ );
and U21648 ( n415, n11504, P1_D_REG_29_ );
and U21649 ( n420, n11504, P1_D_REG_30_ );
xnor U21650 ( ADD_1068_U62, n10861, n10862 );
xnor U21651 ( n10861, P2_ADDR_REG_11_, P1_ADDR_REG_11_ );
nand U21652 ( n1538, n1539, n1541 );
nand U21653 ( n1539, n1477, n1479 );
nand U21654 ( n1541, P1_REG1_REG_11_, n1542 );
nand U21655 ( n1542, n54, n387 );
nand U21656 ( n1536, n1534, n1537 );
nand U21657 ( n1537, P1_REG1_REG_12_, n1532 );
nand U21658 ( n1365, n8530, n8531 );
nand U21659 ( n8531, n11323, P2_IR_REG_6_ );
nor U21660 ( n8530, n8532, n8533 );
nor U21661 ( n8532, n11449, n8537 );
nand U21662 ( n140, n8471, n8472 );
nand U21663 ( n8472, n11409, P1_IR_REG_6_ );
nor U21664 ( n8471, n8473, n8474 );
nor U21665 ( n8473, n11489, n8476 );
nand U21666 ( n1518, n1521, n1522 );
nand U21667 ( n1521, n1524, n1479 );
nand U21668 ( n1522, P1_REG2_REG_11_, n1523 );
nand U21669 ( n1523, n61, n387 );
nor U21670 ( n1507, n377, n1516 );
not U21671 ( n377, n1509 );
nand U21672 ( n1516, n1514, n1517 );
nand U21673 ( n1517, P1_REG2_REG_12_, n1512 );
nor U21674 ( n1719, n1722, n1723 );
nor U21675 ( n1723, n382, n11041 );
nor U21676 ( n1722, n1724, n1726 );
nand U21677 ( n1726, P1_REG2_REG_8_, n1442 );
nor U21678 ( n1811, n1813, n1814 );
nor U21679 ( n1814, n382, n11043 );
nor U21680 ( n1813, n1816, n1817 );
nand U21681 ( n1817, P1_REG1_REG_8_, n1442 );
nand U21682 ( n5848, n5971, n5972 );
nand U21683 ( n5971, P2_REG2_REG_18_, n11287 );
nand U21684 ( n5972, P2_REG1_REG_18_, n11459 );
xnor U21685 ( n1577, n1578, n1579 );
xnor U21686 ( n1579, P1_REG1_REG_15_, n1576 );
xor U21687 ( ADD_1068_U63, n10859, n10860 );
xor U21688 ( n10860, P2_ADDR_REG_10_, P1_ADDR_REG_10_ );
nand U21689 ( n4760, n5309, P2_B_REG );
nor U21690 ( n5309, n5310, n5311 );
nor U21691 ( n5311, n5009, n5312 );
nor U21692 ( n5310, n911, n5313 );
nand U21693 ( n1360, n8541, n8542 );
nand U21694 ( n8542, n11323, P2_IR_REG_5_ );
nor U21695 ( n8541, n8543, n8544 );
nor U21696 ( n8544, n7997, n11451 );
nand U21697 ( n135, n8565, n8566 );
nand U21698 ( n8566, n11409, P1_IR_REG_5_ );
nor U21699 ( n8565, n8567, n8568 );
nor U21700 ( n8568, n8569, n11489 );
nand U21701 ( n1355, n8548, n8549 );
nand U21702 ( n8549, n11323, P2_IR_REG_4_ );
nor U21703 ( n8548, n8550, n8551 );
nor U21704 ( n8550, n11449, n8555 );
nand U21705 ( n130, n8664, n8665 );
nand U21706 ( n8665, n11409, P1_IR_REG_4_ );
nor U21707 ( n8664, n8666, n8667 );
nor U21708 ( n8666, n11489, n8669 );
not U21709 ( n1176, SI_30_ );
nand U21710 ( n1500, n8267, n8268 );
nand U21711 ( n8268, n8253, n8242 );
nand U21712 ( n8267, P2_D_REG_1_, n11461 );
nand U21713 ( n1495, n8278, n8279 );
nand U21714 ( n8279, n8253, n8246 );
nand U21715 ( n8278, P2_D_REG_0_, n11461 );
xnor U21716 ( n1493, n53, n1494 );
xnor U21717 ( n1494, n374, P1_REG1_REG_12_ );
and U21718 ( n1505, n11461, P2_D_REG_2_ );
and U21719 ( n1515, n11461, P2_D_REG_4_ );
and U21720 ( n1525, n11461, P2_D_REG_6_ );
and U21721 ( n1540, n11461, P2_D_REG_9_ );
and U21722 ( n1550, n11461, P2_D_REG_11_ );
and U21723 ( n1560, n11461, P2_D_REG_13_ );
and U21724 ( n1570, n11462, P2_D_REG_15_ );
and U21725 ( n1580, n11462, P2_D_REG_17_ );
and U21726 ( n1590, n11462, P2_D_REG_19_ );
and U21727 ( n1600, n11462, P2_D_REG_21_ );
and U21728 ( n1615, n11462, P2_D_REG_24_ );
and U21729 ( n1625, n11462, P2_D_REG_26_ );
and U21730 ( n1510, n11461, P2_D_REG_3_ );
and U21731 ( n1520, n11461, P2_D_REG_5_ );
and U21732 ( n1535, n11461, P2_D_REG_8_ );
and U21733 ( n1545, n11461, P2_D_REG_10_ );
and U21734 ( n1555, n11461, P2_D_REG_12_ );
and U21735 ( n1565, n11462, P2_D_REG_14_ );
and U21736 ( n1575, n11462, P2_D_REG_16_ );
and U21737 ( n1585, n11462, P2_D_REG_18_ );
and U21738 ( n1595, n11462, P2_D_REG_20_ );
and U21739 ( n1610, n11462, P2_D_REG_23_ );
and U21740 ( n1620, n11462, P2_D_REG_25_ );
and U21741 ( n1630, n11462, P2_D_REG_27_ );
xor U21742 ( n5636, n5637, n5638 );
xnor U21743 ( n5638, n878, P2_REG1_REG_9_ );
xor U21744 ( n1557, n1558, n1559 );
xnor U21745 ( n1559, P1_REG1_REG_14_, n369 );
buf U21746 ( n11322, n8312 );
nor U21747 ( n8312, n11282, P2_IR_REG_31_ );
nand U21748 ( n1350, n8558, n8559 );
nand U21749 ( n8559, n11323, P2_IR_REG_3_ );
nor U21750 ( n8558, n8560, n8561 );
and U21751 ( n8560, n11530, n8064 );
and U21752 ( n1635, n11463, P2_D_REG_28_ );
and U21753 ( n1650, n11463, P2_D_REG_31_ );
and U21754 ( n1640, n11463, P2_D_REG_29_ );
and U21755 ( n1645, n11463, P2_D_REG_30_ );
nand U21756 ( n1457, n1458, n1459 );
nand U21757 ( n1458, n1462, n1442 );
nand U21758 ( n1459, P1_REG1_REG_8_, n1461 );
nand U21759 ( n1461, n56, n389 );
nand U21760 ( n1454, n1453, n1456 );
nand U21761 ( n1456, P1_REG1_REG_9_, n1451 );
nand U21762 ( n1345, n8571, n8572 );
nand U21763 ( n8572, n11323, P2_IR_REG_2_ );
nor U21764 ( n8571, n8573, n8574 );
and U21765 ( n8574, n11530, n8101 );
nand U21766 ( n120, n9044, n9045 );
nand U21767 ( n9045, n11409, P1_IR_REG_2_ );
nor U21768 ( n9044, n9046, n9047 );
nor U21769 ( n9046, n11488, n9049 );
nor U21770 ( n1423, n384, n1432 );
not U21771 ( n384, n1426 );
nand U21772 ( n1432, n1431, n1433 );
nand U21773 ( n1433, P1_REG2_REG_9_, n1428 );
nand U21774 ( n1434, n1437, n1438 );
nand U21775 ( n1437, n1441, n1442 );
nand U21776 ( n1438, P1_REG2_REG_8_, n1439 );
nand U21777 ( n1439, n63, n389 );
nor U21778 ( n1702, n1706, n1707 );
nor U21779 ( n1707, n374, n11049 );
nor U21780 ( n1706, n1708, n1709 );
nand U21781 ( n1709, P1_REG2_REG_11_, n1479 );
nor U21782 ( n1794, n1797, n1798 );
nor U21783 ( n1798, n374, n11051 );
nor U21784 ( n1797, n1799, n1801 );
nand U21785 ( n1801, P1_REG1_REG_11_, n1479 );
xnor U21786 ( ADD_1068_U47, n10892, n10893 );
xnor U21787 ( n10892, P2_ADDR_REG_9_, P1_ADDR_REG_9_ );
buf U21788 ( n11407, n4002 );
nor U21789 ( n4002, n11534, P1_IR_REG_31_ );
nand U21790 ( n1721, P1_REG2_REG_9_, n1436 );
nand U21791 ( n1812, P1_REG1_REG_9_, n1436 );
nand U21792 ( n9562, P1_B_REG, n10451 );
nand U21793 ( n10451, n10452, n10453 );
nand U21794 ( n10453, n10454, n10455 );
nor U21795 ( n10452, n11534, n9375 );
nand U21796 ( n125, n8878, n8879 );
nand U21797 ( n8879, n11409, P1_IR_REG_3_ );
nor U21798 ( n8878, n8880, n8881 );
nor U21799 ( n8881, n8882, n11490 );
xor U21800 ( n5616, n5617, n5618 );
xnor U21801 ( n5618, n876, P2_REG1_REG_8_ );
xnor U21802 ( n1409, n55, n1411 );
xnor U21803 ( n1411, n388, P1_REG1_REG_9_ );
xor U21804 ( ADD_1068_U48, n10890, n10891 );
xor U21805 ( n10891, P2_ADDR_REG_8_, P1_ADDR_REG_8_ );
xnor U21806 ( n1476, n1477, n1478 );
xnor U21807 ( n1478, P1_REG1_REG_11_, n1479 );
nand U21808 ( n1340, n8581, n8582 );
nand U21809 ( n8582, n11323, P2_IR_REG_1_ );
nor U21810 ( n8581, n8583, n8584 );
and U21811 ( n8584, n8130, n8304 );
nand U21812 ( n115, n10498, n10499 );
nand U21813 ( n10499, n11408, P1_IR_REG_1_ );
nor U21814 ( n10498, n10500, n10501 );
and U21815 ( n10501, n10502, n3997 );
nor U21816 ( n1243, P1_IR_REG_0_, n1244 );
nor U21817 ( n1244, n1246, n284 );
nor U21818 ( n1246, P1_REG2_REG_0_, n282 );
nand U21819 ( n9411, n9412, n9413 );
nor U21820 ( n9412, P1_D_REG_4_, P1_D_REG_3_ );
nor U21821 ( n9413, P1_D_REG_6_, P1_D_REG_5_ );
nor U21822 ( n9416, P1_D_REG_17_, P1_D_REG_16_ );
nand U21823 ( n9428, n9429, n9430 );
nor U21824 ( n9429, P1_D_REG_26_, P1_D_REG_25_ );
nor U21825 ( n9430, P1_D_REG_28_, P1_D_REG_27_ );
nor U21826 ( n9433, P1_D_REG_13_, P1_D_REG_12_ );
nor U21827 ( n9415, P1_D_REG_15_, P1_D_REG_14_ );
nand U21828 ( n9419, n9420, n9421 );
nor U21829 ( n9420, P1_D_REG_2_, P1_D_REG_29_ );
nor U21830 ( n9421, P1_D_REG_31_, P1_D_REG_30_ );
nor U21831 ( n9432, P1_D_REG_11_, P1_D_REG_10_ );
nor U21832 ( n9423, P1_D_REG_9_, P1_D_REG_8_ );
xor U21833 ( n5591, n5592, n5593 );
xnor U21834 ( n5593, n874, P2_REG1_REG_7_ );
nand U21835 ( n1703, P1_REG2_REG_13_, n1704 );
nand U21836 ( n1796, P1_REG1_REG_13_, n1704 );
xnor U21837 ( n1394, n56, n1396 );
xnor U21838 ( n1396, n389, P1_REG1_REG_8_ );
xnor U21839 ( ADD_1068_U49, n10888, n10889 );
xnor U21840 ( n10888, P2_ADDR_REG_7_, P1_ADDR_REG_7_ );
nand U21841 ( n8210, n8211, n8212 );
nor U21842 ( n8211, P2_D_REG_4_, P2_D_REG_3_ );
nor U21843 ( n8212, P2_D_REG_6_, P2_D_REG_5_ );
nand U21844 ( n8227, n8228, n8229 );
nor U21845 ( n8228, P2_D_REG_26_, P2_D_REG_25_ );
nor U21846 ( n8229, P2_D_REG_28_, P2_D_REG_27_ );
nor U21847 ( n8215, P2_D_REG_17_, P2_D_REG_16_ );
nor U21848 ( n8232, P2_D_REG_13_, P2_D_REG_12_ );
nor U21849 ( n8214, P2_D_REG_15_, P2_D_REG_14_ );
nand U21850 ( n8218, n8219, n8220 );
nor U21851 ( n8219, P2_D_REG_2_, P2_D_REG_29_ );
nor U21852 ( n8220, P2_D_REG_31_, P2_D_REG_30_ );
nor U21853 ( n8231, P2_D_REG_11_, P2_D_REG_10_ );
nor U21854 ( n8222, P2_D_REG_9_, P2_D_REG_8_ );
nand U21855 ( n110, n10604, n10605 );
nand U21856 ( n10605, P1_IR_REG_0_, n10606 );
nand U21857 ( n10604, n9955, n11534 );
or U21858 ( n10606, n11408, n3997 );
nand U21859 ( n1335, n8588, n8589 );
nand U21860 ( n8589, P2_IR_REG_0_, n8590 );
nand U21861 ( n8588, n8156, n11282 );
or U21862 ( n8590, n11323, n8304 );
xor U21863 ( ADD_1068_U50, n10884, n10885 );
xor U21864 ( n10885, P2_ADDR_REG_6_, P1_ADDR_REG_6_ );
nand U21865 ( n1333, n1334, n64 );
xnor U21866 ( n1334, P1_REG2_REG_6_, n393 );
xor U21867 ( n5535, n5536, n5537 );
xnor U21868 ( n5537, n871, P2_REG1_REG_5_ );
nand U21869 ( n1226, n1318, n1319 );
nand U21870 ( n1318, n1196, n1192 );
nand U21871 ( n1319, P1_REG1_REG_2_, n1320 );
or U21872 ( n1320, n1196, n1192 );
nand U21873 ( n1217, n1299, n1301 );
nand U21874 ( n1299, n1189, n1192 );
nand U21875 ( n1301, P1_REG2_REG_2_, n1302 );
or U21876 ( n1302, n1189, n1192 );
xnor U21877 ( ADD_1068_U51, n10882, n10883 );
xnor U21878 ( n10882, P2_ADDR_REG_5_, P1_ADDR_REG_5_ );
xnor U21879 ( n5870, n907, P2_REG1_REG_19_ );
xnor U21880 ( n5509, n5510, n5511 );
xnor U21881 ( n5511, P2_REG1_REG_4_, n5508 );
nand U21882 ( n1258, n1259, n67 );
xnor U21883 ( n1259, n403, P1_REG2_REG_4_ );
xor U21884 ( ADD_1068_U52, n10880, n10881 );
xor U21885 ( n10881, P2_ADDR_REG_4_, P1_ADDR_REG_4_ );
or U21886 ( n1214, n11257, n1217 );
xor U21887 ( n11257, n407, P1_REG2_REG_3_ );
xnor U21888 ( n1653, n361, P1_REG2_REG_18_ );
xor U21889 ( n5490, n5491, n5492 );
xnor U21890 ( n5492, n864, P2_REG1_REG_3_ );
xnor U21891 ( n5839, P2_REG1_REG_18_, n897 );
xnor U21892 ( ADD_1068_U53, n10878, n10879 );
xnor U21893 ( n10878, P2_ADDR_REG_3_, P1_ADDR_REG_3_ );
xnor U21894 ( n1603, n366, P1_REG1_REG_16_ );
nor U21895 ( n1658, n11533, n11158 );
nor U21896 ( n1609, n11533, n11159 );
nor U21897 ( n1563, P1_STATE_REG, n11160 );
nor U21898 ( n1497, P1_STATE_REG, n11161 );
nor U21899 ( n1464, P1_STATE_REG, n11162 );
nor U21900 ( n1398, P1_STATE_REG, n11163 );
nor U21901 ( n1349, n11533, n11164 );
nor U21902 ( n4040, n11527, n11166 );
nor U21903 ( n4212, n11527, n11167 );
nor U21904 ( n4421, n11527, n11168 );
nor U21905 ( n4113, n11527, n11169 );
nor U21906 ( n4527, n11527, n11170 );
nor U21907 ( n4285, n11527, n11171 );
nor U21908 ( n4491, n11527, n11172 );
nor U21909 ( n4079, n11527, n11173 );
nor U21910 ( n4581, n11527, n11174 );
nor U21911 ( n4154, n11527, n11175 );
nor U21912 ( n4559, n11527, n11176 );
nor U21913 ( n4345, n11527, n11177 );
nor U21914 ( n4367, n11527, n11178 );
nor U21915 ( n4328, n11527, n11179 );
nor U21916 ( n1274, n11533, n11165 );
nor U21917 ( n4717, n11527, n11180 );
xnor U21918 ( n5820, P2_REG1_REG_17_, n5817 );
xnor U21919 ( n1556, P1_REG2_REG_14_, n369 );
xnor U21920 ( n1474, n387, P1_REG2_REG_11_ );
xnor U21921 ( n1408, n388, P1_REG2_REG_9_ );
xnor U21922 ( n1393, n389, P1_REG2_REG_8_ );
xnor U21923 ( n1426, P1_REG2_REG_10_, n1443 );
xnor U21924 ( n1448, P1_REG1_REG_10_, n1443 );
xnor U21925 ( n1492, n374, P1_REG2_REG_12_ );
xnor U21926 ( n5464, n5465, n5466 );
xnor U21927 ( n5466, P2_REG1_REG_2_, n5459 );
xnor U21928 ( n1224, n407, P1_REG1_REG_3_ );
xnor U21929 ( n5567, P2_REG2_REG_6_, n872 );
xnor U21930 ( n5516, n867, P2_REG2_REG_4_ );
xnor U21931 ( n5623, n876, P2_REG2_REG_8_ );
xnor U21932 ( n1343, P1_REG1_REG_6_, n393 );
xnor U21933 ( n5472, n862, P2_REG2_REG_2_ );
xnor U21934 ( n5644, P2_REG2_REG_9_, n5635 );
xnor U21935 ( n5724, P2_REG1_REG_13_, n5721 );
xnor U21936 ( n5543, P2_REG2_REG_5_, n5533 );
xnor U21937 ( n5498, P2_REG2_REG_3_, n5488 );
xnor U21938 ( n5599, P2_REG2_REG_7_, n5586 );
xnor U21939 ( n5703, n886, P2_REG1_REG_12_ );
xor U21940 ( n10900, P1_ADDR_REG_19_, P2_ADDR_REG_19_ );
xor U21941 ( n10804, n10805, n10806 );
nand U21942 ( n10806, P1_REG1_REG_0_, P1_IR_REG_0_ );
nand U21943 ( n10805, n1848, n10807 );
nand U21944 ( n10807, n409, n10973 );
xnor U21945 ( n1272, P1_REG1_REG_4_, n1273 );
xor U21946 ( ADD_1068_U54, n10876, n10877 );
xor U21947 ( n10877, P2_ADDR_REG_2_, P1_ADDR_REG_2_ );
xnor U21948 ( ADD_1068_U5, n10886, n10887 );
xnor U21949 ( n10887, P2_ADDR_REG_1_, n10962 );
xor U21950 ( ADD_1068_U46, P2_ADDR_REG_0_, P1_ADDR_REG_0_ );
xnor U21951 ( U126, P1_RD_REG, P2_RD_REG );
xnor U21952 ( U123, P2_WR_REG, P1_WR_REG );
xnor U21953 ( n5435, n861, P2_REG2_REG_1_ );
xnor U21954 ( n5434, n859, P2_REG1_REG_1_ );
endmodule

