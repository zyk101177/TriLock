
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule

module aes128_ori ( clk, reset, start, state, key, out, out_valid );
input [127:0] state;
input [127:0] key;
output [127:0] out;
input clk, reset, start;
output out_valid;
wire N135, N136, N137, N138, n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, ex_wire30, ex_wire31, ex_wire32, ex_wire33, ex_wire34, ex_wire35, ex_wire36, ex_wire37, ex_wire38, ex_wire39, ex_wire40, ex_wire41, ex_wire42, ex_wire43, ex_wire44, ex_wire45, ex_wire46, ex_wire47, ex_wire48, ex_wire49, ex_wire50, ex_wire51, ex_wire52, ex_wire53, ex_wire54, ex_wire55, ex_wire56, ex_wire57, ex_wire58, ex_wire59, ex_wire60, ex_wire61, ex_wire62, ex_wire63, ex_wire64, ex_wire65, ex_wire66, ex_wire67, ex_wire68, ex_wire69, ex_wire70, ex_wire71, ex_wire72, ex_wire73, ex_wire74, ex_wire75, ex_wire76, ex_wire77, ex_wire78, ex_wire79, ex_wire80, ex_wire81, ex_wire82, ex_wire83, ex_wire84, ex_wire85, ex_wire86, ex_wire87, ex_wire88, ex_wire89, ex_wire90, ex_wire91, ex_wire92, ex_wire93, ex_wire94, ex_wire95, ex_wire96, ex_wire97, ex_wire98, ex_wire99, ex_wire100, ex_wire101, ex_wire102, ex_wire103, ex_wire104, ex_wire105, ex_wire106, ex_wire107, ex_wire108, ex_wire109, ex_wire110, ex_wire111, ex_wire112, ex_wire113, ex_wire114, ex_wire115, ex_wire116, n12,
n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
s9_9_, s9_99_, s9_98_, s9_97_, s9_96_, s9_95_, s9_94_, s9_93_, s9_92_,
s9_91_, s9_90_, s9_8_, s9_89_, s9_88_, s9_87_, s9_86_, s9_85_, s9_84_,
s9_83_, s9_82_, s9_81_, s9_80_, s9_7_, s9_79_, s9_78_, s9_77_, s9_76_,
s9_75_, s9_74_, s9_73_, s9_72_, s9_71_, s9_70_, s9_6_, s9_69_, s9_68_,
s9_67_, s9_66_, s9_65_, s9_64_, s9_63_, s9_62_, s9_61_, s9_60_, s9_5_,
s9_59_, s9_58_, s9_57_, s9_56_, s9_55_, s9_54_, s9_53_, s9_52_,
s9_51_, s9_50_, s9_4_, s9_49_, s9_48_, s9_47_, s9_46_, s9_45_, s9_44_,
s9_43_, s9_42_, s9_41_, s9_40_, s9_3_, s9_39_, s9_38_, s9_37_, s9_36_,
s9_35_, s9_34_, s9_33_, s9_32_, s9_31_, s9_30_, s9_2_, s9_29_, s9_28_,
s9_27_, s9_26_, s9_25_, s9_24_, s9_23_, s9_22_, s9_21_, s9_20_, s9_1_,
s9_19_, s9_18_, s9_17_, s9_16_, s9_15_, s9_14_, s9_13_, s9_12_,
s9_127_, s9_126_, s9_125_, s9_124_, s9_123_, s9_122_, s9_121_,
s9_120_, s9_11_, s9_119_, s9_118_, s9_117_, s9_116_, s9_115_, s9_114_,
s9_113_, s9_112_, s9_111_, s9_110_, s9_10_, s9_109_, s9_108_, s9_107_,
s9_106_, s9_105_, s9_104_, s9_103_, s9_102_, s9_101_, s9_100_, s9_0_,
s8_9_, s8_99_, s8_98_, s8_97_, s8_96_, s8_95_, s8_94_, s8_93_, s8_92_,
s8_91_, s8_90_, s8_8_, s8_89_, s8_88_, s8_87_, s8_86_, s8_85_, s8_84_,
s8_83_, s8_82_, s8_81_, s8_80_, s8_7_, s8_79_, s8_78_, s8_77_, s8_76_,
s8_75_, s8_74_, s8_73_, s8_72_, s8_71_, s8_70_, s8_6_, s8_69_, s8_68_,
s8_67_, s8_66_, s8_65_, s8_64_, s8_63_, s8_62_, s8_61_, s8_60_, s8_5_,
s8_59_, s8_58_, s8_57_, s8_56_, s8_55_, s8_54_, s8_53_, s8_52_,
s8_51_, s8_50_, s8_4_, s8_49_, s8_48_, s8_47_, s8_46_, s8_45_, s8_44_,
s8_43_, s8_42_, s8_41_, s8_40_, s8_3_, s8_39_, s8_38_, s8_37_, s8_36_,
s8_35_, s8_34_, s8_33_, s8_32_, s8_31_, s8_30_, s8_2_, s8_29_, s8_28_,
s8_27_, s8_26_, s8_25_, s8_24_, s8_23_, s8_22_, s8_21_, s8_20_, s8_1_,
s8_19_, s8_18_, s8_17_, s8_16_, s8_15_, s8_14_, s8_13_, s8_12_,
s8_127_, s8_126_, s8_125_, s8_124_, s8_123_, s8_122_, s8_121_,
s8_120_, s8_11_, s8_119_, s8_118_, s8_117_, s8_116_, s8_115_, s8_114_,
s8_113_, s8_112_, s8_111_, s8_110_, s8_10_, s8_109_, s8_108_, s8_107_,
s8_106_, s8_105_, s8_104_, s8_103_, s8_102_, s8_101_, s8_100_, s8_0_,
s7_9_, s7_99_, s7_98_, s7_97_, s7_96_, s7_95_, s7_94_, s7_93_, s7_92_,
s7_91_, s7_90_, s7_8_, s7_89_, s7_88_, s7_87_, s7_86_, s7_85_, s7_84_,
s7_83_, s7_82_, s7_81_, s7_80_, s7_7_, s7_79_, s7_78_, s7_77_, s7_76_,
s7_75_, s7_74_, s7_73_, s7_72_, s7_71_, s7_70_, s7_6_, s7_69_, s7_68_,
s7_67_, s7_66_, s7_65_, s7_64_, s7_63_, s7_62_, s7_61_, s7_60_, s7_5_,
s7_59_, s7_58_, s7_57_, s7_56_, s7_55_, s7_54_, s7_53_, s7_52_,
s7_51_, s7_50_, s7_4_, s7_49_, s7_48_, s7_47_, s7_46_, s7_45_, s7_44_,
s7_43_, s7_42_, s7_41_, s7_40_, s7_3_, s7_39_, s7_38_, s7_37_, s7_36_,
s7_35_, s7_34_, s7_33_, s7_32_, s7_31_, s7_30_, s7_2_, s7_29_, s7_28_,
s7_27_, s7_26_, s7_25_, s7_24_, s7_23_, s7_22_, s7_21_, s7_20_, s7_1_,
s7_19_, s7_18_, s7_17_, s7_16_, s7_15_, s7_14_, s7_13_, s7_12_,
s7_127_, s7_126_, s7_125_, s7_124_, s7_123_, s7_122_, s7_121_,
s7_120_, s7_11_, s7_119_, s7_118_, s7_117_, s7_116_, s7_115_, s7_114_,
s7_113_, s7_112_, s7_111_, s7_110_, s7_10_, s7_109_, s7_108_, s7_107_,
s7_106_, s7_105_, s7_104_, s7_103_, s7_102_, s7_101_, s7_100_, s7_0_,
s6_9_, s6_99_, s6_98_, s6_97_, s6_96_, s6_95_, s6_94_, s6_93_, s6_92_,
s6_91_, s6_90_, s6_8_, s6_89_, s6_88_, s6_87_, s6_86_, s6_85_, s6_84_,
s6_83_, s6_82_, s6_81_, s6_80_, s6_7_, s6_79_, s6_78_, s6_77_, s6_76_,
s6_75_, s6_74_, s6_73_, s6_72_, s6_71_, s6_70_, s6_6_, s6_69_, s6_68_,
s6_67_, s6_66_, s6_65_, s6_64_, s6_63_, s6_62_, s6_61_, s6_60_, s6_5_,
s6_59_, s6_58_, s6_57_, s6_56_, s6_55_, s6_54_, s6_53_, s6_52_,
s6_51_, s6_50_, s6_4_, s6_49_, s6_48_, s6_47_, s6_46_, s6_45_, s6_44_,
s6_43_, s6_42_, s6_41_, s6_40_, s6_3_, s6_39_, s6_38_, s6_37_, s6_36_,
s6_35_, s6_34_, s6_33_, s6_32_, s6_31_, s6_30_, s6_2_, s6_29_, s6_28_,
s6_27_, s6_26_, s6_25_, s6_24_, s6_23_, s6_22_, s6_21_, s6_20_, s6_1_,
s6_19_, s6_18_, s6_17_, s6_16_, s6_15_, s6_14_, s6_13_, s6_12_,
s6_127_, s6_126_, s6_125_, s6_124_, s6_123_, s6_122_, s6_121_,
s6_120_, s6_11_, s6_119_, s6_118_, s6_117_, s6_116_, s6_115_, s6_114_,
s6_113_, s6_112_, s6_111_, s6_110_, s6_10_, s6_109_, s6_108_, s6_107_,
s6_106_, s6_105_, s6_104_, s6_103_, s6_102_, s6_101_, s6_100_, s6_0_,
s5_9_, s5_99_, s5_98_, s5_97_, s5_96_, s5_95_, s5_94_, s5_93_, s5_92_,
s5_91_, s5_90_, s5_8_, s5_89_, s5_88_, s5_87_, s5_86_, s5_85_, s5_84_,
s5_83_, s5_82_, s5_81_, s5_80_, s5_7_, s5_79_, s5_78_, s5_77_, s5_76_,
s5_75_, s5_74_, s5_73_, s5_72_, s5_71_, s5_70_, s5_6_, s5_69_, s5_68_,
s5_67_, s5_66_, s5_65_, s5_64_, s5_63_, s5_62_, s5_61_, s5_60_, s5_5_,
s5_59_, s5_58_, s5_57_, s5_56_, s5_55_, s5_54_, s5_53_, s5_52_,
s5_51_, s5_50_, s5_4_, s5_49_, s5_48_, s5_47_, s5_46_, s5_45_, s5_44_,
s5_43_, s5_42_, s5_41_, s5_40_, s5_3_, s5_39_, s5_38_, s5_37_, s5_36_,
s5_35_, s5_34_, s5_33_, s5_32_, s5_31_, s5_30_, s5_2_, s5_29_, s5_28_,
s5_27_, s5_26_, s5_25_, s5_24_, s5_23_, s5_22_, s5_21_, s5_20_, s5_1_,
s5_19_, s5_18_, s5_17_, s5_16_, s5_15_, s5_14_, s5_13_, s5_12_,
s5_127_, s5_126_, s5_125_, s5_124_, s5_123_, s5_122_, s5_121_,
s5_120_, s5_11_, s5_119_, s5_118_, s5_117_, s5_116_, s5_115_, s5_114_,
s5_113_, s5_112_, s5_111_, s5_110_, s5_10_, s5_109_, s5_108_, s5_107_,
s5_106_, s5_105_, s5_104_, s5_103_, s5_102_, s5_101_, s5_100_, s5_0_,
s4_9_, s4_99_, s4_98_, s4_97_, s4_96_, s4_95_, s4_94_, s4_93_, s4_92_,
s4_91_, s4_90_, s4_8_, s4_89_, s4_88_, s4_87_, s4_86_, s4_85_, s4_84_,
s4_83_, s4_82_, s4_81_, s4_80_, s4_7_, s4_79_, s4_78_, s4_77_, s4_76_,
s4_75_, s4_74_, s4_73_, s4_72_, s4_71_, s4_70_, s4_6_, s4_69_, s4_68_,
s4_67_, s4_66_, s4_65_, s4_64_, s4_63_, s4_62_, s4_61_, s4_60_, s4_5_,
s4_59_, s4_58_, s4_57_, s4_56_, s4_55_, s4_54_, s4_53_, s4_52_,
s4_51_, s4_50_, s4_4_, s4_49_, s4_48_, s4_47_, s4_46_, s4_45_, s4_44_,
s4_43_, s4_42_, s4_41_, s4_40_, s4_3_, s4_39_, s4_38_, s4_37_, s4_36_,
s4_35_, s4_34_, s4_33_, s4_32_, s4_31_, s4_30_, s4_2_, s4_29_, s4_28_,
s4_27_, s4_26_, s4_25_, s4_24_, s4_23_, s4_22_, s4_21_, s4_20_, s4_1_,
s4_19_, s4_18_, s4_17_, s4_16_, s4_15_, s4_14_, s4_13_, s4_12_,
s4_127_, s4_126_, s4_125_, s4_124_, s4_123_, s4_122_, s4_121_,
s4_120_, s4_11_, s4_119_, s4_118_, s4_117_, s4_116_, s4_115_, s4_114_,
s4_113_, s4_112_, s4_111_, s4_110_, s4_10_, s4_109_, s4_108_, s4_107_,
s4_106_, s4_105_, s4_104_, s4_103_, s4_102_, s4_101_, s4_100_, s4_0_,
s3_9_, s3_99_, s3_98_, s3_97_, s3_96_, s3_95_, s3_94_, s3_93_, s3_92_,
s3_91_, s3_90_, s3_8_, s3_89_, s3_88_, s3_87_, s3_86_, s3_85_, s3_84_,
s3_83_, s3_82_, s3_81_, s3_80_, s3_7_, s3_79_, s3_78_, s3_77_, s3_76_,
s3_75_, s3_74_, s3_73_, s3_72_, s3_71_, s3_70_, s3_6_, s3_69_, s3_68_,
s3_67_, s3_66_, s3_65_, s3_64_, s3_63_, s3_62_, s3_61_, s3_60_, s3_5_,
s3_59_, s3_58_, s3_57_, s3_56_, s3_55_, s3_54_, s3_53_, s3_52_,
s3_51_, s3_50_, s3_4_, s3_49_, s3_48_, s3_47_, s3_46_, s3_45_, s3_44_,
s3_43_, s3_42_, s3_41_, s3_40_, s3_3_, s3_39_, s3_38_, s3_37_, s3_36_,
s3_35_, s3_34_, s3_33_, s3_32_, s3_31_, s3_30_, s3_2_, s3_29_, s3_28_,
s3_27_, s3_26_, s3_25_, s3_24_, s3_23_, s3_22_, s3_21_, s3_20_, s3_1_,
s3_19_, s3_18_, s3_17_, s3_16_, s3_15_, s3_14_, s3_13_, s3_12_,
s3_127_, s3_126_, s3_125_, s3_124_, s3_123_, s3_122_, s3_121_,
s3_120_, s3_11_, s3_119_, s3_118_, s3_117_, s3_116_, s3_115_, s3_114_,
s3_113_, s3_112_, s3_111_, s3_110_, s3_10_, s3_109_, s3_108_, s3_107_,
s3_106_, s3_105_, s3_104_, s3_103_, s3_102_, s3_101_, s3_100_, s3_0_,
s2_9_, s2_99_, s2_98_, s2_97_, s2_96_, s2_95_, s2_94_, s2_93_, s2_92_,
s2_91_, s2_90_, s2_8_, s2_89_, s2_88_, s2_87_, s2_86_, s2_85_, s2_84_,
s2_83_, s2_82_, s2_81_, s2_80_, s2_7_, s2_79_, s2_78_, s2_77_, s2_76_,
s2_75_, s2_74_, s2_73_, s2_72_, s2_71_, s2_70_, s2_6_, s2_69_, s2_68_,
s2_67_, s2_66_, s2_65_, s2_64_, s2_63_, s2_62_, s2_61_, s2_60_, s2_5_,
s2_59_, s2_58_, s2_57_, s2_56_, s2_55_, s2_54_, s2_53_, s2_52_,
s2_51_, s2_50_, s2_4_, s2_49_, s2_48_, s2_47_, s2_46_, s2_45_, s2_44_,
s2_43_, s2_42_, s2_41_, s2_40_, s2_3_, s2_39_, s2_38_, s2_37_, s2_36_,
s2_35_, s2_34_, s2_33_, s2_32_, s2_31_, s2_30_, s2_2_, s2_29_, s2_28_,
s2_27_, s2_26_, s2_25_, s2_24_, s2_23_, s2_22_, s2_21_, s2_20_, s2_1_,
s2_19_, s2_18_, s2_17_, s2_16_, s2_15_, s2_14_, s2_13_, s2_12_,
s2_127_, s2_126_, s2_125_, s2_124_, s2_123_, s2_122_, s2_121_,
s2_120_, s2_11_, s2_119_, s2_118_, s2_117_, s2_116_, s2_115_, s2_114_,
s2_113_, s2_112_, s2_111_, s2_110_, s2_10_, s2_109_, s2_108_, s2_107_,
s2_106_, s2_105_, s2_104_, s2_103_, s2_102_, s2_101_, s2_100_, s2_0_,
s1_9_, s1_99_, s1_98_, s1_97_, s1_96_, s1_95_, s1_94_, s1_93_, s1_92_,
s1_91_, s1_90_, s1_8_, s1_89_, s1_88_, s1_87_, s1_86_, s1_85_, s1_84_,
s1_83_, s1_82_, s1_81_, s1_80_, s1_7_, s1_79_, s1_78_, s1_77_, s1_76_,
s1_75_, s1_74_, s1_73_, s1_72_, s1_71_, s1_70_, s1_6_, s1_69_, s1_68_,
s1_67_, s1_66_, s1_65_, s1_64_, s1_63_, s1_62_, s1_61_, s1_60_, s1_5_,
s1_59_, s1_58_, s1_57_, s1_56_, s1_55_, s1_54_, s1_53_, s1_52_,
s1_51_, s1_50_, s1_4_, s1_49_, s1_48_, s1_47_, s1_46_, s1_45_, s1_44_,
s1_43_, s1_42_, s1_41_, s1_40_, s1_3_, s1_39_, s1_38_, s1_37_, s1_36_,
s1_35_, s1_34_, s1_33_, s1_32_, s1_31_, s1_30_, s1_2_, s1_29_, s1_28_,
s1_27_, s1_26_, s1_25_, s1_24_, s1_23_, s1_22_, s1_21_, s1_20_, s1_1_,
s1_19_, s1_18_, s1_17_, s1_16_, s1_15_, s1_14_, s1_13_, s1_12_,
s1_127_, s1_126_, s1_125_, s1_124_, s1_123_, s1_122_, s1_121_,
s1_120_, s1_11_, s1_119_, s1_118_, s1_117_, s1_116_, s1_115_, s1_114_,
s1_113_, s1_112_, s1_111_, s1_110_, s1_10_, s1_109_, s1_108_, s1_107_,
s1_106_, s1_105_, s1_104_, s1_103_, s1_102_, s1_101_, s1_100_, s1_0_,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1589, n1590, n1591,
n1592, n1593;
wire [127:0] s0;
wire [127:0] k0;
wire [4:0] validCounter;
wire [127:0] k1;
wire [127:0] k0b;
wire [127:0] k2;
wire [127:0] k1b;
wire [127:0] k3;
wire [127:0] k2b;
wire [127:0] k4;
wire [127:0] k3b;
wire [127:0] k5;
wire [127:0] k4b;
wire [127:0] k6;
wire [127:0] k5b;
wire [126:0] k7;
wire [127:0] k6b;
wire [127:0] k8;
wire [127:0] k7b;
wire [127:0] k9;
wire [127:0] k8b;
wire [127:0] k9b;
wire [31:0] a1_k4a;
wire [31:0] a1_k3a;
wire [31:0] a1_k2a;
wire [31:0] a1_k1a;
wire [31:0] a1_k0a;
wire [31:0] a1_v3;
wire [31:0] a1_v2;
wire [31:0] a1_v1;
wire [31:0] a2_k4a;
wire [31:0] a2_k3a;
wire [31:0] a2_k2a;
wire [31:0] a2_k1a;
wire [31:0] a2_k0a;
wire [31:0] a2_v3;
wire [31:0] a2_v2;
wire [31:0] a2_v1;
wire [31:0] a3_k4a;
wire [31:0] a3_k3a;
wire [31:0] a3_k2a;
wire [31:0] a3_k1a;
wire [31:0] a3_k0a;
wire [31:0] a3_v3;
wire [31:0] a3_v2;
wire [31:0] a3_v1;
wire [31:0] a4_k4a;
wire [31:0] a4_k3a;
wire [31:0] a4_k2a;
wire [31:0] a4_k1a;
wire [31:0] a4_k0a;
wire [31:0] a4_v3;
wire [31:0] a4_v2;
wire [31:0] a4_v1;
wire [31:0] a5_k4a;
wire [31:0] a5_k3a;
wire [31:0] a5_k2a;
wire [31:0] a5_k1a;
wire [31:0] a5_k0a;
wire [31:0] a5_v3;
wire [31:0] a5_v2;
wire [31:0] a5_v1;
wire [31:0] a6_k4a;
wire [31:0] a6_k3a;
wire [31:0] a6_k2a;
wire [31:0] a6_k1a;
wire [31:0] a6_k0a;
wire [31:0] a6_v3;
wire [31:0] a6_v2;
wire [31:0] a6_v1;
wire [31:0] a7_k4a;
wire [31:0] a7_k3a;
wire [31:0] a7_k2a;
wire [31:0] a7_k1a;
wire [31:0] a7_k0a;
wire [31:0] a7_v3;
wire [31:0] a7_v2;
wire [31:0] a7_v1;
wire [31:0] a8_k4a;
wire [31:0] a8_k3a;
wire [31:0] a8_k2a;
wire [31:0] a8_k1a;
wire [31:0] a8_k0a;
wire [31:0] a8_v3;
wire [31:0] a8_v2;
wire [31:0] a8_v1;
wire [31:0] a9_k4a;
wire [31:0] a9_k3a;
wire [31:0] a9_k2a;
wire [31:0] a9_k1a;
wire [31:0] a9_k0a;
wire [31:0] a9_v3;
wire [31:0] a9_v2;
wire [31:0] a9_v1;
wire [31:0] a10_k4a;
wire [31:0] a10_k3a;
wire [31:0] a10_k2a;
wire [31:0] a10_k1a;
wire [31:0] a10_k0a;
wire [31:0] a10_v3;
wire [31:0] a10_v2;
wire [31:0] a10_v1;

dff a10_k1a_reg_31_ ( clk, n1527_r, a10_k1a[31], a10_v1[31] );
not U_inv0 ( n1527_r, n1527 );
dff a9_k1a_reg_31_ ( clk, n1527_r, a9_k1a[31], a9_v1[31] );
not U_inv1 ( n1527_r, n1527 );
dff a9_k3a_reg_31_ ( clk, n1527_r, a9_k3a[31], a9_v3[31] );
not U_inv2 ( n1527_r, n1527 );
dff a9_out_1_reg_31_ ( clk, n1527_r, k9[31], k8b[31] );
not U_inv3 ( n1527_r, n1527 );
dff a8_k1a_reg_31_ ( clk, n1527_r, a8_k1a[31], a8_v1[31] );
not U_inv4 ( n1527_r, n1527 );
dff a8_k3a_reg_31_ ( clk, n1527_r, a8_k3a[31], a8_v3[31] );
not U_inv5 ( n1527_r, n1527 );
dff a8_out_1_reg_31_ ( clk, n1526_r, k8[31], k7b[31] );
not U_inv6 ( n1526_r, n1526 );
dff a7_k1a_reg_31_ ( clk, n1526_r, a7_k1a[31], a7_v1[31] );
not U_inv7 ( n1526_r, n1526 );
dff a7_k3a_reg_31_ ( clk, n1526_r, a7_k3a[31], a7_v3[31] );
not U_inv8 ( n1526_r, n1526 );
dff a7_out_1_reg_31_ ( clk, n1526_r, k7[31], k6b[31] );
not U_inv9 ( n1526_r, n1526 );
dff a6_k1a_reg_31_ ( clk, n1526_r, a6_k1a[31], a6_v1[31] );
not U_inv10 ( n1526_r, n1526 );
dff a6_k3a_reg_31_ ( clk, n1526_r, a6_k3a[31], a6_v3[31] );
not U_inv11 ( n1526_r, n1526 );
dff a6_out_1_reg_31_ ( clk, n1526_r, k6[31], k5b[31] );
not U_inv12 ( n1526_r, n1526 );
dff a5_k1a_reg_31_ ( clk, n1526_r, a5_k1a[31], a5_v1[31] );
not U_inv13 ( n1526_r, n1526 );
dff a5_k3a_reg_31_ ( clk, n1526_r, a5_k3a[31], a5_v3[31] );
not U_inv14 ( n1526_r, n1526 );
dff a5_out_1_reg_31_ ( clk, n1526_r, k5[31], k4b[31] );
not U_inv15 ( n1526_r, n1526 );
dff a4_k1a_reg_31_ ( clk, n1526_r, a4_k1a[31], a4_v1[31] );
not U_inv16 ( n1526_r, n1526 );
dff a4_k3a_reg_31_ ( clk, n1526_r, a4_k3a[31], a4_v3[31] );
not U_inv17 ( n1526_r, n1526 );
dff a4_out_1_reg_31_ ( clk, n1525_r, k4[31], k3b[31] );
not U_inv18 ( n1525_r, n1525 );
dff a3_k1a_reg_31_ ( clk, n1525_r, a3_k1a[31], a3_v1[31] );
not U_inv19 ( n1525_r, n1525 );
dff a3_k3a_reg_31_ ( clk, n1525_r, a3_k3a[31], a3_v3[31] );
not U_inv20 ( n1525_r, n1525 );
dff a3_out_1_reg_31_ ( clk, n1525_r, k3[31], k2b[31] );
not U_inv21 ( n1525_r, n1525 );
dff a2_k1a_reg_31_ ( clk, n1525_r, a2_k1a[31], a2_v1[31] );
not U_inv22 ( n1525_r, n1525 );
dff a2_k3a_reg_31_ ( clk, n1525_r, a2_k3a[31], a2_v3[31] );
not U_inv23 ( n1525_r, n1525 );
dff a2_out_1_reg_31_ ( clk, n1525_r, k2[31], k1b[31] );
not U_inv24 ( n1525_r, n1525 );
dff a1_k1a_reg_31_ ( clk, n1525_r, a1_k1a[31], a1_v1[31] );
not U_inv25 ( n1525_r, n1525 );
dff a1_k3a_reg_31_ ( clk, n1525_r, a1_k3a[31], a1_v3[31] );
not U_inv26 ( n1525_r, n1525 );
dff a1_out_1_reg_31_ ( clk, n1525_r, k1[31], k0b[31] );
not U_inv27 ( n1525_r, n1525 );
dff k0_reg_0_ ( clk, n1525_r, k0[0], n1282 );
not U_inv28 ( n1525_r, n1525 );
dff start_r_reg ( clk, n1525_r, ex_wire0, start );
not U_inv29 ( n1019, ex_wire0 );
not U_inv30 ( n1525_r, n1525 );
dff s0_reg_127_ ( clk, n1524_r, s0[127], n1281 );
not U_inv31 ( n1524_r, n1524 );
dff s0_reg_126_ ( clk, n1524_r, s0[126], n1280 );
not U_inv32 ( n1524_r, n1524 );
dff s0_reg_125_ ( clk, n1524_r, s0[125], n1279 );
not U_inv33 ( n1524_r, n1524 );
dff s0_reg_124_ ( clk, n1524_r, s0[124], n1278 );
not U_inv34 ( n1524_r, n1524 );
dff s0_reg_123_ ( clk, n1524_r, s0[123], n1277 );
not U_inv35 ( n1524_r, n1524 );
dff s0_reg_122_ ( clk, n1524_r, s0[122], n1276 );
not U_inv36 ( n1524_r, n1524 );
dff s0_reg_121_ ( clk, n1524_r, s0[121], n1275 );
not U_inv37 ( n1524_r, n1524 );
dff s0_reg_120_ ( clk, n1524_r, s0[120], n1274 );
not U_inv38 ( n1524_r, n1524 );
dff s0_reg_119_ ( clk, n1524_r, s0[119], n1273 );
not U_inv39 ( n1524_r, n1524 );
dff s0_reg_118_ ( clk, n1524_r, s0[118], n1272 );
not U_inv40 ( n1524_r, n1524 );
dff s0_reg_117_ ( clk, n1524_r, s0[117], n1271 );
not U_inv41 ( n1524_r, n1524 );
dff s0_reg_116_ ( clk, n1524_r, s0[116], n1270 );
not U_inv42 ( n1524_r, n1524 );
dff s0_reg_115_ ( clk, n1523_r, s0[115], n1269 );
not U_inv43 ( n1523_r, n1523 );
dff s0_reg_114_ ( clk, n1523_r, s0[114], n1268 );
not U_inv44 ( n1523_r, n1523 );
dff s0_reg_113_ ( clk, n1523_r, s0[113], n1267 );
not U_inv45 ( n1523_r, n1523 );
dff s0_reg_112_ ( clk, n1523_r, s0[112], n1266 );
not U_inv46 ( n1523_r, n1523 );
dff s0_reg_111_ ( clk, n1523_r, s0[111], n1265 );
not U_inv47 ( n1523_r, n1523 );
dff s0_reg_110_ ( clk, n1523_r, s0[110], n1264 );
not U_inv48 ( n1523_r, n1523 );
dff s0_reg_109_ ( clk, n1523_r, s0[109], n1263 );
not U_inv49 ( n1523_r, n1523 );
dff s0_reg_108_ ( clk, n1523_r, s0[108], n1262 );
not U_inv50 ( n1523_r, n1523 );
dff s0_reg_107_ ( clk, n1523_r, s0[107], n1261 );
not U_inv51 ( n1523_r, n1523 );
dff s0_reg_106_ ( clk, n1523_r, s0[106], n1260 );
not U_inv52 ( n1523_r, n1523 );
dff s0_reg_105_ ( clk, n1523_r, s0[105], n1259 );
not U_inv53 ( n1523_r, n1523 );
dff s0_reg_104_ ( clk, n1523_r, s0[104], n1258 );
not U_inv54 ( n1523_r, n1523 );
dff s0_reg_103_ ( clk, n1522_r, s0[103], n1257 );
not U_inv55 ( n1522_r, n1522 );
dff s0_reg_102_ ( clk, n1522_r, s0[102], n1256 );
not U_inv56 ( n1522_r, n1522 );
dff s0_reg_101_ ( clk, n1522_r, s0[101], n1255 );
not U_inv57 ( n1522_r, n1522 );
dff s0_reg_100_ ( clk, n1522_r, s0[100], n1254 );
not U_inv58 ( n1522_r, n1522 );
dff s0_reg_99_ ( clk, n1522_r, s0[99], n1253 );
not U_inv59 ( n1522_r, n1522 );
dff s0_reg_98_ ( clk, n1522_r, s0[98], n1252 );
not U_inv60 ( n1522_r, n1522 );
dff s0_reg_97_ ( clk, n1522_r, s0[97], n1251 );
not U_inv61 ( n1522_r, n1522 );
dff s0_reg_96_ ( clk, n1522_r, s0[96], n1250 );
not U_inv62 ( n1522_r, n1522 );
dff s0_reg_95_ ( clk, n1522_r, s0[95], n1249 );
not U_inv63 ( n1522_r, n1522 );
dff s0_reg_94_ ( clk, n1522_r, s0[94], n1248 );
not U_inv64 ( n1522_r, n1522 );
dff s0_reg_93_ ( clk, n1522_r, s0[93], n1247 );
not U_inv65 ( n1522_r, n1522 );
dff s0_reg_92_ ( clk, n1522_r, s0[92], n1246 );
not U_inv66 ( n1522_r, n1522 );
dff s0_reg_91_ ( clk, n1521_r, s0[91], n1245 );
not U_inv67 ( n1521_r, n1521 );
dff s0_reg_90_ ( clk, n1521_r, s0[90], n1244 );
not U_inv68 ( n1521_r, n1521 );
dff s0_reg_89_ ( clk, n1521_r, s0[89], n1243 );
not U_inv69 ( n1521_r, n1521 );
dff s0_reg_88_ ( clk, n1521_r, s0[88], n1242 );
not U_inv70 ( n1521_r, n1521 );
dff s0_reg_87_ ( clk, n1521_r, s0[87], n1241 );
not U_inv71 ( n1521_r, n1521 );
dff s0_reg_86_ ( clk, n1521_r, s0[86], n1240 );
not U_inv72 ( n1521_r, n1521 );
dff s0_reg_85_ ( clk, n1521_r, s0[85], n1239 );
not U_inv73 ( n1521_r, n1521 );
dff s0_reg_84_ ( clk, n1521_r, s0[84], n1238 );
not U_inv74 ( n1521_r, n1521 );
dff s0_reg_83_ ( clk, n1521_r, s0[83], n1237 );
not U_inv75 ( n1521_r, n1521 );
dff s0_reg_82_ ( clk, n1521_r, s0[82], n1236 );
not U_inv76 ( n1521_r, n1521 );
dff s0_reg_81_ ( clk, n1521_r, s0[81], n1235 );
not U_inv77 ( n1521_r, n1521 );
dff s0_reg_80_ ( clk, n1521_r, s0[80], n1234 );
not U_inv78 ( n1521_r, n1521 );
dff s0_reg_79_ ( clk, n1520_r, s0[79], n1233 );
not U_inv79 ( n1520_r, n1520 );
dff s0_reg_78_ ( clk, n1520_r, s0[78], n1232 );
not U_inv80 ( n1520_r, n1520 );
dff s0_reg_77_ ( clk, n1520_r, s0[77], n1231 );
not U_inv81 ( n1520_r, n1520 );
dff s0_reg_76_ ( clk, n1520_r, s0[76], n1230 );
not U_inv82 ( n1520_r, n1520 );
dff s0_reg_75_ ( clk, n1520_r, s0[75], n1229 );
not U_inv83 ( n1520_r, n1520 );
dff s0_reg_74_ ( clk, n1520_r, s0[74], n1228 );
not U_inv84 ( n1520_r, n1520 );
dff s0_reg_73_ ( clk, n1520_r, s0[73], n1227 );
not U_inv85 ( n1520_r, n1520 );
dff s0_reg_72_ ( clk, n1520_r, s0[72], n1226 );
not U_inv86 ( n1520_r, n1520 );
dff s0_reg_71_ ( clk, n1520_r, s0[71], n1225 );
not U_inv87 ( n1520_r, n1520 );
dff s0_reg_70_ ( clk, n1520_r, s0[70], n1224 );
not U_inv88 ( n1520_r, n1520 );
dff s0_reg_69_ ( clk, n1520_r, s0[69], n1223 );
not U_inv89 ( n1520_r, n1520 );
dff s0_reg_68_ ( clk, n1520_r, s0[68], n1222 );
not U_inv90 ( n1520_r, n1520 );
dff s0_reg_67_ ( clk, n1519_r, s0[67], n1221 );
not U_inv91 ( n1519_r, n1519 );
dff s0_reg_66_ ( clk, n1519_r, s0[66], n1220 );
not U_inv92 ( n1519_r, n1519 );
dff s0_reg_65_ ( clk, n1519_r, s0[65], n1219 );
not U_inv93 ( n1519_r, n1519 );
dff s0_reg_64_ ( clk, n1519_r, s0[64], n1218 );
not U_inv94 ( n1519_r, n1519 );
dff s0_reg_63_ ( clk, n1519_r, s0[63], n1217 );
not U_inv95 ( n1519_r, n1519 );
dff s0_reg_62_ ( clk, n1519_r, s0[62], n1216 );
not U_inv96 ( n1519_r, n1519 );
dff s0_reg_61_ ( clk, n1519_r, s0[61], n1215 );
not U_inv97 ( n1519_r, n1519 );
dff s0_reg_60_ ( clk, n1519_r, s0[60], n1214 );
not U_inv98 ( n1519_r, n1519 );
dff s0_reg_59_ ( clk, n1519_r, s0[59], n1213 );
not U_inv99 ( n1519_r, n1519 );
dff s0_reg_58_ ( clk, n1519_r, s0[58], n1212 );
not U_inv100 ( n1519_r, n1519 );
dff s0_reg_57_ ( clk, n1519_r, s0[57], n1211 );
not U_inv101 ( n1519_r, n1519 );
dff s0_reg_56_ ( clk, n1519_r, s0[56], n1210 );
not U_inv102 ( n1519_r, n1519 );
dff s0_reg_55_ ( clk, n1518_r, s0[55], n1209 );
not U_inv103 ( n1518_r, n1518 );
dff s0_reg_54_ ( clk, n1518_r, s0[54], n1208 );
not U_inv104 ( n1518_r, n1518 );
dff s0_reg_53_ ( clk, n1518_r, s0[53], n1207 );
not U_inv105 ( n1518_r, n1518 );
dff s0_reg_52_ ( clk, n1518_r, s0[52], n1206 );
not U_inv106 ( n1518_r, n1518 );
dff s0_reg_51_ ( clk, n1518_r, s0[51], n1205 );
not U_inv107 ( n1518_r, n1518 );
dff s0_reg_50_ ( clk, n1518_r, s0[50], n1204 );
not U_inv108 ( n1518_r, n1518 );
dff s0_reg_49_ ( clk, n1518_r, s0[49], n1203 );
not U_inv109 ( n1518_r, n1518 );
dff s0_reg_48_ ( clk, n1518_r, s0[48], n1202 );
not U_inv110 ( n1518_r, n1518 );
dff s0_reg_47_ ( clk, n1518_r, s0[47], n1201 );
not U_inv111 ( n1518_r, n1518 );
dff s0_reg_46_ ( clk, n1518_r, s0[46], n1200 );
not U_inv112 ( n1518_r, n1518 );
dff s0_reg_45_ ( clk, n1518_r, s0[45], n1199 );
not U_inv113 ( n1518_r, n1518 );
dff s0_reg_44_ ( clk, n1518_r, s0[44], n1198 );
not U_inv114 ( n1518_r, n1518 );
dff s0_reg_43_ ( clk, n1517_r, s0[43], n1197 );
not U_inv115 ( n1517_r, n1517 );
dff s0_reg_42_ ( clk, n1517_r, s0[42], n1196 );
not U_inv116 ( n1517_r, n1517 );
dff s0_reg_41_ ( clk, n1517_r, s0[41], n1195 );
not U_inv117 ( n1517_r, n1517 );
dff s0_reg_40_ ( clk, n1517_r, s0[40], n1194 );
not U_inv118 ( n1517_r, n1517 );
dff s0_reg_39_ ( clk, n1517_r, s0[39], n1193 );
not U_inv119 ( n1517_r, n1517 );
dff s0_reg_38_ ( clk, n1517_r, s0[38], n1192 );
not U_inv120 ( n1517_r, n1517 );
dff s0_reg_37_ ( clk, n1517_r, s0[37], n1191 );
not U_inv121 ( n1517_r, n1517 );
dff s0_reg_36_ ( clk, n1517_r, s0[36], n1190 );
not U_inv122 ( n1517_r, n1517 );
dff s0_reg_35_ ( clk, n1517_r, s0[35], n1189 );
not U_inv123 ( n1517_r, n1517 );
dff s0_reg_34_ ( clk, n1517_r, s0[34], n1188 );
not U_inv124 ( n1517_r, n1517 );
dff s0_reg_33_ ( clk, n1517_r, s0[33], n1187 );
not U_inv125 ( n1517_r, n1517 );
dff s0_reg_32_ ( clk, n1517_r, s0[32], n1186 );
not U_inv126 ( n1517_r, n1517 );
dff s0_reg_31_ ( clk, n1516_r, s0[31], n1185 );
not U_inv127 ( n1516_r, n1516 );
dff s0_reg_30_ ( clk, n1516_r, s0[30], n1184 );
not U_inv128 ( n1516_r, n1516 );
dff s0_reg_29_ ( clk, n1516_r, s0[29], n1183 );
not U_inv129 ( n1516_r, n1516 );
dff s0_reg_28_ ( clk, n1516_r, s0[28], n1182 );
not U_inv130 ( n1516_r, n1516 );
dff s0_reg_27_ ( clk, n1516_r, s0[27], n1181 );
not U_inv131 ( n1516_r, n1516 );
dff s0_reg_26_ ( clk, n1516_r, s0[26], n1180 );
not U_inv132 ( n1516_r, n1516 );
dff s0_reg_25_ ( clk, n1516_r, s0[25], n1179 );
not U_inv133 ( n1516_r, n1516 );
dff s0_reg_24_ ( clk, n1516_r, s0[24], n1178 );
not U_inv134 ( n1516_r, n1516 );
dff s0_reg_23_ ( clk, n1516_r, s0[23], n1177 );
not U_inv135 ( n1516_r, n1516 );
dff s0_reg_22_ ( clk, n1516_r, s0[22], n1176 );
not U_inv136 ( n1516_r, n1516 );
dff s0_reg_21_ ( clk, n1516_r, s0[21], n1175 );
not U_inv137 ( n1516_r, n1516 );
dff s0_reg_20_ ( clk, n1516_r, s0[20], n1174 );
not U_inv138 ( n1516_r, n1516 );
dff s0_reg_19_ ( clk, n1515_r, s0[19], n1173 );
not U_inv139 ( n1515_r, n1515 );
dff s0_reg_18_ ( clk, n1515_r, s0[18], n1172 );
not U_inv140 ( n1515_r, n1515 );
dff s0_reg_17_ ( clk, n1515_r, s0[17], n1171 );
not U_inv141 ( n1515_r, n1515 );
dff s0_reg_16_ ( clk, n1515_r, s0[16], n1170 );
not U_inv142 ( n1515_r, n1515 );
dff s0_reg_15_ ( clk, n1515_r, s0[15], n1169 );
not U_inv143 ( n1515_r, n1515 );
dff s0_reg_14_ ( clk, n1515_r, s0[14], n1168 );
not U_inv144 ( n1515_r, n1515 );
dff s0_reg_13_ ( clk, n1515_r, s0[13], n1167 );
not U_inv145 ( n1515_r, n1515 );
dff s0_reg_12_ ( clk, n1515_r, s0[12], n1166 );
not U_inv146 ( n1515_r, n1515 );
dff s0_reg_11_ ( clk, n1515_r, s0[11], n1165 );
not U_inv147 ( n1515_r, n1515 );
dff s0_reg_10_ ( clk, n1515_r, s0[10], n1164 );
not U_inv148 ( n1515_r, n1515 );
dff s0_reg_9_ ( clk, n1515_r, s0[9], n1163 );
not U_inv149 ( n1515_r, n1515 );
dff s0_reg_8_ ( clk, n1515_r, s0[8], n1162 );
not U_inv150 ( n1515_r, n1515 );
dff s0_reg_7_ ( clk, n1514_r, s0[7], n1161 );
not U_inv151 ( n1514_r, n1514 );
dff s0_reg_6_ ( clk, n1514_r, s0[6], n1160 );
not U_inv152 ( n1514_r, n1514 );
dff s0_reg_5_ ( clk, n1514_r, s0[5], n1159 );
not U_inv153 ( n1514_r, n1514 );
dff s0_reg_4_ ( clk, n1514_r, s0[4], n1158 );
not U_inv154 ( n1514_r, n1514 );
dff s0_reg_3_ ( clk, n1514_r, s0[3], n1157 );
not U_inv155 ( n1514_r, n1514 );
dff s0_reg_2_ ( clk, n1514_r, s0[2], n1156 );
not U_inv156 ( n1514_r, n1514 );
dff s0_reg_1_ ( clk, n1514_r, s0[1], n1155 );
not U_inv157 ( n1514_r, n1514 );
dff s0_reg_0_ ( clk, n1514_r, s0[0], n1154 );
not U_inv158 ( n1514_r, n1514 );
dff k0_reg_127_ ( clk, n1514_r, k0[127], n1153 );
not U_inv159 ( n1018, k0[127] );
not U_inv160 ( n1514_r, n1514 );
dff k0_reg_126_ ( clk, n1514_r, k0[126], n1152 );
not U_inv161 ( n1017, k0[126] );
not U_inv162 ( n1514_r, n1514 );
dff k0_reg_125_ ( clk, n1514_r, k0[125], n1151 );
not U_inv163 ( n1016, k0[125] );
not U_inv164 ( n1514_r, n1514 );
dff k0_reg_124_ ( clk, n1514_r, k0[124], n1150 );
not U_inv165 ( n1015, k0[124] );
not U_inv166 ( n1514_r, n1514 );
dff k0_reg_123_ ( clk, n1513_r, k0[123], n1149 );
not U_inv167 ( n1014, k0[123] );
not U_inv168 ( n1513_r, n1513 );
dff k0_reg_122_ ( clk, n1513_r, k0[122], n1148 );
not U_inv169 ( n1013, k0[122] );
not U_inv170 ( n1513_r, n1513 );
dff k0_reg_121_ ( clk, n1513_r, k0[121], n1147 );
not U_inv171 ( n1012, k0[121] );
not U_inv172 ( n1513_r, n1513 );
dff k0_reg_120_ ( clk, n1513_r, ex_wire1, n1146 );
not U_inv173 ( n1284, ex_wire1 );
not U_inv174 ( n1513_r, n1513 );
dff k0_reg_119_ ( clk, n1513_r, k0[119], n1145 );
not U_inv175 ( n1011, k0[119] );
not U_inv176 ( n1513_r, n1513 );
dff k0_reg_118_ ( clk, n1513_r, k0[118], n1144 );
not U_inv177 ( n1010, k0[118] );
not U_inv178 ( n1513_r, n1513 );
dff k0_reg_117_ ( clk, n1513_r, k0[117], n1143 );
not U_inv179 ( n1009, k0[117] );
not U_inv180 ( n1513_r, n1513 );
dff k0_reg_116_ ( clk, n1513_r, k0[116], n1142 );
not U_inv181 ( n1008, k0[116] );
not U_inv182 ( n1513_r, n1513 );
dff k0_reg_115_ ( clk, n1513_r, k0[115], n1141 );
not U_inv183 ( n1007, k0[115] );
not U_inv184 ( n1513_r, n1513 );
dff k0_reg_114_ ( clk, n1513_r, k0[114], n1140 );
not U_inv185 ( n1006, k0[114] );
not U_inv186 ( n1513_r, n1513 );
dff k0_reg_113_ ( clk, n1513_r, k0[113], n1139 );
not U_inv187 ( n1005, k0[113] );
not U_inv188 ( n1513_r, n1513 );
dff k0_reg_112_ ( clk, n1513_r, k0[112], n1138 );
not U_inv189 ( n1004, k0[112] );
not U_inv190 ( n1513_r, n1513 );
dff k0_reg_111_ ( clk, n1512_r, k0[111], n1137 );
not U_inv191 ( n1003, k0[111] );
not U_inv192 ( n1512_r, n1512 );
dff k0_reg_110_ ( clk, n1512_r, k0[110], n1136 );
not U_inv193 ( n1002, k0[110] );
not U_inv194 ( n1512_r, n1512 );
dff k0_reg_109_ ( clk, n1512_r, k0[109], n1135 );
not U_inv195 ( n1001, k0[109] );
not U_inv196 ( n1512_r, n1512 );
dff k0_reg_108_ ( clk, n1512_r, k0[108], n1134 );
not U_inv197 ( n1000, k0[108] );
not U_inv198 ( n1512_r, n1512 );
dff k0_reg_107_ ( clk, n1512_r, k0[107], n1133 );
not U_inv199 ( n999, k0[107] );
not U_inv200 ( n1512_r, n1512 );
dff k0_reg_106_ ( clk, n1512_r, k0[106], n1132 );
not U_inv201 ( n998, k0[106] );
not U_inv202 ( n1512_r, n1512 );
dff k0_reg_105_ ( clk, n1512_r, k0[105], n1131 );
not U_inv203 ( n997, k0[105] );
not U_inv204 ( n1512_r, n1512 );
dff k0_reg_104_ ( clk, n1512_r, k0[104], n1130 );
not U_inv205 ( n996, k0[104] );
not U_inv206 ( n1512_r, n1512 );
dff k0_reg_103_ ( clk, n1512_r, k0[103], n1129 );
not U_inv207 ( n995, k0[103] );
not U_inv208 ( n1512_r, n1512 );
dff k0_reg_102_ ( clk, n1512_r, k0[102], n1128 );
not U_inv209 ( n994, k0[102] );
not U_inv210 ( n1512_r, n1512 );
dff k0_reg_101_ ( clk, n1512_r, k0[101], n1127 );
not U_inv211 ( n993, k0[101] );
not U_inv212 ( n1512_r, n1512 );
dff k0_reg_100_ ( clk, n1512_r, k0[100], n1126 );
not U_inv213 ( n992, k0[100] );
not U_inv214 ( n1512_r, n1512 );
dff k0_reg_99_ ( clk, n1511_r, k0[99], n1125 );
not U_inv215 ( n991, k0[99] );
not U_inv216 ( n1511_r, n1511 );
dff k0_reg_98_ ( clk, n1511_r, k0[98], n1124 );
not U_inv217 ( n990, k0[98] );
not U_inv218 ( n1511_r, n1511 );
dff k0_reg_97_ ( clk, n1511_r, k0[97], n1123 );
not U_inv219 ( n989, k0[97] );
not U_inv220 ( n1511_r, n1511 );
dff k0_reg_96_ ( clk, n1511_r, k0[96], n1122 );
not U_inv221 ( n988, k0[96] );
not U_inv222 ( n1511_r, n1511 );
dff k0_reg_95_ ( clk, n1511_r, ex_wire2, n1121 );
not U_inv223 ( n987, ex_wire2 );
not U_inv224 ( n1511_r, n1511 );
dff k0_reg_94_ ( clk, n1511_r, ex_wire3, n1120 );
not U_inv225 ( n986, ex_wire3 );
not U_inv226 ( n1511_r, n1511 );
dff k0_reg_93_ ( clk, n1511_r, ex_wire4, n1119 );
not U_inv227 ( n985, ex_wire4 );
not U_inv228 ( n1511_r, n1511 );
dff k0_reg_92_ ( clk, n1511_r, ex_wire5, n1118 );
not U_inv229 ( n984, ex_wire5 );
not U_inv230 ( n1511_r, n1511 );
dff k0_reg_91_ ( clk, n1511_r, ex_wire6, n1117 );
not U_inv231 ( n983, ex_wire6 );
not U_inv232 ( n1511_r, n1511 );
dff k0_reg_90_ ( clk, n1511_r, ex_wire7, n1116 );
not U_inv233 ( n982, ex_wire7 );
not U_inv234 ( n1511_r, n1511 );
dff k0_reg_89_ ( clk, n1511_r, ex_wire8, n1115 );
not U_inv235 ( n981, ex_wire8 );
not U_inv236 ( n1511_r, n1511 );
dff k0_reg_88_ ( clk, n1511_r, ex_wire9, n1114 );
not U_inv237 ( n980, ex_wire9 );
not U_inv238 ( n1511_r, n1511 );
dff k0_reg_87_ ( clk, n1510_r, ex_wire10, n1113 );
not U_inv239 ( n979, ex_wire10 );
not U_inv240 ( n1510_r, n1510 );
dff k0_reg_86_ ( clk, n1510_r, ex_wire11, n1112 );
not U_inv241 ( n978, ex_wire11 );
not U_inv242 ( n1510_r, n1510 );
dff k0_reg_85_ ( clk, n1510_r, ex_wire12, n1111 );
not U_inv243 ( n977, ex_wire12 );
not U_inv244 ( n1510_r, n1510 );
dff k0_reg_84_ ( clk, n1510_r, ex_wire13, n1110 );
not U_inv245 ( n976, ex_wire13 );
not U_inv246 ( n1510_r, n1510 );
dff k0_reg_83_ ( clk, n1510_r, ex_wire14, n1109 );
not U_inv247 ( n975, ex_wire14 );
not U_inv248 ( n1510_r, n1510 );
dff k0_reg_82_ ( clk, n1510_r, ex_wire15, n1108 );
not U_inv249 ( n974, ex_wire15 );
not U_inv250 ( n1510_r, n1510 );
dff k0_reg_81_ ( clk, n1510_r, ex_wire16, n1107 );
not U_inv251 ( n973, ex_wire16 );
not U_inv252 ( n1510_r, n1510 );
dff k0_reg_80_ ( clk, n1510_r, ex_wire17, n1106 );
not U_inv253 ( n972, ex_wire17 );
not U_inv254 ( n1510_r, n1510 );
dff k0_reg_79_ ( clk, n1510_r, ex_wire18, n1105 );
not U_inv255 ( n971, ex_wire18 );
not U_inv256 ( n1510_r, n1510 );
dff k0_reg_78_ ( clk, n1510_r, ex_wire19, n1104 );
not U_inv257 ( n970, ex_wire19 );
not U_inv258 ( n1510_r, n1510 );
dff k0_reg_77_ ( clk, n1510_r, ex_wire20, n1103 );
not U_inv259 ( n969, ex_wire20 );
not U_inv260 ( n1510_r, n1510 );
dff k0_reg_76_ ( clk, n1510_r, ex_wire21, n1102 );
not U_inv261 ( n968, ex_wire21 );
not U_inv262 ( n1510_r, n1510 );
dff k0_reg_75_ ( clk, n1509_r, ex_wire22, n1101 );
not U_inv263 ( n967, ex_wire22 );
not U_inv264 ( n1509_r, n1509 );
dff k0_reg_74_ ( clk, n1509_r, ex_wire23, n1100 );
not U_inv265 ( n966, ex_wire23 );
not U_inv266 ( n1509_r, n1509 );
dff k0_reg_73_ ( clk, n1509_r, ex_wire24, n1099 );
not U_inv267 ( n965, ex_wire24 );
not U_inv268 ( n1509_r, n1509 );
dff k0_reg_72_ ( clk, n1509_r, ex_wire25, n1098 );
not U_inv269 ( n964, ex_wire25 );
not U_inv270 ( n1509_r, n1509 );
dff k0_reg_71_ ( clk, n1509_r, ex_wire26, n1097 );
not U_inv271 ( n963, ex_wire26 );
not U_inv272 ( n1509_r, n1509 );
dff k0_reg_70_ ( clk, n1509_r, ex_wire27, n1096 );
not U_inv273 ( n962, ex_wire27 );
not U_inv274 ( n1509_r, n1509 );
dff k0_reg_69_ ( clk, n1509_r, ex_wire28, n1095 );
not U_inv275 ( n961, ex_wire28 );
not U_inv276 ( n1509_r, n1509 );
dff k0_reg_68_ ( clk, n1509_r, ex_wire29, n1094 );
not U_inv277 ( n960, ex_wire29 );
not U_inv278 ( n1509_r, n1509 );
dff k0_reg_67_ ( clk, n1509_r, ex_wire30, n1093 );
not U_inv279 ( n959, ex_wire30 );
not U_inv280 ( n1509_r, n1509 );
dff k0_reg_66_ ( clk, n1509_r, ex_wire31, n1092 );
not U_inv281 ( n958, ex_wire31 );
not U_inv282 ( n1509_r, n1509 );
dff k0_reg_65_ ( clk, n1509_r, ex_wire32, n1091 );
not U_inv283 ( n957, ex_wire32 );
not U_inv284 ( n1509_r, n1509 );
dff k0_reg_64_ ( clk, n1509_r, ex_wire33, n1090 );
not U_inv285 ( n956, ex_wire33 );
not U_inv286 ( n1509_r, n1509 );
dff k0_reg_63_ ( clk, n1508_r, ex_wire34, n1089 );
not U_inv287 ( n955, ex_wire34 );
not U_inv288 ( n1508_r, n1508 );
dff k0_reg_62_ ( clk, n1508_r, ex_wire35, n1088 );
not U_inv289 ( n954, ex_wire35 );
not U_inv290 ( n1508_r, n1508 );
dff k0_reg_61_ ( clk, n1508_r, ex_wire36, n1087 );
not U_inv291 ( n953, ex_wire36 );
not U_inv292 ( n1508_r, n1508 );
dff k0_reg_60_ ( clk, n1508_r, ex_wire37, n1086 );
not U_inv293 ( n952, ex_wire37 );
not U_inv294 ( n1508_r, n1508 );
dff k0_reg_59_ ( clk, n1508_r, ex_wire38, n1085 );
not U_inv295 ( n951, ex_wire38 );
not U_inv296 ( n1508_r, n1508 );
dff k0_reg_58_ ( clk, n1508_r, ex_wire39, n1084 );
not U_inv297 ( n950, ex_wire39 );
not U_inv298 ( n1508_r, n1508 );
dff k0_reg_57_ ( clk, n1508_r, ex_wire40, n1083 );
not U_inv299 ( n949, ex_wire40 );
not U_inv300 ( n1508_r, n1508 );
dff k0_reg_56_ ( clk, n1508_r, ex_wire41, n1082 );
not U_inv301 ( n948, ex_wire41 );
not U_inv302 ( n1508_r, n1508 );
dff k0_reg_55_ ( clk, n1508_r, ex_wire42, n1081 );
not U_inv303 ( n947, ex_wire42 );
not U_inv304 ( n1508_r, n1508 );
dff k0_reg_54_ ( clk, n1508_r, ex_wire43, n1080 );
not U_inv305 ( n946, ex_wire43 );
not U_inv306 ( n1508_r, n1508 );
dff k0_reg_53_ ( clk, n1508_r, ex_wire44, n1079 );
not U_inv307 ( n945, ex_wire44 );
not U_inv308 ( n1508_r, n1508 );
dff k0_reg_52_ ( clk, n1508_r, ex_wire45, n1078 );
not U_inv309 ( n944, ex_wire45 );
not U_inv310 ( n1508_r, n1508 );
dff k0_reg_51_ ( clk, n1507_r, ex_wire46, n1077 );
not U_inv311 ( n943, ex_wire46 );
not U_inv312 ( n1507_r, n1507 );
dff k0_reg_50_ ( clk, n1507_r, ex_wire47, n1076 );
not U_inv313 ( n942, ex_wire47 );
not U_inv314 ( n1507_r, n1507 );
dff k0_reg_49_ ( clk, n1507_r, ex_wire48, n1075 );
not U_inv315 ( n941, ex_wire48 );
not U_inv316 ( n1507_r, n1507 );
dff k0_reg_48_ ( clk, n1507_r, ex_wire49, n1074 );
not U_inv317 ( n940, ex_wire49 );
not U_inv318 ( n1507_r, n1507 );
dff k0_reg_47_ ( clk, n1507_r, ex_wire50, n1073 );
not U_inv319 ( n939, ex_wire50 );
not U_inv320 ( n1507_r, n1507 );
dff k0_reg_46_ ( clk, n1507_r, ex_wire51, n1072 );
not U_inv321 ( n938, ex_wire51 );
not U_inv322 ( n1507_r, n1507 );
dff k0_reg_45_ ( clk, n1507_r, ex_wire52, n1071 );
not U_inv323 ( n937, ex_wire52 );
not U_inv324 ( n1507_r, n1507 );
dff k0_reg_44_ ( clk, n1507_r, ex_wire53, n1070 );
not U_inv325 ( n936, ex_wire53 );
not U_inv326 ( n1507_r, n1507 );
dff k0_reg_43_ ( clk, n1507_r, ex_wire54, n1069 );
not U_inv327 ( n935, ex_wire54 );
not U_inv328 ( n1507_r, n1507 );
dff k0_reg_42_ ( clk, n1507_r, ex_wire55, n1068 );
not U_inv329 ( n934, ex_wire55 );
not U_inv330 ( n1507_r, n1507 );
dff k0_reg_41_ ( clk, n1507_r, ex_wire56, n1067 );
not U_inv331 ( n933, ex_wire56 );
not U_inv332 ( n1507_r, n1507 );
dff k0_reg_40_ ( clk, n1507_r, ex_wire57, n1066 );
not U_inv333 ( n932, ex_wire57 );
not U_inv334 ( n1507_r, n1507 );
dff k0_reg_39_ ( clk, n1506_r, ex_wire58, n1065 );
not U_inv335 ( n931, ex_wire58 );
not U_inv336 ( n1506_r, n1506 );
dff k0_reg_38_ ( clk, n1506_r, ex_wire59, n1064 );
not U_inv337 ( n930, ex_wire59 );
not U_inv338 ( n1506_r, n1506 );
dff k0_reg_37_ ( clk, n1506_r, ex_wire60, n1063 );
not U_inv339 ( n929, ex_wire60 );
not U_inv340 ( n1506_r, n1506 );
dff k0_reg_36_ ( clk, n1506_r, ex_wire61, n1062 );
not U_inv341 ( n928, ex_wire61 );
not U_inv342 ( n1506_r, n1506 );
dff k0_reg_35_ ( clk, n1506_r, ex_wire62, n1061 );
not U_inv343 ( n927, ex_wire62 );
not U_inv344 ( n1506_r, n1506 );
dff k0_reg_34_ ( clk, n1506_r, ex_wire63, n1060 );
not U_inv345 ( n926, ex_wire63 );
not U_inv346 ( n1506_r, n1506 );
dff k0_reg_33_ ( clk, n1506_r, ex_wire64, n1059 );
not U_inv347 ( n925, ex_wire64 );
not U_inv348 ( n1506_r, n1506 );
dff k0_reg_32_ ( clk, n1506_r, ex_wire65, n1058 );
not U_inv349 ( n924, ex_wire65 );
not U_inv350 ( n1506_r, n1506 );
dff k0_reg_31_ ( clk, n1506_r, k0[31], n1057 );
not U_inv351 ( n1506_r, n1506 );
dff k0_reg_30_ ( clk, n1506_r, k0[30], n1056 );
not U_inv352 ( n1506_r, n1506 );
dff k0_reg_29_ ( clk, n1506_r, k0[29], n1055 );
not U_inv353 ( n1506_r, n1506 );
dff k0_reg_28_ ( clk, n1506_r, k0[28], n1054 );
not U_inv354 ( n1506_r, n1506 );
dff k0_reg_27_ ( clk, n1505_r, k0[27], n1053 );
not U_inv355 ( n1505_r, n1505 );
dff k0_reg_26_ ( clk, n1505_r, k0[26], n1052 );
not U_inv356 ( n1505_r, n1505 );
dff k0_reg_25_ ( clk, n1505_r, k0[25], n1051 );
not U_inv357 ( n1505_r, n1505 );
dff k0_reg_24_ ( clk, n1505_r, k0[24], n1050 );
not U_inv358 ( n1505_r, n1505 );
dff k0_reg_23_ ( clk, n1505_r, k0[23], n1049 );
not U_inv359 ( n1505_r, n1505 );
dff k0_reg_22_ ( clk, n1505_r, k0[22], n1048 );
not U_inv360 ( n1505_r, n1505 );
dff k0_reg_21_ ( clk, n1505_r, k0[21], n1047 );
not U_inv361 ( n1505_r, n1505 );
dff k0_reg_20_ ( clk, n1505_r, k0[20], n1046 );
not U_inv362 ( n1505_r, n1505 );
dff k0_reg_19_ ( clk, n1505_r, k0[19], n1045 );
not U_inv363 ( n1505_r, n1505 );
dff k0_reg_18_ ( clk, n1505_r, k0[18], n1044 );
not U_inv364 ( n1505_r, n1505 );
dff k0_reg_17_ ( clk, n1505_r, k0[17], n1043 );
not U_inv365 ( n1505_r, n1505 );
dff k0_reg_16_ ( clk, n1505_r, k0[16], n1042 );
not U_inv366 ( n1505_r, n1505 );
dff k0_reg_15_ ( clk, n1504_r, k0[15], n1041 );
not U_inv367 ( n1504_r, n1504 );
dff k0_reg_14_ ( clk, n1504_r, k0[14], n1040 );
not U_inv368 ( n1504_r, n1504 );
dff k0_reg_13_ ( clk, n1504_r, k0[13], n1039 );
not U_inv369 ( n1504_r, n1504 );
dff k0_reg_12_ ( clk, n1504_r, k0[12], n1038 );
not U_inv370 ( n1504_r, n1504 );
dff k0_reg_11_ ( clk, n1504_r, k0[11], n1037 );
not U_inv371 ( n1504_r, n1504 );
dff k0_reg_10_ ( clk, n1504_r, k0[10], n1036 );
not U_inv372 ( n1504_r, n1504 );
dff k0_reg_9_ ( clk, n1504_r, k0[9], n1035 );
not U_inv373 ( n1504_r, n1504 );
dff k0_reg_8_ ( clk, n1504_r, k0[8], n1034 );
not U_inv374 ( n1504_r, n1504 );
dff k0_reg_7_ ( clk, n1504_r, k0[7], n1033 );
not U_inv375 ( n1504_r, n1504 );
dff k0_reg_6_ ( clk, n1504_r, k0[6], n1032 );
not U_inv376 ( n1504_r, n1504 );
dff k0_reg_5_ ( clk, n1504_r, k0[5], n1031 );
not U_inv377 ( n1504_r, n1504 );
dff k0_reg_4_ ( clk, n1504_r, k0[4], n1030 );
not U_inv378 ( n1504_r, n1504 );
dff k0_reg_3_ ( clk, n1503_r, k0[3], n1029 );
not U_inv379 ( n1503_r, n1503 );
dff k0_reg_2_ ( clk, n1503_r, k0[2], n1028 );
not U_inv380 ( n1503_r, n1503 );
dff k0_reg_1_ ( clk, n1503_r, k0[1], n1027 );
not U_inv381 ( n1503_r, n1503 );
dff validCounter_reg_0_ ( clk, n1503_r, validCounter[0], n1026 );
not U_inv382 ( n1301, validCounter[0] );
not U_inv383 ( n1503_r, n1503 );
dff validCounter_reg_1_ ( clk, n1503_r, validCounter[1], n1025 );
not U_inv384 ( n1503_r, n1503 );
dff validCounter_reg_2_ ( clk, n1503_r, validCounter[2], n1024 );
not U_inv385 ( n1503_r, n1503 );
dff validCounter_reg_3_ ( clk, n1503_r, validCounter[3], n1023 );
not U_inv386 ( n1020, validCounter[3] );
not U_inv387 ( n1503_r, n1503 );
dff validCounter_reg_4_ ( clk, n1503_r, validCounter[4], n1022 );
not U_inv388 ( n1021, validCounter[4] );
not U_inv389 ( n1503_r, n1503 );
dff a1_k0a_reg_0_ ( clk, n1503_r, a1_k0a[0], k0[96] );
not U_inv390 ( n1503_r, n1503 );
dff a1_out_1_reg_96_ ( clk, n1503_r, k1[96], k0b[96] );
not U_inv391 ( n1503_r, n1503 );
dff a1_k0a_reg_1_ ( clk, n1503_r, a1_k0a[1], k0[97] );
not U_inv392 ( n1503_r, n1503 );
dff a1_out_1_reg_97_ ( clk, n1503_r, k1[97], k0b[97] );
not U_inv393 ( n1503_r, n1503 );
dff a1_k0a_reg_2_ ( clk, n1502_r, a1_k0a[2], k0[98] );
not U_inv394 ( n1502_r, n1502 );
dff a1_out_1_reg_98_ ( clk, n1502_r, k1[98], k0b[98] );
not U_inv395 ( n1502_r, n1502 );
dff a1_k0a_reg_3_ ( clk, n1502_r, a1_k0a[3], k0[99] );
not U_inv396 ( n1502_r, n1502 );
dff a1_out_1_reg_99_ ( clk, n1502_r, k1[99], k0b[99] );
not U_inv397 ( n1502_r, n1502 );
dff a1_k0a_reg_4_ ( clk, n1502_r, a1_k0a[4], k0[100] );
not U_inv398 ( n1502_r, n1502 );
dff a1_out_1_reg_100_ ( clk, n1502_r, k1[100], k0b[100] );
not U_inv399 ( n704, k1[100] );
not U_inv400 ( n1502_r, n1502 );
dff a1_k0a_reg_5_ ( clk, n1502_r, a1_k0a[5], k0[101] );
not U_inv401 ( n1502_r, n1502 );
dff a1_out_1_reg_101_ ( clk, n1502_r, k1[101], k0b[101] );
not U_inv402 ( n705, k1[101] );
not U_inv403 ( n1502_r, n1502 );
dff a1_k0a_reg_6_ ( clk, n1502_r, a1_k0a[6], k0[102] );
not U_inv404 ( n1502_r, n1502 );
dff a1_out_1_reg_102_ ( clk, n1502_r, k1[102], k0b[102] );
not U_inv405 ( n706, k1[102] );
not U_inv406 ( n1502_r, n1502 );
dff a1_k0a_reg_7_ ( clk, n1502_r, a1_k0a[7], k0[103] );
not U_inv407 ( n1502_r, n1502 );
dff a1_out_1_reg_103_ ( clk, n1502_r, k1[103], k0b[103] );
not U_inv408 ( n707, k1[103] );
not U_inv409 ( n1502_r, n1502 );
dff a1_k0a_reg_8_ ( clk, n1501_r, a1_k0a[8], k0[104] );
not U_inv410 ( n1501_r, n1501 );
dff a1_out_1_reg_104_ ( clk, n1501_r, k1[104], k0b[104] );
not U_inv411 ( n708, k1[104] );
not U_inv412 ( n1501_r, n1501 );
dff a1_k0a_reg_9_ ( clk, n1501_r, a1_k0a[9], k0[105] );
not U_inv413 ( n1501_r, n1501 );
dff a1_out_1_reg_105_ ( clk, n1501_r, k1[105], k0b[105] );
not U_inv414 ( n709, k1[105] );
not U_inv415 ( n1501_r, n1501 );
dff a1_k0a_reg_10_ ( clk, n1501_r, a1_k0a[10], k0[106] );
not U_inv416 ( n1501_r, n1501 );
dff a1_out_1_reg_106_ ( clk, n1501_r, k1[106], k0b[106] );
not U_inv417 ( n680, k1[106] );
not U_inv418 ( n1501_r, n1501 );
dff a1_k0a_reg_11_ ( clk, n1501_r, a1_k0a[11], k0[107] );
not U_inv419 ( n1501_r, n1501 );
dff a1_out_1_reg_107_ ( clk, n1501_r, k1[107], k0b[107] );
not U_inv420 ( n681, k1[107] );
not U_inv421 ( n1501_r, n1501 );
dff a1_k0a_reg_12_ ( clk, n1501_r, a1_k0a[12], k0[108] );
not U_inv422 ( n1501_r, n1501 );
dff a1_out_1_reg_108_ ( clk, n1501_r, k1[108], k0b[108] );
not U_inv423 ( n682, k1[108] );
not U_inv424 ( n1501_r, n1501 );
dff a1_k0a_reg_13_ ( clk, n1501_r, a1_k0a[13], k0[109] );
not U_inv425 ( n1501_r, n1501 );
dff a1_out_1_reg_109_ ( clk, n1501_r, k1[109], k0b[109] );
not U_inv426 ( n683, k1[109] );
not U_inv427 ( n1501_r, n1501 );
dff a1_k0a_reg_14_ ( clk, n1500_r, a1_k0a[14], k0[110] );
not U_inv428 ( n1500_r, n1500 );
dff a1_out_1_reg_110_ ( clk, n1500_r, k1[110], k0b[110] );
not U_inv429 ( n684, k1[110] );
not U_inv430 ( n1500_r, n1500 );
dff a1_k0a_reg_15_ ( clk, n1500_r, a1_k0a[15], k0[111] );
not U_inv431 ( n1500_r, n1500 );
dff a1_out_1_reg_111_ ( clk, n1500_r, k1[111], k0b[111] );
not U_inv432 ( n685, k1[111] );
not U_inv433 ( n1500_r, n1500 );
dff a1_k0a_reg_16_ ( clk, n1500_r, a1_k0a[16], k0[112] );
not U_inv434 ( n1500_r, n1500 );
dff a1_out_1_reg_112_ ( clk, n1500_r, k1[112], k0b[112] );
not U_inv435 ( n686, k1[112] );
not U_inv436 ( n1500_r, n1500 );
dff a1_k0a_reg_17_ ( clk, n1500_r, a1_k0a[17], k0[113] );
not U_inv437 ( n1500_r, n1500 );
dff a1_out_1_reg_113_ ( clk, n1500_r, k1[113], k0b[113] );
not U_inv438 ( n687, k1[113] );
not U_inv439 ( n1500_r, n1500 );
dff a1_k0a_reg_18_ ( clk, n1500_r, a1_k0a[18], k0[114] );
not U_inv440 ( n1500_r, n1500 );
dff a1_out_1_reg_114_ ( clk, n1500_r, k1[114], k0b[114] );
not U_inv441 ( n688, k1[114] );
not U_inv442 ( n1500_r, n1500 );
dff a1_k0a_reg_19_ ( clk, n1500_r, a1_k0a[19], k0[115] );
not U_inv443 ( n1500_r, n1500 );
dff a1_out_1_reg_115_ ( clk, n1500_r, k1[115], k0b[115] );
not U_inv444 ( n689, k1[115] );
not U_inv445 ( n1500_r, n1500 );
dff a1_k0a_reg_20_ ( clk, n1499_r, a1_k0a[20], k0[116] );
not U_inv446 ( n1499_r, n1499 );
dff a1_out_1_reg_116_ ( clk, n1499_r, k1[116], k0b[116] );
not U_inv447 ( n691, k1[116] );
not U_inv448 ( n1499_r, n1499 );
dff a1_k0a_reg_21_ ( clk, n1499_r, a1_k0a[21], k0[117] );
not U_inv449 ( n1499_r, n1499 );
dff a1_out_1_reg_117_ ( clk, n1499_r, k1[117], k0b[117] );
not U_inv450 ( n692, k1[117] );
not U_inv451 ( n1499_r, n1499 );
dff a1_k0a_reg_22_ ( clk, n1499_r, a1_k0a[22], k0[118] );
not U_inv452 ( n1499_r, n1499 );
dff a1_out_1_reg_118_ ( clk, n1499_r, k1[118], k0b[118] );
not U_inv453 ( n693, k1[118] );
not U_inv454 ( n1499_r, n1499 );
dff a1_k0a_reg_23_ ( clk, n1499_r, a1_k0a[23], k0[119] );
not U_inv455 ( n1499_r, n1499 );
dff a1_out_1_reg_119_ ( clk, n1499_r, k1[119], k0b[119] );
not U_inv456 ( n694, k1[119] );
not U_inv457 ( n1499_r, n1499 );
dff a1_k0a_reg_24_ ( clk, n1499_r, a1_k0a[24], n1284 );
not U_inv458 ( n1499_r, n1499 );
dff a1_out_1_reg_120_ ( clk, n1499_r, k1[120], k0b[120] );
not U_inv459 ( n695, k1[120] );
not U_inv460 ( n1499_r, n1499 );
dff a1_k0a_reg_25_ ( clk, n1499_r, a1_k0a[25], k0[121] );
not U_inv461 ( n1499_r, n1499 );
dff a1_out_1_reg_121_ ( clk, n1499_r, ex_wire66, k0b[121] );
not U_inv462 ( n1285, ex_wire66 );
not U_inv463 ( n1499_r, n1499 );
dff a1_k0a_reg_26_ ( clk, n1498_r, a1_k0a[26], k0[122] );
not U_inv464 ( n1498_r, n1498 );
dff a1_out_1_reg_122_ ( clk, n1498_r, k1[122], k0b[122] );
not U_inv465 ( n696, k1[122] );
not U_inv466 ( n1498_r, n1498 );
dff a1_k0a_reg_27_ ( clk, n1498_r, a1_k0a[27], k0[123] );
not U_inv467 ( n1498_r, n1498 );
dff a1_out_1_reg_123_ ( clk, n1498_r, k1[123], k0b[123] );
not U_inv468 ( n697, k1[123] );
not U_inv469 ( n1498_r, n1498 );
dff a1_k0a_reg_28_ ( clk, n1498_r, a1_k0a[28], k0[124] );
not U_inv470 ( n1498_r, n1498 );
dff a1_out_1_reg_124_ ( clk, n1498_r, k1[124], k0b[124] );
not U_inv471 ( n698, k1[124] );
not U_inv472 ( n1498_r, n1498 );
dff a1_k0a_reg_29_ ( clk, n1498_r, a1_k0a[29], k0[125] );
not U_inv473 ( n1498_r, n1498 );
dff a1_out_1_reg_125_ ( clk, n1498_r, k1[125], k0b[125] );
not U_inv474 ( n699, k1[125] );
not U_inv475 ( n1498_r, n1498 );
dff a1_k0a_reg_30_ ( clk, n1498_r, a1_k0a[30], k0[126] );
not U_inv476 ( n1498_r, n1498 );
dff a1_out_1_reg_126_ ( clk, n1498_r, k1[126], k0b[126] );
not U_inv477 ( n701, k1[126] );
not U_inv478 ( n1498_r, n1498 );
dff a1_k0a_reg_31_ ( clk, n1498_r, a1_k0a[31], k0[127] );
not U_inv479 ( n1498_r, n1498 );
dff a1_out_1_reg_127_ ( clk, n1498_r, k1[127], k0b[127] );
not U_inv480 ( n702, k1[127] );
not U_inv481 ( n1498_r, n1498 );
dff a1_k3a_reg_0_ ( clk, n1497_r, a1_k3a[0], a1_v3[0] );
not U_inv482 ( n1497_r, n1497 );
dff a1_out_1_reg_0_ ( clk, n1497_r, k1[0], k0b[0] );
not U_inv483 ( n1497_r, n1497 );
dff a1_k3a_reg_1_ ( clk, n1497_r, a1_k3a[1], a1_v3[1] );
not U_inv484 ( n1497_r, n1497 );
dff a1_out_1_reg_1_ ( clk, n1497_r, k1[1], k0b[1] );
not U_inv485 ( n1497_r, n1497 );
dff a1_k3a_reg_2_ ( clk, n1497_r, a1_k3a[2], a1_v3[2] );
not U_inv486 ( n1497_r, n1497 );
dff a1_out_1_reg_2_ ( clk, n1497_r, k1[2], k0b[2] );
not U_inv487 ( n1497_r, n1497 );
dff a1_k3a_reg_3_ ( clk, n1497_r, a1_k3a[3], a1_v3[3] );
not U_inv488 ( n1497_r, n1497 );
dff a1_out_1_reg_3_ ( clk, n1497_r, k1[3], k0b[3] );
not U_inv489 ( n1497_r, n1497 );
dff a1_k3a_reg_4_ ( clk, n1497_r, a1_k3a[4], a1_v3[4] );
not U_inv490 ( n1497_r, n1497 );
dff a1_out_1_reg_4_ ( clk, n1497_r, k1[4], k0b[4] );
not U_inv491 ( n1497_r, n1497 );
dff a1_k3a_reg_5_ ( clk, n1497_r, a1_k3a[5], a1_v3[5] );
not U_inv492 ( n1497_r, n1497 );
dff a1_out_1_reg_5_ ( clk, n1497_r, k1[5], k0b[5] );
not U_inv493 ( n1497_r, n1497 );
dff a1_k3a_reg_6_ ( clk, n1496_r, a1_k3a[6], a1_v3[6] );
not U_inv494 ( n1496_r, n1496 );
dff a1_out_1_reg_6_ ( clk, n1496_r, k1[6], k0b[6] );
not U_inv495 ( n1496_r, n1496 );
dff a1_k3a_reg_7_ ( clk, n1496_r, a1_k3a[7], a1_v3[7] );
not U_inv496 ( n1496_r, n1496 );
dff a1_out_1_reg_7_ ( clk, n1496_r, k1[7], k0b[7] );
not U_inv497 ( n1496_r, n1496 );
dff a1_k3a_reg_8_ ( clk, n1496_r, a1_k3a[8], a1_v3[8] );
not U_inv498 ( n1496_r, n1496 );
dff a1_out_1_reg_8_ ( clk, n1496_r, k1[8], k0b[8] );
not U_inv499 ( n1496_r, n1496 );
dff a1_k3a_reg_9_ ( clk, n1496_r, a1_k3a[9], a1_v3[9] );
not U_inv500 ( n1496_r, n1496 );
dff a1_out_1_reg_9_ ( clk, n1496_r, k1[9], k0b[9] );
not U_inv501 ( n1496_r, n1496 );
dff a1_k3a_reg_10_ ( clk, n1496_r, a1_k3a[10], a1_v3[10] );
not U_inv502 ( n1496_r, n1496 );
dff a1_out_1_reg_10_ ( clk, n1496_r, k1[10], k0b[10] );
not U_inv503 ( n1496_r, n1496 );
dff a1_k3a_reg_11_ ( clk, n1496_r, a1_k3a[11], a1_v3[11] );
not U_inv504 ( n1496_r, n1496 );
dff a1_out_1_reg_11_ ( clk, n1496_r, k1[11], k0b[11] );
not U_inv505 ( n1496_r, n1496 );
dff a1_k3a_reg_12_ ( clk, n1495_r, a1_k3a[12], a1_v3[12] );
not U_inv506 ( n1495_r, n1495 );
dff a1_out_1_reg_12_ ( clk, n1495_r, k1[12], k0b[12] );
not U_inv507 ( n1495_r, n1495 );
dff a1_k3a_reg_13_ ( clk, n1495_r, a1_k3a[13], a1_v3[13] );
not U_inv508 ( n1495_r, n1495 );
dff a1_out_1_reg_13_ ( clk, n1495_r, k1[13], k0b[13] );
not U_inv509 ( n1495_r, n1495 );
dff a1_k3a_reg_14_ ( clk, n1495_r, a1_k3a[14], a1_v3[14] );
not U_inv510 ( n1495_r, n1495 );
dff a1_out_1_reg_14_ ( clk, n1495_r, k1[14], k0b[14] );
not U_inv511 ( n1495_r, n1495 );
dff a1_k3a_reg_15_ ( clk, n1495_r, a1_k3a[15], a1_v3[15] );
not U_inv512 ( n1495_r, n1495 );
dff a1_out_1_reg_15_ ( clk, n1495_r, k1[15], k0b[15] );
not U_inv513 ( n1495_r, n1495 );
dff a1_k3a_reg_16_ ( clk, n1495_r, a1_k3a[16], a1_v3[16] );
not U_inv514 ( n1495_r, n1495 );
dff a1_out_1_reg_16_ ( clk, n1495_r, k1[16], k0b[16] );
not U_inv515 ( n1495_r, n1495 );
dff a1_k3a_reg_17_ ( clk, n1495_r, a1_k3a[17], a1_v3[17] );
not U_inv516 ( n1495_r, n1495 );
dff a1_out_1_reg_17_ ( clk, n1495_r, k1[17], k0b[17] );
not U_inv517 ( n1495_r, n1495 );
dff a1_k3a_reg_18_ ( clk, n1494_r, a1_k3a[18], a1_v3[18] );
not U_inv518 ( n1494_r, n1494 );
dff a1_out_1_reg_18_ ( clk, n1494_r, k1[18], k0b[18] );
not U_inv519 ( n1494_r, n1494 );
dff a1_k3a_reg_19_ ( clk, n1494_r, a1_k3a[19], a1_v3[19] );
not U_inv520 ( n1494_r, n1494 );
dff a1_out_1_reg_19_ ( clk, n1494_r, k1[19], k0b[19] );
not U_inv521 ( n1494_r, n1494 );
dff a1_k3a_reg_20_ ( clk, n1494_r, a1_k3a[20], a1_v3[20] );
not U_inv522 ( n1494_r, n1494 );
dff a1_out_1_reg_20_ ( clk, n1494_r, k1[20], k0b[20] );
not U_inv523 ( n1494_r, n1494 );
dff a1_k3a_reg_21_ ( clk, n1494_r, a1_k3a[21], a1_v3[21] );
not U_inv524 ( n1494_r, n1494 );
dff a1_out_1_reg_21_ ( clk, n1494_r, k1[21], k0b[21] );
not U_inv525 ( n1494_r, n1494 );
dff a1_k3a_reg_22_ ( clk, n1494_r, a1_k3a[22], a1_v3[22] );
not U_inv526 ( n1494_r, n1494 );
dff a1_out_1_reg_22_ ( clk, n1494_r, k1[22], k0b[22] );
not U_inv527 ( n1494_r, n1494 );
dff a1_k3a_reg_23_ ( clk, n1494_r, a1_k3a[23], a1_v3[23] );
not U_inv528 ( n1494_r, n1494 );
dff a1_out_1_reg_23_ ( clk, n1494_r, k1[23], k0b[23] );
not U_inv529 ( n1494_r, n1494 );
dff a1_k3a_reg_24_ ( clk, n1493_r, a1_k3a[24], a1_v3[24] );
not U_inv530 ( n1493_r, n1493 );
dff a1_out_1_reg_24_ ( clk, n1493_r, k1[24], k0b[24] );
not U_inv531 ( n1493_r, n1493 );
dff a1_k3a_reg_25_ ( clk, n1493_r, a1_k3a[25], a1_v3[25] );
not U_inv532 ( n1493_r, n1493 );
dff a1_out_1_reg_25_ ( clk, n1493_r, k1[25], k0b[25] );
not U_inv533 ( n1493_r, n1493 );
dff a1_k3a_reg_26_ ( clk, n1493_r, a1_k3a[26], a1_v3[26] );
not U_inv534 ( n1493_r, n1493 );
dff a1_out_1_reg_26_ ( clk, n1493_r, k1[26], k0b[26] );
not U_inv535 ( n1493_r, n1493 );
dff a1_k3a_reg_27_ ( clk, n1493_r, a1_k3a[27], a1_v3[27] );
not U_inv536 ( n1493_r, n1493 );
dff a1_out_1_reg_27_ ( clk, n1493_r, k1[27], k0b[27] );
not U_inv537 ( n1493_r, n1493 );
dff a1_k3a_reg_28_ ( clk, n1493_r, a1_k3a[28], a1_v3[28] );
not U_inv538 ( n1493_r, n1493 );
dff a1_out_1_reg_28_ ( clk, n1493_r, k1[28], k0b[28] );
not U_inv539 ( n1493_r, n1493 );
dff a1_k3a_reg_29_ ( clk, n1493_r, a1_k3a[29], a1_v3[29] );
not U_inv540 ( n1493_r, n1493 );
dff a1_out_1_reg_29_ ( clk, n1493_r, k1[29], k0b[29] );
not U_inv541 ( n1493_r, n1493 );
dff a1_k3a_reg_30_ ( clk, n1492_r, a1_k3a[30], a1_v3[30] );
not U_inv542 ( n1492_r, n1492 );
dff a1_out_1_reg_30_ ( clk, n1492_r, k1[30], k0b[30] );
not U_inv543 ( n1492_r, n1492 );
dff a1_k2a_reg_0_ ( clk, n1492_r, a1_k2a[0], a1_v2[0] );
not U_inv544 ( n1492_r, n1492 );
dff a1_out_1_reg_32_ ( clk, n1492_r, k1[32], k0b[32] );
not U_inv545 ( n1492_r, n1492 );
dff a1_k2a_reg_1_ ( clk, n1492_r, a1_k2a[1], a1_v2[1] );
not U_inv546 ( n1492_r, n1492 );
dff a1_out_1_reg_33_ ( clk, n1492_r, k1[33], k0b[33] );
not U_inv547 ( n1492_r, n1492 );
dff a1_k2a_reg_2_ ( clk, n1492_r, a1_k2a[2], a1_v2[2] );
not U_inv548 ( n1492_r, n1492 );
dff a1_out_1_reg_34_ ( clk, n1492_r, k1[34], k0b[34] );
not U_inv549 ( n1492_r, n1492 );
dff a1_k2a_reg_3_ ( clk, n1492_r, a1_k2a[3], a1_v2[3] );
not U_inv550 ( n1492_r, n1492 );
dff a1_out_1_reg_35_ ( clk, n1492_r, k1[35], k0b[35] );
not U_inv551 ( n1492_r, n1492 );
dff a1_k2a_reg_4_ ( clk, n1492_r, a1_k2a[4], a1_v2[4] );
not U_inv552 ( n1492_r, n1492 );
dff a1_out_1_reg_36_ ( clk, n1492_r, k1[36], k0b[36] );
not U_inv553 ( n1492_r, n1492 );
dff a1_k2a_reg_5_ ( clk, n1491_r, a1_k2a[5], a1_v2[5] );
not U_inv554 ( n1491_r, n1491 );
dff a1_out_1_reg_37_ ( clk, n1491_r, k1[37], k0b[37] );
not U_inv555 ( n1491_r, n1491 );
dff a1_k2a_reg_6_ ( clk, n1491_r, a1_k2a[6], a1_v2[6] );
not U_inv556 ( n1491_r, n1491 );
dff a1_out_1_reg_38_ ( clk, n1491_r, k1[38], k0b[38] );
not U_inv557 ( n1491_r, n1491 );
dff a1_k2a_reg_7_ ( clk, n1491_r, a1_k2a[7], a1_v2[7] );
not U_inv558 ( n1491_r, n1491 );
dff a1_out_1_reg_39_ ( clk, n1491_r, k1[39], k0b[39] );
not U_inv559 ( n1491_r, n1491 );
dff a1_k2a_reg_8_ ( clk, n1491_r, a1_k2a[8], a1_v2[8] );
not U_inv560 ( n1491_r, n1491 );
dff a1_out_1_reg_40_ ( clk, n1491_r, k1[40], k0b[40] );
not U_inv561 ( n1491_r, n1491 );
dff a1_k2a_reg_9_ ( clk, n1491_r, a1_k2a[9], a1_v2[9] );
not U_inv562 ( n1491_r, n1491 );
dff a1_out_1_reg_41_ ( clk, n1491_r, k1[41], k0b[41] );
not U_inv563 ( n1491_r, n1491 );
dff a1_k2a_reg_10_ ( clk, n1491_r, a1_k2a[10], a1_v2[10] );
not U_inv564 ( n1491_r, n1491 );
dff a1_out_1_reg_42_ ( clk, n1491_r, k1[42], k0b[42] );
not U_inv565 ( n1491_r, n1491 );
dff a1_k2a_reg_11_ ( clk, n1490_r, a1_k2a[11], a1_v2[11] );
not U_inv566 ( n1490_r, n1490 );
dff a1_out_1_reg_43_ ( clk, n1490_r, k1[43], k0b[43] );
not U_inv567 ( n1490_r, n1490 );
dff a1_k2a_reg_12_ ( clk, n1490_r, a1_k2a[12], a1_v2[12] );
not U_inv568 ( n1490_r, n1490 );
dff a1_out_1_reg_44_ ( clk, n1490_r, k1[44], k0b[44] );
not U_inv569 ( n1490_r, n1490 );
dff a1_k2a_reg_13_ ( clk, n1490_r, a1_k2a[13], a1_v2[13] );
not U_inv570 ( n1490_r, n1490 );
dff a1_out_1_reg_45_ ( clk, n1490_r, k1[45], k0b[45] );
not U_inv571 ( n1490_r, n1490 );
dff a1_k2a_reg_14_ ( clk, n1490_r, a1_k2a[14], a1_v2[14] );
not U_inv572 ( n1490_r, n1490 );
dff a1_out_1_reg_46_ ( clk, n1490_r, k1[46], k0b[46] );
not U_inv573 ( n1490_r, n1490 );
dff a1_k2a_reg_15_ ( clk, n1490_r, a1_k2a[15], a1_v2[15] );
not U_inv574 ( n1490_r, n1490 );
dff a1_out_1_reg_47_ ( clk, n1490_r, k1[47], k0b[47] );
not U_inv575 ( n1490_r, n1490 );
dff a1_k2a_reg_16_ ( clk, n1490_r, a1_k2a[16], a1_v2[16] );
not U_inv576 ( n1490_r, n1490 );
dff a1_out_1_reg_48_ ( clk, n1490_r, k1[48], k0b[48] );
not U_inv577 ( n1490_r, n1490 );
dff a1_k2a_reg_17_ ( clk, n1489_r, a1_k2a[17], a1_v2[17] );
not U_inv578 ( n1489_r, n1489 );
dff a1_out_1_reg_49_ ( clk, n1489_r, k1[49], k0b[49] );
not U_inv579 ( n1489_r, n1489 );
dff a1_k2a_reg_18_ ( clk, n1489_r, a1_k2a[18], a1_v2[18] );
not U_inv580 ( n1489_r, n1489 );
dff a1_out_1_reg_50_ ( clk, n1489_r, k1[50], k0b[50] );
not U_inv581 ( n1489_r, n1489 );
dff a1_k2a_reg_19_ ( clk, n1489_r, a1_k2a[19], a1_v2[19] );
not U_inv582 ( n1489_r, n1489 );
dff a1_out_1_reg_51_ ( clk, n1489_r, k1[51], k0b[51] );
not U_inv583 ( n1489_r, n1489 );
dff a1_k2a_reg_20_ ( clk, n1489_r, a1_k2a[20], a1_v2[20] );
not U_inv584 ( n1489_r, n1489 );
dff a1_out_1_reg_52_ ( clk, n1489_r, k1[52], k0b[52] );
not U_inv585 ( n1489_r, n1489 );
dff a1_k2a_reg_21_ ( clk, n1489_r, a1_k2a[21], a1_v2[21] );
not U_inv586 ( n1489_r, n1489 );
dff a1_out_1_reg_53_ ( clk, n1489_r, k1[53], k0b[53] );
not U_inv587 ( n1489_r, n1489 );
dff a1_k2a_reg_22_ ( clk, n1489_r, a1_k2a[22], a1_v2[22] );
not U_inv588 ( n1489_r, n1489 );
dff a1_out_1_reg_54_ ( clk, n1489_r, k1[54], k0b[54] );
not U_inv589 ( n1489_r, n1489 );
dff a1_k2a_reg_23_ ( clk, n1488_r, a1_k2a[23], a1_v2[23] );
not U_inv590 ( n1488_r, n1488 );
dff a1_out_1_reg_55_ ( clk, n1488_r, k1[55], k0b[55] );
not U_inv591 ( n1488_r, n1488 );
dff a1_k2a_reg_24_ ( clk, n1488_r, a1_k2a[24], a1_v2[24] );
not U_inv592 ( n1488_r, n1488 );
dff a1_out_1_reg_56_ ( clk, n1488_r, k1[56], k0b[56] );
not U_inv593 ( n1488_r, n1488 );
dff a1_k2a_reg_25_ ( clk, n1488_r, a1_k2a[25], a1_v2[25] );
not U_inv594 ( n1488_r, n1488 );
dff a1_out_1_reg_57_ ( clk, n1488_r, k1[57], k0b[57] );
not U_inv595 ( n1488_r, n1488 );
dff a1_k2a_reg_26_ ( clk, n1488_r, a1_k2a[26], a1_v2[26] );
not U_inv596 ( n1488_r, n1488 );
dff a1_out_1_reg_58_ ( clk, n1488_r, k1[58], k0b[58] );
not U_inv597 ( n1488_r, n1488 );
dff a1_k2a_reg_27_ ( clk, n1488_r, a1_k2a[27], a1_v2[27] );
not U_inv598 ( n1488_r, n1488 );
dff a1_out_1_reg_59_ ( clk, n1488_r, k1[59], k0b[59] );
not U_inv599 ( n1488_r, n1488 );
dff a1_k2a_reg_28_ ( clk, n1488_r, a1_k2a[28], a1_v2[28] );
not U_inv600 ( n1488_r, n1488 );
dff a1_out_1_reg_60_ ( clk, n1488_r, k1[60], k0b[60] );
not U_inv601 ( n1488_r, n1488 );
dff a1_k2a_reg_29_ ( clk, n1487_r, a1_k2a[29], a1_v2[29] );
not U_inv602 ( n1487_r, n1487 );
dff a1_out_1_reg_61_ ( clk, n1487_r, k1[61], k0b[61] );
not U_inv603 ( n1487_r, n1487 );
dff a1_k2a_reg_30_ ( clk, n1487_r, a1_k2a[30], a1_v2[30] );
not U_inv604 ( n1487_r, n1487 );
dff a1_out_1_reg_62_ ( clk, n1487_r, k1[62], k0b[62] );
not U_inv605 ( n1487_r, n1487 );
dff a1_k2a_reg_31_ ( clk, n1487_r, a1_k2a[31], a1_v2[31] );
not U_inv606 ( n1487_r, n1487 );
dff a1_out_1_reg_63_ ( clk, n1487_r, k1[63], k0b[63] );
not U_inv607 ( n1487_r, n1487 );
dff a1_k1a_reg_0_ ( clk, n1487_r, a1_k1a[0], a1_v1[0] );
not U_inv608 ( n1487_r, n1487 );
dff a1_out_1_reg_64_ ( clk, n1487_r, ex_wire67, k0b[64] );
not U_inv609 ( n679, ex_wire67 );
not U_inv610 ( n1487_r, n1487 );
dff a1_k1a_reg_1_ ( clk, n1487_r, a1_k1a[1], a1_v1[1] );
not U_inv611 ( n1487_r, n1487 );
dff a1_out_1_reg_65_ ( clk, n1487_r, ex_wire68, k0b[65] );
not U_inv612 ( n690, ex_wire68 );
not U_inv613 ( n1487_r, n1487 );
dff a1_k1a_reg_2_ ( clk, n1487_r, a1_k1a[2], a1_v1[2] );
not U_inv614 ( n1487_r, n1487 );
dff a1_out_1_reg_66_ ( clk, n1487_r, ex_wire69, k0b[66] );
not U_inv615 ( n700, ex_wire69 );
not U_inv616 ( n1487_r, n1487 );
dff a1_k1a_reg_3_ ( clk, n1486_r, a1_k1a[3], a1_v1[3] );
not U_inv617 ( n1486_r, n1486 );
dff a1_out_1_reg_67_ ( clk, n1486_r, ex_wire70, k0b[67] );
not U_inv618 ( n703, ex_wire70 );
not U_inv619 ( n1486_r, n1486 );
dff a1_k1a_reg_4_ ( clk, n1486_r, a1_k1a[4], a1_v1[4] );
not U_inv620 ( n1486_r, n1486 );
dff a1_out_1_reg_68_ ( clk, n1486_r, k1[68], k0b[68] );
not U_inv621 ( n1486_r, n1486 );
dff a1_k1a_reg_5_ ( clk, n1486_r, a1_k1a[5], a1_v1[5] );
not U_inv622 ( n1486_r, n1486 );
dff a1_out_1_reg_69_ ( clk, n1486_r, k1[69], k0b[69] );
not U_inv623 ( n1486_r, n1486 );
dff a1_k1a_reg_6_ ( clk, n1486_r, a1_k1a[6], a1_v1[6] );
not U_inv624 ( n1486_r, n1486 );
dff a1_out_1_reg_70_ ( clk, n1486_r, k1[70], k0b[70] );
not U_inv625 ( n1486_r, n1486 );
dff a1_k1a_reg_7_ ( clk, n1486_r, a1_k1a[7], a1_v1[7] );
not U_inv626 ( n1486_r, n1486 );
dff a1_out_1_reg_71_ ( clk, n1486_r, k1[71], k0b[71] );
not U_inv627 ( n1486_r, n1486 );
dff a1_k1a_reg_8_ ( clk, n1486_r, a1_k1a[8], a1_v1[8] );
not U_inv628 ( n1486_r, n1486 );
dff a1_out_1_reg_72_ ( clk, n1486_r, k1[72], k0b[72] );
not U_inv629 ( n1486_r, n1486 );
dff a1_k1a_reg_9_ ( clk, n1485_r, a1_k1a[9], a1_v1[9] );
not U_inv630 ( n1485_r, n1485 );
dff a1_out_1_reg_73_ ( clk, n1485_r, k1[73], k0b[73] );
not U_inv631 ( n1485_r, n1485 );
dff a1_k1a_reg_10_ ( clk, n1485_r, a1_k1a[10], a1_v1[10] );
not U_inv632 ( n1485_r, n1485 );
dff a1_out_1_reg_74_ ( clk, n1485_r, k1[74], k0b[74] );
not U_inv633 ( n1485_r, n1485 );
dff a1_k1a_reg_11_ ( clk, n1485_r, a1_k1a[11], a1_v1[11] );
not U_inv634 ( n1485_r, n1485 );
dff a1_out_1_reg_75_ ( clk, n1485_r, k1[75], k0b[75] );
not U_inv635 ( n1485_r, n1485 );
dff a1_k1a_reg_12_ ( clk, n1485_r, a1_k1a[12], a1_v1[12] );
not U_inv636 ( n1485_r, n1485 );
dff a1_out_1_reg_76_ ( clk, n1485_r, k1[76], k0b[76] );
not U_inv637 ( n1485_r, n1485 );
dff a1_k1a_reg_13_ ( clk, n1485_r, a1_k1a[13], a1_v1[13] );
not U_inv638 ( n1485_r, n1485 );
dff a1_out_1_reg_77_ ( clk, n1485_r, k1[77], k0b[77] );
not U_inv639 ( n1485_r, n1485 );
dff a1_k1a_reg_14_ ( clk, n1485_r, a1_k1a[14], a1_v1[14] );
not U_inv640 ( n1485_r, n1485 );
dff a1_out_1_reg_78_ ( clk, n1485_r, k1[78], k0b[78] );
not U_inv641 ( n1485_r, n1485 );
dff a1_k1a_reg_15_ ( clk, n1484_r, a1_k1a[15], a1_v1[15] );
not U_inv642 ( n1484_r, n1484 );
dff a1_out_1_reg_79_ ( clk, n1484_r, k1[79], k0b[79] );
not U_inv643 ( n1484_r, n1484 );
dff a1_k1a_reg_16_ ( clk, n1484_r, a1_k1a[16], a1_v1[16] );
not U_inv644 ( n1484_r, n1484 );
dff a1_out_1_reg_80_ ( clk, n1484_r, k1[80], k0b[80] );
not U_inv645 ( n1484_r, n1484 );
dff a1_k1a_reg_17_ ( clk, n1484_r, a1_k1a[17], a1_v1[17] );
not U_inv646 ( n1484_r, n1484 );
dff a1_out_1_reg_81_ ( clk, n1484_r, k1[81], k0b[81] );
not U_inv647 ( n1484_r, n1484 );
dff a1_k1a_reg_18_ ( clk, n1484_r, a1_k1a[18], a1_v1[18] );
not U_inv648 ( n1484_r, n1484 );
dff a1_out_1_reg_82_ ( clk, n1484_r, k1[82], k0b[82] );
not U_inv649 ( n1484_r, n1484 );
dff a1_k1a_reg_19_ ( clk, n1484_r, a1_k1a[19], a1_v1[19] );
not U_inv650 ( n1484_r, n1484 );
dff a1_out_1_reg_83_ ( clk, n1484_r, k1[83], k0b[83] );
not U_inv651 ( n1484_r, n1484 );
dff a1_k1a_reg_20_ ( clk, n1484_r, a1_k1a[20], a1_v1[20] );
not U_inv652 ( n1484_r, n1484 );
dff a1_out_1_reg_84_ ( clk, n1484_r, k1[84], k0b[84] );
not U_inv653 ( n1484_r, n1484 );
dff a1_k1a_reg_21_ ( clk, n1483_r, a1_k1a[21], a1_v1[21] );
not U_inv654 ( n1483_r, n1483 );
dff a1_out_1_reg_85_ ( clk, n1483_r, k1[85], k0b[85] );
not U_inv655 ( n1483_r, n1483 );
dff a1_k1a_reg_22_ ( clk, n1483_r, a1_k1a[22], a1_v1[22] );
not U_inv656 ( n1483_r, n1483 );
dff a1_out_1_reg_86_ ( clk, n1483_r, k1[86], k0b[86] );
not U_inv657 ( n1483_r, n1483 );
dff a1_k1a_reg_23_ ( clk, n1483_r, a1_k1a[23], a1_v1[23] );
not U_inv658 ( n1483_r, n1483 );
dff a1_out_1_reg_87_ ( clk, n1483_r, k1[87], k0b[87] );
not U_inv659 ( n1483_r, n1483 );
dff a1_k1a_reg_24_ ( clk, n1483_r, a1_k1a[24], a1_v1[24] );
not U_inv660 ( n1483_r, n1483 );
dff a1_out_1_reg_88_ ( clk, n1483_r, k1[88], k0b[88] );
not U_inv661 ( n1483_r, n1483 );
dff a1_k1a_reg_25_ ( clk, n1483_r, a1_k1a[25], a1_v1[25] );
not U_inv662 ( n1483_r, n1483 );
dff a1_out_1_reg_89_ ( clk, n1483_r, k1[89], k0b[89] );
not U_inv663 ( n1483_r, n1483 );
dff a1_k1a_reg_26_ ( clk, n1483_r, a1_k1a[26], a1_v1[26] );
not U_inv664 ( n1483_r, n1483 );
dff a1_out_1_reg_90_ ( clk, n1483_r, k1[90], k0b[90] );
not U_inv665 ( n1483_r, n1483 );
dff a1_k1a_reg_27_ ( clk, n1482_r, a1_k1a[27], a1_v1[27] );
not U_inv666 ( n1482_r, n1482 );
dff a1_out_1_reg_91_ ( clk, n1482_r, k1[91], k0b[91] );
not U_inv667 ( n1482_r, n1482 );
dff a1_k1a_reg_28_ ( clk, n1482_r, a1_k1a[28], a1_v1[28] );
not U_inv668 ( n1482_r, n1482 );
dff a1_out_1_reg_92_ ( clk, n1482_r, k1[92], k0b[92] );
not U_inv669 ( n1482_r, n1482 );
dff a1_k1a_reg_29_ ( clk, n1482_r, a1_k1a[29], a1_v1[29] );
not U_inv670 ( n1482_r, n1482 );
dff a1_out_1_reg_93_ ( clk, n1482_r, k1[93], k0b[93] );
not U_inv671 ( n1482_r, n1482 );
dff a1_k1a_reg_30_ ( clk, n1482_r, a1_k1a[30], a1_v1[30] );
not U_inv672 ( n1482_r, n1482 );
dff a1_out_1_reg_94_ ( clk, n1482_r, k1[94], k0b[94] );
not U_inv673 ( n1482_r, n1482 );
dff a1_out_1_reg_95_ ( clk, n1482_r, k1[95], k0b[95] );
not U_inv674 ( n1482_r, n1482 );
dff a2_k0a_reg_0_ ( clk, n1482_r, a2_k0a[0], k1[96] );
not U_inv675 ( n1482_r, n1482 );
dff a2_out_1_reg_96_ ( clk, n1482_r, k2[96], k1b[96] );
not U_inv676 ( n1482_r, n1482 );
dff a2_k0a_reg_1_ ( clk, n1482_r, a2_k0a[1], k1[97] );
not U_inv677 ( n1482_r, n1482 );
dff a2_out_1_reg_97_ ( clk, n1481_r, k2[97], k1b[97] );
not U_inv678 ( n1481_r, n1481 );
dff a2_k0a_reg_2_ ( clk, n1481_r, a2_k0a[2], k1[98] );
not U_inv679 ( n1481_r, n1481 );
dff a2_out_1_reg_98_ ( clk, n1481_r, k2[98], k1b[98] );
not U_inv680 ( n1481_r, n1481 );
dff a2_k0a_reg_3_ ( clk, n1481_r, a2_k0a[3], k1[99] );
not U_inv681 ( n1481_r, n1481 );
dff a2_out_1_reg_99_ ( clk, n1481_r, k2[99], k1b[99] );
not U_inv682 ( n1481_r, n1481 );
dff a2_k0a_reg_4_ ( clk, n1481_r, a2_k0a[4], k1[100] );
not U_inv683 ( n1481_r, n1481 );
dff a2_out_1_reg_100_ ( clk, n1481_r, k2[100], k1b[100] );
not U_inv684 ( n735, k2[100] );
not U_inv685 ( n1481_r, n1481 );
dff a2_k0a_reg_5_ ( clk, n1481_r, a2_k0a[5], k1[101] );
not U_inv686 ( n1481_r, n1481 );
dff a2_out_1_reg_101_ ( clk, n1481_r, k2[101], k1b[101] );
not U_inv687 ( n736, k2[101] );
not U_inv688 ( n1481_r, n1481 );
dff a2_k0a_reg_6_ ( clk, n1481_r, a2_k0a[6], k1[102] );
not U_inv689 ( n1481_r, n1481 );
dff a2_out_1_reg_102_ ( clk, n1481_r, k2[102], k1b[102] );
not U_inv690 ( n737, k2[102] );
not U_inv691 ( n1481_r, n1481 );
dff a2_k0a_reg_7_ ( clk, n1481_r, a2_k0a[7], k1[103] );
not U_inv692 ( n1481_r, n1481 );
dff a2_out_1_reg_103_ ( clk, n1480_r, k2[103], k1b[103] );
not U_inv693 ( n738, k2[103] );
not U_inv694 ( n1480_r, n1480 );
dff a2_k0a_reg_8_ ( clk, n1480_r, a2_k0a[8], k1[104] );
not U_inv695 ( n1480_r, n1480 );
dff a2_out_1_reg_104_ ( clk, n1480_r, k2[104], k1b[104] );
not U_inv696 ( n739, k2[104] );
not U_inv697 ( n1480_r, n1480 );
dff a2_k0a_reg_9_ ( clk, n1480_r, a2_k0a[9], k1[105] );
not U_inv698 ( n1480_r, n1480 );
dff a2_out_1_reg_105_ ( clk, n1480_r, k2[105], k1b[105] );
not U_inv699 ( n740, k2[105] );
not U_inv700 ( n1480_r, n1480 );
dff a2_k0a_reg_10_ ( clk, n1480_r, a2_k0a[10], k1[106] );
not U_inv701 ( n1480_r, n1480 );
dff a2_out_1_reg_106_ ( clk, n1480_r, k2[106], k1b[106] );
not U_inv702 ( n711, k2[106] );
not U_inv703 ( n1480_r, n1480 );
dff a2_k0a_reg_11_ ( clk, n1480_r, a2_k0a[11], k1[107] );
not U_inv704 ( n1480_r, n1480 );
dff a2_out_1_reg_107_ ( clk, n1480_r, k2[107], k1b[107] );
not U_inv705 ( n712, k2[107] );
not U_inv706 ( n1480_r, n1480 );
dff a2_k0a_reg_12_ ( clk, n1480_r, a2_k0a[12], k1[108] );
not U_inv707 ( n1480_r, n1480 );
dff a2_out_1_reg_108_ ( clk, n1480_r, k2[108], k1b[108] );
not U_inv708 ( n713, k2[108] );
not U_inv709 ( n1480_r, n1480 );
dff a2_k0a_reg_13_ ( clk, n1480_r, a2_k0a[13], k1[109] );
not U_inv710 ( n1480_r, n1480 );
dff a2_out_1_reg_109_ ( clk, n1479_r, k2[109], k1b[109] );
not U_inv711 ( n714, k2[109] );
not U_inv712 ( n1479_r, n1479 );
dff a2_k0a_reg_14_ ( clk, n1479_r, a2_k0a[14], k1[110] );
not U_inv713 ( n1479_r, n1479 );
dff a2_out_1_reg_110_ ( clk, n1479_r, k2[110], k1b[110] );
not U_inv714 ( n715, k2[110] );
not U_inv715 ( n1479_r, n1479 );
dff a2_k0a_reg_15_ ( clk, n1479_r, a2_k0a[15], k1[111] );
not U_inv716 ( n1479_r, n1479 );
dff a2_out_1_reg_111_ ( clk, n1479_r, k2[111], k1b[111] );
not U_inv717 ( n716, k2[111] );
not U_inv718 ( n1479_r, n1479 );
dff a2_k0a_reg_16_ ( clk, n1479_r, a2_k0a[16], k1[112] );
not U_inv719 ( n1479_r, n1479 );
dff a2_out_1_reg_112_ ( clk, n1479_r, k2[112], k1b[112] );
not U_inv720 ( n717, k2[112] );
not U_inv721 ( n1479_r, n1479 );
dff a2_k0a_reg_17_ ( clk, n1479_r, a2_k0a[17], k1[113] );
not U_inv722 ( n1479_r, n1479 );
dff a2_out_1_reg_113_ ( clk, n1479_r, k2[113], k1b[113] );
not U_inv723 ( n718, k2[113] );
not U_inv724 ( n1479_r, n1479 );
dff a2_k0a_reg_18_ ( clk, n1479_r, a2_k0a[18], k1[114] );
not U_inv725 ( n1479_r, n1479 );
dff a2_out_1_reg_114_ ( clk, n1479_r, k2[114], k1b[114] );
not U_inv726 ( n719, k2[114] );
not U_inv727 ( n1479_r, n1479 );
dff a2_k0a_reg_19_ ( clk, n1479_r, a2_k0a[19], k1[115] );
not U_inv728 ( n1479_r, n1479 );
dff a2_out_1_reg_115_ ( clk, n1478_r, k2[115], k1b[115] );
not U_inv729 ( n720, k2[115] );
not U_inv730 ( n1478_r, n1478 );
dff a2_k0a_reg_20_ ( clk, n1478_r, a2_k0a[20], k1[116] );
not U_inv731 ( n1478_r, n1478 );
dff a2_out_1_reg_116_ ( clk, n1478_r, k2[116], k1b[116] );
not U_inv732 ( n722, k2[116] );
not U_inv733 ( n1478_r, n1478 );
dff a2_k0a_reg_21_ ( clk, n1478_r, a2_k0a[21], k1[117] );
not U_inv734 ( n1478_r, n1478 );
dff a2_out_1_reg_117_ ( clk, n1478_r, k2[117], k1b[117] );
not U_inv735 ( n723, k2[117] );
not U_inv736 ( n1478_r, n1478 );
dff a2_k0a_reg_22_ ( clk, n1478_r, a2_k0a[22], k1[118] );
not U_inv737 ( n1478_r, n1478 );
dff a2_out_1_reg_118_ ( clk, n1478_r, k2[118], k1b[118] );
not U_inv738 ( n724, k2[118] );
not U_inv739 ( n1478_r, n1478 );
dff a2_k0a_reg_23_ ( clk, n1478_r, a2_k0a[23], k1[119] );
not U_inv740 ( n1478_r, n1478 );
dff a2_out_1_reg_119_ ( clk, n1478_r, k2[119], k1b[119] );
not U_inv741 ( n725, k2[119] );
not U_inv742 ( n1478_r, n1478 );
dff a2_k0a_reg_24_ ( clk, n1478_r, a2_k0a[24], k1[120] );
not U_inv743 ( n1478_r, n1478 );
dff a2_out_1_reg_120_ ( clk, n1478_r, k2[120], k1b[120] );
not U_inv744 ( n726, k2[120] );
not U_inv745 ( n1478_r, n1478 );
dff a2_k0a_reg_25_ ( clk, n1478_r, a2_k0a[25], n1285 );
not U_inv746 ( n1478_r, n1478 );
dff a2_out_1_reg_121_ ( clk, n1477_r, k2[121], k1b[121] );
not U_inv747 ( n727, k2[121] );
not U_inv748 ( n1477_r, n1477 );
dff a2_k0a_reg_26_ ( clk, n1477_r, a2_k0a[26], k1[122] );
not U_inv749 ( n1477_r, n1477 );
dff a2_out_1_reg_122_ ( clk, n1477_r, ex_wire71, k1b[122] );
not U_inv750 ( n1286, ex_wire71 );
not U_inv751 ( n1477_r, n1477 );
dff a2_k0a_reg_27_ ( clk, n1477_r, a2_k0a[27], k1[123] );
not U_inv752 ( n1477_r, n1477 );
dff a2_out_1_reg_123_ ( clk, n1477_r, k2[123], k1b[123] );
not U_inv753 ( n728, k2[123] );
not U_inv754 ( n1477_r, n1477 );
dff a2_k0a_reg_28_ ( clk, n1477_r, a2_k0a[28], k1[124] );
not U_inv755 ( n1477_r, n1477 );
dff a2_out_1_reg_124_ ( clk, n1477_r, k2[124], k1b[124] );
not U_inv756 ( n729, k2[124] );
not U_inv757 ( n1477_r, n1477 );
dff a2_k0a_reg_29_ ( clk, n1477_r, a2_k0a[29], k1[125] );
not U_inv758 ( n1477_r, n1477 );
dff a2_out_1_reg_125_ ( clk, n1477_r, k2[125], k1b[125] );
not U_inv759 ( n730, k2[125] );
not U_inv760 ( n1477_r, n1477 );
dff a2_k0a_reg_30_ ( clk, n1477_r, a2_k0a[30], k1[126] );
not U_inv761 ( n1477_r, n1477 );
dff a2_out_1_reg_126_ ( clk, n1477_r, k2[126], k1b[126] );
not U_inv762 ( n732, k2[126] );
not U_inv763 ( n1477_r, n1477 );
dff a2_k0a_reg_31_ ( clk, n1477_r, a2_k0a[31], k1[127] );
not U_inv764 ( n1477_r, n1477 );
dff a2_out_1_reg_127_ ( clk, n1476_r, k2[127], k1b[127] );
not U_inv765 ( n733, k2[127] );
not U_inv766 ( n1476_r, n1476 );
dff a2_k3a_reg_0_ ( clk, n1476_r, a2_k3a[0], a2_v3[0] );
not U_inv767 ( n1476_r, n1476 );
dff a2_out_1_reg_0_ ( clk, n1476_r, k2[0], k1b[0] );
not U_inv768 ( n1476_r, n1476 );
dff a2_k3a_reg_1_ ( clk, n1476_r, a2_k3a[1], a2_v3[1] );
not U_inv769 ( n1476_r, n1476 );
dff a2_out_1_reg_1_ ( clk, n1476_r, k2[1], k1b[1] );
not U_inv770 ( n1476_r, n1476 );
dff a2_k3a_reg_2_ ( clk, n1476_r, a2_k3a[2], a2_v3[2] );
not U_inv771 ( n1476_r, n1476 );
dff a2_out_1_reg_2_ ( clk, n1476_r, k2[2], k1b[2] );
not U_inv772 ( n1476_r, n1476 );
dff a2_k3a_reg_3_ ( clk, n1476_r, a2_k3a[3], a2_v3[3] );
not U_inv773 ( n1476_r, n1476 );
dff a2_out_1_reg_3_ ( clk, n1476_r, k2[3], k1b[3] );
not U_inv774 ( n1476_r, n1476 );
dff a2_k3a_reg_4_ ( clk, n1476_r, a2_k3a[4], a2_v3[4] );
not U_inv775 ( n1476_r, n1476 );
dff a2_out_1_reg_4_ ( clk, n1476_r, k2[4], k1b[4] );
not U_inv776 ( n1476_r, n1476 );
dff a2_k3a_reg_5_ ( clk, n1476_r, a2_k3a[5], a2_v3[5] );
not U_inv777 ( n1476_r, n1476 );
dff a2_out_1_reg_5_ ( clk, n1475_r, k2[5], k1b[5] );
not U_inv778 ( n1475_r, n1475 );
dff a2_k3a_reg_6_ ( clk, n1475_r, a2_k3a[6], a2_v3[6] );
not U_inv779 ( n1475_r, n1475 );
dff a2_out_1_reg_6_ ( clk, n1475_r, k2[6], k1b[6] );
not U_inv780 ( n1475_r, n1475 );
dff a2_k3a_reg_7_ ( clk, n1475_r, a2_k3a[7], a2_v3[7] );
not U_inv781 ( n1475_r, n1475 );
dff a2_out_1_reg_7_ ( clk, n1475_r, k2[7], k1b[7] );
not U_inv782 ( n1475_r, n1475 );
dff a2_k3a_reg_8_ ( clk, n1475_r, a2_k3a[8], a2_v3[8] );
not U_inv783 ( n1475_r, n1475 );
dff a2_out_1_reg_8_ ( clk, n1475_r, k2[8], k1b[8] );
not U_inv784 ( n1475_r, n1475 );
dff a2_k3a_reg_9_ ( clk, n1475_r, a2_k3a[9], a2_v3[9] );
not U_inv785 ( n1475_r, n1475 );
dff a2_out_1_reg_9_ ( clk, n1475_r, k2[9], k1b[9] );
not U_inv786 ( n1475_r, n1475 );
dff a2_k3a_reg_10_ ( clk, n1475_r, a2_k3a[10], a2_v3[10] );
not U_inv787 ( n1475_r, n1475 );
dff a2_out_1_reg_10_ ( clk, n1475_r, k2[10], k1b[10] );
not U_inv788 ( n1475_r, n1475 );
dff a2_k3a_reg_11_ ( clk, n1475_r, a2_k3a[11], a2_v3[11] );
not U_inv789 ( n1475_r, n1475 );
dff a2_out_1_reg_11_ ( clk, n1474_r, k2[11], k1b[11] );
not U_inv790 ( n1474_r, n1474 );
dff a2_k3a_reg_12_ ( clk, n1474_r, a2_k3a[12], a2_v3[12] );
not U_inv791 ( n1474_r, n1474 );
dff a2_out_1_reg_12_ ( clk, n1474_r, k2[12], k1b[12] );
not U_inv792 ( n1474_r, n1474 );
dff a2_k3a_reg_13_ ( clk, n1474_r, a2_k3a[13], a2_v3[13] );
not U_inv793 ( n1474_r, n1474 );
dff a2_out_1_reg_13_ ( clk, n1474_r, k2[13], k1b[13] );
not U_inv794 ( n1474_r, n1474 );
dff a2_k3a_reg_14_ ( clk, n1474_r, a2_k3a[14], a2_v3[14] );
not U_inv795 ( n1474_r, n1474 );
dff a2_out_1_reg_14_ ( clk, n1474_r, k2[14], k1b[14] );
not U_inv796 ( n1474_r, n1474 );
dff a2_k3a_reg_15_ ( clk, n1474_r, a2_k3a[15], a2_v3[15] );
not U_inv797 ( n1474_r, n1474 );
dff a2_out_1_reg_15_ ( clk, n1474_r, k2[15], k1b[15] );
not U_inv798 ( n1474_r, n1474 );
dff a2_k3a_reg_16_ ( clk, n1474_r, a2_k3a[16], a2_v3[16] );
not U_inv799 ( n1474_r, n1474 );
dff a2_out_1_reg_16_ ( clk, n1474_r, k2[16], k1b[16] );
not U_inv800 ( n1474_r, n1474 );
dff a2_k3a_reg_17_ ( clk, n1474_r, a2_k3a[17], a2_v3[17] );
not U_inv801 ( n1474_r, n1474 );
dff a2_out_1_reg_17_ ( clk, n1473_r, k2[17], k1b[17] );
not U_inv802 ( n1473_r, n1473 );
dff a2_k3a_reg_18_ ( clk, n1473_r, a2_k3a[18], a2_v3[18] );
not U_inv803 ( n1473_r, n1473 );
dff a2_out_1_reg_18_ ( clk, n1473_r, k2[18], k1b[18] );
not U_inv804 ( n1473_r, n1473 );
dff a2_k3a_reg_19_ ( clk, n1473_r, a2_k3a[19], a2_v3[19] );
not U_inv805 ( n1473_r, n1473 );
dff a2_out_1_reg_19_ ( clk, n1473_r, k2[19], k1b[19] );
not U_inv806 ( n1473_r, n1473 );
dff a2_k3a_reg_20_ ( clk, n1473_r, a2_k3a[20], a2_v3[20] );
not U_inv807 ( n1473_r, n1473 );
dff a2_out_1_reg_20_ ( clk, n1473_r, k2[20], k1b[20] );
not U_inv808 ( n1473_r, n1473 );
dff a2_k3a_reg_21_ ( clk, n1473_r, a2_k3a[21], a2_v3[21] );
not U_inv809 ( n1473_r, n1473 );
dff a2_out_1_reg_21_ ( clk, n1473_r, k2[21], k1b[21] );
not U_inv810 ( n1473_r, n1473 );
dff a2_k3a_reg_22_ ( clk, n1473_r, a2_k3a[22], a2_v3[22] );
not U_inv811 ( n1473_r, n1473 );
dff a2_out_1_reg_22_ ( clk, n1473_r, k2[22], k1b[22] );
not U_inv812 ( n1473_r, n1473 );
dff a2_k3a_reg_23_ ( clk, n1473_r, a2_k3a[23], a2_v3[23] );
not U_inv813 ( n1473_r, n1473 );
dff a2_out_1_reg_23_ ( clk, n1472_r, k2[23], k1b[23] );
not U_inv814 ( n1472_r, n1472 );
dff a2_k3a_reg_24_ ( clk, n1472_r, a2_k3a[24], a2_v3[24] );
not U_inv815 ( n1472_r, n1472 );
dff a2_out_1_reg_24_ ( clk, n1472_r, k2[24], k1b[24] );
not U_inv816 ( n1472_r, n1472 );
dff a2_k3a_reg_25_ ( clk, n1472_r, a2_k3a[25], a2_v3[25] );
not U_inv817 ( n1472_r, n1472 );
dff a2_out_1_reg_25_ ( clk, n1472_r, k2[25], k1b[25] );
not U_inv818 ( n1472_r, n1472 );
dff a2_k3a_reg_26_ ( clk, n1472_r, a2_k3a[26], a2_v3[26] );
not U_inv819 ( n1472_r, n1472 );
dff a2_out_1_reg_26_ ( clk, n1472_r, k2[26], k1b[26] );
not U_inv820 ( n1472_r, n1472 );
dff a2_k3a_reg_27_ ( clk, n1472_r, a2_k3a[27], a2_v3[27] );
not U_inv821 ( n1472_r, n1472 );
dff a2_out_1_reg_27_ ( clk, n1472_r, k2[27], k1b[27] );
not U_inv822 ( n1472_r, n1472 );
dff a2_k3a_reg_28_ ( clk, n1472_r, a2_k3a[28], a2_v3[28] );
not U_inv823 ( n1472_r, n1472 );
dff a2_out_1_reg_28_ ( clk, n1472_r, k2[28], k1b[28] );
not U_inv824 ( n1472_r, n1472 );
dff a2_k3a_reg_29_ ( clk, n1472_r, a2_k3a[29], a2_v3[29] );
not U_inv825 ( n1472_r, n1472 );
dff a2_out_1_reg_29_ ( clk, n1471_r, k2[29], k1b[29] );
not U_inv826 ( n1471_r, n1471 );
dff a2_k3a_reg_30_ ( clk, n1471_r, a2_k3a[30], a2_v3[30] );
not U_inv827 ( n1471_r, n1471 );
dff a2_out_1_reg_30_ ( clk, n1471_r, k2[30], k1b[30] );
not U_inv828 ( n1471_r, n1471 );
dff a2_k2a_reg_0_ ( clk, n1471_r, a2_k2a[0], a2_v2[0] );
not U_inv829 ( n1471_r, n1471 );
dff a2_out_1_reg_32_ ( clk, n1471_r, k2[32], k1b[32] );
not U_inv830 ( n1471_r, n1471 );
dff a2_k2a_reg_1_ ( clk, n1471_r, a2_k2a[1], a2_v2[1] );
not U_inv831 ( n1471_r, n1471 );
dff a2_out_1_reg_33_ ( clk, n1471_r, k2[33], k1b[33] );
not U_inv832 ( n1471_r, n1471 );
dff a2_k2a_reg_2_ ( clk, n1471_r, a2_k2a[2], a2_v2[2] );
not U_inv833 ( n1471_r, n1471 );
dff a2_out_1_reg_34_ ( clk, n1471_r, k2[34], k1b[34] );
not U_inv834 ( n1471_r, n1471 );
dff a2_k2a_reg_3_ ( clk, n1471_r, a2_k2a[3], a2_v2[3] );
not U_inv835 ( n1471_r, n1471 );
dff a2_out_1_reg_35_ ( clk, n1471_r, k2[35], k1b[35] );
not U_inv836 ( n1471_r, n1471 );
dff a2_k2a_reg_4_ ( clk, n1471_r, a2_k2a[4], a2_v2[4] );
not U_inv837 ( n1471_r, n1471 );
dff a2_out_1_reg_36_ ( clk, n1470_r, k2[36], k1b[36] );
not U_inv838 ( n1470_r, n1470 );
dff a2_k2a_reg_5_ ( clk, n1470_r, a2_k2a[5], a2_v2[5] );
not U_inv839 ( n1470_r, n1470 );
dff a2_out_1_reg_37_ ( clk, n1470_r, k2[37], k1b[37] );
not U_inv840 ( n1470_r, n1470 );
dff a2_k2a_reg_6_ ( clk, n1470_r, a2_k2a[6], a2_v2[6] );
not U_inv841 ( n1470_r, n1470 );
dff a2_out_1_reg_38_ ( clk, n1470_r, k2[38], k1b[38] );
not U_inv842 ( n1470_r, n1470 );
dff a2_k2a_reg_7_ ( clk, n1470_r, a2_k2a[7], a2_v2[7] );
not U_inv843 ( n1470_r, n1470 );
dff a2_out_1_reg_39_ ( clk, n1470_r, k2[39], k1b[39] );
not U_inv844 ( n1470_r, n1470 );
dff a2_k2a_reg_8_ ( clk, n1470_r, a2_k2a[8], a2_v2[8] );
not U_inv845 ( n1470_r, n1470 );
dff a2_out_1_reg_40_ ( clk, n1470_r, k2[40], k1b[40] );
not U_inv846 ( n1470_r, n1470 );
dff a2_k2a_reg_9_ ( clk, n1470_r, a2_k2a[9], a2_v2[9] );
not U_inv847 ( n1470_r, n1470 );
dff a2_out_1_reg_41_ ( clk, n1470_r, k2[41], k1b[41] );
not U_inv848 ( n1470_r, n1470 );
dff a2_k2a_reg_10_ ( clk, n1470_r, a2_k2a[10], a2_v2[10] );
not U_inv849 ( n1470_r, n1470 );
dff a2_out_1_reg_42_ ( clk, n1469_r, k2[42], k1b[42] );
not U_inv850 ( n1469_r, n1469 );
dff a2_k2a_reg_11_ ( clk, n1469_r, a2_k2a[11], a2_v2[11] );
not U_inv851 ( n1469_r, n1469 );
dff a2_out_1_reg_43_ ( clk, n1469_r, k2[43], k1b[43] );
not U_inv852 ( n1469_r, n1469 );
dff a2_k2a_reg_12_ ( clk, n1469_r, a2_k2a[12], a2_v2[12] );
not U_inv853 ( n1469_r, n1469 );
dff a2_out_1_reg_44_ ( clk, n1469_r, k2[44], k1b[44] );
not U_inv854 ( n1469_r, n1469 );
dff a2_k2a_reg_13_ ( clk, n1469_r, a2_k2a[13], a2_v2[13] );
not U_inv855 ( n1469_r, n1469 );
dff a2_out_1_reg_45_ ( clk, n1469_r, k2[45], k1b[45] );
not U_inv856 ( n1469_r, n1469 );
dff a2_k2a_reg_14_ ( clk, n1469_r, a2_k2a[14], a2_v2[14] );
not U_inv857 ( n1469_r, n1469 );
dff a2_out_1_reg_46_ ( clk, n1469_r, k2[46], k1b[46] );
not U_inv858 ( n1469_r, n1469 );
dff a2_k2a_reg_15_ ( clk, n1469_r, a2_k2a[15], a2_v2[15] );
not U_inv859 ( n1469_r, n1469 );
dff a2_out_1_reg_47_ ( clk, n1469_r, k2[47], k1b[47] );
not U_inv860 ( n1469_r, n1469 );
dff a2_k2a_reg_16_ ( clk, n1469_r, a2_k2a[16], a2_v2[16] );
not U_inv861 ( n1469_r, n1469 );
dff a2_out_1_reg_48_ ( clk, n1468_r, k2[48], k1b[48] );
not U_inv862 ( n1468_r, n1468 );
dff a2_k2a_reg_17_ ( clk, n1468_r, a2_k2a[17], a2_v2[17] );
not U_inv863 ( n1468_r, n1468 );
dff a2_out_1_reg_49_ ( clk, n1468_r, k2[49], k1b[49] );
not U_inv864 ( n1468_r, n1468 );
dff a2_k2a_reg_18_ ( clk, n1468_r, a2_k2a[18], a2_v2[18] );
not U_inv865 ( n1468_r, n1468 );
dff a2_out_1_reg_50_ ( clk, n1468_r, k2[50], k1b[50] );
not U_inv866 ( n1468_r, n1468 );
dff a2_k2a_reg_19_ ( clk, n1468_r, a2_k2a[19], a2_v2[19] );
not U_inv867 ( n1468_r, n1468 );
dff a2_out_1_reg_51_ ( clk, n1468_r, k2[51], k1b[51] );
not U_inv868 ( n1468_r, n1468 );
dff a2_k2a_reg_20_ ( clk, n1468_r, a2_k2a[20], a2_v2[20] );
not U_inv869 ( n1468_r, n1468 );
dff a2_out_1_reg_52_ ( clk, n1468_r, k2[52], k1b[52] );
not U_inv870 ( n1468_r, n1468 );
dff a2_k2a_reg_21_ ( clk, n1468_r, a2_k2a[21], a2_v2[21] );
not U_inv871 ( n1468_r, n1468 );
dff a2_out_1_reg_53_ ( clk, n1468_r, k2[53], k1b[53] );
not U_inv872 ( n1468_r, n1468 );
dff a2_k2a_reg_22_ ( clk, n1468_r, a2_k2a[22], a2_v2[22] );
not U_inv873 ( n1468_r, n1468 );
dff a2_out_1_reg_54_ ( clk, n1467_r, k2[54], k1b[54] );
not U_inv874 ( n1467_r, n1467 );
dff a2_k2a_reg_23_ ( clk, n1467_r, a2_k2a[23], a2_v2[23] );
not U_inv875 ( n1467_r, n1467 );
dff a2_out_1_reg_55_ ( clk, n1467_r, k2[55], k1b[55] );
not U_inv876 ( n1467_r, n1467 );
dff a2_k2a_reg_24_ ( clk, n1467_r, a2_k2a[24], a2_v2[24] );
not U_inv877 ( n1467_r, n1467 );
dff a2_out_1_reg_56_ ( clk, n1467_r, k2[56], k1b[56] );
not U_inv878 ( n1467_r, n1467 );
dff a2_k2a_reg_25_ ( clk, n1467_r, a2_k2a[25], a2_v2[25] );
not U_inv879 ( n1467_r, n1467 );
dff a2_out_1_reg_57_ ( clk, n1467_r, k2[57], k1b[57] );
not U_inv880 ( n1467_r, n1467 );
dff a2_k2a_reg_26_ ( clk, n1467_r, a2_k2a[26], a2_v2[26] );
not U_inv881 ( n1467_r, n1467 );
dff a2_out_1_reg_58_ ( clk, n1467_r, k2[58], k1b[58] );
not U_inv882 ( n1467_r, n1467 );
dff a2_k2a_reg_27_ ( clk, n1467_r, a2_k2a[27], a2_v2[27] );
not U_inv883 ( n1467_r, n1467 );
dff a2_out_1_reg_59_ ( clk, n1467_r, k2[59], k1b[59] );
not U_inv884 ( n1467_r, n1467 );
dff a2_k2a_reg_28_ ( clk, n1467_r, a2_k2a[28], a2_v2[28] );
not U_inv885 ( n1467_r, n1467 );
dff a2_out_1_reg_60_ ( clk, n1466_r, k2[60], k1b[60] );
not U_inv886 ( n1466_r, n1466 );
dff a2_k2a_reg_29_ ( clk, n1466_r, a2_k2a[29], a2_v2[29] );
not U_inv887 ( n1466_r, n1466 );
dff a2_out_1_reg_61_ ( clk, n1466_r, k2[61], k1b[61] );
not U_inv888 ( n1466_r, n1466 );
dff a2_k2a_reg_30_ ( clk, n1466_r, a2_k2a[30], a2_v2[30] );
not U_inv889 ( n1466_r, n1466 );
dff a2_out_1_reg_62_ ( clk, n1466_r, k2[62], k1b[62] );
not U_inv890 ( n1466_r, n1466 );
dff a2_k2a_reg_31_ ( clk, n1466_r, a2_k2a[31], a2_v2[31] );
not U_inv891 ( n1466_r, n1466 );
dff a2_out_1_reg_63_ ( clk, n1466_r, k2[63], k1b[63] );
not U_inv892 ( n1466_r, n1466 );
dff a2_k1a_reg_0_ ( clk, n1466_r, a2_k1a[0], a2_v1[0] );
not U_inv893 ( n1466_r, n1466 );
dff a2_out_1_reg_64_ ( clk, n1466_r, ex_wire72, k1b[64] );
not U_inv894 ( n710, ex_wire72 );
not U_inv895 ( n1466_r, n1466 );
dff a2_k1a_reg_1_ ( clk, n1466_r, a2_k1a[1], a2_v1[1] );
not U_inv896 ( n1466_r, n1466 );
dff a2_out_1_reg_65_ ( clk, n1466_r, ex_wire73, k1b[65] );
not U_inv897 ( n721, ex_wire73 );
not U_inv898 ( n1466_r, n1466 );
dff a2_k1a_reg_2_ ( clk, n1466_r, a2_k1a[2], a2_v1[2] );
not U_inv899 ( n1466_r, n1466 );
dff a2_out_1_reg_66_ ( clk, n1465_r, ex_wire74, k1b[66] );
not U_inv900 ( n731, ex_wire74 );
not U_inv901 ( n1465_r, n1465 );
dff a2_k1a_reg_3_ ( clk, n1465_r, a2_k1a[3], a2_v1[3] );
not U_inv902 ( n1465_r, n1465 );
dff a2_out_1_reg_67_ ( clk, n1465_r, ex_wire75, k1b[67] );
not U_inv903 ( n734, ex_wire75 );
not U_inv904 ( n1465_r, n1465 );
dff a2_k1a_reg_4_ ( clk, n1465_r, a2_k1a[4], a2_v1[4] );
not U_inv905 ( n1465_r, n1465 );
dff a2_out_1_reg_68_ ( clk, n1465_r, k2[68], k1b[68] );
not U_inv906 ( n1465_r, n1465 );
dff a2_k1a_reg_5_ ( clk, n1465_r, a2_k1a[5], a2_v1[5] );
not U_inv907 ( n1465_r, n1465 );
dff a2_out_1_reg_69_ ( clk, n1465_r, k2[69], k1b[69] );
not U_inv908 ( n1465_r, n1465 );
dff a2_k1a_reg_6_ ( clk, n1465_r, a2_k1a[6], a2_v1[6] );
not U_inv909 ( n1465_r, n1465 );
dff a2_out_1_reg_70_ ( clk, n1465_r, k2[70], k1b[70] );
not U_inv910 ( n1465_r, n1465 );
dff a2_k1a_reg_7_ ( clk, n1465_r, a2_k1a[7], a2_v1[7] );
not U_inv911 ( n1465_r, n1465 );
dff a2_out_1_reg_71_ ( clk, n1465_r, k2[71], k1b[71] );
not U_inv912 ( n1465_r, n1465 );
dff a2_k1a_reg_8_ ( clk, n1465_r, a2_k1a[8], a2_v1[8] );
not U_inv913 ( n1465_r, n1465 );
dff a2_out_1_reg_72_ ( clk, n1464_r, k2[72], k1b[72] );
not U_inv914 ( n1464_r, n1464 );
dff a2_k1a_reg_9_ ( clk, n1464_r, a2_k1a[9], a2_v1[9] );
not U_inv915 ( n1464_r, n1464 );
dff a2_out_1_reg_73_ ( clk, n1464_r, k2[73], k1b[73] );
not U_inv916 ( n1464_r, n1464 );
dff a2_k1a_reg_10_ ( clk, n1464_r, a2_k1a[10], a2_v1[10] );
not U_inv917 ( n1464_r, n1464 );
dff a2_out_1_reg_74_ ( clk, n1464_r, k2[74], k1b[74] );
not U_inv918 ( n1464_r, n1464 );
dff a2_k1a_reg_11_ ( clk, n1464_r, a2_k1a[11], a2_v1[11] );
not U_inv919 ( n1464_r, n1464 );
dff a2_out_1_reg_75_ ( clk, n1464_r, k2[75], k1b[75] );
not U_inv920 ( n1464_r, n1464 );
dff a2_k1a_reg_12_ ( clk, n1464_r, a2_k1a[12], a2_v1[12] );
not U_inv921 ( n1464_r, n1464 );
dff a2_out_1_reg_76_ ( clk, n1464_r, k2[76], k1b[76] );
not U_inv922 ( n1464_r, n1464 );
dff a2_k1a_reg_13_ ( clk, n1464_r, a2_k1a[13], a2_v1[13] );
not U_inv923 ( n1464_r, n1464 );
dff a2_out_1_reg_77_ ( clk, n1464_r, k2[77], k1b[77] );
not U_inv924 ( n1464_r, n1464 );
dff a2_k1a_reg_14_ ( clk, n1464_r, a2_k1a[14], a2_v1[14] );
not U_inv925 ( n1464_r, n1464 );
dff a2_out_1_reg_78_ ( clk, n1463_r, k2[78], k1b[78] );
not U_inv926 ( n1463_r, n1463 );
dff a2_k1a_reg_15_ ( clk, n1463_r, a2_k1a[15], a2_v1[15] );
not U_inv927 ( n1463_r, n1463 );
dff a2_out_1_reg_79_ ( clk, n1463_r, k2[79], k1b[79] );
not U_inv928 ( n1463_r, n1463 );
dff a2_k1a_reg_16_ ( clk, n1463_r, a2_k1a[16], a2_v1[16] );
not U_inv929 ( n1463_r, n1463 );
dff a2_out_1_reg_80_ ( clk, n1463_r, k2[80], k1b[80] );
not U_inv930 ( n1463_r, n1463 );
dff a2_k1a_reg_17_ ( clk, n1463_r, a2_k1a[17], a2_v1[17] );
not U_inv931 ( n1463_r, n1463 );
dff a2_out_1_reg_81_ ( clk, n1463_r, k2[81], k1b[81] );
not U_inv932 ( n1463_r, n1463 );
dff a2_k1a_reg_18_ ( clk, n1463_r, a2_k1a[18], a2_v1[18] );
not U_inv933 ( n1463_r, n1463 );
dff a2_out_1_reg_82_ ( clk, n1463_r, k2[82], k1b[82] );
not U_inv934 ( n1463_r, n1463 );
dff a2_k1a_reg_19_ ( clk, n1463_r, a2_k1a[19], a2_v1[19] );
not U_inv935 ( n1463_r, n1463 );
dff a2_out_1_reg_83_ ( clk, n1463_r, k2[83], k1b[83] );
not U_inv936 ( n1463_r, n1463 );
dff a2_k1a_reg_20_ ( clk, n1463_r, a2_k1a[20], a2_v1[20] );
not U_inv937 ( n1463_r, n1463 );
dff a2_out_1_reg_84_ ( clk, n1462_r, k2[84], k1b[84] );
not U_inv938 ( n1462_r, n1462 );
dff a2_k1a_reg_21_ ( clk, n1462_r, a2_k1a[21], a2_v1[21] );
not U_inv939 ( n1462_r, n1462 );
dff a2_out_1_reg_85_ ( clk, n1462_r, k2[85], k1b[85] );
not U_inv940 ( n1462_r, n1462 );
dff a2_k1a_reg_22_ ( clk, n1462_r, a2_k1a[22], a2_v1[22] );
not U_inv941 ( n1462_r, n1462 );
dff a2_out_1_reg_86_ ( clk, n1462_r, k2[86], k1b[86] );
not U_inv942 ( n1462_r, n1462 );
dff a2_k1a_reg_23_ ( clk, n1462_r, a2_k1a[23], a2_v1[23] );
not U_inv943 ( n1462_r, n1462 );
dff a2_out_1_reg_87_ ( clk, n1462_r, k2[87], k1b[87] );
not U_inv944 ( n1462_r, n1462 );
dff a2_k1a_reg_24_ ( clk, n1462_r, a2_k1a[24], a2_v1[24] );
not U_inv945 ( n1462_r, n1462 );
dff a2_out_1_reg_88_ ( clk, n1462_r, k2[88], k1b[88] );
not U_inv946 ( n1462_r, n1462 );
dff a2_k1a_reg_25_ ( clk, n1462_r, a2_k1a[25], a2_v1[25] );
not U_inv947 ( n1462_r, n1462 );
dff a2_out_1_reg_89_ ( clk, n1462_r, k2[89], k1b[89] );
not U_inv948 ( n1462_r, n1462 );
dff a2_k1a_reg_26_ ( clk, n1462_r, a2_k1a[26], a2_v1[26] );
not U_inv949 ( n1462_r, n1462 );
dff a2_out_1_reg_90_ ( clk, n1461_r, k2[90], k1b[90] );
not U_inv950 ( n1461_r, n1461 );
dff a2_k1a_reg_27_ ( clk, n1461_r, a2_k1a[27], a2_v1[27] );
not U_inv951 ( n1461_r, n1461 );
dff a2_out_1_reg_91_ ( clk, n1461_r, k2[91], k1b[91] );
not U_inv952 ( n1461_r, n1461 );
dff a2_k1a_reg_28_ ( clk, n1461_r, a2_k1a[28], a2_v1[28] );
not U_inv953 ( n1461_r, n1461 );
dff a2_out_1_reg_92_ ( clk, n1461_r, k2[92], k1b[92] );
not U_inv954 ( n1461_r, n1461 );
dff a2_k1a_reg_29_ ( clk, n1461_r, a2_k1a[29], a2_v1[29] );
not U_inv955 ( n1461_r, n1461 );
dff a2_out_1_reg_93_ ( clk, n1461_r, k2[93], k1b[93] );
not U_inv956 ( n1461_r, n1461 );
dff a2_k1a_reg_30_ ( clk, n1461_r, a2_k1a[30], a2_v1[30] );
not U_inv957 ( n1461_r, n1461 );
dff a2_out_1_reg_94_ ( clk, n1461_r, k2[94], k1b[94] );
not U_inv958 ( n1461_r, n1461 );
dff a2_out_1_reg_95_ ( clk, n1461_r, k2[95], k1b[95] );
not U_inv959 ( n1461_r, n1461 );
dff a3_k0a_reg_0_ ( clk, n1461_r, a3_k0a[0], k2[96] );
not U_inv960 ( n1461_r, n1461 );
dff a3_out_1_reg_96_ ( clk, n1461_r, k3[96], k2b[96] );
not U_inv961 ( n1461_r, n1461 );
dff a3_k0a_reg_1_ ( clk, n1460_r, a3_k0a[1], k2[97] );
not U_inv962 ( n1460_r, n1460 );
dff a3_out_1_reg_97_ ( clk, n1460_r, k3[97], k2b[97] );
not U_inv963 ( n1460_r, n1460 );
dff a3_k0a_reg_2_ ( clk, n1460_r, a3_k0a[2], k2[98] );
not U_inv964 ( n1460_r, n1460 );
dff a3_out_1_reg_98_ ( clk, n1460_r, k3[98], k2b[98] );
not U_inv965 ( n1460_r, n1460 );
dff a3_k0a_reg_3_ ( clk, n1460_r, a3_k0a[3], k2[99] );
not U_inv966 ( n1460_r, n1460 );
dff a3_out_1_reg_99_ ( clk, n1460_r, k3[99], k2b[99] );
not U_inv967 ( n1460_r, n1460 );
dff a3_k0a_reg_4_ ( clk, n1460_r, a3_k0a[4], k2[100] );
not U_inv968 ( n1460_r, n1460 );
dff a3_out_1_reg_100_ ( clk, n1460_r, k3[100], k2b[100] );
not U_inv969 ( n766, k3[100] );
not U_inv970 ( n1460_r, n1460 );
dff a3_k0a_reg_5_ ( clk, n1460_r, a3_k0a[5], k2[101] );
not U_inv971 ( n1460_r, n1460 );
dff a3_out_1_reg_101_ ( clk, n1460_r, k3[101], k2b[101] );
not U_inv972 ( n767, k3[101] );
not U_inv973 ( n1460_r, n1460 );
dff a3_k0a_reg_6_ ( clk, n1460_r, a3_k0a[6], k2[102] );
not U_inv974 ( n1460_r, n1460 );
dff a3_out_1_reg_102_ ( clk, n1460_r, k3[102], k2b[102] );
not U_inv975 ( n768, k3[102] );
not U_inv976 ( n1460_r, n1460 );
dff a3_k0a_reg_7_ ( clk, n1459_r, a3_k0a[7], k2[103] );
not U_inv977 ( n1459_r, n1459 );
dff a3_out_1_reg_103_ ( clk, n1459_r, k3[103], k2b[103] );
not U_inv978 ( n769, k3[103] );
not U_inv979 ( n1459_r, n1459 );
dff a3_k0a_reg_8_ ( clk, n1459_r, a3_k0a[8], k2[104] );
not U_inv980 ( n1459_r, n1459 );
dff a3_out_1_reg_104_ ( clk, n1459_r, k3[104], k2b[104] );
not U_inv981 ( n770, k3[104] );
not U_inv982 ( n1459_r, n1459 );
dff a3_k0a_reg_9_ ( clk, n1459_r, a3_k0a[9], k2[105] );
not U_inv983 ( n1459_r, n1459 );
dff a3_out_1_reg_105_ ( clk, n1459_r, k3[105], k2b[105] );
not U_inv984 ( n771, k3[105] );
not U_inv985 ( n1459_r, n1459 );
dff a3_k0a_reg_10_ ( clk, n1459_r, a3_k0a[10], k2[106] );
not U_inv986 ( n1459_r, n1459 );
dff a3_out_1_reg_106_ ( clk, n1459_r, k3[106], k2b[106] );
not U_inv987 ( n742, k3[106] );
not U_inv988 ( n1459_r, n1459 );
dff a3_k0a_reg_11_ ( clk, n1459_r, a3_k0a[11], k2[107] );
not U_inv989 ( n1459_r, n1459 );
dff a3_out_1_reg_107_ ( clk, n1459_r, k3[107], k2b[107] );
not U_inv990 ( n743, k3[107] );
not U_inv991 ( n1459_r, n1459 );
dff a3_k0a_reg_12_ ( clk, n1459_r, a3_k0a[12], k2[108] );
not U_inv992 ( n1459_r, n1459 );
dff a3_out_1_reg_108_ ( clk, n1459_r, k3[108], k2b[108] );
not U_inv993 ( n744, k3[108] );
not U_inv994 ( n1459_r, n1459 );
dff a3_k0a_reg_13_ ( clk, n1458_r, a3_k0a[13], k2[109] );
not U_inv995 ( n1458_r, n1458 );
dff a3_out_1_reg_109_ ( clk, n1458_r, k3[109], k2b[109] );
not U_inv996 ( n745, k3[109] );
not U_inv997 ( n1458_r, n1458 );
dff a3_k0a_reg_14_ ( clk, n1458_r, a3_k0a[14], k2[110] );
not U_inv998 ( n1458_r, n1458 );
dff a3_out_1_reg_110_ ( clk, n1458_r, k3[110], k2b[110] );
not U_inv999 ( n746, k3[110] );
not U_inv1000 ( n1458_r, n1458 );
dff a3_k0a_reg_15_ ( clk, n1458_r, a3_k0a[15], k2[111] );
not U_inv1001 ( n1458_r, n1458 );
dff a3_out_1_reg_111_ ( clk, n1458_r, k3[111], k2b[111] );
not U_inv1002 ( n747, k3[111] );
not U_inv1003 ( n1458_r, n1458 );
dff a3_k0a_reg_16_ ( clk, n1458_r, a3_k0a[16], k2[112] );
not U_inv1004 ( n1458_r, n1458 );
dff a3_out_1_reg_112_ ( clk, n1458_r, k3[112], k2b[112] );
not U_inv1005 ( n748, k3[112] );
not U_inv1006 ( n1458_r, n1458 );
dff a3_k0a_reg_17_ ( clk, n1458_r, a3_k0a[17], k2[113] );
not U_inv1007 ( n1458_r, n1458 );
dff a3_out_1_reg_113_ ( clk, n1458_r, k3[113], k2b[113] );
not U_inv1008 ( n749, k3[113] );
not U_inv1009 ( n1458_r, n1458 );
dff a3_k0a_reg_18_ ( clk, n1458_r, a3_k0a[18], k2[114] );
not U_inv1010 ( n1458_r, n1458 );
dff a3_out_1_reg_114_ ( clk, n1458_r, k3[114], k2b[114] );
not U_inv1011 ( n750, k3[114] );
not U_inv1012 ( n1458_r, n1458 );
dff a3_k0a_reg_19_ ( clk, n1457_r, a3_k0a[19], k2[115] );
not U_inv1013 ( n1457_r, n1457 );
dff a3_out_1_reg_115_ ( clk, n1457_r, k3[115], k2b[115] );
not U_inv1014 ( n751, k3[115] );
not U_inv1015 ( n1457_r, n1457 );
dff a3_k0a_reg_20_ ( clk, n1457_r, a3_k0a[20], k2[116] );
not U_inv1016 ( n1457_r, n1457 );
dff a3_out_1_reg_116_ ( clk, n1457_r, k3[116], k2b[116] );
not U_inv1017 ( n753, k3[116] );
not U_inv1018 ( n1457_r, n1457 );
dff a3_k0a_reg_21_ ( clk, n1457_r, a3_k0a[21], k2[117] );
not U_inv1019 ( n1457_r, n1457 );
dff a3_out_1_reg_117_ ( clk, n1457_r, k3[117], k2b[117] );
not U_inv1020 ( n754, k3[117] );
not U_inv1021 ( n1457_r, n1457 );
dff a3_k0a_reg_22_ ( clk, n1457_r, a3_k0a[22], k2[118] );
not U_inv1022 ( n1457_r, n1457 );
dff a3_out_1_reg_118_ ( clk, n1457_r, k3[118], k2b[118] );
not U_inv1023 ( n755, k3[118] );
not U_inv1024 ( n1457_r, n1457 );
dff a3_k0a_reg_23_ ( clk, n1457_r, a3_k0a[23], k2[119] );
not U_inv1025 ( n1457_r, n1457 );
dff a3_out_1_reg_119_ ( clk, n1457_r, k3[119], k2b[119] );
not U_inv1026 ( n756, k3[119] );
not U_inv1027 ( n1457_r, n1457 );
dff a3_k0a_reg_24_ ( clk, n1457_r, a3_k0a[24], k2[120] );
not U_inv1028 ( n1457_r, n1457 );
dff a3_out_1_reg_120_ ( clk, n1457_r, k3[120], k2b[120] );
not U_inv1029 ( n757, k3[120] );
not U_inv1030 ( n1457_r, n1457 );
dff a3_k0a_reg_25_ ( clk, n1456_r, a3_k0a[25], k2[121] );
not U_inv1031 ( n1456_r, n1456 );
dff a3_out_1_reg_121_ ( clk, n1456_r, k3[121], k2b[121] );
not U_inv1032 ( n758, k3[121] );
not U_inv1033 ( n1456_r, n1456 );
dff a3_k0a_reg_26_ ( clk, n1456_r, a3_k0a[26], n1286 );
not U_inv1034 ( n1456_r, n1456 );
dff a3_out_1_reg_122_ ( clk, n1456_r, k3[122], k2b[122] );
not U_inv1035 ( n759, k3[122] );
not U_inv1036 ( n1456_r, n1456 );
dff a3_k0a_reg_27_ ( clk, n1456_r, a3_k0a[27], k2[123] );
not U_inv1037 ( n1456_r, n1456 );
dff a3_out_1_reg_123_ ( clk, n1456_r, ex_wire76, k2b[123] );
not U_inv1038 ( n1287, ex_wire76 );
not U_inv1039 ( n1456_r, n1456 );
dff a3_k0a_reg_28_ ( clk, n1456_r, a3_k0a[28], k2[124] );
not U_inv1040 ( n1456_r, n1456 );
dff a3_out_1_reg_124_ ( clk, n1456_r, k3[124], k2b[124] );
not U_inv1041 ( n760, k3[124] );
not U_inv1042 ( n1456_r, n1456 );
dff a3_k0a_reg_29_ ( clk, n1456_r, a3_k0a[29], k2[125] );
not U_inv1043 ( n1456_r, n1456 );
dff a3_out_1_reg_125_ ( clk, n1456_r, k3[125], k2b[125] );
not U_inv1044 ( n761, k3[125] );
not U_inv1045 ( n1456_r, n1456 );
dff a3_k0a_reg_30_ ( clk, n1456_r, a3_k0a[30], k2[126] );
not U_inv1046 ( n1456_r, n1456 );
dff a3_out_1_reg_126_ ( clk, n1456_r, k3[126], k2b[126] );
not U_inv1047 ( n763, k3[126] );
not U_inv1048 ( n1456_r, n1456 );
dff a3_k0a_reg_31_ ( clk, n1455_r, a3_k0a[31], k2[127] );
not U_inv1049 ( n1455_r, n1455 );
dff a3_out_1_reg_127_ ( clk, n1455_r, k3[127], k2b[127] );
not U_inv1050 ( n764, k3[127] );
not U_inv1051 ( n1455_r, n1455 );
dff a3_k3a_reg_0_ ( clk, n1455_r, a3_k3a[0], a3_v3[0] );
not U_inv1052 ( n1455_r, n1455 );
dff a3_out_1_reg_0_ ( clk, n1455_r, k3[0], k2b[0] );
not U_inv1053 ( n1455_r, n1455 );
dff a3_k3a_reg_1_ ( clk, n1455_r, a3_k3a[1], a3_v3[1] );
not U_inv1054 ( n1455_r, n1455 );
dff a3_out_1_reg_1_ ( clk, n1455_r, k3[1], k2b[1] );
not U_inv1055 ( n1455_r, n1455 );
dff a3_k3a_reg_2_ ( clk, n1455_r, a3_k3a[2], a3_v3[2] );
not U_inv1056 ( n1455_r, n1455 );
dff a3_out_1_reg_2_ ( clk, n1455_r, k3[2], k2b[2] );
not U_inv1057 ( n1455_r, n1455 );
dff a3_k3a_reg_3_ ( clk, n1455_r, a3_k3a[3], a3_v3[3] );
not U_inv1058 ( n1455_r, n1455 );
dff a3_out_1_reg_3_ ( clk, n1455_r, k3[3], k2b[3] );
not U_inv1059 ( n1455_r, n1455 );
dff a3_k3a_reg_4_ ( clk, n1455_r, a3_k3a[4], a3_v3[4] );
not U_inv1060 ( n1455_r, n1455 );
dff a3_out_1_reg_4_ ( clk, n1455_r, k3[4], k2b[4] );
not U_inv1061 ( n1455_r, n1455 );
dff a3_k3a_reg_5_ ( clk, n1454_r, a3_k3a[5], a3_v3[5] );
not U_inv1062 ( n1454_r, n1454 );
dff a3_out_1_reg_5_ ( clk, n1454_r, k3[5], k2b[5] );
not U_inv1063 ( n1454_r, n1454 );
dff a3_k3a_reg_6_ ( clk, n1454_r, a3_k3a[6], a3_v3[6] );
not U_inv1064 ( n1454_r, n1454 );
dff a3_out_1_reg_6_ ( clk, n1454_r, k3[6], k2b[6] );
not U_inv1065 ( n1454_r, n1454 );
dff a3_k3a_reg_7_ ( clk, n1454_r, a3_k3a[7], a3_v3[7] );
not U_inv1066 ( n1454_r, n1454 );
dff a3_out_1_reg_7_ ( clk, n1454_r, k3[7], k2b[7] );
not U_inv1067 ( n1454_r, n1454 );
dff a3_k3a_reg_8_ ( clk, n1454_r, a3_k3a[8], a3_v3[8] );
not U_inv1068 ( n1454_r, n1454 );
dff a3_out_1_reg_8_ ( clk, n1454_r, k3[8], k2b[8] );
not U_inv1069 ( n1454_r, n1454 );
dff a3_k3a_reg_9_ ( clk, n1454_r, a3_k3a[9], a3_v3[9] );
not U_inv1070 ( n1454_r, n1454 );
dff a3_out_1_reg_9_ ( clk, n1454_r, k3[9], k2b[9] );
not U_inv1071 ( n1454_r, n1454 );
dff a3_k3a_reg_10_ ( clk, n1454_r, a3_k3a[10], a3_v3[10] );
not U_inv1072 ( n1454_r, n1454 );
dff a3_out_1_reg_10_ ( clk, n1454_r, k3[10], k2b[10] );
not U_inv1073 ( n1454_r, n1454 );
dff a3_k3a_reg_11_ ( clk, n1453_r, a3_k3a[11], a3_v3[11] );
not U_inv1074 ( n1453_r, n1453 );
dff a3_out_1_reg_11_ ( clk, n1453_r, k3[11], k2b[11] );
not U_inv1075 ( n1453_r, n1453 );
dff a3_k3a_reg_12_ ( clk, n1453_r, a3_k3a[12], a3_v3[12] );
not U_inv1076 ( n1453_r, n1453 );
dff a3_out_1_reg_12_ ( clk, n1453_r, k3[12], k2b[12] );
not U_inv1077 ( n1453_r, n1453 );
dff a3_k3a_reg_13_ ( clk, n1453_r, a3_k3a[13], a3_v3[13] );
not U_inv1078 ( n1453_r, n1453 );
dff a3_out_1_reg_13_ ( clk, n1453_r, k3[13], k2b[13] );
not U_inv1079 ( n1453_r, n1453 );
dff a3_k3a_reg_14_ ( clk, n1453_r, a3_k3a[14], a3_v3[14] );
not U_inv1080 ( n1453_r, n1453 );
dff a3_out_1_reg_14_ ( clk, n1453_r, k3[14], k2b[14] );
not U_inv1081 ( n1453_r, n1453 );
dff a3_k3a_reg_15_ ( clk, n1453_r, a3_k3a[15], a3_v3[15] );
not U_inv1082 ( n1453_r, n1453 );
dff a3_out_1_reg_15_ ( clk, n1453_r, k3[15], k2b[15] );
not U_inv1083 ( n1453_r, n1453 );
dff a3_k3a_reg_16_ ( clk, n1453_r, a3_k3a[16], a3_v3[16] );
not U_inv1084 ( n1453_r, n1453 );
dff a3_out_1_reg_16_ ( clk, n1453_r, k3[16], k2b[16] );
not U_inv1085 ( n1453_r, n1453 );
dff a3_k3a_reg_17_ ( clk, n1452_r, a3_k3a[17], a3_v3[17] );
not U_inv1086 ( n1452_r, n1452 );
dff a3_out_1_reg_17_ ( clk, n1452_r, k3[17], k2b[17] );
not U_inv1087 ( n1452_r, n1452 );
dff a3_k3a_reg_18_ ( clk, n1452_r, a3_k3a[18], a3_v3[18] );
not U_inv1088 ( n1452_r, n1452 );
dff a3_out_1_reg_18_ ( clk, n1452_r, k3[18], k2b[18] );
not U_inv1089 ( n1452_r, n1452 );
dff a3_k3a_reg_19_ ( clk, n1452_r, a3_k3a[19], a3_v3[19] );
not U_inv1090 ( n1452_r, n1452 );
dff a3_out_1_reg_19_ ( clk, n1452_r, k3[19], k2b[19] );
not U_inv1091 ( n1452_r, n1452 );
dff a3_k3a_reg_20_ ( clk, n1452_r, a3_k3a[20], a3_v3[20] );
not U_inv1092 ( n1452_r, n1452 );
dff a3_out_1_reg_20_ ( clk, n1452_r, k3[20], k2b[20] );
not U_inv1093 ( n1452_r, n1452 );
dff a3_k3a_reg_21_ ( clk, n1452_r, a3_k3a[21], a3_v3[21] );
not U_inv1094 ( n1452_r, n1452 );
dff a3_out_1_reg_21_ ( clk, n1452_r, k3[21], k2b[21] );
not U_inv1095 ( n1452_r, n1452 );
dff a3_k3a_reg_22_ ( clk, n1452_r, a3_k3a[22], a3_v3[22] );
not U_inv1096 ( n1452_r, n1452 );
dff a3_out_1_reg_22_ ( clk, n1452_r, k3[22], k2b[22] );
not U_inv1097 ( n1452_r, n1452 );
dff a3_k3a_reg_23_ ( clk, n1451_r, a3_k3a[23], a3_v3[23] );
not U_inv1098 ( n1451_r, n1451 );
dff a3_out_1_reg_23_ ( clk, n1451_r, k3[23], k2b[23] );
not U_inv1099 ( n1451_r, n1451 );
dff a3_k3a_reg_24_ ( clk, n1451_r, a3_k3a[24], a3_v3[24] );
not U_inv1100 ( n1451_r, n1451 );
dff a3_out_1_reg_24_ ( clk, n1451_r, k3[24], k2b[24] );
not U_inv1101 ( n1451_r, n1451 );
dff a3_k3a_reg_25_ ( clk, n1451_r, a3_k3a[25], a3_v3[25] );
not U_inv1102 ( n1451_r, n1451 );
dff a3_out_1_reg_25_ ( clk, n1451_r, k3[25], k2b[25] );
not U_inv1103 ( n1451_r, n1451 );
dff a3_k3a_reg_26_ ( clk, n1451_r, a3_k3a[26], a3_v3[26] );
not U_inv1104 ( n1451_r, n1451 );
dff a3_out_1_reg_26_ ( clk, n1451_r, k3[26], k2b[26] );
not U_inv1105 ( n1451_r, n1451 );
dff a3_k3a_reg_27_ ( clk, n1451_r, a3_k3a[27], a3_v3[27] );
not U_inv1106 ( n1451_r, n1451 );
dff a3_out_1_reg_27_ ( clk, n1451_r, k3[27], k2b[27] );
not U_inv1107 ( n1451_r, n1451 );
dff a3_k3a_reg_28_ ( clk, n1451_r, a3_k3a[28], a3_v3[28] );
not U_inv1108 ( n1451_r, n1451 );
dff a3_out_1_reg_28_ ( clk, n1451_r, k3[28], k2b[28] );
not U_inv1109 ( n1451_r, n1451 );
dff a3_k3a_reg_29_ ( clk, n1450_r, a3_k3a[29], a3_v3[29] );
not U_inv1110 ( n1450_r, n1450 );
dff a3_out_1_reg_29_ ( clk, n1450_r, k3[29], k2b[29] );
not U_inv1111 ( n1450_r, n1450 );
dff a3_k3a_reg_30_ ( clk, n1450_r, a3_k3a[30], a3_v3[30] );
not U_inv1112 ( n1450_r, n1450 );
dff a3_out_1_reg_30_ ( clk, n1450_r, k3[30], k2b[30] );
not U_inv1113 ( n1450_r, n1450 );
dff a3_k2a_reg_0_ ( clk, n1450_r, a3_k2a[0], a3_v2[0] );
not U_inv1114 ( n1450_r, n1450 );
dff a3_out_1_reg_32_ ( clk, n1450_r, k3[32], k2b[32] );
not U_inv1115 ( n1450_r, n1450 );
dff a3_k2a_reg_1_ ( clk, n1450_r, a3_k2a[1], a3_v2[1] );
not U_inv1116 ( n1450_r, n1450 );
dff a3_out_1_reg_33_ ( clk, n1450_r, k3[33], k2b[33] );
not U_inv1117 ( n1450_r, n1450 );
dff a3_k2a_reg_2_ ( clk, n1450_r, a3_k2a[2], a3_v2[2] );
not U_inv1118 ( n1450_r, n1450 );
dff a3_out_1_reg_34_ ( clk, n1450_r, k3[34], k2b[34] );
not U_inv1119 ( n1450_r, n1450 );
dff a3_k2a_reg_3_ ( clk, n1450_r, a3_k2a[3], a3_v2[3] );
not U_inv1120 ( n1450_r, n1450 );
dff a3_out_1_reg_35_ ( clk, n1450_r, k3[35], k2b[35] );
not U_inv1121 ( n1450_r, n1450 );
dff a3_k2a_reg_4_ ( clk, n1449_r, a3_k2a[4], a3_v2[4] );
not U_inv1122 ( n1449_r, n1449 );
dff a3_out_1_reg_36_ ( clk, n1449_r, k3[36], k2b[36] );
not U_inv1123 ( n1449_r, n1449 );
dff a3_k2a_reg_5_ ( clk, n1449_r, a3_k2a[5], a3_v2[5] );
not U_inv1124 ( n1449_r, n1449 );
dff a3_out_1_reg_37_ ( clk, n1449_r, k3[37], k2b[37] );
not U_inv1125 ( n1449_r, n1449 );
dff a3_k2a_reg_6_ ( clk, n1449_r, a3_k2a[6], a3_v2[6] );
not U_inv1126 ( n1449_r, n1449 );
dff a3_out_1_reg_38_ ( clk, n1449_r, k3[38], k2b[38] );
not U_inv1127 ( n1449_r, n1449 );
dff a3_k2a_reg_7_ ( clk, n1449_r, a3_k2a[7], a3_v2[7] );
not U_inv1128 ( n1449_r, n1449 );
dff a3_out_1_reg_39_ ( clk, n1449_r, k3[39], k2b[39] );
not U_inv1129 ( n1449_r, n1449 );
dff a3_k2a_reg_8_ ( clk, n1449_r, a3_k2a[8], a3_v2[8] );
not U_inv1130 ( n1449_r, n1449 );
dff a3_out_1_reg_40_ ( clk, n1449_r, k3[40], k2b[40] );
not U_inv1131 ( n1449_r, n1449 );
dff a3_k2a_reg_9_ ( clk, n1449_r, a3_k2a[9], a3_v2[9] );
not U_inv1132 ( n1449_r, n1449 );
dff a3_out_1_reg_41_ ( clk, n1449_r, k3[41], k2b[41] );
not U_inv1133 ( n1449_r, n1449 );
dff a3_k2a_reg_10_ ( clk, n1448_r, a3_k2a[10], a3_v2[10] );
not U_inv1134 ( n1448_r, n1448 );
dff a3_out_1_reg_42_ ( clk, n1448_r, k3[42], k2b[42] );
not U_inv1135 ( n1448_r, n1448 );
dff a3_k2a_reg_11_ ( clk, n1448_r, a3_k2a[11], a3_v2[11] );
not U_inv1136 ( n1448_r, n1448 );
dff a3_out_1_reg_43_ ( clk, n1448_r, k3[43], k2b[43] );
not U_inv1137 ( n1448_r, n1448 );
dff a3_k2a_reg_12_ ( clk, n1448_r, a3_k2a[12], a3_v2[12] );
not U_inv1138 ( n1448_r, n1448 );
dff a3_out_1_reg_44_ ( clk, n1448_r, k3[44], k2b[44] );
not U_inv1139 ( n1448_r, n1448 );
dff a3_k2a_reg_13_ ( clk, n1448_r, a3_k2a[13], a3_v2[13] );
not U_inv1140 ( n1448_r, n1448 );
dff a3_out_1_reg_45_ ( clk, n1448_r, k3[45], k2b[45] );
not U_inv1141 ( n1448_r, n1448 );
dff a3_k2a_reg_14_ ( clk, n1448_r, a3_k2a[14], a3_v2[14] );
not U_inv1142 ( n1448_r, n1448 );
dff a3_out_1_reg_46_ ( clk, n1448_r, k3[46], k2b[46] );
not U_inv1143 ( n1448_r, n1448 );
dff a3_k2a_reg_15_ ( clk, n1448_r, a3_k2a[15], a3_v2[15] );
not U_inv1144 ( n1448_r, n1448 );
dff a3_out_1_reg_47_ ( clk, n1448_r, k3[47], k2b[47] );
not U_inv1145 ( n1448_r, n1448 );
dff a3_k2a_reg_16_ ( clk, n1447_r, a3_k2a[16], a3_v2[16] );
not U_inv1146 ( n1447_r, n1447 );
dff a3_out_1_reg_48_ ( clk, n1447_r, k3[48], k2b[48] );
not U_inv1147 ( n1447_r, n1447 );
dff a3_k2a_reg_17_ ( clk, n1447_r, a3_k2a[17], a3_v2[17] );
not U_inv1148 ( n1447_r, n1447 );
dff a3_out_1_reg_49_ ( clk, n1447_r, k3[49], k2b[49] );
not U_inv1149 ( n1447_r, n1447 );
dff a3_k2a_reg_18_ ( clk, n1447_r, a3_k2a[18], a3_v2[18] );
not U_inv1150 ( n1447_r, n1447 );
dff a3_out_1_reg_50_ ( clk, n1447_r, k3[50], k2b[50] );
not U_inv1151 ( n1447_r, n1447 );
dff a3_k2a_reg_19_ ( clk, n1447_r, a3_k2a[19], a3_v2[19] );
not U_inv1152 ( n1447_r, n1447 );
dff a3_out_1_reg_51_ ( clk, n1447_r, k3[51], k2b[51] );
not U_inv1153 ( n1447_r, n1447 );
dff a3_k2a_reg_20_ ( clk, n1447_r, a3_k2a[20], a3_v2[20] );
not U_inv1154 ( n1447_r, n1447 );
dff a3_out_1_reg_52_ ( clk, n1447_r, k3[52], k2b[52] );
not U_inv1155 ( n1447_r, n1447 );
dff a3_k2a_reg_21_ ( clk, n1447_r, a3_k2a[21], a3_v2[21] );
not U_inv1156 ( n1447_r, n1447 );
dff a3_out_1_reg_53_ ( clk, n1447_r, k3[53], k2b[53] );
not U_inv1157 ( n1447_r, n1447 );
dff a3_k2a_reg_22_ ( clk, n1446_r, a3_k2a[22], a3_v2[22] );
not U_inv1158 ( n1446_r, n1446 );
dff a3_out_1_reg_54_ ( clk, n1446_r, k3[54], k2b[54] );
not U_inv1159 ( n1446_r, n1446 );
dff a3_k2a_reg_23_ ( clk, n1446_r, a3_k2a[23], a3_v2[23] );
not U_inv1160 ( n1446_r, n1446 );
dff a3_out_1_reg_55_ ( clk, n1446_r, k3[55], k2b[55] );
not U_inv1161 ( n1446_r, n1446 );
dff a3_k2a_reg_24_ ( clk, n1446_r, a3_k2a[24], a3_v2[24] );
not U_inv1162 ( n1446_r, n1446 );
dff a3_out_1_reg_56_ ( clk, n1446_r, k3[56], k2b[56] );
not U_inv1163 ( n1446_r, n1446 );
dff a3_k2a_reg_25_ ( clk, n1446_r, a3_k2a[25], a3_v2[25] );
not U_inv1164 ( n1446_r, n1446 );
dff a3_out_1_reg_57_ ( clk, n1446_r, k3[57], k2b[57] );
not U_inv1165 ( n1446_r, n1446 );
dff a3_k2a_reg_26_ ( clk, n1446_r, a3_k2a[26], a3_v2[26] );
not U_inv1166 ( n1446_r, n1446 );
dff a3_out_1_reg_58_ ( clk, n1446_r, k3[58], k2b[58] );
not U_inv1167 ( n1446_r, n1446 );
dff a3_k2a_reg_27_ ( clk, n1446_r, a3_k2a[27], a3_v2[27] );
not U_inv1168 ( n1446_r, n1446 );
dff a3_out_1_reg_59_ ( clk, n1446_r, k3[59], k2b[59] );
not U_inv1169 ( n1446_r, n1446 );
dff a3_k2a_reg_28_ ( clk, n1445_r, a3_k2a[28], a3_v2[28] );
not U_inv1170 ( n1445_r, n1445 );
dff a3_out_1_reg_60_ ( clk, n1445_r, k3[60], k2b[60] );
not U_inv1171 ( n1445_r, n1445 );
dff a3_k2a_reg_29_ ( clk, n1445_r, a3_k2a[29], a3_v2[29] );
not U_inv1172 ( n1445_r, n1445 );
dff a3_out_1_reg_61_ ( clk, n1445_r, k3[61], k2b[61] );
not U_inv1173 ( n1445_r, n1445 );
dff a3_k2a_reg_30_ ( clk, n1445_r, a3_k2a[30], a3_v2[30] );
not U_inv1174 ( n1445_r, n1445 );
dff a3_out_1_reg_62_ ( clk, n1445_r, k3[62], k2b[62] );
not U_inv1175 ( n1445_r, n1445 );
dff a3_k2a_reg_31_ ( clk, n1445_r, a3_k2a[31], a3_v2[31] );
not U_inv1176 ( n1445_r, n1445 );
dff a3_out_1_reg_63_ ( clk, n1445_r, k3[63], k2b[63] );
not U_inv1177 ( n1445_r, n1445 );
dff a3_k1a_reg_0_ ( clk, n1445_r, a3_k1a[0], a3_v1[0] );
not U_inv1178 ( n1445_r, n1445 );
dff a3_out_1_reg_64_ ( clk, n1445_r, ex_wire77, k2b[64] );
not U_inv1179 ( n741, ex_wire77 );
not U_inv1180 ( n1445_r, n1445 );
dff a3_k1a_reg_1_ ( clk, n1445_r, a3_k1a[1], a3_v1[1] );
not U_inv1181 ( n1445_r, n1445 );
dff a3_out_1_reg_65_ ( clk, n1445_r, ex_wire78, k2b[65] );
not U_inv1182 ( n752, ex_wire78 );
not U_inv1183 ( n1445_r, n1445 );
dff a3_k1a_reg_2_ ( clk, n1444_r, a3_k1a[2], a3_v1[2] );
not U_inv1184 ( n1444_r, n1444 );
dff a3_out_1_reg_66_ ( clk, n1444_r, ex_wire79, k2b[66] );
not U_inv1185 ( n762, ex_wire79 );
not U_inv1186 ( n1444_r, n1444 );
dff a3_k1a_reg_3_ ( clk, n1444_r, a3_k1a[3], a3_v1[3] );
not U_inv1187 ( n1444_r, n1444 );
dff a3_out_1_reg_67_ ( clk, n1444_r, ex_wire80, k2b[67] );
not U_inv1188 ( n765, ex_wire80 );
not U_inv1189 ( n1444_r, n1444 );
dff a3_k1a_reg_4_ ( clk, n1444_r, a3_k1a[4], a3_v1[4] );
not U_inv1190 ( n1444_r, n1444 );
dff a3_out_1_reg_68_ ( clk, n1444_r, k3[68], k2b[68] );
not U_inv1191 ( n1444_r, n1444 );
dff a3_k1a_reg_5_ ( clk, n1444_r, a3_k1a[5], a3_v1[5] );
not U_inv1192 ( n1444_r, n1444 );
dff a3_out_1_reg_69_ ( clk, n1444_r, k3[69], k2b[69] );
not U_inv1193 ( n1444_r, n1444 );
dff a3_k1a_reg_6_ ( clk, n1444_r, a3_k1a[6], a3_v1[6] );
not U_inv1194 ( n1444_r, n1444 );
dff a3_out_1_reg_70_ ( clk, n1444_r, k3[70], k2b[70] );
not U_inv1195 ( n1444_r, n1444 );
dff a3_k1a_reg_7_ ( clk, n1444_r, a3_k1a[7], a3_v1[7] );
not U_inv1196 ( n1444_r, n1444 );
dff a3_out_1_reg_71_ ( clk, n1444_r, k3[71], k2b[71] );
not U_inv1197 ( n1444_r, n1444 );
dff a3_k1a_reg_8_ ( clk, n1443_r, a3_k1a[8], a3_v1[8] );
not U_inv1198 ( n1443_r, n1443 );
dff a3_out_1_reg_72_ ( clk, n1443_r, k3[72], k2b[72] );
not U_inv1199 ( n1443_r, n1443 );
dff a3_k1a_reg_9_ ( clk, n1443_r, a3_k1a[9], a3_v1[9] );
not U_inv1200 ( n1443_r, n1443 );
dff a3_out_1_reg_73_ ( clk, n1443_r, k3[73], k2b[73] );
not U_inv1201 ( n1443_r, n1443 );
dff a3_k1a_reg_10_ ( clk, n1443_r, a3_k1a[10], a3_v1[10] );
not U_inv1202 ( n1443_r, n1443 );
dff a3_out_1_reg_74_ ( clk, n1443_r, k3[74], k2b[74] );
not U_inv1203 ( n1443_r, n1443 );
dff a3_k1a_reg_11_ ( clk, n1443_r, a3_k1a[11], a3_v1[11] );
not U_inv1204 ( n1443_r, n1443 );
dff a3_out_1_reg_75_ ( clk, n1443_r, k3[75], k2b[75] );
not U_inv1205 ( n1443_r, n1443 );
dff a3_k1a_reg_12_ ( clk, n1443_r, a3_k1a[12], a3_v1[12] );
not U_inv1206 ( n1443_r, n1443 );
dff a3_out_1_reg_76_ ( clk, n1443_r, k3[76], k2b[76] );
not U_inv1207 ( n1443_r, n1443 );
dff a3_k1a_reg_13_ ( clk, n1443_r, a3_k1a[13], a3_v1[13] );
not U_inv1208 ( n1443_r, n1443 );
dff a3_out_1_reg_77_ ( clk, n1443_r, k3[77], k2b[77] );
not U_inv1209 ( n1443_r, n1443 );
dff a3_k1a_reg_14_ ( clk, n1442_r, a3_k1a[14], a3_v1[14] );
not U_inv1210 ( n1442_r, n1442 );
dff a3_out_1_reg_78_ ( clk, n1442_r, k3[78], k2b[78] );
not U_inv1211 ( n1442_r, n1442 );
dff a3_k1a_reg_15_ ( clk, n1442_r, a3_k1a[15], a3_v1[15] );
not U_inv1212 ( n1442_r, n1442 );
dff a3_out_1_reg_79_ ( clk, n1442_r, k3[79], k2b[79] );
not U_inv1213 ( n1442_r, n1442 );
dff a3_k1a_reg_16_ ( clk, n1442_r, a3_k1a[16], a3_v1[16] );
not U_inv1214 ( n1442_r, n1442 );
dff a3_out_1_reg_80_ ( clk, n1442_r, k3[80], k2b[80] );
not U_inv1215 ( n1442_r, n1442 );
dff a3_k1a_reg_17_ ( clk, n1442_r, a3_k1a[17], a3_v1[17] );
not U_inv1216 ( n1442_r, n1442 );
dff a3_out_1_reg_81_ ( clk, n1442_r, k3[81], k2b[81] );
not U_inv1217 ( n1442_r, n1442 );
dff a3_k1a_reg_18_ ( clk, n1442_r, a3_k1a[18], a3_v1[18] );
not U_inv1218 ( n1442_r, n1442 );
dff a3_out_1_reg_82_ ( clk, n1442_r, k3[82], k2b[82] );
not U_inv1219 ( n1442_r, n1442 );
dff a3_k1a_reg_19_ ( clk, n1442_r, a3_k1a[19], a3_v1[19] );
not U_inv1220 ( n1442_r, n1442 );
dff a3_out_1_reg_83_ ( clk, n1442_r, k3[83], k2b[83] );
not U_inv1221 ( n1442_r, n1442 );
dff a3_k1a_reg_20_ ( clk, n1441_r, a3_k1a[20], a3_v1[20] );
not U_inv1222 ( n1441_r, n1441 );
dff a3_out_1_reg_84_ ( clk, n1441_r, k3[84], k2b[84] );
not U_inv1223 ( n1441_r, n1441 );
dff a3_k1a_reg_21_ ( clk, n1441_r, a3_k1a[21], a3_v1[21] );
not U_inv1224 ( n1441_r, n1441 );
dff a3_out_1_reg_85_ ( clk, n1441_r, k3[85], k2b[85] );
not U_inv1225 ( n1441_r, n1441 );
dff a3_k1a_reg_22_ ( clk, n1441_r, a3_k1a[22], a3_v1[22] );
not U_inv1226 ( n1441_r, n1441 );
dff a3_out_1_reg_86_ ( clk, n1441_r, k3[86], k2b[86] );
not U_inv1227 ( n1441_r, n1441 );
dff a3_k1a_reg_23_ ( clk, n1441_r, a3_k1a[23], a3_v1[23] );
not U_inv1228 ( n1441_r, n1441 );
dff a3_out_1_reg_87_ ( clk, n1441_r, k3[87], k2b[87] );
not U_inv1229 ( n1441_r, n1441 );
dff a3_k1a_reg_24_ ( clk, n1441_r, a3_k1a[24], a3_v1[24] );
not U_inv1230 ( n1441_r, n1441 );
dff a3_out_1_reg_88_ ( clk, n1441_r, k3[88], k2b[88] );
not U_inv1231 ( n1441_r, n1441 );
dff a3_k1a_reg_25_ ( clk, n1441_r, a3_k1a[25], a3_v1[25] );
not U_inv1232 ( n1441_r, n1441 );
dff a3_out_1_reg_89_ ( clk, n1441_r, k3[89], k2b[89] );
not U_inv1233 ( n1441_r, n1441 );
dff a3_k1a_reg_26_ ( clk, n1440_r, a3_k1a[26], a3_v1[26] );
not U_inv1234 ( n1440_r, n1440 );
dff a3_out_1_reg_90_ ( clk, n1440_r, k3[90], k2b[90] );
not U_inv1235 ( n1440_r, n1440 );
dff a3_k1a_reg_27_ ( clk, n1440_r, a3_k1a[27], a3_v1[27] );
not U_inv1236 ( n1440_r, n1440 );
dff a3_out_1_reg_91_ ( clk, n1440_r, k3[91], k2b[91] );
not U_inv1237 ( n1440_r, n1440 );
dff a3_k1a_reg_28_ ( clk, n1440_r, a3_k1a[28], a3_v1[28] );
not U_inv1238 ( n1440_r, n1440 );
dff a3_out_1_reg_92_ ( clk, n1440_r, k3[92], k2b[92] );
not U_inv1239 ( n1440_r, n1440 );
dff a3_k1a_reg_29_ ( clk, n1440_r, a3_k1a[29], a3_v1[29] );
not U_inv1240 ( n1440_r, n1440 );
dff a3_out_1_reg_93_ ( clk, n1440_r, k3[93], k2b[93] );
not U_inv1241 ( n1440_r, n1440 );
dff a3_k1a_reg_30_ ( clk, n1440_r, a3_k1a[30], a3_v1[30] );
not U_inv1242 ( n1440_r, n1440 );
dff a3_out_1_reg_94_ ( clk, n1440_r, k3[94], k2b[94] );
not U_inv1243 ( n1440_r, n1440 );
dff a3_out_1_reg_95_ ( clk, n1440_r, k3[95], k2b[95] );
not U_inv1244 ( n1440_r, n1440 );
dff a4_k0a_reg_0_ ( clk, n1440_r, a4_k0a[0], k3[96] );
not U_inv1245 ( n1440_r, n1440 );
dff a4_out_1_reg_96_ ( clk, n1439_r, k4[96], k3b[96] );
not U_inv1246 ( n1439_r, n1439 );
dff a4_k0a_reg_1_ ( clk, n1439_r, a4_k0a[1], k3[97] );
not U_inv1247 ( n1439_r, n1439 );
dff a4_out_1_reg_97_ ( clk, n1439_r, k4[97], k3b[97] );
not U_inv1248 ( n1439_r, n1439 );
dff a4_k0a_reg_2_ ( clk, n1439_r, a4_k0a[2], k3[98] );
not U_inv1249 ( n1439_r, n1439 );
dff a4_out_1_reg_98_ ( clk, n1439_r, k4[98], k3b[98] );
not U_inv1250 ( n1439_r, n1439 );
dff a4_k0a_reg_3_ ( clk, n1439_r, a4_k0a[3], k3[99] );
not U_inv1251 ( n1439_r, n1439 );
dff a4_out_1_reg_99_ ( clk, n1439_r, k4[99], k3b[99] );
not U_inv1252 ( n1439_r, n1439 );
dff a4_k0a_reg_4_ ( clk, n1439_r, a4_k0a[4], k3[100] );
not U_inv1253 ( n1439_r, n1439 );
dff a4_out_1_reg_100_ ( clk, n1439_r, k4[100], k3b[100] );
not U_inv1254 ( n797, k4[100] );
not U_inv1255 ( n1439_r, n1439 );
dff a4_k0a_reg_5_ ( clk, n1439_r, a4_k0a[5], k3[101] );
not U_inv1256 ( n1439_r, n1439 );
dff a4_out_1_reg_101_ ( clk, n1439_r, k4[101], k3b[101] );
not U_inv1257 ( n798, k4[101] );
not U_inv1258 ( n1439_r, n1439 );
dff a4_k0a_reg_6_ ( clk, n1439_r, a4_k0a[6], k3[102] );
not U_inv1259 ( n1439_r, n1439 );
dff a4_out_1_reg_102_ ( clk, n1438_r, k4[102], k3b[102] );
not U_inv1260 ( n799, k4[102] );
not U_inv1261 ( n1438_r, n1438 );
dff a4_k0a_reg_7_ ( clk, n1438_r, a4_k0a[7], k3[103] );
not U_inv1262 ( n1438_r, n1438 );
dff a4_out_1_reg_103_ ( clk, n1438_r, k4[103], k3b[103] );
not U_inv1263 ( n800, k4[103] );
not U_inv1264 ( n1438_r, n1438 );
dff a4_k0a_reg_8_ ( clk, n1438_r, a4_k0a[8], k3[104] );
not U_inv1265 ( n1438_r, n1438 );
dff a4_out_1_reg_104_ ( clk, n1438_r, k4[104], k3b[104] );
not U_inv1266 ( n801, k4[104] );
not U_inv1267 ( n1438_r, n1438 );
dff a4_k0a_reg_9_ ( clk, n1438_r, a4_k0a[9], k3[105] );
not U_inv1268 ( n1438_r, n1438 );
dff a4_out_1_reg_105_ ( clk, n1438_r, k4[105], k3b[105] );
not U_inv1269 ( n802, k4[105] );
not U_inv1270 ( n1438_r, n1438 );
dff a4_k0a_reg_10_ ( clk, n1438_r, a4_k0a[10], k3[106] );
not U_inv1271 ( n1438_r, n1438 );
dff a4_out_1_reg_106_ ( clk, n1438_r, k4[106], k3b[106] );
not U_inv1272 ( n773, k4[106] );
not U_inv1273 ( n1438_r, n1438 );
dff a4_k0a_reg_11_ ( clk, n1438_r, a4_k0a[11], k3[107] );
not U_inv1274 ( n1438_r, n1438 );
dff a4_out_1_reg_107_ ( clk, n1438_r, k4[107], k3b[107] );
not U_inv1275 ( n774, k4[107] );
not U_inv1276 ( n1438_r, n1438 );
dff a4_k0a_reg_12_ ( clk, n1438_r, a4_k0a[12], k3[108] );
not U_inv1277 ( n1438_r, n1438 );
dff a4_out_1_reg_108_ ( clk, n1437_r, k4[108], k3b[108] );
not U_inv1278 ( n775, k4[108] );
not U_inv1279 ( n1437_r, n1437 );
dff a4_k0a_reg_13_ ( clk, n1437_r, a4_k0a[13], k3[109] );
not U_inv1280 ( n1437_r, n1437 );
dff a4_out_1_reg_109_ ( clk, n1437_r, k4[109], k3b[109] );
not U_inv1281 ( n776, k4[109] );
not U_inv1282 ( n1437_r, n1437 );
dff a4_k0a_reg_14_ ( clk, n1437_r, a4_k0a[14], k3[110] );
not U_inv1283 ( n1437_r, n1437 );
dff a4_out_1_reg_110_ ( clk, n1437_r, k4[110], k3b[110] );
not U_inv1284 ( n777, k4[110] );
not U_inv1285 ( n1437_r, n1437 );
dff a4_k0a_reg_15_ ( clk, n1437_r, a4_k0a[15], k3[111] );
not U_inv1286 ( n1437_r, n1437 );
dff a4_out_1_reg_111_ ( clk, n1437_r, k4[111], k3b[111] );
not U_inv1287 ( n778, k4[111] );
not U_inv1288 ( n1437_r, n1437 );
dff a4_k0a_reg_16_ ( clk, n1437_r, a4_k0a[16], k3[112] );
not U_inv1289 ( n1437_r, n1437 );
dff a4_out_1_reg_112_ ( clk, n1437_r, k4[112], k3b[112] );
not U_inv1290 ( n779, k4[112] );
not U_inv1291 ( n1437_r, n1437 );
dff a4_k0a_reg_17_ ( clk, n1437_r, a4_k0a[17], k3[113] );
not U_inv1292 ( n1437_r, n1437 );
dff a4_out_1_reg_113_ ( clk, n1437_r, k4[113], k3b[113] );
not U_inv1293 ( n780, k4[113] );
not U_inv1294 ( n1437_r, n1437 );
dff a4_k0a_reg_18_ ( clk, n1437_r, a4_k0a[18], k3[114] );
not U_inv1295 ( n1437_r, n1437 );
dff a4_out_1_reg_114_ ( clk, n1436_r, k4[114], k3b[114] );
not U_inv1296 ( n781, k4[114] );
not U_inv1297 ( n1436_r, n1436 );
dff a4_k0a_reg_19_ ( clk, n1436_r, a4_k0a[19], k3[115] );
not U_inv1298 ( n1436_r, n1436 );
dff a4_out_1_reg_115_ ( clk, n1436_r, k4[115], k3b[115] );
not U_inv1299 ( n782, k4[115] );
not U_inv1300 ( n1436_r, n1436 );
dff a4_k0a_reg_20_ ( clk, n1436_r, a4_k0a[20], k3[116] );
not U_inv1301 ( n1436_r, n1436 );
dff a4_out_1_reg_116_ ( clk, n1436_r, k4[116], k3b[116] );
not U_inv1302 ( n784, k4[116] );
not U_inv1303 ( n1436_r, n1436 );
dff a4_k0a_reg_21_ ( clk, n1436_r, a4_k0a[21], k3[117] );
not U_inv1304 ( n1436_r, n1436 );
dff a4_out_1_reg_117_ ( clk, n1436_r, k4[117], k3b[117] );
not U_inv1305 ( n785, k4[117] );
not U_inv1306 ( n1436_r, n1436 );
dff a4_k0a_reg_22_ ( clk, n1436_r, a4_k0a[22], k3[118] );
not U_inv1307 ( n1436_r, n1436 );
dff a4_out_1_reg_118_ ( clk, n1436_r, k4[118], k3b[118] );
not U_inv1308 ( n786, k4[118] );
not U_inv1309 ( n1436_r, n1436 );
dff a4_k0a_reg_23_ ( clk, n1436_r, a4_k0a[23], k3[119] );
not U_inv1310 ( n1436_r, n1436 );
dff a4_out_1_reg_119_ ( clk, n1436_r, k4[119], k3b[119] );
not U_inv1311 ( n787, k4[119] );
not U_inv1312 ( n1436_r, n1436 );
dff a4_k0a_reg_24_ ( clk, n1436_r, a4_k0a[24], k3[120] );
not U_inv1313 ( n1436_r, n1436 );
dff a4_out_1_reg_120_ ( clk, n1435_r, k4[120], k3b[120] );
not U_inv1314 ( n788, k4[120] );
not U_inv1315 ( n1435_r, n1435 );
dff a4_k0a_reg_25_ ( clk, n1435_r, a4_k0a[25], k3[121] );
not U_inv1316 ( n1435_r, n1435 );
dff a4_out_1_reg_121_ ( clk, n1435_r, k4[121], k3b[121] );
not U_inv1317 ( n789, k4[121] );
not U_inv1318 ( n1435_r, n1435 );
dff a4_k0a_reg_26_ ( clk, n1435_r, a4_k0a[26], k3[122] );
not U_inv1319 ( n1435_r, n1435 );
dff a4_out_1_reg_122_ ( clk, n1435_r, k4[122], k3b[122] );
not U_inv1320 ( n790, k4[122] );
not U_inv1321 ( n1435_r, n1435 );
dff a4_k0a_reg_27_ ( clk, n1435_r, a4_k0a[27], n1287 );
not U_inv1322 ( n1435_r, n1435 );
dff a4_out_1_reg_123_ ( clk, n1435_r, k4[123], k3b[123] );
not U_inv1323 ( n791, k4[123] );
not U_inv1324 ( n1435_r, n1435 );
dff a4_k0a_reg_28_ ( clk, n1435_r, a4_k0a[28], k3[124] );
not U_inv1325 ( n1435_r, n1435 );
dff a4_out_1_reg_124_ ( clk, n1435_r, ex_wire81, k3b[124] );
not U_inv1326 ( n1288, ex_wire81 );
not U_inv1327 ( n1435_r, n1435 );
dff a4_k0a_reg_29_ ( clk, n1435_r, a4_k0a[29], k3[125] );
not U_inv1328 ( n1435_r, n1435 );
dff a4_out_1_reg_125_ ( clk, n1435_r, k4[125], k3b[125] );
not U_inv1329 ( n792, k4[125] );
not U_inv1330 ( n1435_r, n1435 );
dff a4_k0a_reg_30_ ( clk, n1435_r, a4_k0a[30], k3[126] );
not U_inv1331 ( n1435_r, n1435 );
dff a4_out_1_reg_126_ ( clk, n1434_r, k4[126], k3b[126] );
not U_inv1332 ( n794, k4[126] );
not U_inv1333 ( n1434_r, n1434 );
dff a4_k0a_reg_31_ ( clk, n1434_r, a4_k0a[31], k3[127] );
not U_inv1334 ( n1434_r, n1434 );
dff a4_out_1_reg_127_ ( clk, n1434_r, k4[127], k3b[127] );
not U_inv1335 ( n795, k4[127] );
not U_inv1336 ( n1434_r, n1434 );
dff a4_k3a_reg_0_ ( clk, n1434_r, a4_k3a[0], a4_v3[0] );
not U_inv1337 ( n1434_r, n1434 );
dff a4_out_1_reg_0_ ( clk, n1434_r, k4[0], k3b[0] );
not U_inv1338 ( n1434_r, n1434 );
dff a4_k3a_reg_1_ ( clk, n1434_r, a4_k3a[1], a4_v3[1] );
not U_inv1339 ( n1434_r, n1434 );
dff a4_out_1_reg_1_ ( clk, n1434_r, k4[1], k3b[1] );
not U_inv1340 ( n1434_r, n1434 );
dff a4_k3a_reg_2_ ( clk, n1434_r, a4_k3a[2], a4_v3[2] );
not U_inv1341 ( n1434_r, n1434 );
dff a4_out_1_reg_2_ ( clk, n1434_r, k4[2], k3b[2] );
not U_inv1342 ( n1434_r, n1434 );
dff a4_k3a_reg_3_ ( clk, n1434_r, a4_k3a[3], a4_v3[3] );
not U_inv1343 ( n1434_r, n1434 );
dff a4_out_1_reg_3_ ( clk, n1434_r, k4[3], k3b[3] );
not U_inv1344 ( n1434_r, n1434 );
dff a4_k3a_reg_4_ ( clk, n1434_r, a4_k3a[4], a4_v3[4] );
not U_inv1345 ( n1434_r, n1434 );
dff a4_out_1_reg_4_ ( clk, n1433_r, k4[4], k3b[4] );
not U_inv1346 ( n1433_r, n1433 );
dff a4_k3a_reg_5_ ( clk, n1433_r, a4_k3a[5], a4_v3[5] );
not U_inv1347 ( n1433_r, n1433 );
dff a4_out_1_reg_5_ ( clk, n1433_r, k4[5], k3b[5] );
not U_inv1348 ( n1433_r, n1433 );
dff a4_k3a_reg_6_ ( clk, n1433_r, a4_k3a[6], a4_v3[6] );
not U_inv1349 ( n1433_r, n1433 );
dff a4_out_1_reg_6_ ( clk, n1433_r, k4[6], k3b[6] );
not U_inv1350 ( n1433_r, n1433 );
dff a4_k3a_reg_7_ ( clk, n1433_r, a4_k3a[7], a4_v3[7] );
not U_inv1351 ( n1433_r, n1433 );
dff a4_out_1_reg_7_ ( clk, n1433_r, k4[7], k3b[7] );
not U_inv1352 ( n1433_r, n1433 );
dff a4_k3a_reg_8_ ( clk, n1433_r, a4_k3a[8], a4_v3[8] );
not U_inv1353 ( n1433_r, n1433 );
dff a4_out_1_reg_8_ ( clk, n1433_r, k4[8], k3b[8] );
not U_inv1354 ( n1433_r, n1433 );
dff a4_k3a_reg_9_ ( clk, n1433_r, a4_k3a[9], a4_v3[9] );
not U_inv1355 ( n1433_r, n1433 );
dff a4_out_1_reg_9_ ( clk, n1433_r, k4[9], k3b[9] );
not U_inv1356 ( n1433_r, n1433 );
dff a4_k3a_reg_10_ ( clk, n1433_r, a4_k3a[10], a4_v3[10] );
not U_inv1357 ( n1433_r, n1433 );
dff a4_out_1_reg_10_ ( clk, n1432_r, k4[10], k3b[10] );
not U_inv1358 ( n1432_r, n1432 );
dff a4_k3a_reg_11_ ( clk, n1432_r, a4_k3a[11], a4_v3[11] );
not U_inv1359 ( n1432_r, n1432 );
dff a4_out_1_reg_11_ ( clk, n1432_r, k4[11], k3b[11] );
not U_inv1360 ( n1432_r, n1432 );
dff a4_k3a_reg_12_ ( clk, n1432_r, a4_k3a[12], a4_v3[12] );
not U_inv1361 ( n1432_r, n1432 );
dff a4_out_1_reg_12_ ( clk, n1432_r, k4[12], k3b[12] );
not U_inv1362 ( n1432_r, n1432 );
dff a4_k3a_reg_13_ ( clk, n1432_r, a4_k3a[13], a4_v3[13] );
not U_inv1363 ( n1432_r, n1432 );
dff a4_out_1_reg_13_ ( clk, n1432_r, k4[13], k3b[13] );
not U_inv1364 ( n1432_r, n1432 );
dff a4_k3a_reg_14_ ( clk, n1432_r, a4_k3a[14], a4_v3[14] );
not U_inv1365 ( n1432_r, n1432 );
dff a4_out_1_reg_14_ ( clk, n1432_r, k4[14], k3b[14] );
not U_inv1366 ( n1432_r, n1432 );
dff a4_k3a_reg_15_ ( clk, n1432_r, a4_k3a[15], a4_v3[15] );
not U_inv1367 ( n1432_r, n1432 );
dff a4_out_1_reg_15_ ( clk, n1432_r, k4[15], k3b[15] );
not U_inv1368 ( n1432_r, n1432 );
dff a4_k3a_reg_16_ ( clk, n1432_r, a4_k3a[16], a4_v3[16] );
not U_inv1369 ( n1432_r, n1432 );
dff a4_out_1_reg_16_ ( clk, n1431_r, k4[16], k3b[16] );
not U_inv1370 ( n1431_r, n1431 );
dff a4_k3a_reg_17_ ( clk, n1431_r, a4_k3a[17], a4_v3[17] );
not U_inv1371 ( n1431_r, n1431 );
dff a4_out_1_reg_17_ ( clk, n1431_r, k4[17], k3b[17] );
not U_inv1372 ( n1431_r, n1431 );
dff a4_k3a_reg_18_ ( clk, n1431_r, a4_k3a[18], a4_v3[18] );
not U_inv1373 ( n1431_r, n1431 );
dff a4_out_1_reg_18_ ( clk, n1431_r, k4[18], k3b[18] );
not U_inv1374 ( n1431_r, n1431 );
dff a4_k3a_reg_19_ ( clk, n1431_r, a4_k3a[19], a4_v3[19] );
not U_inv1375 ( n1431_r, n1431 );
dff a4_out_1_reg_19_ ( clk, n1431_r, k4[19], k3b[19] );
not U_inv1376 ( n1431_r, n1431 );
dff a4_k3a_reg_20_ ( clk, n1431_r, a4_k3a[20], a4_v3[20] );
not U_inv1377 ( n1431_r, n1431 );
dff a4_out_1_reg_20_ ( clk, n1431_r, k4[20], k3b[20] );
not U_inv1378 ( n1431_r, n1431 );
dff a4_k3a_reg_21_ ( clk, n1431_r, a4_k3a[21], a4_v3[21] );
not U_inv1379 ( n1431_r, n1431 );
dff a4_out_1_reg_21_ ( clk, n1431_r, k4[21], k3b[21] );
not U_inv1380 ( n1431_r, n1431 );
dff a4_k3a_reg_22_ ( clk, n1431_r, a4_k3a[22], a4_v3[22] );
not U_inv1381 ( n1431_r, n1431 );
dff a4_out_1_reg_22_ ( clk, n1430_r, k4[22], k3b[22] );
not U_inv1382 ( n1430_r, n1430 );
dff a4_k3a_reg_23_ ( clk, n1430_r, a4_k3a[23], a4_v3[23] );
not U_inv1383 ( n1430_r, n1430 );
dff a4_out_1_reg_23_ ( clk, n1430_r, k4[23], k3b[23] );
not U_inv1384 ( n1430_r, n1430 );
dff a4_k3a_reg_24_ ( clk, n1430_r, a4_k3a[24], a4_v3[24] );
not U_inv1385 ( n1430_r, n1430 );
dff a4_out_1_reg_24_ ( clk, n1430_r, k4[24], k3b[24] );
not U_inv1386 ( n1430_r, n1430 );
dff a4_k3a_reg_25_ ( clk, n1430_r, a4_k3a[25], a4_v3[25] );
not U_inv1387 ( n1430_r, n1430 );
dff a4_out_1_reg_25_ ( clk, n1430_r, k4[25], k3b[25] );
not U_inv1388 ( n1430_r, n1430 );
dff a4_k3a_reg_26_ ( clk, n1430_r, a4_k3a[26], a4_v3[26] );
not U_inv1389 ( n1430_r, n1430 );
dff a4_out_1_reg_26_ ( clk, n1430_r, k4[26], k3b[26] );
not U_inv1390 ( n1430_r, n1430 );
dff a4_k3a_reg_27_ ( clk, n1430_r, a4_k3a[27], a4_v3[27] );
not U_inv1391 ( n1430_r, n1430 );
dff a4_out_1_reg_27_ ( clk, n1430_r, k4[27], k3b[27] );
not U_inv1392 ( n1430_r, n1430 );
dff a4_k3a_reg_28_ ( clk, n1430_r, a4_k3a[28], a4_v3[28] );
not U_inv1393 ( n1430_r, n1430 );
dff a4_out_1_reg_28_ ( clk, n1429_r, k4[28], k3b[28] );
not U_inv1394 ( n1429_r, n1429 );
dff a4_k3a_reg_29_ ( clk, n1429_r, a4_k3a[29], a4_v3[29] );
not U_inv1395 ( n1429_r, n1429 );
dff a4_out_1_reg_29_ ( clk, n1429_r, k4[29], k3b[29] );
not U_inv1396 ( n1429_r, n1429 );
dff a4_k3a_reg_30_ ( clk, n1429_r, a4_k3a[30], a4_v3[30] );
not U_inv1397 ( n1429_r, n1429 );
dff a4_out_1_reg_30_ ( clk, n1429_r, k4[30], k3b[30] );
not U_inv1398 ( n1429_r, n1429 );
dff a4_k2a_reg_0_ ( clk, n1429_r, a4_k2a[0], a4_v2[0] );
not U_inv1399 ( n1429_r, n1429 );
dff a4_out_1_reg_32_ ( clk, n1429_r, k4[32], k3b[32] );
not U_inv1400 ( n1429_r, n1429 );
dff a4_k2a_reg_1_ ( clk, n1429_r, a4_k2a[1], a4_v2[1] );
not U_inv1401 ( n1429_r, n1429 );
dff a4_out_1_reg_33_ ( clk, n1429_r, k4[33], k3b[33] );
not U_inv1402 ( n1429_r, n1429 );
dff a4_k2a_reg_2_ ( clk, n1429_r, a4_k2a[2], a4_v2[2] );
not U_inv1403 ( n1429_r, n1429 );
dff a4_out_1_reg_34_ ( clk, n1429_r, k4[34], k3b[34] );
not U_inv1404 ( n1429_r, n1429 );
dff a4_k2a_reg_3_ ( clk, n1429_r, a4_k2a[3], a4_v2[3] );
not U_inv1405 ( n1429_r, n1429 );
dff a4_out_1_reg_35_ ( clk, n1428_r, k4[35], k3b[35] );
not U_inv1406 ( n1428_r, n1428 );
dff a4_k2a_reg_4_ ( clk, n1428_r, a4_k2a[4], a4_v2[4] );
not U_inv1407 ( n1428_r, n1428 );
dff a4_out_1_reg_36_ ( clk, n1428_r, k4[36], k3b[36] );
not U_inv1408 ( n1428_r, n1428 );
dff a4_k2a_reg_5_ ( clk, n1428_r, a4_k2a[5], a4_v2[5] );
not U_inv1409 ( n1428_r, n1428 );
dff a4_out_1_reg_37_ ( clk, n1428_r, k4[37], k3b[37] );
not U_inv1410 ( n1428_r, n1428 );
dff a4_k2a_reg_6_ ( clk, n1428_r, a4_k2a[6], a4_v2[6] );
not U_inv1411 ( n1428_r, n1428 );
dff a4_out_1_reg_38_ ( clk, n1428_r, k4[38], k3b[38] );
not U_inv1412 ( n1428_r, n1428 );
dff a4_k2a_reg_7_ ( clk, n1428_r, a4_k2a[7], a4_v2[7] );
not U_inv1413 ( n1428_r, n1428 );
dff a4_out_1_reg_39_ ( clk, n1428_r, k4[39], k3b[39] );
not U_inv1414 ( n1428_r, n1428 );
dff a4_k2a_reg_8_ ( clk, n1428_r, a4_k2a[8], a4_v2[8] );
not U_inv1415 ( n1428_r, n1428 );
dff a4_out_1_reg_40_ ( clk, n1428_r, k4[40], k3b[40] );
not U_inv1416 ( n1428_r, n1428 );
dff a4_k2a_reg_9_ ( clk, n1428_r, a4_k2a[9], a4_v2[9] );
not U_inv1417 ( n1428_r, n1428 );
dff a4_out_1_reg_41_ ( clk, n1427_r, k4[41], k3b[41] );
not U_inv1418 ( n1427_r, n1427 );
dff a4_k2a_reg_10_ ( clk, n1427_r, a4_k2a[10], a4_v2[10] );
not U_inv1419 ( n1427_r, n1427 );
dff a4_out_1_reg_42_ ( clk, n1427_r, k4[42], k3b[42] );
not U_inv1420 ( n1427_r, n1427 );
dff a4_k2a_reg_11_ ( clk, n1427_r, a4_k2a[11], a4_v2[11] );
not U_inv1421 ( n1427_r, n1427 );
dff a4_out_1_reg_43_ ( clk, n1427_r, k4[43], k3b[43] );
not U_inv1422 ( n1427_r, n1427 );
dff a4_k2a_reg_12_ ( clk, n1427_r, a4_k2a[12], a4_v2[12] );
not U_inv1423 ( n1427_r, n1427 );
dff a4_out_1_reg_44_ ( clk, n1427_r, k4[44], k3b[44] );
not U_inv1424 ( n1427_r, n1427 );
dff a4_k2a_reg_13_ ( clk, n1427_r, a4_k2a[13], a4_v2[13] );
not U_inv1425 ( n1427_r, n1427 );
dff a4_out_1_reg_45_ ( clk, n1427_r, k4[45], k3b[45] );
not U_inv1426 ( n1427_r, n1427 );
dff a4_k2a_reg_14_ ( clk, n1427_r, a4_k2a[14], a4_v2[14] );
not U_inv1427 ( n1427_r, n1427 );
dff a4_out_1_reg_46_ ( clk, n1427_r, k4[46], k3b[46] );
not U_inv1428 ( n1427_r, n1427 );
dff a4_k2a_reg_15_ ( clk, n1427_r, a4_k2a[15], a4_v2[15] );
not U_inv1429 ( n1427_r, n1427 );
dff a4_out_1_reg_47_ ( clk, n1426_r, k4[47], k3b[47] );
not U_inv1430 ( n1426_r, n1426 );
dff a4_k2a_reg_16_ ( clk, n1426_r, a4_k2a[16], a4_v2[16] );
not U_inv1431 ( n1426_r, n1426 );
dff a4_out_1_reg_48_ ( clk, n1426_r, k4[48], k3b[48] );
not U_inv1432 ( n1426_r, n1426 );
dff a4_k2a_reg_17_ ( clk, n1426_r, a4_k2a[17], a4_v2[17] );
not U_inv1433 ( n1426_r, n1426 );
dff a4_out_1_reg_49_ ( clk, n1426_r, k4[49], k3b[49] );
not U_inv1434 ( n1426_r, n1426 );
dff a4_k2a_reg_18_ ( clk, n1426_r, a4_k2a[18], a4_v2[18] );
not U_inv1435 ( n1426_r, n1426 );
dff a4_out_1_reg_50_ ( clk, n1426_r, k4[50], k3b[50] );
not U_inv1436 ( n1426_r, n1426 );
dff a4_k2a_reg_19_ ( clk, n1426_r, a4_k2a[19], a4_v2[19] );
not U_inv1437 ( n1426_r, n1426 );
dff a4_out_1_reg_51_ ( clk, n1426_r, k4[51], k3b[51] );
not U_inv1438 ( n1426_r, n1426 );
dff a4_k2a_reg_20_ ( clk, n1426_r, a4_k2a[20], a4_v2[20] );
not U_inv1439 ( n1426_r, n1426 );
dff a4_out_1_reg_52_ ( clk, n1426_r, k4[52], k3b[52] );
not U_inv1440 ( n1426_r, n1426 );
dff a4_k2a_reg_21_ ( clk, n1426_r, a4_k2a[21], a4_v2[21] );
not U_inv1441 ( n1426_r, n1426 );
dff a4_out_1_reg_53_ ( clk, n1425_r, k4[53], k3b[53] );
not U_inv1442 ( n1425_r, n1425 );
dff a4_k2a_reg_22_ ( clk, n1425_r, a4_k2a[22], a4_v2[22] );
not U_inv1443 ( n1425_r, n1425 );
dff a4_out_1_reg_54_ ( clk, n1425_r, k4[54], k3b[54] );
not U_inv1444 ( n1425_r, n1425 );
dff a4_k2a_reg_23_ ( clk, n1425_r, a4_k2a[23], a4_v2[23] );
not U_inv1445 ( n1425_r, n1425 );
dff a4_out_1_reg_55_ ( clk, n1425_r, k4[55], k3b[55] );
not U_inv1446 ( n1425_r, n1425 );
dff a4_k2a_reg_24_ ( clk, n1425_r, a4_k2a[24], a4_v2[24] );
not U_inv1447 ( n1425_r, n1425 );
dff a4_out_1_reg_56_ ( clk, n1425_r, k4[56], k3b[56] );
not U_inv1448 ( n1425_r, n1425 );
dff a4_k2a_reg_25_ ( clk, n1425_r, a4_k2a[25], a4_v2[25] );
not U_inv1449 ( n1425_r, n1425 );
dff a4_out_1_reg_57_ ( clk, n1425_r, k4[57], k3b[57] );
not U_inv1450 ( n1425_r, n1425 );
dff a4_k2a_reg_26_ ( clk, n1425_r, a4_k2a[26], a4_v2[26] );
not U_inv1451 ( n1425_r, n1425 );
dff a4_out_1_reg_58_ ( clk, n1425_r, k4[58], k3b[58] );
not U_inv1452 ( n1425_r, n1425 );
dff a4_k2a_reg_27_ ( clk, n1425_r, a4_k2a[27], a4_v2[27] );
not U_inv1453 ( n1425_r, n1425 );
dff a4_out_1_reg_59_ ( clk, n1424_r, k4[59], k3b[59] );
not U_inv1454 ( n1424_r, n1424 );
dff a4_k2a_reg_28_ ( clk, n1424_r, a4_k2a[28], a4_v2[28] );
not U_inv1455 ( n1424_r, n1424 );
dff a4_out_1_reg_60_ ( clk, n1424_r, k4[60], k3b[60] );
not U_inv1456 ( n1424_r, n1424 );
dff a4_k2a_reg_29_ ( clk, n1424_r, a4_k2a[29], a4_v2[29] );
not U_inv1457 ( n1424_r, n1424 );
dff a4_out_1_reg_61_ ( clk, n1424_r, k4[61], k3b[61] );
not U_inv1458 ( n1424_r, n1424 );
dff a4_k2a_reg_30_ ( clk, n1424_r, a4_k2a[30], a4_v2[30] );
not U_inv1459 ( n1424_r, n1424 );
dff a4_out_1_reg_62_ ( clk, n1424_r, k4[62], k3b[62] );
not U_inv1460 ( n1424_r, n1424 );
dff a4_k2a_reg_31_ ( clk, n1424_r, a4_k2a[31], a4_v2[31] );
not U_inv1461 ( n1424_r, n1424 );
dff a4_out_1_reg_63_ ( clk, n1424_r, k4[63], k3b[63] );
not U_inv1462 ( n1424_r, n1424 );
dff a4_k1a_reg_0_ ( clk, n1424_r, a4_k1a[0], a4_v1[0] );
not U_inv1463 ( n1424_r, n1424 );
dff a4_out_1_reg_64_ ( clk, n1424_r, ex_wire82, k3b[64] );
not U_inv1464 ( n772, ex_wire82 );
not U_inv1465 ( n1424_r, n1424 );
dff a4_k1a_reg_1_ ( clk, n1424_r, a4_k1a[1], a4_v1[1] );
not U_inv1466 ( n1424_r, n1424 );
dff a4_out_1_reg_65_ ( clk, n1423_r, ex_wire83, k3b[65] );
not U_inv1467 ( n783, ex_wire83 );
not U_inv1468 ( n1423_r, n1423 );
dff a4_k1a_reg_2_ ( clk, n1423_r, a4_k1a[2], a4_v1[2] );
not U_inv1469 ( n1423_r, n1423 );
dff a4_out_1_reg_66_ ( clk, n1423_r, ex_wire84, k3b[66] );
not U_inv1470 ( n793, ex_wire84 );
not U_inv1471 ( n1423_r, n1423 );
dff a4_k1a_reg_3_ ( clk, n1423_r, a4_k1a[3], a4_v1[3] );
not U_inv1472 ( n1423_r, n1423 );
dff a4_out_1_reg_67_ ( clk, n1423_r, ex_wire85, k3b[67] );
not U_inv1473 ( n796, ex_wire85 );
not U_inv1474 ( n1423_r, n1423 );
dff a4_k1a_reg_4_ ( clk, n1423_r, a4_k1a[4], a4_v1[4] );
not U_inv1475 ( n1423_r, n1423 );
dff a4_out_1_reg_68_ ( clk, n1423_r, k4[68], k3b[68] );
not U_inv1476 ( n1423_r, n1423 );
dff a4_k1a_reg_5_ ( clk, n1423_r, a4_k1a[5], a4_v1[5] );
not U_inv1477 ( n1423_r, n1423 );
dff a4_out_1_reg_69_ ( clk, n1423_r, k4[69], k3b[69] );
not U_inv1478 ( n1423_r, n1423 );
dff a4_k1a_reg_6_ ( clk, n1423_r, a4_k1a[6], a4_v1[6] );
not U_inv1479 ( n1423_r, n1423 );
dff a4_out_1_reg_70_ ( clk, n1423_r, k4[70], k3b[70] );
not U_inv1480 ( n1423_r, n1423 );
dff a4_k1a_reg_7_ ( clk, n1423_r, a4_k1a[7], a4_v1[7] );
not U_inv1481 ( n1423_r, n1423 );
dff a4_out_1_reg_71_ ( clk, n1422_r, k4[71], k3b[71] );
not U_inv1482 ( n1422_r, n1422 );
dff a4_k1a_reg_8_ ( clk, n1422_r, a4_k1a[8], a4_v1[8] );
not U_inv1483 ( n1422_r, n1422 );
dff a4_out_1_reg_72_ ( clk, n1422_r, k4[72], k3b[72] );
not U_inv1484 ( n1422_r, n1422 );
dff a4_k1a_reg_9_ ( clk, n1422_r, a4_k1a[9], a4_v1[9] );
not U_inv1485 ( n1422_r, n1422 );
dff a4_out_1_reg_73_ ( clk, n1422_r, k4[73], k3b[73] );
not U_inv1486 ( n1422_r, n1422 );
dff a4_k1a_reg_10_ ( clk, n1422_r, a4_k1a[10], a4_v1[10] );
not U_inv1487 ( n1422_r, n1422 );
dff a4_out_1_reg_74_ ( clk, n1422_r, k4[74], k3b[74] );
not U_inv1488 ( n1422_r, n1422 );
dff a4_k1a_reg_11_ ( clk, n1422_r, a4_k1a[11], a4_v1[11] );
not U_inv1489 ( n1422_r, n1422 );
dff a4_out_1_reg_75_ ( clk, n1422_r, k4[75], k3b[75] );
not U_inv1490 ( n1422_r, n1422 );
dff a4_k1a_reg_12_ ( clk, n1422_r, a4_k1a[12], a4_v1[12] );
not U_inv1491 ( n1422_r, n1422 );
dff a4_out_1_reg_76_ ( clk, n1422_r, k4[76], k3b[76] );
not U_inv1492 ( n1422_r, n1422 );
dff a4_k1a_reg_13_ ( clk, n1422_r, a4_k1a[13], a4_v1[13] );
not U_inv1493 ( n1422_r, n1422 );
dff a4_out_1_reg_77_ ( clk, n1421_r, k4[77], k3b[77] );
not U_inv1494 ( n1421_r, n1421 );
dff a4_k1a_reg_14_ ( clk, n1421_r, a4_k1a[14], a4_v1[14] );
not U_inv1495 ( n1421_r, n1421 );
dff a4_out_1_reg_78_ ( clk, n1421_r, k4[78], k3b[78] );
not U_inv1496 ( n1421_r, n1421 );
dff a4_k1a_reg_15_ ( clk, n1421_r, a4_k1a[15], a4_v1[15] );
not U_inv1497 ( n1421_r, n1421 );
dff a4_out_1_reg_79_ ( clk, n1421_r, k4[79], k3b[79] );
not U_inv1498 ( n1421_r, n1421 );
dff a4_k1a_reg_16_ ( clk, n1421_r, a4_k1a[16], a4_v1[16] );
not U_inv1499 ( n1421_r, n1421 );
dff a4_out_1_reg_80_ ( clk, n1421_r, k4[80], k3b[80] );
not U_inv1500 ( n1421_r, n1421 );
dff a4_k1a_reg_17_ ( clk, n1421_r, a4_k1a[17], a4_v1[17] );
not U_inv1501 ( n1421_r, n1421 );
dff a4_out_1_reg_81_ ( clk, n1421_r, k4[81], k3b[81] );
not U_inv1502 ( n1421_r, n1421 );
dff a4_k1a_reg_18_ ( clk, n1421_r, a4_k1a[18], a4_v1[18] );
not U_inv1503 ( n1421_r, n1421 );
dff a4_out_1_reg_82_ ( clk, n1421_r, k4[82], k3b[82] );
not U_inv1504 ( n1421_r, n1421 );
dff a4_k1a_reg_19_ ( clk, n1421_r, a4_k1a[19], a4_v1[19] );
not U_inv1505 ( n1421_r, n1421 );
dff a4_out_1_reg_83_ ( clk, n1420_r, k4[83], k3b[83] );
not U_inv1506 ( n1420_r, n1420 );
dff a4_k1a_reg_20_ ( clk, n1420_r, a4_k1a[20], a4_v1[20] );
not U_inv1507 ( n1420_r, n1420 );
dff a4_out_1_reg_84_ ( clk, n1420_r, k4[84], k3b[84] );
not U_inv1508 ( n1420_r, n1420 );
dff a4_k1a_reg_21_ ( clk, n1420_r, a4_k1a[21], a4_v1[21] );
not U_inv1509 ( n1420_r, n1420 );
dff a4_out_1_reg_85_ ( clk, n1420_r, k4[85], k3b[85] );
not U_inv1510 ( n1420_r, n1420 );
dff a4_k1a_reg_22_ ( clk, n1420_r, a4_k1a[22], a4_v1[22] );
not U_inv1511 ( n1420_r, n1420 );
dff a4_out_1_reg_86_ ( clk, n1420_r, k4[86], k3b[86] );
not U_inv1512 ( n1420_r, n1420 );
dff a4_k1a_reg_23_ ( clk, n1420_r, a4_k1a[23], a4_v1[23] );
not U_inv1513 ( n1420_r, n1420 );
dff a4_out_1_reg_87_ ( clk, n1420_r, k4[87], k3b[87] );
not U_inv1514 ( n1420_r, n1420 );
dff a4_k1a_reg_24_ ( clk, n1420_r, a4_k1a[24], a4_v1[24] );
not U_inv1515 ( n1420_r, n1420 );
dff a4_out_1_reg_88_ ( clk, n1420_r, k4[88], k3b[88] );
not U_inv1516 ( n1420_r, n1420 );
dff a4_k1a_reg_25_ ( clk, n1420_r, a4_k1a[25], a4_v1[25] );
not U_inv1517 ( n1420_r, n1420 );
dff a4_out_1_reg_89_ ( clk, n1419_r, k4[89], k3b[89] );
not U_inv1518 ( n1419_r, n1419 );
dff a4_k1a_reg_26_ ( clk, n1419_r, a4_k1a[26], a4_v1[26] );
not U_inv1519 ( n1419_r, n1419 );
dff a4_out_1_reg_90_ ( clk, n1419_r, k4[90], k3b[90] );
not U_inv1520 ( n1419_r, n1419 );
dff a4_k1a_reg_27_ ( clk, n1419_r, a4_k1a[27], a4_v1[27] );
not U_inv1521 ( n1419_r, n1419 );
dff a4_out_1_reg_91_ ( clk, n1419_r, k4[91], k3b[91] );
not U_inv1522 ( n1419_r, n1419 );
dff a4_k1a_reg_28_ ( clk, n1419_r, a4_k1a[28], a4_v1[28] );
not U_inv1523 ( n1419_r, n1419 );
dff a4_out_1_reg_92_ ( clk, n1419_r, k4[92], k3b[92] );
not U_inv1524 ( n1419_r, n1419 );
dff a4_k1a_reg_29_ ( clk, n1419_r, a4_k1a[29], a4_v1[29] );
not U_inv1525 ( n1419_r, n1419 );
dff a4_out_1_reg_93_ ( clk, n1419_r, k4[93], k3b[93] );
not U_inv1526 ( n1419_r, n1419 );
dff a4_k1a_reg_30_ ( clk, n1419_r, a4_k1a[30], a4_v1[30] );
not U_inv1527 ( n1419_r, n1419 );
dff a4_out_1_reg_94_ ( clk, n1419_r, k4[94], k3b[94] );
not U_inv1528 ( n1419_r, n1419 );
dff a4_out_1_reg_95_ ( clk, n1419_r, k4[95], k3b[95] );
not U_inv1529 ( n1419_r, n1419 );
dff a5_k0a_reg_0_ ( clk, n1418_r, a5_k0a[0], k4[96] );
not U_inv1530 ( n1418_r, n1418 );
dff a5_out_1_reg_96_ ( clk, n1418_r, k5[96], k4b[96] );
not U_inv1531 ( n1418_r, n1418 );
dff a5_k0a_reg_1_ ( clk, n1418_r, a5_k0a[1], k4[97] );
not U_inv1532 ( n1418_r, n1418 );
dff a5_out_1_reg_97_ ( clk, n1418_r, k5[97], k4b[97] );
not U_inv1533 ( n1418_r, n1418 );
dff a5_k0a_reg_2_ ( clk, n1418_r, a5_k0a[2], k4[98] );
not U_inv1534 ( n1418_r, n1418 );
dff a5_out_1_reg_98_ ( clk, n1418_r, k5[98], k4b[98] );
not U_inv1535 ( n1418_r, n1418 );
dff a5_k0a_reg_3_ ( clk, n1418_r, a5_k0a[3], k4[99] );
not U_inv1536 ( n1418_r, n1418 );
dff a5_out_1_reg_99_ ( clk, n1418_r, k5[99], k4b[99] );
not U_inv1537 ( n1418_r, n1418 );
dff a5_k0a_reg_4_ ( clk, n1418_r, a5_k0a[4], k4[100] );
not U_inv1538 ( n1418_r, n1418 );
dff a5_out_1_reg_100_ ( clk, n1418_r, k5[100], k4b[100] );
not U_inv1539 ( n828, k5[100] );
not U_inv1540 ( n1418_r, n1418 );
dff a5_k0a_reg_5_ ( clk, n1418_r, a5_k0a[5], k4[101] );
not U_inv1541 ( n1418_r, n1418 );
dff a5_out_1_reg_101_ ( clk, n1418_r, k5[101], k4b[101] );
not U_inv1542 ( n829, k5[101] );
not U_inv1543 ( n1418_r, n1418 );
dff a5_k0a_reg_6_ ( clk, n1417_r, a5_k0a[6], k4[102] );
not U_inv1544 ( n1417_r, n1417 );
dff a5_out_1_reg_102_ ( clk, n1417_r, k5[102], k4b[102] );
not U_inv1545 ( n830, k5[102] );
not U_inv1546 ( n1417_r, n1417 );
dff a5_k0a_reg_7_ ( clk, n1417_r, a5_k0a[7], k4[103] );
not U_inv1547 ( n1417_r, n1417 );
dff a5_out_1_reg_103_ ( clk, n1417_r, k5[103], k4b[103] );
not U_inv1548 ( n831, k5[103] );
not U_inv1549 ( n1417_r, n1417 );
dff a5_k0a_reg_8_ ( clk, n1417_r, a5_k0a[8], k4[104] );
not U_inv1550 ( n1417_r, n1417 );
dff a5_out_1_reg_104_ ( clk, n1417_r, k5[104], k4b[104] );
not U_inv1551 ( n832, k5[104] );
not U_inv1552 ( n1417_r, n1417 );
dff a5_k0a_reg_9_ ( clk, n1417_r, a5_k0a[9], k4[105] );
not U_inv1553 ( n1417_r, n1417 );
dff a5_out_1_reg_105_ ( clk, n1417_r, k5[105], k4b[105] );
not U_inv1554 ( n833, k5[105] );
not U_inv1555 ( n1417_r, n1417 );
dff a5_k0a_reg_10_ ( clk, n1417_r, a5_k0a[10], k4[106] );
not U_inv1556 ( n1417_r, n1417 );
dff a5_out_1_reg_106_ ( clk, n1417_r, k5[106], k4b[106] );
not U_inv1557 ( n804, k5[106] );
not U_inv1558 ( n1417_r, n1417 );
dff a5_k0a_reg_11_ ( clk, n1417_r, a5_k0a[11], k4[107] );
not U_inv1559 ( n1417_r, n1417 );
dff a5_out_1_reg_107_ ( clk, n1417_r, k5[107], k4b[107] );
not U_inv1560 ( n805, k5[107] );
not U_inv1561 ( n1417_r, n1417 );
dff a5_k0a_reg_12_ ( clk, n1416_r, a5_k0a[12], k4[108] );
not U_inv1562 ( n1416_r, n1416 );
dff a5_out_1_reg_108_ ( clk, n1416_r, k5[108], k4b[108] );
not U_inv1563 ( n806, k5[108] );
not U_inv1564 ( n1416_r, n1416 );
dff a5_k0a_reg_13_ ( clk, n1416_r, a5_k0a[13], k4[109] );
not U_inv1565 ( n1416_r, n1416 );
dff a5_out_1_reg_109_ ( clk, n1416_r, k5[109], k4b[109] );
not U_inv1566 ( n807, k5[109] );
not U_inv1567 ( n1416_r, n1416 );
dff a5_k0a_reg_14_ ( clk, n1416_r, a5_k0a[14], k4[110] );
not U_inv1568 ( n1416_r, n1416 );
dff a5_out_1_reg_110_ ( clk, n1416_r, k5[110], k4b[110] );
not U_inv1569 ( n808, k5[110] );
not U_inv1570 ( n1416_r, n1416 );
dff a5_k0a_reg_15_ ( clk, n1416_r, a5_k0a[15], k4[111] );
not U_inv1571 ( n1416_r, n1416 );
dff a5_out_1_reg_111_ ( clk, n1416_r, k5[111], k4b[111] );
not U_inv1572 ( n809, k5[111] );
not U_inv1573 ( n1416_r, n1416 );
dff a5_k0a_reg_16_ ( clk, n1416_r, a5_k0a[16], k4[112] );
not U_inv1574 ( n1416_r, n1416 );
dff a5_out_1_reg_112_ ( clk, n1416_r, k5[112], k4b[112] );
not U_inv1575 ( n810, k5[112] );
not U_inv1576 ( n1416_r, n1416 );
dff a5_k0a_reg_17_ ( clk, n1416_r, a5_k0a[17], k4[113] );
not U_inv1577 ( n1416_r, n1416 );
dff a5_out_1_reg_113_ ( clk, n1416_r, k5[113], k4b[113] );
not U_inv1578 ( n811, k5[113] );
not U_inv1579 ( n1416_r, n1416 );
dff a5_k0a_reg_18_ ( clk, n1415_r, a5_k0a[18], k4[114] );
not U_inv1580 ( n1415_r, n1415 );
dff a5_out_1_reg_114_ ( clk, n1415_r, k5[114], k4b[114] );
not U_inv1581 ( n812, k5[114] );
not U_inv1582 ( n1415_r, n1415 );
dff a5_k0a_reg_19_ ( clk, n1415_r, a5_k0a[19], k4[115] );
not U_inv1583 ( n1415_r, n1415 );
dff a5_out_1_reg_115_ ( clk, n1415_r, k5[115], k4b[115] );
not U_inv1584 ( n813, k5[115] );
not U_inv1585 ( n1415_r, n1415 );
dff a5_k0a_reg_20_ ( clk, n1415_r, a5_k0a[20], k4[116] );
not U_inv1586 ( n1415_r, n1415 );
dff a5_out_1_reg_116_ ( clk, n1415_r, k5[116], k4b[116] );
not U_inv1587 ( n815, k5[116] );
not U_inv1588 ( n1415_r, n1415 );
dff a5_k0a_reg_21_ ( clk, n1415_r, a5_k0a[21], k4[117] );
not U_inv1589 ( n1415_r, n1415 );
dff a5_out_1_reg_117_ ( clk, n1415_r, k5[117], k4b[117] );
not U_inv1590 ( n816, k5[117] );
not U_inv1591 ( n1415_r, n1415 );
dff a5_k0a_reg_22_ ( clk, n1415_r, a5_k0a[22], k4[118] );
not U_inv1592 ( n1415_r, n1415 );
dff a5_out_1_reg_118_ ( clk, n1415_r, k5[118], k4b[118] );
not U_inv1593 ( n817, k5[118] );
not U_inv1594 ( n1415_r, n1415 );
dff a5_k0a_reg_23_ ( clk, n1415_r, a5_k0a[23], k4[119] );
not U_inv1595 ( n1415_r, n1415 );
dff a5_out_1_reg_119_ ( clk, n1415_r, k5[119], k4b[119] );
not U_inv1596 ( n818, k5[119] );
not U_inv1597 ( n1415_r, n1415 );
dff a5_k0a_reg_24_ ( clk, n1414_r, a5_k0a[24], k4[120] );
not U_inv1598 ( n1414_r, n1414 );
dff a5_out_1_reg_120_ ( clk, n1414_r, k5[120], k4b[120] );
not U_inv1599 ( n819, k5[120] );
not U_inv1600 ( n1414_r, n1414 );
dff a5_k0a_reg_25_ ( clk, n1414_r, a5_k0a[25], k4[121] );
not U_inv1601 ( n1414_r, n1414 );
dff a5_out_1_reg_121_ ( clk, n1414_r, k5[121], k4b[121] );
not U_inv1602 ( n820, k5[121] );
not U_inv1603 ( n1414_r, n1414 );
dff a5_k0a_reg_26_ ( clk, n1414_r, a5_k0a[26], k4[122] );
not U_inv1604 ( n1414_r, n1414 );
dff a5_out_1_reg_122_ ( clk, n1414_r, k5[122], k4b[122] );
not U_inv1605 ( n821, k5[122] );
not U_inv1606 ( n1414_r, n1414 );
dff a5_k0a_reg_27_ ( clk, n1414_r, a5_k0a[27], k4[123] );
not U_inv1607 ( n1414_r, n1414 );
dff a5_out_1_reg_123_ ( clk, n1414_r, k5[123], k4b[123] );
not U_inv1608 ( n822, k5[123] );
not U_inv1609 ( n1414_r, n1414 );
dff a5_k0a_reg_28_ ( clk, n1414_r, a5_k0a[28], n1288 );
not U_inv1610 ( n1414_r, n1414 );
dff a5_out_1_reg_124_ ( clk, n1414_r, k5[124], k4b[124] );
not U_inv1611 ( n823, k5[124] );
not U_inv1612 ( n1414_r, n1414 );
dff a5_k0a_reg_29_ ( clk, n1414_r, a5_k0a[29], k4[125] );
not U_inv1613 ( n1414_r, n1414 );
dff a5_out_1_reg_125_ ( clk, n1414_r, ex_wire86, k4b[125] );
not U_inv1614 ( n1289, ex_wire86 );
not U_inv1615 ( n1414_r, n1414 );
dff a5_k0a_reg_30_ ( clk, n1413_r, a5_k0a[30], k4[126] );
not U_inv1616 ( n1413_r, n1413 );
dff a5_out_1_reg_126_ ( clk, n1413_r, k5[126], k4b[126] );
not U_inv1617 ( n825, k5[126] );
not U_inv1618 ( n1413_r, n1413 );
dff a5_k0a_reg_31_ ( clk, n1413_r, a5_k0a[31], k4[127] );
not U_inv1619 ( n1413_r, n1413 );
dff a5_out_1_reg_127_ ( clk, n1413_r, k5[127], k4b[127] );
not U_inv1620 ( n826, k5[127] );
not U_inv1621 ( n1413_r, n1413 );
dff a5_k3a_reg_0_ ( clk, n1413_r, a5_k3a[0], a5_v3[0] );
not U_inv1622 ( n1413_r, n1413 );
dff a5_out_1_reg_0_ ( clk, n1413_r, k5[0], k4b[0] );
not U_inv1623 ( n1413_r, n1413 );
dff a5_k3a_reg_1_ ( clk, n1413_r, a5_k3a[1], a5_v3[1] );
not U_inv1624 ( n1413_r, n1413 );
dff a5_out_1_reg_1_ ( clk, n1413_r, k5[1], k4b[1] );
not U_inv1625 ( n1413_r, n1413 );
dff a5_k3a_reg_2_ ( clk, n1413_r, a5_k3a[2], a5_v3[2] );
not U_inv1626 ( n1413_r, n1413 );
dff a5_out_1_reg_2_ ( clk, n1413_r, k5[2], k4b[2] );
not U_inv1627 ( n1413_r, n1413 );
dff a5_k3a_reg_3_ ( clk, n1413_r, a5_k3a[3], a5_v3[3] );
not U_inv1628 ( n1413_r, n1413 );
dff a5_out_1_reg_3_ ( clk, n1413_r, k5[3], k4b[3] );
not U_inv1629 ( n1413_r, n1413 );
dff a5_k3a_reg_4_ ( clk, n1412_r, a5_k3a[4], a5_v3[4] );
not U_inv1630 ( n1412_r, n1412 );
dff a5_out_1_reg_4_ ( clk, n1412_r, k5[4], k4b[4] );
not U_inv1631 ( n1412_r, n1412 );
dff a5_k3a_reg_5_ ( clk, n1412_r, a5_k3a[5], a5_v3[5] );
not U_inv1632 ( n1412_r, n1412 );
dff a5_out_1_reg_5_ ( clk, n1412_r, k5[5], k4b[5] );
not U_inv1633 ( n1412_r, n1412 );
dff a5_k3a_reg_6_ ( clk, n1412_r, a5_k3a[6], a5_v3[6] );
not U_inv1634 ( n1412_r, n1412 );
dff a5_out_1_reg_6_ ( clk, n1412_r, k5[6], k4b[6] );
not U_inv1635 ( n1412_r, n1412 );
dff a5_k3a_reg_7_ ( clk, n1412_r, a5_k3a[7], a5_v3[7] );
not U_inv1636 ( n1412_r, n1412 );
dff a5_out_1_reg_7_ ( clk, n1412_r, k5[7], k4b[7] );
not U_inv1637 ( n1412_r, n1412 );
dff a5_k3a_reg_8_ ( clk, n1412_r, a5_k3a[8], a5_v3[8] );
not U_inv1638 ( n1412_r, n1412 );
dff a5_out_1_reg_8_ ( clk, n1412_r, k5[8], k4b[8] );
not U_inv1639 ( n1412_r, n1412 );
dff a5_k3a_reg_9_ ( clk, n1412_r, a5_k3a[9], a5_v3[9] );
not U_inv1640 ( n1412_r, n1412 );
dff a5_out_1_reg_9_ ( clk, n1412_r, k5[9], k4b[9] );
not U_inv1641 ( n1412_r, n1412 );
dff a5_k3a_reg_10_ ( clk, n1411_r, a5_k3a[10], a5_v3[10] );
not U_inv1642 ( n1411_r, n1411 );
dff a5_out_1_reg_10_ ( clk, n1411_r, k5[10], k4b[10] );
not U_inv1643 ( n1411_r, n1411 );
dff a5_k3a_reg_11_ ( clk, n1411_r, a5_k3a[11], a5_v3[11] );
not U_inv1644 ( n1411_r, n1411 );
dff a5_out_1_reg_11_ ( clk, n1411_r, k5[11], k4b[11] );
not U_inv1645 ( n1411_r, n1411 );
dff a5_k3a_reg_12_ ( clk, n1411_r, a5_k3a[12], a5_v3[12] );
not U_inv1646 ( n1411_r, n1411 );
dff a5_out_1_reg_12_ ( clk, n1411_r, k5[12], k4b[12] );
not U_inv1647 ( n1411_r, n1411 );
dff a5_k3a_reg_13_ ( clk, n1411_r, a5_k3a[13], a5_v3[13] );
not U_inv1648 ( n1411_r, n1411 );
dff a5_out_1_reg_13_ ( clk, n1411_r, k5[13], k4b[13] );
not U_inv1649 ( n1411_r, n1411 );
dff a5_k3a_reg_14_ ( clk, n1411_r, a5_k3a[14], a5_v3[14] );
not U_inv1650 ( n1411_r, n1411 );
dff a5_out_1_reg_14_ ( clk, n1411_r, k5[14], k4b[14] );
not U_inv1651 ( n1411_r, n1411 );
dff a5_k3a_reg_15_ ( clk, n1411_r, a5_k3a[15], a5_v3[15] );
not U_inv1652 ( n1411_r, n1411 );
dff a5_out_1_reg_15_ ( clk, n1411_r, k5[15], k4b[15] );
not U_inv1653 ( n1411_r, n1411 );
dff a5_k3a_reg_16_ ( clk, n1410_r, a5_k3a[16], a5_v3[16] );
not U_inv1654 ( n1410_r, n1410 );
dff a5_out_1_reg_16_ ( clk, n1410_r, k5[16], k4b[16] );
not U_inv1655 ( n1410_r, n1410 );
dff a5_k3a_reg_17_ ( clk, n1410_r, a5_k3a[17], a5_v3[17] );
not U_inv1656 ( n1410_r, n1410 );
dff a5_out_1_reg_17_ ( clk, n1410_r, k5[17], k4b[17] );
not U_inv1657 ( n1410_r, n1410 );
dff a5_k3a_reg_18_ ( clk, n1410_r, a5_k3a[18], a5_v3[18] );
not U_inv1658 ( n1410_r, n1410 );
dff a5_out_1_reg_18_ ( clk, n1410_r, k5[18], k4b[18] );
not U_inv1659 ( n1410_r, n1410 );
dff a5_k3a_reg_19_ ( clk, n1410_r, a5_k3a[19], a5_v3[19] );
not U_inv1660 ( n1410_r, n1410 );
dff a5_out_1_reg_19_ ( clk, n1410_r, k5[19], k4b[19] );
not U_inv1661 ( n1410_r, n1410 );
dff a5_k3a_reg_20_ ( clk, n1410_r, a5_k3a[20], a5_v3[20] );
not U_inv1662 ( n1410_r, n1410 );
dff a5_out_1_reg_20_ ( clk, n1410_r, k5[20], k4b[20] );
not U_inv1663 ( n1410_r, n1410 );
dff a5_k3a_reg_21_ ( clk, n1410_r, a5_k3a[21], a5_v3[21] );
not U_inv1664 ( n1410_r, n1410 );
dff a5_out_1_reg_21_ ( clk, n1410_r, k5[21], k4b[21] );
not U_inv1665 ( n1410_r, n1410 );
dff a5_k3a_reg_22_ ( clk, n1409_r, a5_k3a[22], a5_v3[22] );
not U_inv1666 ( n1409_r, n1409 );
dff a5_out_1_reg_22_ ( clk, n1409_r, k5[22], k4b[22] );
not U_inv1667 ( n1409_r, n1409 );
dff a5_k3a_reg_23_ ( clk, n1409_r, a5_k3a[23], a5_v3[23] );
not U_inv1668 ( n1409_r, n1409 );
dff a5_out_1_reg_23_ ( clk, n1409_r, k5[23], k4b[23] );
not U_inv1669 ( n1409_r, n1409 );
dff a5_k3a_reg_24_ ( clk, n1409_r, a5_k3a[24], a5_v3[24] );
not U_inv1670 ( n1409_r, n1409 );
dff a5_out_1_reg_24_ ( clk, n1409_r, k5[24], k4b[24] );
not U_inv1671 ( n1409_r, n1409 );
dff a5_k3a_reg_25_ ( clk, n1409_r, a5_k3a[25], a5_v3[25] );
not U_inv1672 ( n1409_r, n1409 );
dff a5_out_1_reg_25_ ( clk, n1409_r, k5[25], k4b[25] );
not U_inv1673 ( n1409_r, n1409 );
dff a5_k3a_reg_26_ ( clk, n1409_r, a5_k3a[26], a5_v3[26] );
not U_inv1674 ( n1409_r, n1409 );
dff a5_out_1_reg_26_ ( clk, n1409_r, k5[26], k4b[26] );
not U_inv1675 ( n1409_r, n1409 );
dff a5_k3a_reg_27_ ( clk, n1409_r, a5_k3a[27], a5_v3[27] );
not U_inv1676 ( n1409_r, n1409 );
dff a5_out_1_reg_27_ ( clk, n1409_r, k5[27], k4b[27] );
not U_inv1677 ( n1409_r, n1409 );
dff a5_k3a_reg_28_ ( clk, n1408_r, a5_k3a[28], a5_v3[28] );
not U_inv1678 ( n1408_r, n1408 );
dff a5_out_1_reg_28_ ( clk, n1408_r, k5[28], k4b[28] );
not U_inv1679 ( n1408_r, n1408 );
dff a5_k3a_reg_29_ ( clk, n1408_r, a5_k3a[29], a5_v3[29] );
not U_inv1680 ( n1408_r, n1408 );
dff a5_out_1_reg_29_ ( clk, n1408_r, k5[29], k4b[29] );
not U_inv1681 ( n1408_r, n1408 );
dff a5_k3a_reg_30_ ( clk, n1408_r, a5_k3a[30], a5_v3[30] );
not U_inv1682 ( n1408_r, n1408 );
dff a5_out_1_reg_30_ ( clk, n1408_r, k5[30], k4b[30] );
not U_inv1683 ( n1408_r, n1408 );
dff a5_k2a_reg_0_ ( clk, n1408_r, a5_k2a[0], a5_v2[0] );
not U_inv1684 ( n1408_r, n1408 );
dff a5_out_1_reg_32_ ( clk, n1408_r, k5[32], k4b[32] );
not U_inv1685 ( n1408_r, n1408 );
dff a5_k2a_reg_1_ ( clk, n1408_r, a5_k2a[1], a5_v2[1] );
not U_inv1686 ( n1408_r, n1408 );
dff a5_out_1_reg_33_ ( clk, n1408_r, k5[33], k4b[33] );
not U_inv1687 ( n1408_r, n1408 );
dff a5_k2a_reg_2_ ( clk, n1408_r, a5_k2a[2], a5_v2[2] );
not U_inv1688 ( n1408_r, n1408 );
dff a5_out_1_reg_34_ ( clk, n1408_r, k5[34], k4b[34] );
not U_inv1689 ( n1408_r, n1408 );
dff a5_k2a_reg_3_ ( clk, n1407_r, a5_k2a[3], a5_v2[3] );
not U_inv1690 ( n1407_r, n1407 );
dff a5_out_1_reg_35_ ( clk, n1407_r, k5[35], k4b[35] );
not U_inv1691 ( n1407_r, n1407 );
dff a5_k2a_reg_4_ ( clk, n1407_r, a5_k2a[4], a5_v2[4] );
not U_inv1692 ( n1407_r, n1407 );
dff a5_out_1_reg_36_ ( clk, n1407_r, k5[36], k4b[36] );
not U_inv1693 ( n1407_r, n1407 );
dff a5_k2a_reg_5_ ( clk, n1407_r, a5_k2a[5], a5_v2[5] );
not U_inv1694 ( n1407_r, n1407 );
dff a5_out_1_reg_37_ ( clk, n1407_r, k5[37], k4b[37] );
not U_inv1695 ( n1407_r, n1407 );
dff a5_k2a_reg_6_ ( clk, n1407_r, a5_k2a[6], a5_v2[6] );
not U_inv1696 ( n1407_r, n1407 );
dff a5_out_1_reg_38_ ( clk, n1407_r, k5[38], k4b[38] );
not U_inv1697 ( n1407_r, n1407 );
dff a5_k2a_reg_7_ ( clk, n1407_r, a5_k2a[7], a5_v2[7] );
not U_inv1698 ( n1407_r, n1407 );
dff a5_out_1_reg_39_ ( clk, n1407_r, k5[39], k4b[39] );
not U_inv1699 ( n1407_r, n1407 );
dff a5_k2a_reg_8_ ( clk, n1407_r, a5_k2a[8], a5_v2[8] );
not U_inv1700 ( n1407_r, n1407 );
dff a5_out_1_reg_40_ ( clk, n1407_r, k5[40], k4b[40] );
not U_inv1701 ( n1407_r, n1407 );
dff a5_k2a_reg_9_ ( clk, n1406_r, a5_k2a[9], a5_v2[9] );
not U_inv1702 ( n1406_r, n1406 );
dff a5_out_1_reg_41_ ( clk, n1406_r, k5[41], k4b[41] );
not U_inv1703 ( n1406_r, n1406 );
dff a5_k2a_reg_10_ ( clk, n1406_r, a5_k2a[10], a5_v2[10] );
not U_inv1704 ( n1406_r, n1406 );
dff a5_out_1_reg_42_ ( clk, n1406_r, k5[42], k4b[42] );
not U_inv1705 ( n1406_r, n1406 );
dff a5_k2a_reg_11_ ( clk, n1406_r, a5_k2a[11], a5_v2[11] );
not U_inv1706 ( n1406_r, n1406 );
dff a5_out_1_reg_43_ ( clk, n1406_r, k5[43], k4b[43] );
not U_inv1707 ( n1406_r, n1406 );
dff a5_k2a_reg_12_ ( clk, n1406_r, a5_k2a[12], a5_v2[12] );
not U_inv1708 ( n1406_r, n1406 );
dff a5_out_1_reg_44_ ( clk, n1406_r, k5[44], k4b[44] );
not U_inv1709 ( n1406_r, n1406 );
dff a5_k2a_reg_13_ ( clk, n1406_r, a5_k2a[13], a5_v2[13] );
not U_inv1710 ( n1406_r, n1406 );
dff a5_out_1_reg_45_ ( clk, n1406_r, k5[45], k4b[45] );
not U_inv1711 ( n1406_r, n1406 );
dff a5_k2a_reg_14_ ( clk, n1406_r, a5_k2a[14], a5_v2[14] );
not U_inv1712 ( n1406_r, n1406 );
dff a5_out_1_reg_46_ ( clk, n1406_r, k5[46], k4b[46] );
not U_inv1713 ( n1406_r, n1406 );
dff a5_k2a_reg_15_ ( clk, n1405_r, a5_k2a[15], a5_v2[15] );
not U_inv1714 ( n1405_r, n1405 );
dff a5_out_1_reg_47_ ( clk, n1405_r, k5[47], k4b[47] );
not U_inv1715 ( n1405_r, n1405 );
dff a5_k2a_reg_16_ ( clk, n1405_r, a5_k2a[16], a5_v2[16] );
not U_inv1716 ( n1405_r, n1405 );
dff a5_out_1_reg_48_ ( clk, n1405_r, k5[48], k4b[48] );
not U_inv1717 ( n1405_r, n1405 );
dff a5_k2a_reg_17_ ( clk, n1405_r, a5_k2a[17], a5_v2[17] );
not U_inv1718 ( n1405_r, n1405 );
dff a5_out_1_reg_49_ ( clk, n1405_r, k5[49], k4b[49] );
not U_inv1719 ( n1405_r, n1405 );
dff a5_k2a_reg_18_ ( clk, n1405_r, a5_k2a[18], a5_v2[18] );
not U_inv1720 ( n1405_r, n1405 );
dff a5_out_1_reg_50_ ( clk, n1405_r, k5[50], k4b[50] );
not U_inv1721 ( n1405_r, n1405 );
dff a5_k2a_reg_19_ ( clk, n1405_r, a5_k2a[19], a5_v2[19] );
not U_inv1722 ( n1405_r, n1405 );
dff a5_out_1_reg_51_ ( clk, n1405_r, k5[51], k4b[51] );
not U_inv1723 ( n1405_r, n1405 );
dff a5_k2a_reg_20_ ( clk, n1405_r, a5_k2a[20], a5_v2[20] );
not U_inv1724 ( n1405_r, n1405 );
dff a5_out_1_reg_52_ ( clk, n1405_r, k5[52], k4b[52] );
not U_inv1725 ( n1405_r, n1405 );
dff a5_k2a_reg_21_ ( clk, n1404_r, a5_k2a[21], a5_v2[21] );
not U_inv1726 ( n1404_r, n1404 );
dff a5_out_1_reg_53_ ( clk, n1404_r, k5[53], k4b[53] );
not U_inv1727 ( n1404_r, n1404 );
dff a5_k2a_reg_22_ ( clk, n1404_r, a5_k2a[22], a5_v2[22] );
not U_inv1728 ( n1404_r, n1404 );
dff a5_out_1_reg_54_ ( clk, n1404_r, k5[54], k4b[54] );
not U_inv1729 ( n1404_r, n1404 );
dff a5_k2a_reg_23_ ( clk, n1404_r, a5_k2a[23], a5_v2[23] );
not U_inv1730 ( n1404_r, n1404 );
dff a5_out_1_reg_55_ ( clk, n1404_r, k5[55], k4b[55] );
not U_inv1731 ( n1404_r, n1404 );
dff a5_k2a_reg_24_ ( clk, n1404_r, a5_k2a[24], a5_v2[24] );
not U_inv1732 ( n1404_r, n1404 );
dff a5_out_1_reg_56_ ( clk, n1404_r, k5[56], k4b[56] );
not U_inv1733 ( n1404_r, n1404 );
dff a5_k2a_reg_25_ ( clk, n1404_r, a5_k2a[25], a5_v2[25] );
not U_inv1734 ( n1404_r, n1404 );
dff a5_out_1_reg_57_ ( clk, n1404_r, k5[57], k4b[57] );
not U_inv1735 ( n1404_r, n1404 );
dff a5_k2a_reg_26_ ( clk, n1404_r, a5_k2a[26], a5_v2[26] );
not U_inv1736 ( n1404_r, n1404 );
dff a5_out_1_reg_58_ ( clk, n1404_r, k5[58], k4b[58] );
not U_inv1737 ( n1404_r, n1404 );
dff a5_k2a_reg_27_ ( clk, n1403_r, a5_k2a[27], a5_v2[27] );
not U_inv1738 ( n1403_r, n1403 );
dff a5_out_1_reg_59_ ( clk, n1403_r, k5[59], k4b[59] );
not U_inv1739 ( n1403_r, n1403 );
dff a5_k2a_reg_28_ ( clk, n1403_r, a5_k2a[28], a5_v2[28] );
not U_inv1740 ( n1403_r, n1403 );
dff a5_out_1_reg_60_ ( clk, n1403_r, k5[60], k4b[60] );
not U_inv1741 ( n1403_r, n1403 );
dff a5_k2a_reg_29_ ( clk, n1403_r, a5_k2a[29], a5_v2[29] );
not U_inv1742 ( n1403_r, n1403 );
dff a5_out_1_reg_61_ ( clk, n1403_r, k5[61], k4b[61] );
not U_inv1743 ( n1403_r, n1403 );
dff a5_k2a_reg_30_ ( clk, n1403_r, a5_k2a[30], a5_v2[30] );
not U_inv1744 ( n1403_r, n1403 );
dff a5_out_1_reg_62_ ( clk, n1403_r, k5[62], k4b[62] );
not U_inv1745 ( n1403_r, n1403 );
dff a5_k2a_reg_31_ ( clk, n1403_r, a5_k2a[31], a5_v2[31] );
not U_inv1746 ( n1403_r, n1403 );
dff a5_out_1_reg_63_ ( clk, n1403_r, k5[63], k4b[63] );
not U_inv1747 ( n1403_r, n1403 );
dff a5_k1a_reg_0_ ( clk, n1403_r, a5_k1a[0], a5_v1[0] );
not U_inv1748 ( n1403_r, n1403 );
dff a5_out_1_reg_64_ ( clk, n1403_r, ex_wire87, k4b[64] );
not U_inv1749 ( n803, ex_wire87 );
not U_inv1750 ( n1403_r, n1403 );
dff a5_k1a_reg_1_ ( clk, n1402_r, a5_k1a[1], a5_v1[1] );
not U_inv1751 ( n1402_r, n1402 );
dff a5_out_1_reg_65_ ( clk, n1402_r, ex_wire88, k4b[65] );
not U_inv1752 ( n814, ex_wire88 );
not U_inv1753 ( n1402_r, n1402 );
dff a5_k1a_reg_2_ ( clk, n1402_r, a5_k1a[2], a5_v1[2] );
not U_inv1754 ( n1402_r, n1402 );
dff a5_out_1_reg_66_ ( clk, n1402_r, ex_wire89, k4b[66] );
not U_inv1755 ( n824, ex_wire89 );
not U_inv1756 ( n1402_r, n1402 );
dff a5_k1a_reg_3_ ( clk, n1402_r, a5_k1a[3], a5_v1[3] );
not U_inv1757 ( n1402_r, n1402 );
dff a5_out_1_reg_67_ ( clk, n1402_r, ex_wire90, k4b[67] );
not U_inv1758 ( n827, ex_wire90 );
not U_inv1759 ( n1402_r, n1402 );
dff a5_k1a_reg_4_ ( clk, n1402_r, a5_k1a[4], a5_v1[4] );
not U_inv1760 ( n1402_r, n1402 );
dff a5_out_1_reg_68_ ( clk, n1402_r, k5[68], k4b[68] );
not U_inv1761 ( n1402_r, n1402 );
dff a5_k1a_reg_5_ ( clk, n1402_r, a5_k1a[5], a5_v1[5] );
not U_inv1762 ( n1402_r, n1402 );
dff a5_out_1_reg_69_ ( clk, n1402_r, k5[69], k4b[69] );
not U_inv1763 ( n1402_r, n1402 );
dff a5_k1a_reg_6_ ( clk, n1402_r, a5_k1a[6], a5_v1[6] );
not U_inv1764 ( n1402_r, n1402 );
dff a5_out_1_reg_70_ ( clk, n1402_r, k5[70], k4b[70] );
not U_inv1765 ( n1402_r, n1402 );
dff a5_k1a_reg_7_ ( clk, n1401_r, a5_k1a[7], a5_v1[7] );
not U_inv1766 ( n1401_r, n1401 );
dff a5_out_1_reg_71_ ( clk, n1401_r, k5[71], k4b[71] );
not U_inv1767 ( n1401_r, n1401 );
dff a5_k1a_reg_8_ ( clk, n1401_r, a5_k1a[8], a5_v1[8] );
not U_inv1768 ( n1401_r, n1401 );
dff a5_out_1_reg_72_ ( clk, n1401_r, k5[72], k4b[72] );
not U_inv1769 ( n1401_r, n1401 );
dff a5_k1a_reg_9_ ( clk, n1401_r, a5_k1a[9], a5_v1[9] );
not U_inv1770 ( n1401_r, n1401 );
dff a5_out_1_reg_73_ ( clk, n1401_r, k5[73], k4b[73] );
not U_inv1771 ( n1401_r, n1401 );
dff a5_k1a_reg_10_ ( clk, n1401_r, a5_k1a[10], a5_v1[10] );
not U_inv1772 ( n1401_r, n1401 );
dff a5_out_1_reg_74_ ( clk, n1401_r, k5[74], k4b[74] );
not U_inv1773 ( n1401_r, n1401 );
dff a5_k1a_reg_11_ ( clk, n1401_r, a5_k1a[11], a5_v1[11] );
not U_inv1774 ( n1401_r, n1401 );
dff a5_out_1_reg_75_ ( clk, n1401_r, k5[75], k4b[75] );
not U_inv1775 ( n1401_r, n1401 );
dff a5_k1a_reg_12_ ( clk, n1401_r, a5_k1a[12], a5_v1[12] );
not U_inv1776 ( n1401_r, n1401 );
dff a5_out_1_reg_76_ ( clk, n1401_r, k5[76], k4b[76] );
not U_inv1777 ( n1401_r, n1401 );
dff a5_k1a_reg_13_ ( clk, n1400_r, a5_k1a[13], a5_v1[13] );
not U_inv1778 ( n1400_r, n1400 );
dff a5_out_1_reg_77_ ( clk, n1400_r, k5[77], k4b[77] );
not U_inv1779 ( n1400_r, n1400 );
dff a5_k1a_reg_14_ ( clk, n1400_r, a5_k1a[14], a5_v1[14] );
not U_inv1780 ( n1400_r, n1400 );
dff a5_out_1_reg_78_ ( clk, n1400_r, k5[78], k4b[78] );
not U_inv1781 ( n1400_r, n1400 );
dff a5_k1a_reg_15_ ( clk, n1400_r, a5_k1a[15], a5_v1[15] );
not U_inv1782 ( n1400_r, n1400 );
dff a5_out_1_reg_79_ ( clk, n1400_r, k5[79], k4b[79] );
not U_inv1783 ( n1400_r, n1400 );
dff a5_k1a_reg_16_ ( clk, n1400_r, a5_k1a[16], a5_v1[16] );
not U_inv1784 ( n1400_r, n1400 );
dff a5_out_1_reg_80_ ( clk, n1400_r, k5[80], k4b[80] );
not U_inv1785 ( n1400_r, n1400 );
dff a5_k1a_reg_17_ ( clk, n1400_r, a5_k1a[17], a5_v1[17] );
not U_inv1786 ( n1400_r, n1400 );
dff a5_out_1_reg_81_ ( clk, n1400_r, k5[81], k4b[81] );
not U_inv1787 ( n1400_r, n1400 );
dff a5_k1a_reg_18_ ( clk, n1400_r, a5_k1a[18], a5_v1[18] );
not U_inv1788 ( n1400_r, n1400 );
dff a5_out_1_reg_82_ ( clk, n1400_r, k5[82], k4b[82] );
not U_inv1789 ( n1400_r, n1400 );
dff a5_k1a_reg_19_ ( clk, n1399_r, a5_k1a[19], a5_v1[19] );
not U_inv1790 ( n1399_r, n1399 );
dff a5_out_1_reg_83_ ( clk, n1399_r, k5[83], k4b[83] );
not U_inv1791 ( n1399_r, n1399 );
dff a5_k1a_reg_20_ ( clk, n1399_r, a5_k1a[20], a5_v1[20] );
not U_inv1792 ( n1399_r, n1399 );
dff a5_out_1_reg_84_ ( clk, n1399_r, k5[84], k4b[84] );
not U_inv1793 ( n1399_r, n1399 );
dff a5_k1a_reg_21_ ( clk, n1399_r, a5_k1a[21], a5_v1[21] );
not U_inv1794 ( n1399_r, n1399 );
dff a5_out_1_reg_85_ ( clk, n1399_r, k5[85], k4b[85] );
not U_inv1795 ( n1399_r, n1399 );
dff a5_k1a_reg_22_ ( clk, n1399_r, a5_k1a[22], a5_v1[22] );
not U_inv1796 ( n1399_r, n1399 );
dff a5_out_1_reg_86_ ( clk, n1399_r, k5[86], k4b[86] );
not U_inv1797 ( n1399_r, n1399 );
dff a5_k1a_reg_23_ ( clk, n1399_r, a5_k1a[23], a5_v1[23] );
not U_inv1798 ( n1399_r, n1399 );
dff a5_out_1_reg_87_ ( clk, n1399_r, k5[87], k4b[87] );
not U_inv1799 ( n1399_r, n1399 );
dff a5_k1a_reg_24_ ( clk, n1399_r, a5_k1a[24], a5_v1[24] );
not U_inv1800 ( n1399_r, n1399 );
dff a5_out_1_reg_88_ ( clk, n1399_r, k5[88], k4b[88] );
not U_inv1801 ( n1399_r, n1399 );
dff a5_k1a_reg_25_ ( clk, n1398_r, a5_k1a[25], a5_v1[25] );
not U_inv1802 ( n1398_r, n1398 );
dff a5_out_1_reg_89_ ( clk, n1398_r, k5[89], k4b[89] );
not U_inv1803 ( n1398_r, n1398 );
dff a5_k1a_reg_26_ ( clk, n1398_r, a5_k1a[26], a5_v1[26] );
not U_inv1804 ( n1398_r, n1398 );
dff a5_out_1_reg_90_ ( clk, n1398_r, k5[90], k4b[90] );
not U_inv1805 ( n1398_r, n1398 );
dff a5_k1a_reg_27_ ( clk, n1398_r, a5_k1a[27], a5_v1[27] );
not U_inv1806 ( n1398_r, n1398 );
dff a5_out_1_reg_91_ ( clk, n1398_r, k5[91], k4b[91] );
not U_inv1807 ( n1398_r, n1398 );
dff a5_k1a_reg_28_ ( clk, n1398_r, a5_k1a[28], a5_v1[28] );
not U_inv1808 ( n1398_r, n1398 );
dff a5_out_1_reg_92_ ( clk, n1398_r, k5[92], k4b[92] );
not U_inv1809 ( n1398_r, n1398 );
dff a5_k1a_reg_29_ ( clk, n1398_r, a5_k1a[29], a5_v1[29] );
not U_inv1810 ( n1398_r, n1398 );
dff a5_out_1_reg_93_ ( clk, n1398_r, k5[93], k4b[93] );
not U_inv1811 ( n1398_r, n1398 );
dff a5_k1a_reg_30_ ( clk, n1398_r, a5_k1a[30], a5_v1[30] );
not U_inv1812 ( n1398_r, n1398 );
dff a5_out_1_reg_94_ ( clk, n1398_r, k5[94], k4b[94] );
not U_inv1813 ( n1398_r, n1398 );
dff a5_out_1_reg_95_ ( clk, n1397_r, k5[95], k4b[95] );
not U_inv1814 ( n1397_r, n1397 );
dff a6_k0a_reg_0_ ( clk, n1397_r, a6_k0a[0], k5[96] );
not U_inv1815 ( n1397_r, n1397 );
dff a6_out_1_reg_96_ ( clk, n1397_r, k6[96], k5b[96] );
not U_inv1816 ( n1397_r, n1397 );
dff a6_k0a_reg_1_ ( clk, n1397_r, a6_k0a[1], k5[97] );
not U_inv1817 ( n1397_r, n1397 );
dff a6_out_1_reg_97_ ( clk, n1397_r, k6[97], k5b[97] );
not U_inv1818 ( n1397_r, n1397 );
dff a6_k0a_reg_2_ ( clk, n1397_r, a6_k0a[2], k5[98] );
not U_inv1819 ( n1397_r, n1397 );
dff a6_out_1_reg_98_ ( clk, n1397_r, k6[98], k5b[98] );
not U_inv1820 ( n1397_r, n1397 );
dff a6_k0a_reg_3_ ( clk, n1397_r, a6_k0a[3], k5[99] );
not U_inv1821 ( n1397_r, n1397 );
dff a6_out_1_reg_99_ ( clk, n1397_r, k6[99], k5b[99] );
not U_inv1822 ( n1397_r, n1397 );
dff a6_k0a_reg_4_ ( clk, n1397_r, a6_k0a[4], k5[100] );
not U_inv1823 ( n1397_r, n1397 );
dff a6_out_1_reg_100_ ( clk, n1397_r, k6[100], k5b[100] );
not U_inv1824 ( n859, k6[100] );
not U_inv1825 ( n1397_r, n1397 );
dff a6_k0a_reg_5_ ( clk, n1397_r, a6_k0a[5], k5[101] );
not U_inv1826 ( n1397_r, n1397 );
dff a6_out_1_reg_101_ ( clk, n1396_r, k6[101], k5b[101] );
not U_inv1827 ( n860, k6[101] );
not U_inv1828 ( n1396_r, n1396 );
dff a6_k0a_reg_6_ ( clk, n1396_r, a6_k0a[6], k5[102] );
not U_inv1829 ( n1396_r, n1396 );
dff a6_out_1_reg_102_ ( clk, n1396_r, k6[102], k5b[102] );
not U_inv1830 ( n861, k6[102] );
not U_inv1831 ( n1396_r, n1396 );
dff a6_k0a_reg_7_ ( clk, n1396_r, a6_k0a[7], k5[103] );
not U_inv1832 ( n1396_r, n1396 );
dff a6_out_1_reg_103_ ( clk, n1396_r, k6[103], k5b[103] );
not U_inv1833 ( n862, k6[103] );
not U_inv1834 ( n1396_r, n1396 );
dff a6_k0a_reg_8_ ( clk, n1396_r, a6_k0a[8], k5[104] );
not U_inv1835 ( n1396_r, n1396 );
dff a6_out_1_reg_104_ ( clk, n1396_r, k6[104], k5b[104] );
not U_inv1836 ( n863, k6[104] );
not U_inv1837 ( n1396_r, n1396 );
dff a6_k0a_reg_9_ ( clk, n1396_r, a6_k0a[9], k5[105] );
not U_inv1838 ( n1396_r, n1396 );
dff a6_out_1_reg_105_ ( clk, n1396_r, k6[105], k5b[105] );
not U_inv1839 ( n864, k6[105] );
not U_inv1840 ( n1396_r, n1396 );
dff a6_k0a_reg_10_ ( clk, n1396_r, a6_k0a[10], k5[106] );
not U_inv1841 ( n1396_r, n1396 );
dff a6_out_1_reg_106_ ( clk, n1396_r, k6[106], k5b[106] );
not U_inv1842 ( n835, k6[106] );
not U_inv1843 ( n1396_r, n1396 );
dff a6_k0a_reg_11_ ( clk, n1396_r, a6_k0a[11], k5[107] );
not U_inv1844 ( n1396_r, n1396 );
dff a6_out_1_reg_107_ ( clk, n1395_r, k6[107], k5b[107] );
not U_inv1845 ( n836, k6[107] );
not U_inv1846 ( n1395_r, n1395 );
dff a6_k0a_reg_12_ ( clk, n1395_r, a6_k0a[12], k5[108] );
not U_inv1847 ( n1395_r, n1395 );
dff a6_out_1_reg_108_ ( clk, n1395_r, k6[108], k5b[108] );
not U_inv1848 ( n837, k6[108] );
not U_inv1849 ( n1395_r, n1395 );
dff a6_k0a_reg_13_ ( clk, n1395_r, a6_k0a[13], k5[109] );
not U_inv1850 ( n1395_r, n1395 );
dff a6_out_1_reg_109_ ( clk, n1395_r, k6[109], k5b[109] );
not U_inv1851 ( n838, k6[109] );
not U_inv1852 ( n1395_r, n1395 );
dff a6_k0a_reg_14_ ( clk, n1395_r, a6_k0a[14], k5[110] );
not U_inv1853 ( n1395_r, n1395 );
dff a6_out_1_reg_110_ ( clk, n1395_r, k6[110], k5b[110] );
not U_inv1854 ( n839, k6[110] );
not U_inv1855 ( n1395_r, n1395 );
dff a6_k0a_reg_15_ ( clk, n1395_r, a6_k0a[15], k5[111] );
not U_inv1856 ( n1395_r, n1395 );
dff a6_out_1_reg_111_ ( clk, n1395_r, k6[111], k5b[111] );
not U_inv1857 ( n840, k6[111] );
not U_inv1858 ( n1395_r, n1395 );
dff a6_k0a_reg_16_ ( clk, n1395_r, a6_k0a[16], k5[112] );
not U_inv1859 ( n1395_r, n1395 );
dff a6_out_1_reg_112_ ( clk, n1395_r, k6[112], k5b[112] );
not U_inv1860 ( n841, k6[112] );
not U_inv1861 ( n1395_r, n1395 );
dff a6_k0a_reg_17_ ( clk, n1395_r, a6_k0a[17], k5[113] );
not U_inv1862 ( n1395_r, n1395 );
dff a6_out_1_reg_113_ ( clk, n1394_r, k6[113], k5b[113] );
not U_inv1863 ( n842, k6[113] );
not U_inv1864 ( n1394_r, n1394 );
dff a6_k0a_reg_18_ ( clk, n1394_r, a6_k0a[18], k5[114] );
not U_inv1865 ( n1394_r, n1394 );
dff a6_out_1_reg_114_ ( clk, n1394_r, k6[114], k5b[114] );
not U_inv1866 ( n843, k6[114] );
not U_inv1867 ( n1394_r, n1394 );
dff a6_k0a_reg_19_ ( clk, n1394_r, a6_k0a[19], k5[115] );
not U_inv1868 ( n1394_r, n1394 );
dff a6_out_1_reg_115_ ( clk, n1394_r, k6[115], k5b[115] );
not U_inv1869 ( n844, k6[115] );
not U_inv1870 ( n1394_r, n1394 );
dff a6_k0a_reg_20_ ( clk, n1394_r, a6_k0a[20], k5[116] );
not U_inv1871 ( n1394_r, n1394 );
dff a6_out_1_reg_116_ ( clk, n1394_r, k6[116], k5b[116] );
not U_inv1872 ( n846, k6[116] );
not U_inv1873 ( n1394_r, n1394 );
dff a6_k0a_reg_21_ ( clk, n1394_r, a6_k0a[21], k5[117] );
not U_inv1874 ( n1394_r, n1394 );
dff a6_out_1_reg_117_ ( clk, n1394_r, k6[117], k5b[117] );
not U_inv1875 ( n847, k6[117] );
not U_inv1876 ( n1394_r, n1394 );
dff a6_k0a_reg_22_ ( clk, n1394_r, a6_k0a[22], k5[118] );
not U_inv1877 ( n1394_r, n1394 );
dff a6_out_1_reg_118_ ( clk, n1394_r, k6[118], k5b[118] );
not U_inv1878 ( n848, k6[118] );
not U_inv1879 ( n1394_r, n1394 );
dff a6_k0a_reg_23_ ( clk, n1394_r, a6_k0a[23], k5[119] );
not U_inv1880 ( n1394_r, n1394 );
dff a6_out_1_reg_119_ ( clk, n1393_r, k6[119], k5b[119] );
not U_inv1881 ( n849, k6[119] );
not U_inv1882 ( n1393_r, n1393 );
dff a6_k0a_reg_24_ ( clk, n1393_r, a6_k0a[24], k5[120] );
not U_inv1883 ( n1393_r, n1393 );
dff a6_out_1_reg_120_ ( clk, n1393_r, k6[120], k5b[120] );
not U_inv1884 ( n850, k6[120] );
not U_inv1885 ( n1393_r, n1393 );
dff a6_k0a_reg_25_ ( clk, n1393_r, a6_k0a[25], k5[121] );
not U_inv1886 ( n1393_r, n1393 );
dff a6_out_1_reg_121_ ( clk, n1393_r, k6[121], k5b[121] );
not U_inv1887 ( n851, k6[121] );
not U_inv1888 ( n1393_r, n1393 );
dff a6_k0a_reg_26_ ( clk, n1393_r, a6_k0a[26], k5[122] );
not U_inv1889 ( n1393_r, n1393 );
dff a6_out_1_reg_122_ ( clk, n1393_r, k6[122], k5b[122] );
not U_inv1890 ( n852, k6[122] );
not U_inv1891 ( n1393_r, n1393 );
dff a6_k0a_reg_27_ ( clk, n1393_r, a6_k0a[27], k5[123] );
not U_inv1892 ( n1393_r, n1393 );
dff a6_out_1_reg_123_ ( clk, n1393_r, k6[123], k5b[123] );
not U_inv1893 ( n853, k6[123] );
not U_inv1894 ( n1393_r, n1393 );
dff a6_k0a_reg_28_ ( clk, n1393_r, a6_k0a[28], k5[124] );
not U_inv1895 ( n1393_r, n1393 );
dff a6_out_1_reg_124_ ( clk, n1393_r, k6[124], k5b[124] );
not U_inv1896 ( n854, k6[124] );
not U_inv1897 ( n1393_r, n1393 );
dff a6_k0a_reg_29_ ( clk, n1393_r, a6_k0a[29], n1289 );
not U_inv1898 ( n1393_r, n1393 );
dff a6_out_1_reg_125_ ( clk, n1392_r, k6[125], k5b[125] );
not U_inv1899 ( n855, k6[125] );
not U_inv1900 ( n1392_r, n1392 );
dff a6_k0a_reg_30_ ( clk, n1392_r, a6_k0a[30], k5[126] );
not U_inv1901 ( n1392_r, n1392 );
dff a6_out_1_reg_126_ ( clk, n1392_r, ex_wire91, k5b[126] );
not U_inv1902 ( n1290, ex_wire91 );
not U_inv1903 ( n1392_r, n1392 );
dff a6_k0a_reg_31_ ( clk, n1392_r, a6_k0a[31], k5[127] );
not U_inv1904 ( n1392_r, n1392 );
dff a6_out_1_reg_127_ ( clk, n1392_r, k6[127], k5b[127] );
not U_inv1905 ( n857, k6[127] );
not U_inv1906 ( n1392_r, n1392 );
dff a6_k3a_reg_0_ ( clk, n1392_r, a6_k3a[0], a6_v3[0] );
not U_inv1907 ( n1392_r, n1392 );
dff a6_out_1_reg_0_ ( clk, n1392_r, k6[0], k5b[0] );
not U_inv1908 ( n1392_r, n1392 );
dff a6_k3a_reg_1_ ( clk, n1392_r, a6_k3a[1], a6_v3[1] );
not U_inv1909 ( n1392_r, n1392 );
dff a6_out_1_reg_1_ ( clk, n1392_r, k6[1], k5b[1] );
not U_inv1910 ( n1392_r, n1392 );
dff a6_k3a_reg_2_ ( clk, n1392_r, a6_k3a[2], a6_v3[2] );
not U_inv1911 ( n1392_r, n1392 );
dff a6_out_1_reg_2_ ( clk, n1392_r, k6[2], k5b[2] );
not U_inv1912 ( n1392_r, n1392 );
dff a6_k3a_reg_3_ ( clk, n1392_r, a6_k3a[3], a6_v3[3] );
not U_inv1913 ( n1392_r, n1392 );
dff a6_out_1_reg_3_ ( clk, n1391_r, k6[3], k5b[3] );
not U_inv1914 ( n1391_r, n1391 );
dff a6_k3a_reg_4_ ( clk, n1391_r, a6_k3a[4], a6_v3[4] );
not U_inv1915 ( n1391_r, n1391 );
dff a6_out_1_reg_4_ ( clk, n1391_r, k6[4], k5b[4] );
not U_inv1916 ( n1391_r, n1391 );
dff a6_k3a_reg_5_ ( clk, n1391_r, a6_k3a[5], a6_v3[5] );
not U_inv1917 ( n1391_r, n1391 );
dff a6_out_1_reg_5_ ( clk, n1391_r, k6[5], k5b[5] );
not U_inv1918 ( n1391_r, n1391 );
dff a6_k3a_reg_6_ ( clk, n1391_r, a6_k3a[6], a6_v3[6] );
not U_inv1919 ( n1391_r, n1391 );
dff a6_out_1_reg_6_ ( clk, n1391_r, k6[6], k5b[6] );
not U_inv1920 ( n1391_r, n1391 );
dff a6_k3a_reg_7_ ( clk, n1391_r, a6_k3a[7], a6_v3[7] );
not U_inv1921 ( n1391_r, n1391 );
dff a6_out_1_reg_7_ ( clk, n1391_r, k6[7], k5b[7] );
not U_inv1922 ( n1391_r, n1391 );
dff a6_k3a_reg_8_ ( clk, n1391_r, a6_k3a[8], a6_v3[8] );
not U_inv1923 ( n1391_r, n1391 );
dff a6_out_1_reg_8_ ( clk, n1391_r, k6[8], k5b[8] );
not U_inv1924 ( n1391_r, n1391 );
dff a6_k3a_reg_9_ ( clk, n1391_r, a6_k3a[9], a6_v3[9] );
not U_inv1925 ( n1391_r, n1391 );
dff a6_out_1_reg_9_ ( clk, n1390_r, k6[9], k5b[9] );
not U_inv1926 ( n1390_r, n1390 );
dff a6_k3a_reg_10_ ( clk, n1390_r, a6_k3a[10], a6_v3[10] );
not U_inv1927 ( n1390_r, n1390 );
dff a6_out_1_reg_10_ ( clk, n1390_r, k6[10], k5b[10] );
not U_inv1928 ( n1390_r, n1390 );
dff a6_k3a_reg_11_ ( clk, n1390_r, a6_k3a[11], a6_v3[11] );
not U_inv1929 ( n1390_r, n1390 );
dff a6_out_1_reg_11_ ( clk, n1390_r, k6[11], k5b[11] );
not U_inv1930 ( n1390_r, n1390 );
dff a6_k3a_reg_12_ ( clk, n1390_r, a6_k3a[12], a6_v3[12] );
not U_inv1931 ( n1390_r, n1390 );
dff a6_out_1_reg_12_ ( clk, n1390_r, k6[12], k5b[12] );
not U_inv1932 ( n1390_r, n1390 );
dff a6_k3a_reg_13_ ( clk, n1390_r, a6_k3a[13], a6_v3[13] );
not U_inv1933 ( n1390_r, n1390 );
dff a6_out_1_reg_13_ ( clk, n1390_r, k6[13], k5b[13] );
not U_inv1934 ( n1390_r, n1390 );
dff a6_k3a_reg_14_ ( clk, n1390_r, a6_k3a[14], a6_v3[14] );
not U_inv1935 ( n1390_r, n1390 );
dff a6_out_1_reg_14_ ( clk, n1390_r, k6[14], k5b[14] );
not U_inv1936 ( n1390_r, n1390 );
dff a6_k3a_reg_15_ ( clk, n1390_r, a6_k3a[15], a6_v3[15] );
not U_inv1937 ( n1390_r, n1390 );
dff a6_out_1_reg_15_ ( clk, n1389_r, k6[15], k5b[15] );
not U_inv1938 ( n1389_r, n1389 );
dff a6_k3a_reg_16_ ( clk, n1389_r, a6_k3a[16], a6_v3[16] );
not U_inv1939 ( n1389_r, n1389 );
dff a6_out_1_reg_16_ ( clk, n1389_r, k6[16], k5b[16] );
not U_inv1940 ( n1389_r, n1389 );
dff a6_k3a_reg_17_ ( clk, n1389_r, a6_k3a[17], a6_v3[17] );
not U_inv1941 ( n1389_r, n1389 );
dff a6_out_1_reg_17_ ( clk, n1389_r, k6[17], k5b[17] );
not U_inv1942 ( n1389_r, n1389 );
dff a6_k3a_reg_18_ ( clk, n1389_r, a6_k3a[18], a6_v3[18] );
not U_inv1943 ( n1389_r, n1389 );
dff a6_out_1_reg_18_ ( clk, n1389_r, k6[18], k5b[18] );
not U_inv1944 ( n1389_r, n1389 );
dff a6_k3a_reg_19_ ( clk, n1389_r, a6_k3a[19], a6_v3[19] );
not U_inv1945 ( n1389_r, n1389 );
dff a6_out_1_reg_19_ ( clk, n1389_r, k6[19], k5b[19] );
not U_inv1946 ( n1389_r, n1389 );
dff a6_k3a_reg_20_ ( clk, n1389_r, a6_k3a[20], a6_v3[20] );
not U_inv1947 ( n1389_r, n1389 );
dff a6_out_1_reg_20_ ( clk, n1389_r, k6[20], k5b[20] );
not U_inv1948 ( n1389_r, n1389 );
dff a6_k3a_reg_21_ ( clk, n1389_r, a6_k3a[21], a6_v3[21] );
not U_inv1949 ( n1389_r, n1389 );
dff a6_out_1_reg_21_ ( clk, n1388_r, k6[21], k5b[21] );
not U_inv1950 ( n1388_r, n1388 );
dff a6_k3a_reg_22_ ( clk, n1388_r, a6_k3a[22], a6_v3[22] );
not U_inv1951 ( n1388_r, n1388 );
dff a6_out_1_reg_22_ ( clk, n1388_r, k6[22], k5b[22] );
not U_inv1952 ( n1388_r, n1388 );
dff a6_k3a_reg_23_ ( clk, n1388_r, a6_k3a[23], a6_v3[23] );
not U_inv1953 ( n1388_r, n1388 );
dff a6_out_1_reg_23_ ( clk, n1388_r, k6[23], k5b[23] );
not U_inv1954 ( n1388_r, n1388 );
dff a6_k3a_reg_24_ ( clk, n1388_r, a6_k3a[24], a6_v3[24] );
not U_inv1955 ( n1388_r, n1388 );
dff a6_out_1_reg_24_ ( clk, n1388_r, k6[24], k5b[24] );
not U_inv1956 ( n1388_r, n1388 );
dff a6_k3a_reg_25_ ( clk, n1388_r, a6_k3a[25], a6_v3[25] );
not U_inv1957 ( n1388_r, n1388 );
dff a6_out_1_reg_25_ ( clk, n1388_r, k6[25], k5b[25] );
not U_inv1958 ( n1388_r, n1388 );
dff a6_k3a_reg_26_ ( clk, n1388_r, a6_k3a[26], a6_v3[26] );
not U_inv1959 ( n1388_r, n1388 );
dff a6_out_1_reg_26_ ( clk, n1388_r, k6[26], k5b[26] );
not U_inv1960 ( n1388_r, n1388 );
dff a6_k3a_reg_27_ ( clk, n1388_r, a6_k3a[27], a6_v3[27] );
not U_inv1961 ( n1388_r, n1388 );
dff a6_out_1_reg_27_ ( clk, n1387_r, k6[27], k5b[27] );
not U_inv1962 ( n1387_r, n1387 );
dff a6_k3a_reg_28_ ( clk, n1387_r, a6_k3a[28], a6_v3[28] );
not U_inv1963 ( n1387_r, n1387 );
dff a6_out_1_reg_28_ ( clk, n1387_r, k6[28], k5b[28] );
not U_inv1964 ( n1387_r, n1387 );
dff a6_k3a_reg_29_ ( clk, n1387_r, a6_k3a[29], a6_v3[29] );
not U_inv1965 ( n1387_r, n1387 );
dff a6_out_1_reg_29_ ( clk, n1387_r, k6[29], k5b[29] );
not U_inv1966 ( n1387_r, n1387 );
dff a6_k3a_reg_30_ ( clk, n1387_r, a6_k3a[30], a6_v3[30] );
not U_inv1967 ( n1387_r, n1387 );
dff a6_out_1_reg_30_ ( clk, n1387_r, k6[30], k5b[30] );
not U_inv1968 ( n1387_r, n1387 );
dff a6_k2a_reg_0_ ( clk, n1387_r, a6_k2a[0], a6_v2[0] );
not U_inv1969 ( n1387_r, n1387 );
dff a6_out_1_reg_32_ ( clk, n1387_r, k6[32], k5b[32] );
not U_inv1970 ( n1387_r, n1387 );
dff a6_k2a_reg_1_ ( clk, n1387_r, a6_k2a[1], a6_v2[1] );
not U_inv1971 ( n1387_r, n1387 );
dff a6_out_1_reg_33_ ( clk, n1387_r, k6[33], k5b[33] );
not U_inv1972 ( n1387_r, n1387 );
dff a6_k2a_reg_2_ ( clk, n1387_r, a6_k2a[2], a6_v2[2] );
not U_inv1973 ( n1387_r, n1387 );
dff a6_out_1_reg_34_ ( clk, n1386_r, k6[34], k5b[34] );
not U_inv1974 ( n1386_r, n1386 );
dff a6_k2a_reg_3_ ( clk, n1386_r, a6_k2a[3], a6_v2[3] );
not U_inv1975 ( n1386_r, n1386 );
dff a6_out_1_reg_35_ ( clk, n1386_r, k6[35], k5b[35] );
not U_inv1976 ( n1386_r, n1386 );
dff a6_k2a_reg_4_ ( clk, n1386_r, a6_k2a[4], a6_v2[4] );
not U_inv1977 ( n1386_r, n1386 );
dff a6_out_1_reg_36_ ( clk, n1386_r, k6[36], k5b[36] );
not U_inv1978 ( n1386_r, n1386 );
dff a6_k2a_reg_5_ ( clk, n1386_r, a6_k2a[5], a6_v2[5] );
not U_inv1979 ( n1386_r, n1386 );
dff a6_out_1_reg_37_ ( clk, n1386_r, k6[37], k5b[37] );
not U_inv1980 ( n1386_r, n1386 );
dff a6_k2a_reg_6_ ( clk, n1386_r, a6_k2a[6], a6_v2[6] );
not U_inv1981 ( n1386_r, n1386 );
dff a6_out_1_reg_38_ ( clk, n1386_r, k6[38], k5b[38] );
not U_inv1982 ( n1386_r, n1386 );
dff a6_k2a_reg_7_ ( clk, n1386_r, a6_k2a[7], a6_v2[7] );
not U_inv1983 ( n1386_r, n1386 );
dff a6_out_1_reg_39_ ( clk, n1386_r, k6[39], k5b[39] );
not U_inv1984 ( n1386_r, n1386 );
dff a6_k2a_reg_8_ ( clk, n1386_r, a6_k2a[8], a6_v2[8] );
not U_inv1985 ( n1386_r, n1386 );
dff a6_out_1_reg_40_ ( clk, n1385_r, k6[40], k5b[40] );
not U_inv1986 ( n1385_r, n1385 );
dff a6_k2a_reg_9_ ( clk, n1385_r, a6_k2a[9], a6_v2[9] );
not U_inv1987 ( n1385_r, n1385 );
dff a6_out_1_reg_41_ ( clk, n1385_r, k6[41], k5b[41] );
not U_inv1988 ( n1385_r, n1385 );
dff a6_k2a_reg_10_ ( clk, n1385_r, a6_k2a[10], a6_v2[10] );
not U_inv1989 ( n1385_r, n1385 );
dff a6_out_1_reg_42_ ( clk, n1385_r, k6[42], k5b[42] );
not U_inv1990 ( n1385_r, n1385 );
dff a6_k2a_reg_11_ ( clk, n1385_r, a6_k2a[11], a6_v2[11] );
not U_inv1991 ( n1385_r, n1385 );
dff a6_out_1_reg_43_ ( clk, n1385_r, k6[43], k5b[43] );
not U_inv1992 ( n1385_r, n1385 );
dff a6_k2a_reg_12_ ( clk, n1385_r, a6_k2a[12], a6_v2[12] );
not U_inv1993 ( n1385_r, n1385 );
dff a6_out_1_reg_44_ ( clk, n1385_r, k6[44], k5b[44] );
not U_inv1994 ( n1385_r, n1385 );
dff a6_k2a_reg_13_ ( clk, n1385_r, a6_k2a[13], a6_v2[13] );
not U_inv1995 ( n1385_r, n1385 );
dff a6_out_1_reg_45_ ( clk, n1385_r, k6[45], k5b[45] );
not U_inv1996 ( n1385_r, n1385 );
dff a6_k2a_reg_14_ ( clk, n1385_r, a6_k2a[14], a6_v2[14] );
not U_inv1997 ( n1385_r, n1385 );
dff a6_out_1_reg_46_ ( clk, n1384_r, k6[46], k5b[46] );
not U_inv1998 ( n1384_r, n1384 );
dff a6_k2a_reg_15_ ( clk, n1384_r, a6_k2a[15], a6_v2[15] );
not U_inv1999 ( n1384_r, n1384 );
dff a6_out_1_reg_47_ ( clk, n1384_r, k6[47], k5b[47] );
not U_inv2000 ( n1384_r, n1384 );
dff a6_k2a_reg_16_ ( clk, n1384_r, a6_k2a[16], a6_v2[16] );
not U_inv2001 ( n1384_r, n1384 );
dff a6_out_1_reg_48_ ( clk, n1384_r, k6[48], k5b[48] );
not U_inv2002 ( n1384_r, n1384 );
dff a6_k2a_reg_17_ ( clk, n1384_r, a6_k2a[17], a6_v2[17] );
not U_inv2003 ( n1384_r, n1384 );
dff a6_out_1_reg_49_ ( clk, n1384_r, k6[49], k5b[49] );
not U_inv2004 ( n1384_r, n1384 );
dff a6_k2a_reg_18_ ( clk, n1384_r, a6_k2a[18], a6_v2[18] );
not U_inv2005 ( n1384_r, n1384 );
dff a6_out_1_reg_50_ ( clk, n1384_r, k6[50], k5b[50] );
not U_inv2006 ( n1384_r, n1384 );
dff a6_k2a_reg_19_ ( clk, n1384_r, a6_k2a[19], a6_v2[19] );
not U_inv2007 ( n1384_r, n1384 );
dff a6_out_1_reg_51_ ( clk, n1384_r, k6[51], k5b[51] );
not U_inv2008 ( n1384_r, n1384 );
dff a6_k2a_reg_20_ ( clk, n1384_r, a6_k2a[20], a6_v2[20] );
not U_inv2009 ( n1384_r, n1384 );
dff a6_out_1_reg_52_ ( clk, n1383_r, k6[52], k5b[52] );
not U_inv2010 ( n1383_r, n1383 );
dff a6_k2a_reg_21_ ( clk, n1383_r, a6_k2a[21], a6_v2[21] );
not U_inv2011 ( n1383_r, n1383 );
dff a6_out_1_reg_53_ ( clk, n1383_r, k6[53], k5b[53] );
not U_inv2012 ( n1383_r, n1383 );
dff a6_k2a_reg_22_ ( clk, n1383_r, a6_k2a[22], a6_v2[22] );
not U_inv2013 ( n1383_r, n1383 );
dff a6_out_1_reg_54_ ( clk, n1383_r, k6[54], k5b[54] );
not U_inv2014 ( n1383_r, n1383 );
dff a6_k2a_reg_23_ ( clk, n1383_r, a6_k2a[23], a6_v2[23] );
not U_inv2015 ( n1383_r, n1383 );
dff a6_out_1_reg_55_ ( clk, n1383_r, k6[55], k5b[55] );
not U_inv2016 ( n1383_r, n1383 );
dff a6_k2a_reg_24_ ( clk, n1383_r, a6_k2a[24], a6_v2[24] );
not U_inv2017 ( n1383_r, n1383 );
dff a6_out_1_reg_56_ ( clk, n1383_r, k6[56], k5b[56] );
not U_inv2018 ( n1383_r, n1383 );
dff a6_k2a_reg_25_ ( clk, n1383_r, a6_k2a[25], a6_v2[25] );
not U_inv2019 ( n1383_r, n1383 );
dff a6_out_1_reg_57_ ( clk, n1383_r, k6[57], k5b[57] );
not U_inv2020 ( n1383_r, n1383 );
dff a6_k2a_reg_26_ ( clk, n1383_r, a6_k2a[26], a6_v2[26] );
not U_inv2021 ( n1383_r, n1383 );
dff a6_out_1_reg_58_ ( clk, n1382_r, k6[58], k5b[58] );
not U_inv2022 ( n1382_r, n1382 );
dff a6_k2a_reg_27_ ( clk, n1382_r, a6_k2a[27], a6_v2[27] );
not U_inv2023 ( n1382_r, n1382 );
dff a6_out_1_reg_59_ ( clk, n1382_r, k6[59], k5b[59] );
not U_inv2024 ( n1382_r, n1382 );
dff a6_k2a_reg_28_ ( clk, n1382_r, a6_k2a[28], a6_v2[28] );
not U_inv2025 ( n1382_r, n1382 );
dff a6_out_1_reg_60_ ( clk, n1382_r, k6[60], k5b[60] );
not U_inv2026 ( n1382_r, n1382 );
dff a6_k2a_reg_29_ ( clk, n1382_r, a6_k2a[29], a6_v2[29] );
not U_inv2027 ( n1382_r, n1382 );
dff a6_out_1_reg_61_ ( clk, n1382_r, k6[61], k5b[61] );
not U_inv2028 ( n1382_r, n1382 );
dff a6_k2a_reg_30_ ( clk, n1382_r, a6_k2a[30], a6_v2[30] );
not U_inv2029 ( n1382_r, n1382 );
dff a6_out_1_reg_62_ ( clk, n1382_r, k6[62], k5b[62] );
not U_inv2030 ( n1382_r, n1382 );
dff a6_k2a_reg_31_ ( clk, n1382_r, a6_k2a[31], a6_v2[31] );
not U_inv2031 ( n1382_r, n1382 );
dff a6_out_1_reg_63_ ( clk, n1382_r, k6[63], k5b[63] );
not U_inv2032 ( n1382_r, n1382 );
dff a6_k1a_reg_0_ ( clk, n1382_r, a6_k1a[0], a6_v1[0] );
not U_inv2033 ( n1382_r, n1382 );
dff a6_out_1_reg_64_ ( clk, n1381_r, ex_wire92, k5b[64] );
not U_inv2034 ( n834, ex_wire92 );
not U_inv2035 ( n1381_r, n1381 );
dff a6_k1a_reg_1_ ( clk, n1381_r, a6_k1a[1], a6_v1[1] );
not U_inv2036 ( n1381_r, n1381 );
dff a6_out_1_reg_65_ ( clk, n1381_r, ex_wire93, k5b[65] );
not U_inv2037 ( n845, ex_wire93 );
not U_inv2038 ( n1381_r, n1381 );
dff a6_k1a_reg_2_ ( clk, n1381_r, a6_k1a[2], a6_v1[2] );
not U_inv2039 ( n1381_r, n1381 );
dff a6_out_1_reg_66_ ( clk, n1381_r, ex_wire94, k5b[66] );
not U_inv2040 ( n856, ex_wire94 );
not U_inv2041 ( n1381_r, n1381 );
dff a6_k1a_reg_3_ ( clk, n1381_r, a6_k1a[3], a6_v1[3] );
not U_inv2042 ( n1381_r, n1381 );
dff a6_out_1_reg_67_ ( clk, n1381_r, ex_wire95, k5b[67] );
not U_inv2043 ( n858, ex_wire95 );
not U_inv2044 ( n1381_r, n1381 );
dff a6_k1a_reg_4_ ( clk, n1381_r, a6_k1a[4], a6_v1[4] );
not U_inv2045 ( n1381_r, n1381 );
dff a6_out_1_reg_68_ ( clk, n1381_r, k6[68], k5b[68] );
not U_inv2046 ( n1381_r, n1381 );
dff a6_k1a_reg_5_ ( clk, n1381_r, a6_k1a[5], a6_v1[5] );
not U_inv2047 ( n1381_r, n1381 );
dff a6_out_1_reg_69_ ( clk, n1381_r, k6[69], k5b[69] );
not U_inv2048 ( n1381_r, n1381 );
dff a6_k1a_reg_6_ ( clk, n1381_r, a6_k1a[6], a6_v1[6] );
not U_inv2049 ( n1381_r, n1381 );
dff a6_out_1_reg_70_ ( clk, n1380_r, k6[70], k5b[70] );
not U_inv2050 ( n1380_r, n1380 );
dff a6_k1a_reg_7_ ( clk, n1380_r, a6_k1a[7], a6_v1[7] );
not U_inv2051 ( n1380_r, n1380 );
dff a6_out_1_reg_71_ ( clk, n1380_r, k6[71], k5b[71] );
not U_inv2052 ( n1380_r, n1380 );
dff a6_k1a_reg_8_ ( clk, n1380_r, a6_k1a[8], a6_v1[8] );
not U_inv2053 ( n1380_r, n1380 );
dff a6_out_1_reg_72_ ( clk, n1380_r, k6[72], k5b[72] );
not U_inv2054 ( n1380_r, n1380 );
dff a6_k1a_reg_9_ ( clk, n1380_r, a6_k1a[9], a6_v1[9] );
not U_inv2055 ( n1380_r, n1380 );
dff a6_out_1_reg_73_ ( clk, n1380_r, k6[73], k5b[73] );
not U_inv2056 ( n1380_r, n1380 );
dff a6_k1a_reg_10_ ( clk, n1380_r, a6_k1a[10], a6_v1[10] );
not U_inv2057 ( n1380_r, n1380 );
dff a6_out_1_reg_74_ ( clk, n1380_r, k6[74], k5b[74] );
not U_inv2058 ( n1380_r, n1380 );
dff a6_k1a_reg_11_ ( clk, n1380_r, a6_k1a[11], a6_v1[11] );
not U_inv2059 ( n1380_r, n1380 );
dff a6_out_1_reg_75_ ( clk, n1380_r, k6[75], k5b[75] );
not U_inv2060 ( n1380_r, n1380 );
dff a6_k1a_reg_12_ ( clk, n1380_r, a6_k1a[12], a6_v1[12] );
not U_inv2061 ( n1380_r, n1380 );
dff a6_out_1_reg_76_ ( clk, n1379_r, k6[76], k5b[76] );
not U_inv2062 ( n1379_r, n1379 );
dff a6_k1a_reg_13_ ( clk, n1379_r, a6_k1a[13], a6_v1[13] );
not U_inv2063 ( n1379_r, n1379 );
dff a6_out_1_reg_77_ ( clk, n1379_r, k6[77], k5b[77] );
not U_inv2064 ( n1379_r, n1379 );
dff a6_k1a_reg_14_ ( clk, n1379_r, a6_k1a[14], a6_v1[14] );
not U_inv2065 ( n1379_r, n1379 );
dff a6_out_1_reg_78_ ( clk, n1379_r, k6[78], k5b[78] );
not U_inv2066 ( n1379_r, n1379 );
dff a6_k1a_reg_15_ ( clk, n1379_r, a6_k1a[15], a6_v1[15] );
not U_inv2067 ( n1379_r, n1379 );
dff a6_out_1_reg_79_ ( clk, n1379_r, k6[79], k5b[79] );
not U_inv2068 ( n1379_r, n1379 );
dff a6_k1a_reg_16_ ( clk, n1379_r, a6_k1a[16], a6_v1[16] );
not U_inv2069 ( n1379_r, n1379 );
dff a6_out_1_reg_80_ ( clk, n1379_r, k6[80], k5b[80] );
not U_inv2070 ( n1379_r, n1379 );
dff a6_k1a_reg_17_ ( clk, n1379_r, a6_k1a[17], a6_v1[17] );
not U_inv2071 ( n1379_r, n1379 );
dff a6_out_1_reg_81_ ( clk, n1379_r, k6[81], k5b[81] );
not U_inv2072 ( n1379_r, n1379 );
dff a6_k1a_reg_18_ ( clk, n1379_r, a6_k1a[18], a6_v1[18] );
not U_inv2073 ( n1379_r, n1379 );
dff a6_out_1_reg_82_ ( clk, n1378_r, k6[82], k5b[82] );
not U_inv2074 ( n1378_r, n1378 );
dff a6_k1a_reg_19_ ( clk, n1378_r, a6_k1a[19], a6_v1[19] );
not U_inv2075 ( n1378_r, n1378 );
dff a6_out_1_reg_83_ ( clk, n1378_r, k6[83], k5b[83] );
not U_inv2076 ( n1378_r, n1378 );
dff a6_k1a_reg_20_ ( clk, n1378_r, a6_k1a[20], a6_v1[20] );
not U_inv2077 ( n1378_r, n1378 );
dff a6_out_1_reg_84_ ( clk, n1378_r, k6[84], k5b[84] );
not U_inv2078 ( n1378_r, n1378 );
dff a6_k1a_reg_21_ ( clk, n1378_r, a6_k1a[21], a6_v1[21] );
not U_inv2079 ( n1378_r, n1378 );
dff a6_out_1_reg_85_ ( clk, n1378_r, k6[85], k5b[85] );
not U_inv2080 ( n1378_r, n1378 );
dff a6_k1a_reg_22_ ( clk, n1378_r, a6_k1a[22], a6_v1[22] );
not U_inv2081 ( n1378_r, n1378 );
dff a6_out_1_reg_86_ ( clk, n1378_r, k6[86], k5b[86] );
not U_inv2082 ( n1378_r, n1378 );
dff a6_k1a_reg_23_ ( clk, n1378_r, a6_k1a[23], a6_v1[23] );
not U_inv2083 ( n1378_r, n1378 );
dff a6_out_1_reg_87_ ( clk, n1378_r, k6[87], k5b[87] );
not U_inv2084 ( n1378_r, n1378 );
dff a6_k1a_reg_24_ ( clk, n1378_r, a6_k1a[24], a6_v1[24] );
not U_inv2085 ( n1378_r, n1378 );
dff a6_out_1_reg_88_ ( clk, n1377_r, k6[88], k5b[88] );
not U_inv2086 ( n1377_r, n1377 );
dff a6_k1a_reg_25_ ( clk, n1377_r, a6_k1a[25], a6_v1[25] );
not U_inv2087 ( n1377_r, n1377 );
dff a6_out_1_reg_89_ ( clk, n1377_r, k6[89], k5b[89] );
not U_inv2088 ( n1377_r, n1377 );
dff a6_k1a_reg_26_ ( clk, n1377_r, a6_k1a[26], a6_v1[26] );
not U_inv2089 ( n1377_r, n1377 );
dff a6_out_1_reg_90_ ( clk, n1377_r, k6[90], k5b[90] );
not U_inv2090 ( n1377_r, n1377 );
dff a6_k1a_reg_27_ ( clk, n1377_r, a6_k1a[27], a6_v1[27] );
not U_inv2091 ( n1377_r, n1377 );
dff a6_out_1_reg_91_ ( clk, n1377_r, k6[91], k5b[91] );
not U_inv2092 ( n1377_r, n1377 );
dff a6_k1a_reg_28_ ( clk, n1377_r, a6_k1a[28], a6_v1[28] );
not U_inv2093 ( n1377_r, n1377 );
dff a6_out_1_reg_92_ ( clk, n1377_r, k6[92], k5b[92] );
not U_inv2094 ( n1377_r, n1377 );
dff a6_k1a_reg_29_ ( clk, n1377_r, a6_k1a[29], a6_v1[29] );
not U_inv2095 ( n1377_r, n1377 );
dff a6_out_1_reg_93_ ( clk, n1377_r, k6[93], k5b[93] );
not U_inv2096 ( n1377_r, n1377 );
dff a6_k1a_reg_30_ ( clk, n1377_r, a6_k1a[30], a6_v1[30] );
not U_inv2097 ( n1377_r, n1377 );
dff a6_out_1_reg_94_ ( clk, n1376_r, k6[94], k5b[94] );
not U_inv2098 ( n1376_r, n1376 );
dff a6_out_1_reg_95_ ( clk, n1376_r, k6[95], k5b[95] );
not U_inv2099 ( n1376_r, n1376 );
dff a7_k0a_reg_0_ ( clk, n1376_r, a7_k0a[0], k6[96] );
not U_inv2100 ( n1376_r, n1376 );
dff a7_out_1_reg_96_ ( clk, n1376_r, k7[96], k6b[96] );
not U_inv2101 ( n1376_r, n1376 );
dff a7_k0a_reg_1_ ( clk, n1376_r, a7_k0a[1], k6[97] );
not U_inv2102 ( n1376_r, n1376 );
dff a7_out_1_reg_97_ ( clk, n1376_r, k7[97], k6b[97] );
not U_inv2103 ( n1376_r, n1376 );
dff a7_k0a_reg_2_ ( clk, n1376_r, a7_k0a[2], k6[98] );
not U_inv2104 ( n1376_r, n1376 );
dff a7_out_1_reg_98_ ( clk, n1376_r, k7[98], k6b[98] );
not U_inv2105 ( n1376_r, n1376 );
dff a7_k0a_reg_3_ ( clk, n1376_r, a7_k0a[3], k6[99] );
not U_inv2106 ( n1376_r, n1376 );
dff a7_out_1_reg_99_ ( clk, n1376_r, k7[99], k6b[99] );
not U_inv2107 ( n1376_r, n1376 );
dff a7_k0a_reg_4_ ( clk, n1376_r, a7_k0a[4], k6[100] );
not U_inv2108 ( n1376_r, n1376 );
dff a7_out_1_reg_100_ ( clk, n1376_r, k7[100], k6b[100] );
not U_inv2109 ( n890, k7[100] );
not U_inv2110 ( n1376_r, n1376 );
dff a7_k0a_reg_5_ ( clk, n1375_r, a7_k0a[5], k6[101] );
not U_inv2111 ( n1375_r, n1375 );
dff a7_out_1_reg_101_ ( clk, n1375_r, k7[101], k6b[101] );
not U_inv2112 ( n891, k7[101] );
not U_inv2113 ( n1375_r, n1375 );
dff a7_k0a_reg_6_ ( clk, n1375_r, a7_k0a[6], k6[102] );
not U_inv2114 ( n1375_r, n1375 );
dff a7_out_1_reg_102_ ( clk, n1375_r, k7[102], k6b[102] );
not U_inv2115 ( n892, k7[102] );
not U_inv2116 ( n1375_r, n1375 );
dff a7_k0a_reg_7_ ( clk, n1375_r, a7_k0a[7], k6[103] );
not U_inv2117 ( n1375_r, n1375 );
dff a7_out_1_reg_103_ ( clk, n1375_r, k7[103], k6b[103] );
not U_inv2118 ( n893, k7[103] );
not U_inv2119 ( n1375_r, n1375 );
dff a7_k0a_reg_8_ ( clk, n1375_r, a7_k0a[8], k6[104] );
not U_inv2120 ( n1375_r, n1375 );
dff a7_out_1_reg_104_ ( clk, n1375_r, k7[104], k6b[104] );
not U_inv2121 ( n894, k7[104] );
not U_inv2122 ( n1375_r, n1375 );
dff a7_k0a_reg_9_ ( clk, n1375_r, a7_k0a[9], k6[105] );
not U_inv2123 ( n1375_r, n1375 );
dff a7_out_1_reg_105_ ( clk, n1375_r, k7[105], k6b[105] );
not U_inv2124 ( n895, k7[105] );
not U_inv2125 ( n1375_r, n1375 );
dff a7_k0a_reg_10_ ( clk, n1375_r, a7_k0a[10], k6[106] );
not U_inv2126 ( n1375_r, n1375 );
dff a7_out_1_reg_106_ ( clk, n1375_r, k7[106], k6b[106] );
not U_inv2127 ( n866, k7[106] );
not U_inv2128 ( n1375_r, n1375 );
dff a7_k0a_reg_11_ ( clk, n1374_r, a7_k0a[11], k6[107] );
not U_inv2129 ( n1374_r, n1374 );
dff a7_out_1_reg_107_ ( clk, n1374_r, k7[107], k6b[107] );
not U_inv2130 ( n867, k7[107] );
not U_inv2131 ( n1374_r, n1374 );
dff a7_k0a_reg_12_ ( clk, n1374_r, a7_k0a[12], k6[108] );
not U_inv2132 ( n1374_r, n1374 );
dff a7_out_1_reg_108_ ( clk, n1374_r, k7[108], k6b[108] );
not U_inv2133 ( n868, k7[108] );
not U_inv2134 ( n1374_r, n1374 );
dff a7_k0a_reg_13_ ( clk, n1374_r, a7_k0a[13], k6[109] );
not U_inv2135 ( n1374_r, n1374 );
dff a7_out_1_reg_109_ ( clk, n1374_r, k7[109], k6b[109] );
not U_inv2136 ( n869, k7[109] );
not U_inv2137 ( n1374_r, n1374 );
dff a7_k0a_reg_14_ ( clk, n1374_r, a7_k0a[14], k6[110] );
not U_inv2138 ( n1374_r, n1374 );
dff a7_out_1_reg_110_ ( clk, n1374_r, k7[110], k6b[110] );
not U_inv2139 ( n870, k7[110] );
not U_inv2140 ( n1374_r, n1374 );
dff a7_k0a_reg_15_ ( clk, n1374_r, a7_k0a[15], k6[111] );
not U_inv2141 ( n1374_r, n1374 );
dff a7_out_1_reg_111_ ( clk, n1374_r, k7[111], k6b[111] );
not U_inv2142 ( n871, k7[111] );
not U_inv2143 ( n1374_r, n1374 );
dff a7_k0a_reg_16_ ( clk, n1374_r, a7_k0a[16], k6[112] );
not U_inv2144 ( n1374_r, n1374 );
dff a7_out_1_reg_112_ ( clk, n1374_r, k7[112], k6b[112] );
not U_inv2145 ( n872, k7[112] );
not U_inv2146 ( n1374_r, n1374 );
dff a7_k0a_reg_17_ ( clk, n1373_r, a7_k0a[17], k6[113] );
not U_inv2147 ( n1373_r, n1373 );
dff a7_out_1_reg_113_ ( clk, n1373_r, k7[113], k6b[113] );
not U_inv2148 ( n873, k7[113] );
not U_inv2149 ( n1373_r, n1373 );
dff a7_k0a_reg_18_ ( clk, n1373_r, a7_k0a[18], k6[114] );
not U_inv2150 ( n1373_r, n1373 );
dff a7_out_1_reg_114_ ( clk, n1373_r, k7[114], k6b[114] );
not U_inv2151 ( n874, k7[114] );
not U_inv2152 ( n1373_r, n1373 );
dff a7_k0a_reg_19_ ( clk, n1373_r, a7_k0a[19], k6[115] );
not U_inv2153 ( n1373_r, n1373 );
dff a7_out_1_reg_115_ ( clk, n1373_r, k7[115], k6b[115] );
not U_inv2154 ( n875, k7[115] );
not U_inv2155 ( n1373_r, n1373 );
dff a7_k0a_reg_20_ ( clk, n1373_r, a7_k0a[20], k6[116] );
not U_inv2156 ( n1373_r, n1373 );
dff a7_out_1_reg_116_ ( clk, n1373_r, k7[116], k6b[116] );
not U_inv2157 ( n877, k7[116] );
not U_inv2158 ( n1373_r, n1373 );
dff a7_k0a_reg_21_ ( clk, n1373_r, a7_k0a[21], k6[117] );
not U_inv2159 ( n1373_r, n1373 );
dff a7_out_1_reg_117_ ( clk, n1373_r, k7[117], k6b[117] );
not U_inv2160 ( n878, k7[117] );
not U_inv2161 ( n1373_r, n1373 );
dff a7_k0a_reg_22_ ( clk, n1373_r, a7_k0a[22], k6[118] );
not U_inv2162 ( n1373_r, n1373 );
dff a7_out_1_reg_118_ ( clk, n1373_r, k7[118], k6b[118] );
not U_inv2163 ( n879, k7[118] );
not U_inv2164 ( n1373_r, n1373 );
dff a7_k0a_reg_23_ ( clk, n1372_r, a7_k0a[23], k6[119] );
not U_inv2165 ( n1372_r, n1372 );
dff a7_out_1_reg_119_ ( clk, n1372_r, k7[119], k6b[119] );
not U_inv2166 ( n880, k7[119] );
not U_inv2167 ( n1372_r, n1372 );
dff a7_k0a_reg_24_ ( clk, n1372_r, a7_k0a[24], k6[120] );
not U_inv2168 ( n1372_r, n1372 );
dff a7_out_1_reg_120_ ( clk, n1372_r, k7[120], k6b[120] );
not U_inv2169 ( n881, k7[120] );
not U_inv2170 ( n1372_r, n1372 );
dff a7_k0a_reg_25_ ( clk, n1372_r, a7_k0a[25], k6[121] );
not U_inv2171 ( n1372_r, n1372 );
dff a7_out_1_reg_121_ ( clk, n1372_r, k7[121], k6b[121] );
not U_inv2172 ( n882, k7[121] );
not U_inv2173 ( n1372_r, n1372 );
dff a7_k0a_reg_26_ ( clk, n1372_r, a7_k0a[26], k6[122] );
not U_inv2174 ( n1372_r, n1372 );
dff a7_out_1_reg_122_ ( clk, n1372_r, k7[122], k6b[122] );
not U_inv2175 ( n883, k7[122] );
not U_inv2176 ( n1372_r, n1372 );
dff a7_k0a_reg_27_ ( clk, n1372_r, a7_k0a[27], k6[123] );
not U_inv2177 ( n1372_r, n1372 );
dff a7_out_1_reg_123_ ( clk, n1372_r, k7[123], k6b[123] );
not U_inv2178 ( n884, k7[123] );
not U_inv2179 ( n1372_r, n1372 );
dff a7_k0a_reg_28_ ( clk, n1372_r, a7_k0a[28], k6[124] );
not U_inv2180 ( n1372_r, n1372 );
dff a7_out_1_reg_124_ ( clk, n1372_r, k7[124], k6b[124] );
not U_inv2181 ( n885, k7[124] );
not U_inv2182 ( n1372_r, n1372 );
dff a7_k0a_reg_29_ ( clk, n1371_r, a7_k0a[29], k6[125] );
not U_inv2183 ( n1371_r, n1371 );
dff a7_out_1_reg_125_ ( clk, n1371_r, k7[125], k6b[125] );
not U_inv2184 ( n886, k7[125] );
not U_inv2185 ( n1371_r, n1371 );
dff a7_k0a_reg_30_ ( clk, n1371_r, a7_k0a[30], n1290 );
not U_inv2186 ( n1371_r, n1371 );
dff a7_out_1_reg_126_ ( clk, n1371_r, k7[126], k6b[126] );
not U_inv2187 ( n888, k7[126] );
not U_inv2188 ( n1371_r, n1371 );
dff a7_k0a_reg_31_ ( clk, n1371_r, a7_k0a[31], k6[127] );
not U_inv2189 ( n1371_r, n1371 );
dff a7_out_1_reg_127_ ( clk, n1371_r, ex_wire96, k6b[127] );
not U_inv2190 ( n1291, ex_wire96 );
not U_inv2191 ( n1371_r, n1371 );
dff a7_k3a_reg_0_ ( clk, n1371_r, a7_k3a[0], a7_v3[0] );
not U_inv2192 ( n1371_r, n1371 );
dff a7_out_1_reg_0_ ( clk, n1371_r, k7[0], k6b[0] );
not U_inv2193 ( n1371_r, n1371 );
dff a7_k3a_reg_1_ ( clk, n1371_r, a7_k3a[1], a7_v3[1] );
not U_inv2194 ( n1371_r, n1371 );
dff a7_out_1_reg_1_ ( clk, n1371_r, k7[1], k6b[1] );
not U_inv2195 ( n1371_r, n1371 );
dff a7_k3a_reg_2_ ( clk, n1371_r, a7_k3a[2], a7_v3[2] );
not U_inv2196 ( n1371_r, n1371 );
dff a7_out_1_reg_2_ ( clk, n1371_r, k7[2], k6b[2] );
not U_inv2197 ( n1371_r, n1371 );
dff a7_k3a_reg_3_ ( clk, n1370_r, a7_k3a[3], a7_v3[3] );
not U_inv2198 ( n1370_r, n1370 );
dff a7_out_1_reg_3_ ( clk, n1370_r, k7[3], k6b[3] );
not U_inv2199 ( n1370_r, n1370 );
dff a7_k3a_reg_4_ ( clk, n1370_r, a7_k3a[4], a7_v3[4] );
not U_inv2200 ( n1370_r, n1370 );
dff a7_out_1_reg_4_ ( clk, n1370_r, k7[4], k6b[4] );
not U_inv2201 ( n1370_r, n1370 );
dff a7_k3a_reg_5_ ( clk, n1370_r, a7_k3a[5], a7_v3[5] );
not U_inv2202 ( n1370_r, n1370 );
dff a7_out_1_reg_5_ ( clk, n1370_r, k7[5], k6b[5] );
not U_inv2203 ( n1370_r, n1370 );
dff a7_k3a_reg_6_ ( clk, n1370_r, a7_k3a[6], a7_v3[6] );
not U_inv2204 ( n1370_r, n1370 );
dff a7_out_1_reg_6_ ( clk, n1370_r, k7[6], k6b[6] );
not U_inv2205 ( n1370_r, n1370 );
dff a7_k3a_reg_7_ ( clk, n1370_r, a7_k3a[7], a7_v3[7] );
not U_inv2206 ( n1370_r, n1370 );
dff a7_out_1_reg_7_ ( clk, n1370_r, k7[7], k6b[7] );
not U_inv2207 ( n1370_r, n1370 );
dff a7_k3a_reg_8_ ( clk, n1370_r, a7_k3a[8], a7_v3[8] );
not U_inv2208 ( n1370_r, n1370 );
dff a7_out_1_reg_8_ ( clk, n1370_r, k7[8], k6b[8] );
not U_inv2209 ( n1370_r, n1370 );
dff a7_k3a_reg_9_ ( clk, n1369_r, a7_k3a[9], a7_v3[9] );
not U_inv2210 ( n1369_r, n1369 );
dff a7_out_1_reg_9_ ( clk, n1369_r, k7[9], k6b[9] );
not U_inv2211 ( n1369_r, n1369 );
dff a7_k3a_reg_10_ ( clk, n1369_r, a7_k3a[10], a7_v3[10] );
not U_inv2212 ( n1369_r, n1369 );
dff a7_out_1_reg_10_ ( clk, n1369_r, k7[10], k6b[10] );
not U_inv2213 ( n1369_r, n1369 );
dff a7_k3a_reg_11_ ( clk, n1369_r, a7_k3a[11], a7_v3[11] );
not U_inv2214 ( n1369_r, n1369 );
dff a7_out_1_reg_11_ ( clk, n1369_r, k7[11], k6b[11] );
not U_inv2215 ( n1369_r, n1369 );
dff a7_k3a_reg_12_ ( clk, n1369_r, a7_k3a[12], a7_v3[12] );
not U_inv2216 ( n1369_r, n1369 );
dff a7_out_1_reg_12_ ( clk, n1369_r, k7[12], k6b[12] );
not U_inv2217 ( n1369_r, n1369 );
dff a7_k3a_reg_13_ ( clk, n1369_r, a7_k3a[13], a7_v3[13] );
not U_inv2218 ( n1369_r, n1369 );
dff a7_out_1_reg_13_ ( clk, n1369_r, k7[13], k6b[13] );
not U_inv2219 ( n1369_r, n1369 );
dff a7_k3a_reg_14_ ( clk, n1369_r, a7_k3a[14], a7_v3[14] );
not U_inv2220 ( n1369_r, n1369 );
dff a7_out_1_reg_14_ ( clk, n1369_r, k7[14], k6b[14] );
not U_inv2221 ( n1369_r, n1369 );
dff a7_k3a_reg_15_ ( clk, n1368_r, a7_k3a[15], a7_v3[15] );
not U_inv2222 ( n1368_r, n1368 );
dff a7_out_1_reg_15_ ( clk, n1368_r, k7[15], k6b[15] );
not U_inv2223 ( n1368_r, n1368 );
dff a7_k3a_reg_16_ ( clk, n1368_r, a7_k3a[16], a7_v3[16] );
not U_inv2224 ( n1368_r, n1368 );
dff a7_out_1_reg_16_ ( clk, n1368_r, k7[16], k6b[16] );
not U_inv2225 ( n1368_r, n1368 );
dff a7_k3a_reg_17_ ( clk, n1368_r, a7_k3a[17], a7_v3[17] );
not U_inv2226 ( n1368_r, n1368 );
dff a7_out_1_reg_17_ ( clk, n1368_r, k7[17], k6b[17] );
not U_inv2227 ( n1368_r, n1368 );
dff a7_k3a_reg_18_ ( clk, n1368_r, a7_k3a[18], a7_v3[18] );
not U_inv2228 ( n1368_r, n1368 );
dff a7_out_1_reg_18_ ( clk, n1368_r, k7[18], k6b[18] );
not U_inv2229 ( n1368_r, n1368 );
dff a7_k3a_reg_19_ ( clk, n1368_r, a7_k3a[19], a7_v3[19] );
not U_inv2230 ( n1368_r, n1368 );
dff a7_out_1_reg_19_ ( clk, n1368_r, k7[19], k6b[19] );
not U_inv2231 ( n1368_r, n1368 );
dff a7_k3a_reg_20_ ( clk, n1368_r, a7_k3a[20], a7_v3[20] );
not U_inv2232 ( n1368_r, n1368 );
dff a7_out_1_reg_20_ ( clk, n1368_r, k7[20], k6b[20] );
not U_inv2233 ( n1368_r, n1368 );
dff a7_k3a_reg_21_ ( clk, n1367_r, a7_k3a[21], a7_v3[21] );
not U_inv2234 ( n1367_r, n1367 );
dff a7_out_1_reg_21_ ( clk, n1367_r, k7[21], k6b[21] );
not U_inv2235 ( n1367_r, n1367 );
dff a7_k3a_reg_22_ ( clk, n1367_r, a7_k3a[22], a7_v3[22] );
not U_inv2236 ( n1367_r, n1367 );
dff a7_out_1_reg_22_ ( clk, n1367_r, k7[22], k6b[22] );
not U_inv2237 ( n1367_r, n1367 );
dff a7_k3a_reg_23_ ( clk, n1367_r, a7_k3a[23], a7_v3[23] );
not U_inv2238 ( n1367_r, n1367 );
dff a7_out_1_reg_23_ ( clk, n1367_r, k7[23], k6b[23] );
not U_inv2239 ( n1367_r, n1367 );
dff a7_k3a_reg_24_ ( clk, n1367_r, a7_k3a[24], a7_v3[24] );
not U_inv2240 ( n1367_r, n1367 );
dff a7_out_1_reg_24_ ( clk, n1367_r, k7[24], k6b[24] );
not U_inv2241 ( n1367_r, n1367 );
dff a7_k3a_reg_25_ ( clk, n1367_r, a7_k3a[25], a7_v3[25] );
not U_inv2242 ( n1367_r, n1367 );
dff a7_out_1_reg_25_ ( clk, n1367_r, k7[25], k6b[25] );
not U_inv2243 ( n1367_r, n1367 );
dff a7_k3a_reg_26_ ( clk, n1367_r, a7_k3a[26], a7_v3[26] );
not U_inv2244 ( n1367_r, n1367 );
dff a7_out_1_reg_26_ ( clk, n1367_r, k7[26], k6b[26] );
not U_inv2245 ( n1367_r, n1367 );
dff a7_k3a_reg_27_ ( clk, n1366_r, a7_k3a[27], a7_v3[27] );
not U_inv2246 ( n1366_r, n1366 );
dff a7_out_1_reg_27_ ( clk, n1366_r, k7[27], k6b[27] );
not U_inv2247 ( n1366_r, n1366 );
dff a7_k3a_reg_28_ ( clk, n1366_r, a7_k3a[28], a7_v3[28] );
not U_inv2248 ( n1366_r, n1366 );
dff a7_out_1_reg_28_ ( clk, n1366_r, k7[28], k6b[28] );
not U_inv2249 ( n1366_r, n1366 );
dff a7_k3a_reg_29_ ( clk, n1366_r, a7_k3a[29], a7_v3[29] );
not U_inv2250 ( n1366_r, n1366 );
dff a7_out_1_reg_29_ ( clk, n1366_r, k7[29], k6b[29] );
not U_inv2251 ( n1366_r, n1366 );
dff a7_k3a_reg_30_ ( clk, n1366_r, a7_k3a[30], a7_v3[30] );
not U_inv2252 ( n1366_r, n1366 );
dff a7_out_1_reg_30_ ( clk, n1366_r, k7[30], k6b[30] );
not U_inv2253 ( n1366_r, n1366 );
dff a7_k2a_reg_0_ ( clk, n1366_r, a7_k2a[0], a7_v2[0] );
not U_inv2254 ( n1366_r, n1366 );
dff a7_out_1_reg_32_ ( clk, n1366_r, k7[32], k6b[32] );
not U_inv2255 ( n1366_r, n1366 );
dff a7_k2a_reg_1_ ( clk, n1366_r, a7_k2a[1], a7_v2[1] );
not U_inv2256 ( n1366_r, n1366 );
dff a7_out_1_reg_33_ ( clk, n1366_r, k7[33], k6b[33] );
not U_inv2257 ( n1366_r, n1366 );
dff a7_k2a_reg_2_ ( clk, n1365_r, a7_k2a[2], a7_v2[2] );
not U_inv2258 ( n1365_r, n1365 );
dff a7_out_1_reg_34_ ( clk, n1365_r, k7[34], k6b[34] );
not U_inv2259 ( n1365_r, n1365 );
dff a7_k2a_reg_3_ ( clk, n1365_r, a7_k2a[3], a7_v2[3] );
not U_inv2260 ( n1365_r, n1365 );
dff a7_out_1_reg_35_ ( clk, n1365_r, k7[35], k6b[35] );
not U_inv2261 ( n1365_r, n1365 );
dff a7_k2a_reg_4_ ( clk, n1365_r, a7_k2a[4], a7_v2[4] );
not U_inv2262 ( n1365_r, n1365 );
dff a7_out_1_reg_36_ ( clk, n1365_r, k7[36], k6b[36] );
not U_inv2263 ( n1365_r, n1365 );
dff a7_k2a_reg_5_ ( clk, n1365_r, a7_k2a[5], a7_v2[5] );
not U_inv2264 ( n1365_r, n1365 );
dff a7_out_1_reg_37_ ( clk, n1365_r, k7[37], k6b[37] );
not U_inv2265 ( n1365_r, n1365 );
dff a7_k2a_reg_6_ ( clk, n1365_r, a7_k2a[6], a7_v2[6] );
not U_inv2266 ( n1365_r, n1365 );
dff a7_out_1_reg_38_ ( clk, n1365_r, k7[38], k6b[38] );
not U_inv2267 ( n1365_r, n1365 );
dff a7_k2a_reg_7_ ( clk, n1365_r, a7_k2a[7], a7_v2[7] );
not U_inv2268 ( n1365_r, n1365 );
dff a7_out_1_reg_39_ ( clk, n1365_r, k7[39], k6b[39] );
not U_inv2269 ( n1365_r, n1365 );
dff a7_k2a_reg_8_ ( clk, n1364_r, a7_k2a[8], a7_v2[8] );
not U_inv2270 ( n1364_r, n1364 );
dff a7_out_1_reg_40_ ( clk, n1364_r, k7[40], k6b[40] );
not U_inv2271 ( n1364_r, n1364 );
dff a7_k2a_reg_9_ ( clk, n1364_r, a7_k2a[9], a7_v2[9] );
not U_inv2272 ( n1364_r, n1364 );
dff a7_out_1_reg_41_ ( clk, n1364_r, k7[41], k6b[41] );
not U_inv2273 ( n1364_r, n1364 );
dff a7_k2a_reg_10_ ( clk, n1364_r, a7_k2a[10], a7_v2[10] );
not U_inv2274 ( n1364_r, n1364 );
dff a7_out_1_reg_42_ ( clk, n1364_r, k7[42], k6b[42] );
not U_inv2275 ( n1364_r, n1364 );
dff a7_k2a_reg_11_ ( clk, n1364_r, a7_k2a[11], a7_v2[11] );
not U_inv2276 ( n1364_r, n1364 );
dff a7_out_1_reg_43_ ( clk, n1364_r, k7[43], k6b[43] );
not U_inv2277 ( n1364_r, n1364 );
dff a7_k2a_reg_12_ ( clk, n1364_r, a7_k2a[12], a7_v2[12] );
not U_inv2278 ( n1364_r, n1364 );
dff a7_out_1_reg_44_ ( clk, n1364_r, k7[44], k6b[44] );
not U_inv2279 ( n1364_r, n1364 );
dff a7_k2a_reg_13_ ( clk, n1364_r, a7_k2a[13], a7_v2[13] );
not U_inv2280 ( n1364_r, n1364 );
dff a7_out_1_reg_45_ ( clk, n1364_r, k7[45], k6b[45] );
not U_inv2281 ( n1364_r, n1364 );
dff a7_k2a_reg_14_ ( clk, n1363_r, a7_k2a[14], a7_v2[14] );
not U_inv2282 ( n1363_r, n1363 );
dff a7_out_1_reg_46_ ( clk, n1363_r, k7[46], k6b[46] );
not U_inv2283 ( n1363_r, n1363 );
dff a7_k2a_reg_15_ ( clk, n1363_r, a7_k2a[15], a7_v2[15] );
not U_inv2284 ( n1363_r, n1363 );
dff a7_out_1_reg_47_ ( clk, n1363_r, k7[47], k6b[47] );
not U_inv2285 ( n1363_r, n1363 );
dff a7_k2a_reg_16_ ( clk, n1363_r, a7_k2a[16], a7_v2[16] );
not U_inv2286 ( n1363_r, n1363 );
dff a7_out_1_reg_48_ ( clk, n1363_r, k7[48], k6b[48] );
not U_inv2287 ( n1363_r, n1363 );
dff a7_k2a_reg_17_ ( clk, n1363_r, a7_k2a[17], a7_v2[17] );
not U_inv2288 ( n1363_r, n1363 );
dff a7_out_1_reg_49_ ( clk, n1363_r, k7[49], k6b[49] );
not U_inv2289 ( n1363_r, n1363 );
dff a7_k2a_reg_18_ ( clk, n1363_r, a7_k2a[18], a7_v2[18] );
not U_inv2290 ( n1363_r, n1363 );
dff a7_out_1_reg_50_ ( clk, n1363_r, k7[50], k6b[50] );
not U_inv2291 ( n1363_r, n1363 );
dff a7_k2a_reg_19_ ( clk, n1363_r, a7_k2a[19], a7_v2[19] );
not U_inv2292 ( n1363_r, n1363 );
dff a7_out_1_reg_51_ ( clk, n1363_r, k7[51], k6b[51] );
not U_inv2293 ( n1363_r, n1363 );
dff a7_k2a_reg_20_ ( clk, n1362_r, a7_k2a[20], a7_v2[20] );
not U_inv2294 ( n1362_r, n1362 );
dff a7_out_1_reg_52_ ( clk, n1362_r, k7[52], k6b[52] );
not U_inv2295 ( n1362_r, n1362 );
dff a7_k2a_reg_21_ ( clk, n1362_r, a7_k2a[21], a7_v2[21] );
not U_inv2296 ( n1362_r, n1362 );
dff a7_out_1_reg_53_ ( clk, n1362_r, k7[53], k6b[53] );
not U_inv2297 ( n1362_r, n1362 );
dff a7_k2a_reg_22_ ( clk, n1362_r, a7_k2a[22], a7_v2[22] );
not U_inv2298 ( n1362_r, n1362 );
dff a7_out_1_reg_54_ ( clk, n1362_r, k7[54], k6b[54] );
not U_inv2299 ( n1362_r, n1362 );
dff a7_k2a_reg_23_ ( clk, n1362_r, a7_k2a[23], a7_v2[23] );
not U_inv2300 ( n1362_r, n1362 );
dff a7_out_1_reg_55_ ( clk, n1362_r, k7[55], k6b[55] );
not U_inv2301 ( n1362_r, n1362 );
dff a7_k2a_reg_24_ ( clk, n1362_r, a7_k2a[24], a7_v2[24] );
not U_inv2302 ( n1362_r, n1362 );
dff a7_out_1_reg_56_ ( clk, n1362_r, k7[56], k6b[56] );
not U_inv2303 ( n1362_r, n1362 );
dff a7_k2a_reg_25_ ( clk, n1362_r, a7_k2a[25], a7_v2[25] );
not U_inv2304 ( n1362_r, n1362 );
dff a7_out_1_reg_57_ ( clk, n1362_r, k7[57], k6b[57] );
not U_inv2305 ( n1362_r, n1362 );
dff a7_k2a_reg_26_ ( clk, n1361_r, a7_k2a[26], a7_v2[26] );
not U_inv2306 ( n1361_r, n1361 );
dff a7_out_1_reg_58_ ( clk, n1361_r, k7[58], k6b[58] );
not U_inv2307 ( n1361_r, n1361 );
dff a7_k2a_reg_27_ ( clk, n1361_r, a7_k2a[27], a7_v2[27] );
not U_inv2308 ( n1361_r, n1361 );
dff a7_out_1_reg_59_ ( clk, n1361_r, k7[59], k6b[59] );
not U_inv2309 ( n1361_r, n1361 );
dff a7_k2a_reg_28_ ( clk, n1361_r, a7_k2a[28], a7_v2[28] );
not U_inv2310 ( n1361_r, n1361 );
dff a7_out_1_reg_60_ ( clk, n1361_r, k7[60], k6b[60] );
not U_inv2311 ( n1361_r, n1361 );
dff a7_k2a_reg_29_ ( clk, n1361_r, a7_k2a[29], a7_v2[29] );
not U_inv2312 ( n1361_r, n1361 );
dff a7_out_1_reg_61_ ( clk, n1361_r, k7[61], k6b[61] );
not U_inv2313 ( n1361_r, n1361 );
dff a7_k2a_reg_30_ ( clk, n1361_r, a7_k2a[30], a7_v2[30] );
not U_inv2314 ( n1361_r, n1361 );
dff a7_out_1_reg_62_ ( clk, n1361_r, k7[62], k6b[62] );
not U_inv2315 ( n1361_r, n1361 );
dff a7_k2a_reg_31_ ( clk, n1361_r, a7_k2a[31], a7_v2[31] );
not U_inv2316 ( n1361_r, n1361 );
dff a7_out_1_reg_63_ ( clk, n1361_r, k7[63], k6b[63] );
not U_inv2317 ( n1361_r, n1361 );
dff a7_k1a_reg_0_ ( clk, n1360_r, a7_k1a[0], a7_v1[0] );
not U_inv2318 ( n1360_r, n1360 );
dff a7_out_1_reg_64_ ( clk, n1360_r, ex_wire97, k6b[64] );
not U_inv2319 ( n865, ex_wire97 );
not U_inv2320 ( n1360_r, n1360 );
dff a7_k1a_reg_1_ ( clk, n1360_r, a7_k1a[1], a7_v1[1] );
not U_inv2321 ( n1360_r, n1360 );
dff a7_out_1_reg_65_ ( clk, n1360_r, ex_wire98, k6b[65] );
not U_inv2322 ( n876, ex_wire98 );
not U_inv2323 ( n1360_r, n1360 );
dff a7_k1a_reg_2_ ( clk, n1360_r, a7_k1a[2], a7_v1[2] );
not U_inv2324 ( n1360_r, n1360 );
dff a7_out_1_reg_66_ ( clk, n1360_r, ex_wire99, k6b[66] );
not U_inv2325 ( n887, ex_wire99 );
not U_inv2326 ( n1360_r, n1360 );
dff a7_k1a_reg_3_ ( clk, n1360_r, a7_k1a[3], a7_v1[3] );
not U_inv2327 ( n1360_r, n1360 );
dff a7_out_1_reg_67_ ( clk, n1360_r, ex_wire100, k6b[67] );
not U_inv2328 ( n889, ex_wire100 );
not U_inv2329 ( n1360_r, n1360 );
dff a7_k1a_reg_4_ ( clk, n1360_r, a7_k1a[4], a7_v1[4] );
not U_inv2330 ( n1360_r, n1360 );
dff a7_out_1_reg_68_ ( clk, n1360_r, k7[68], k6b[68] );
not U_inv2331 ( n1360_r, n1360 );
dff a7_k1a_reg_5_ ( clk, n1360_r, a7_k1a[5], a7_v1[5] );
not U_inv2332 ( n1360_r, n1360 );
dff a7_out_1_reg_69_ ( clk, n1360_r, k7[69], k6b[69] );
not U_inv2333 ( n1360_r, n1360 );
dff a7_k1a_reg_6_ ( clk, n1359_r, a7_k1a[6], a7_v1[6] );
not U_inv2334 ( n1359_r, n1359 );
dff a7_out_1_reg_70_ ( clk, n1359_r, k7[70], k6b[70] );
not U_inv2335 ( n1359_r, n1359 );
dff a7_k1a_reg_7_ ( clk, n1359_r, a7_k1a[7], a7_v1[7] );
not U_inv2336 ( n1359_r, n1359 );
dff a7_out_1_reg_71_ ( clk, n1359_r, k7[71], k6b[71] );
not U_inv2337 ( n1359_r, n1359 );
dff a7_k1a_reg_8_ ( clk, n1359_r, a7_k1a[8], a7_v1[8] );
not U_inv2338 ( n1359_r, n1359 );
dff a7_out_1_reg_72_ ( clk, n1359_r, k7[72], k6b[72] );
not U_inv2339 ( n1359_r, n1359 );
dff a7_k1a_reg_9_ ( clk, n1359_r, a7_k1a[9], a7_v1[9] );
not U_inv2340 ( n1359_r, n1359 );
dff a7_out_1_reg_73_ ( clk, n1359_r, k7[73], k6b[73] );
not U_inv2341 ( n1359_r, n1359 );
dff a7_k1a_reg_10_ ( clk, n1359_r, a7_k1a[10], a7_v1[10] );
not U_inv2342 ( n1359_r, n1359 );
dff a7_out_1_reg_74_ ( clk, n1359_r, k7[74], k6b[74] );
not U_inv2343 ( n1359_r, n1359 );
dff a7_k1a_reg_11_ ( clk, n1359_r, a7_k1a[11], a7_v1[11] );
not U_inv2344 ( n1359_r, n1359 );
dff a7_out_1_reg_75_ ( clk, n1359_r, k7[75], k6b[75] );
not U_inv2345 ( n1359_r, n1359 );
dff a7_k1a_reg_12_ ( clk, n1358_r, a7_k1a[12], a7_v1[12] );
not U_inv2346 ( n1358_r, n1358 );
dff a7_out_1_reg_76_ ( clk, n1358_r, k7[76], k6b[76] );
not U_inv2347 ( n1358_r, n1358 );
dff a7_k1a_reg_13_ ( clk, n1358_r, a7_k1a[13], a7_v1[13] );
not U_inv2348 ( n1358_r, n1358 );
dff a7_out_1_reg_77_ ( clk, n1358_r, k7[77], k6b[77] );
not U_inv2349 ( n1358_r, n1358 );
dff a7_k1a_reg_14_ ( clk, n1358_r, a7_k1a[14], a7_v1[14] );
not U_inv2350 ( n1358_r, n1358 );
dff a7_out_1_reg_78_ ( clk, n1358_r, k7[78], k6b[78] );
not U_inv2351 ( n1358_r, n1358 );
dff a7_k1a_reg_15_ ( clk, n1358_r, a7_k1a[15], a7_v1[15] );
not U_inv2352 ( n1358_r, n1358 );
dff a7_out_1_reg_79_ ( clk, n1358_r, k7[79], k6b[79] );
not U_inv2353 ( n1358_r, n1358 );
dff a7_k1a_reg_16_ ( clk, n1358_r, a7_k1a[16], a7_v1[16] );
not U_inv2354 ( n1358_r, n1358 );
dff a7_out_1_reg_80_ ( clk, n1358_r, k7[80], k6b[80] );
not U_inv2355 ( n1358_r, n1358 );
dff a7_k1a_reg_17_ ( clk, n1358_r, a7_k1a[17], a7_v1[17] );
not U_inv2356 ( n1358_r, n1358 );
dff a7_out_1_reg_81_ ( clk, n1358_r, k7[81], k6b[81] );
not U_inv2357 ( n1358_r, n1358 );
dff a7_k1a_reg_18_ ( clk, n1357_r, a7_k1a[18], a7_v1[18] );
not U_inv2358 ( n1357_r, n1357 );
dff a7_out_1_reg_82_ ( clk, n1357_r, k7[82], k6b[82] );
not U_inv2359 ( n1357_r, n1357 );
dff a7_k1a_reg_19_ ( clk, n1357_r, a7_k1a[19], a7_v1[19] );
not U_inv2360 ( n1357_r, n1357 );
dff a7_out_1_reg_83_ ( clk, n1357_r, k7[83], k6b[83] );
not U_inv2361 ( n1357_r, n1357 );
dff a7_k1a_reg_20_ ( clk, n1357_r, a7_k1a[20], a7_v1[20] );
not U_inv2362 ( n1357_r, n1357 );
dff a7_out_1_reg_84_ ( clk, n1357_r, k7[84], k6b[84] );
not U_inv2363 ( n1357_r, n1357 );
dff a7_k1a_reg_21_ ( clk, n1357_r, a7_k1a[21], a7_v1[21] );
not U_inv2364 ( n1357_r, n1357 );
dff a7_out_1_reg_85_ ( clk, n1357_r, k7[85], k6b[85] );
not U_inv2365 ( n1357_r, n1357 );
dff a7_k1a_reg_22_ ( clk, n1357_r, a7_k1a[22], a7_v1[22] );
not U_inv2366 ( n1357_r, n1357 );
dff a7_out_1_reg_86_ ( clk, n1357_r, k7[86], k6b[86] );
not U_inv2367 ( n1357_r, n1357 );
dff a7_k1a_reg_23_ ( clk, n1357_r, a7_k1a[23], a7_v1[23] );
not U_inv2368 ( n1357_r, n1357 );
dff a7_out_1_reg_87_ ( clk, n1357_r, k7[87], k6b[87] );
not U_inv2369 ( n1357_r, n1357 );
dff a7_k1a_reg_24_ ( clk, n1356_r, a7_k1a[24], a7_v1[24] );
not U_inv2370 ( n1356_r, n1356 );
dff a7_out_1_reg_88_ ( clk, n1356_r, k7[88], k6b[88] );
not U_inv2371 ( n1356_r, n1356 );
dff a7_k1a_reg_25_ ( clk, n1356_r, a7_k1a[25], a7_v1[25] );
not U_inv2372 ( n1356_r, n1356 );
dff a7_out_1_reg_89_ ( clk, n1356_r, k7[89], k6b[89] );
not U_inv2373 ( n1356_r, n1356 );
dff a7_k1a_reg_26_ ( clk, n1356_r, a7_k1a[26], a7_v1[26] );
not U_inv2374 ( n1356_r, n1356 );
dff a7_out_1_reg_90_ ( clk, n1356_r, k7[90], k6b[90] );
not U_inv2375 ( n1356_r, n1356 );
dff a7_k1a_reg_27_ ( clk, n1356_r, a7_k1a[27], a7_v1[27] );
not U_inv2376 ( n1356_r, n1356 );
dff a7_out_1_reg_91_ ( clk, n1356_r, k7[91], k6b[91] );
not U_inv2377 ( n1356_r, n1356 );
dff a7_k1a_reg_28_ ( clk, n1356_r, a7_k1a[28], a7_v1[28] );
not U_inv2378 ( n1356_r, n1356 );
dff a7_out_1_reg_92_ ( clk, n1356_r, k7[92], k6b[92] );
not U_inv2379 ( n1356_r, n1356 );
dff a7_k1a_reg_29_ ( clk, n1356_r, a7_k1a[29], a7_v1[29] );
not U_inv2380 ( n1356_r, n1356 );
dff a7_out_1_reg_93_ ( clk, n1356_r, k7[93], k6b[93] );
not U_inv2381 ( n1356_r, n1356 );
dff a7_k1a_reg_30_ ( clk, n1355_r, a7_k1a[30], a7_v1[30] );
not U_inv2382 ( n1355_r, n1355 );
dff a7_out_1_reg_94_ ( clk, n1355_r, k7[94], k6b[94] );
not U_inv2383 ( n1355_r, n1355 );
dff a7_out_1_reg_95_ ( clk, n1355_r, k7[95], k6b[95] );
not U_inv2384 ( n1355_r, n1355 );
dff a8_k0a_reg_0_ ( clk, n1355_r, a8_k0a[0], k7[96] );
not U_inv2385 ( n1355_r, n1355 );
dff a8_out_1_reg_96_ ( clk, n1355_r, k8[96], k7b[96] );
not U_inv2386 ( n1355_r, n1355 );
dff a8_k0a_reg_1_ ( clk, n1355_r, a8_k0a[1], k7[97] );
not U_inv2387 ( n1355_r, n1355 );
dff a8_out_1_reg_97_ ( clk, n1355_r, k8[97], k7b[97] );
not U_inv2388 ( n1355_r, n1355 );
dff a8_k0a_reg_2_ ( clk, n1355_r, a8_k0a[2], k7[98] );
not U_inv2389 ( n1355_r, n1355 );
dff a8_out_1_reg_98_ ( clk, n1355_r, k8[98], k7b[98] );
not U_inv2390 ( n1355_r, n1355 );
dff a8_k0a_reg_3_ ( clk, n1355_r, a8_k0a[3], k7[99] );
not U_inv2391 ( n1355_r, n1355 );
dff a8_out_1_reg_99_ ( clk, n1355_r, k8[99], k7b[99] );
not U_inv2392 ( n1355_r, n1355 );
dff a8_k0a_reg_4_ ( clk, n1355_r, a8_k0a[4], k7[100] );
not U_inv2393 ( n1355_r, n1355 );
dff a8_out_1_reg_100_ ( clk, n1354_r, k8[100], k7b[100] );
not U_inv2394 ( n918, k8[100] );
not U_inv2395 ( n1354_r, n1354 );
dff a8_k0a_reg_5_ ( clk, n1354_r, a8_k0a[5], k7[101] );
not U_inv2396 ( n1354_r, n1354 );
dff a8_out_1_reg_101_ ( clk, n1354_r, k8[101], k7b[101] );
not U_inv2397 ( n919, k8[101] );
not U_inv2398 ( n1354_r, n1354 );
dff a8_k0a_reg_6_ ( clk, n1354_r, a8_k0a[6], k7[102] );
not U_inv2399 ( n1354_r, n1354 );
dff a8_out_1_reg_102_ ( clk, n1354_r, k8[102], k7b[102] );
not U_inv2400 ( n920, k8[102] );
not U_inv2401 ( n1354_r, n1354 );
dff a8_k0a_reg_7_ ( clk, n1354_r, a8_k0a[7], k7[103] );
not U_inv2402 ( n1354_r, n1354 );
dff a8_out_1_reg_103_ ( clk, n1354_r, k8[103], k7b[103] );
not U_inv2403 ( n921, k8[103] );
not U_inv2404 ( n1354_r, n1354 );
dff a8_k0a_reg_8_ ( clk, n1354_r, a8_k0a[8], k7[104] );
not U_inv2405 ( n1354_r, n1354 );
dff a8_out_1_reg_104_ ( clk, n1354_r, k8[104], k7b[104] );
not U_inv2406 ( n922, k8[104] );
not U_inv2407 ( n1354_r, n1354 );
dff a8_k0a_reg_9_ ( clk, n1354_r, a8_k0a[9], k7[105] );
not U_inv2408 ( n1354_r, n1354 );
dff a8_out_1_reg_105_ ( clk, n1354_r, k8[105], k7b[105] );
not U_inv2409 ( n923, k8[105] );
not U_inv2410 ( n1354_r, n1354 );
dff a8_k0a_reg_10_ ( clk, n1354_r, a8_k0a[10], k7[106] );
not U_inv2411 ( n1354_r, n1354 );
dff a8_out_1_reg_106_ ( clk, n1353_r, k8[106], k7b[106] );
not U_inv2412 ( n897, k8[106] );
not U_inv2413 ( n1353_r, n1353 );
dff a8_k0a_reg_11_ ( clk, n1353_r, a8_k0a[11], k7[107] );
not U_inv2414 ( n1353_r, n1353 );
dff a8_out_1_reg_107_ ( clk, n1353_r, k8[107], k7b[107] );
not U_inv2415 ( n898, k8[107] );
not U_inv2416 ( n1353_r, n1353 );
dff a8_k0a_reg_12_ ( clk, n1353_r, a8_k0a[12], k7[108] );
not U_inv2417 ( n1353_r, n1353 );
dff a8_out_1_reg_108_ ( clk, n1353_r, k8[108], k7b[108] );
not U_inv2418 ( n899, k8[108] );
not U_inv2419 ( n1353_r, n1353 );
dff a8_k0a_reg_13_ ( clk, n1353_r, a8_k0a[13], k7[109] );
not U_inv2420 ( n1353_r, n1353 );
dff a8_out_1_reg_109_ ( clk, n1353_r, k8[109], k7b[109] );
not U_inv2421 ( n900, k8[109] );
not U_inv2422 ( n1353_r, n1353 );
dff a8_k0a_reg_14_ ( clk, n1353_r, a8_k0a[14], k7[110] );
not U_inv2423 ( n1353_r, n1353 );
dff a8_out_1_reg_110_ ( clk, n1353_r, k8[110], k7b[110] );
not U_inv2424 ( n901, k8[110] );
not U_inv2425 ( n1353_r, n1353 );
dff a8_k0a_reg_15_ ( clk, n1353_r, a8_k0a[15], k7[111] );
not U_inv2426 ( n1353_r, n1353 );
dff a8_out_1_reg_111_ ( clk, n1353_r, k8[111], k7b[111] );
not U_inv2427 ( n902, k8[111] );
not U_inv2428 ( n1353_r, n1353 );
dff a8_k0a_reg_16_ ( clk, n1353_r, a8_k0a[16], k7[112] );
not U_inv2429 ( n1353_r, n1353 );
dff a8_out_1_reg_112_ ( clk, n1352_r, k8[112], k7b[112] );
not U_inv2430 ( n903, k8[112] );
not U_inv2431 ( n1352_r, n1352 );
dff a8_k0a_reg_17_ ( clk, n1352_r, a8_k0a[17], k7[113] );
not U_inv2432 ( n1352_r, n1352 );
dff a8_out_1_reg_113_ ( clk, n1352_r, k8[113], k7b[113] );
not U_inv2433 ( n904, k8[113] );
not U_inv2434 ( n1352_r, n1352 );
dff a8_k0a_reg_18_ ( clk, n1352_r, a8_k0a[18], k7[114] );
not U_inv2435 ( n1352_r, n1352 );
dff a8_out_1_reg_114_ ( clk, n1352_r, k8[114], k7b[114] );
not U_inv2436 ( n905, k8[114] );
not U_inv2437 ( n1352_r, n1352 );
dff a8_k0a_reg_19_ ( clk, n1352_r, a8_k0a[19], k7[115] );
not U_inv2438 ( n1352_r, n1352 );
dff a8_out_1_reg_115_ ( clk, n1352_r, k8[115], k7b[115] );
not U_inv2439 ( n906, k8[115] );
not U_inv2440 ( n1352_r, n1352 );
dff a8_k0a_reg_20_ ( clk, n1352_r, a8_k0a[20], k7[116] );
not U_inv2441 ( n1352_r, n1352 );
dff a8_out_1_reg_116_ ( clk, n1352_r, k8[116], k7b[116] );
not U_inv2442 ( n908, k8[116] );
not U_inv2443 ( n1352_r, n1352 );
dff a8_k0a_reg_21_ ( clk, n1352_r, a8_k0a[21], k7[117] );
not U_inv2444 ( n1352_r, n1352 );
dff a8_out_1_reg_117_ ( clk, n1352_r, k8[117], k7b[117] );
not U_inv2445 ( n909, k8[117] );
not U_inv2446 ( n1352_r, n1352 );
dff a8_k0a_reg_22_ ( clk, n1352_r, a8_k0a[22], k7[118] );
not U_inv2447 ( n1352_r, n1352 );
dff a8_out_1_reg_118_ ( clk, n1351_r, k8[118], k7b[118] );
not U_inv2448 ( n910, k8[118] );
not U_inv2449 ( n1351_r, n1351 );
dff a8_k0a_reg_23_ ( clk, n1351_r, a8_k0a[23], k7[119] );
not U_inv2450 ( n1351_r, n1351 );
dff a8_out_1_reg_119_ ( clk, n1351_r, k8[119], k7b[119] );
not U_inv2451 ( n911, k8[119] );
not U_inv2452 ( n1351_r, n1351 );
dff a8_k0a_reg_24_ ( clk, n1351_r, a8_k0a[24], k7[120] );
not U_inv2453 ( n1351_r, n1351 );
dff a8_out_1_reg_120_ ( clk, n1351_r, ex_wire101, k7b[120] );
not U_inv2454 ( n1292, ex_wire101 );
not U_inv2455 ( n1351_r, n1351 );
dff a8_k0a_reg_25_ ( clk, n1351_r, a8_k0a[25], k7[121] );
not U_inv2456 ( n1351_r, n1351 );
dff a8_out_1_reg_121_ ( clk, n1351_r, ex_wire102, k7b[121] );
not U_inv2457 ( n1293, ex_wire102 );
not U_inv2458 ( n1351_r, n1351 );
dff a8_k0a_reg_26_ ( clk, n1351_r, a8_k0a[26], k7[122] );
not U_inv2459 ( n1351_r, n1351 );
dff a8_out_1_reg_122_ ( clk, n1351_r, k8[122], k7b[122] );
not U_inv2460 ( n912, k8[122] );
not U_inv2461 ( n1351_r, n1351 );
dff a8_k0a_reg_27_ ( clk, n1351_r, a8_k0a[27], k7[123] );
not U_inv2462 ( n1351_r, n1351 );
dff a8_out_1_reg_123_ ( clk, n1351_r, ex_wire103, k7b[123] );
not U_inv2463 ( n1294, ex_wire103 );
not U_inv2464 ( n1351_r, n1351 );
dff a8_k0a_reg_28_ ( clk, n1351_r, a8_k0a[28], k7[124] );
not U_inv2465 ( n1351_r, n1351 );
dff a8_out_1_reg_124_ ( clk, n1350_r, ex_wire104, k7b[124] );
not U_inv2466 ( n1295, ex_wire104 );
not U_inv2467 ( n1350_r, n1350 );
dff a8_k0a_reg_29_ ( clk, n1350_r, a8_k0a[29], k7[125] );
not U_inv2468 ( n1350_r, n1350 );
dff a8_out_1_reg_125_ ( clk, n1350_r, k8[125], k7b[125] );
not U_inv2469 ( n913, k8[125] );
not U_inv2470 ( n1350_r, n1350 );
dff a8_k0a_reg_30_ ( clk, n1350_r, a8_k0a[30], k7[126] );
not U_inv2471 ( n1350_r, n1350 );
dff a8_out_1_reg_126_ ( clk, n1350_r, k8[126], k7b[126] );
not U_inv2472 ( n915, k8[126] );
not U_inv2473 ( n1350_r, n1350 );
dff a8_k0a_reg_31_ ( clk, n1350_r, a8_k0a[31], n1291 );
not U_inv2474 ( n1350_r, n1350 );
dff a8_out_1_reg_127_ ( clk, n1350_r, k8[127], k7b[127] );
not U_inv2475 ( n916, k8[127] );
not U_inv2476 ( n1350_r, n1350 );
dff a8_k3a_reg_0_ ( clk, n1350_r, a8_k3a[0], a8_v3[0] );
not U_inv2477 ( n1350_r, n1350 );
dff a8_out_1_reg_0_ ( clk, n1350_r, k8[0], k7b[0] );
not U_inv2478 ( n1350_r, n1350 );
dff a8_k3a_reg_1_ ( clk, n1350_r, a8_k3a[1], a8_v3[1] );
not U_inv2479 ( n1350_r, n1350 );
dff a8_out_1_reg_1_ ( clk, n1350_r, k8[1], k7b[1] );
not U_inv2480 ( n1350_r, n1350 );
dff a8_k3a_reg_2_ ( clk, n1350_r, a8_k3a[2], a8_v3[2] );
not U_inv2481 ( n1350_r, n1350 );
dff a8_out_1_reg_2_ ( clk, n1349_r, k8[2], k7b[2] );
not U_inv2482 ( n1349_r, n1349 );
dff a8_k3a_reg_3_ ( clk, n1349_r, a8_k3a[3], a8_v3[3] );
not U_inv2483 ( n1349_r, n1349 );
dff a8_out_1_reg_3_ ( clk, n1349_r, k8[3], k7b[3] );
not U_inv2484 ( n1349_r, n1349 );
dff a8_k3a_reg_4_ ( clk, n1349_r, a8_k3a[4], a8_v3[4] );
not U_inv2485 ( n1349_r, n1349 );
dff a8_out_1_reg_4_ ( clk, n1349_r, k8[4], k7b[4] );
not U_inv2486 ( n1349_r, n1349 );
dff a8_k3a_reg_5_ ( clk, n1349_r, a8_k3a[5], a8_v3[5] );
not U_inv2487 ( n1349_r, n1349 );
dff a8_out_1_reg_5_ ( clk, n1349_r, k8[5], k7b[5] );
not U_inv2488 ( n1349_r, n1349 );
dff a8_k3a_reg_6_ ( clk, n1349_r, a8_k3a[6], a8_v3[6] );
not U_inv2489 ( n1349_r, n1349 );
dff a8_out_1_reg_6_ ( clk, n1349_r, k8[6], k7b[6] );
not U_inv2490 ( n1349_r, n1349 );
dff a8_k3a_reg_7_ ( clk, n1349_r, a8_k3a[7], a8_v3[7] );
not U_inv2491 ( n1349_r, n1349 );
dff a8_out_1_reg_7_ ( clk, n1349_r, k8[7], k7b[7] );
not U_inv2492 ( n1349_r, n1349 );
dff a8_k3a_reg_8_ ( clk, n1349_r, a8_k3a[8], a8_v3[8] );
not U_inv2493 ( n1349_r, n1349 );
dff a8_out_1_reg_8_ ( clk, n1348_r, k8[8], k7b[8] );
not U_inv2494 ( n1348_r, n1348 );
dff a8_k3a_reg_9_ ( clk, n1348_r, a8_k3a[9], a8_v3[9] );
not U_inv2495 ( n1348_r, n1348 );
dff a8_out_1_reg_9_ ( clk, n1348_r, k8[9], k7b[9] );
not U_inv2496 ( n1348_r, n1348 );
dff a8_k3a_reg_10_ ( clk, n1348_r, a8_k3a[10], a8_v3[10] );
not U_inv2497 ( n1348_r, n1348 );
dff a8_out_1_reg_10_ ( clk, n1348_r, k8[10], k7b[10] );
not U_inv2498 ( n1348_r, n1348 );
dff a8_k3a_reg_11_ ( clk, n1348_r, a8_k3a[11], a8_v3[11] );
not U_inv2499 ( n1348_r, n1348 );
dff a8_out_1_reg_11_ ( clk, n1348_r, k8[11], k7b[11] );
not U_inv2500 ( n1348_r, n1348 );
dff a8_k3a_reg_12_ ( clk, n1348_r, a8_k3a[12], a8_v3[12] );
not U_inv2501 ( n1348_r, n1348 );
dff a8_out_1_reg_12_ ( clk, n1348_r, k8[12], k7b[12] );
not U_inv2502 ( n1348_r, n1348 );
dff a8_k3a_reg_13_ ( clk, n1348_r, a8_k3a[13], a8_v3[13] );
not U_inv2503 ( n1348_r, n1348 );
dff a8_out_1_reg_13_ ( clk, n1348_r, k8[13], k7b[13] );
not U_inv2504 ( n1348_r, n1348 );
dff a8_k3a_reg_14_ ( clk, n1348_r, a8_k3a[14], a8_v3[14] );
not U_inv2505 ( n1348_r, n1348 );
dff a8_out_1_reg_14_ ( clk, n1347_r, k8[14], k7b[14] );
not U_inv2506 ( n1347_r, n1347 );
dff a8_k3a_reg_15_ ( clk, n1347_r, a8_k3a[15], a8_v3[15] );
not U_inv2507 ( n1347_r, n1347 );
dff a8_out_1_reg_15_ ( clk, n1347_r, k8[15], k7b[15] );
not U_inv2508 ( n1347_r, n1347 );
dff a8_k3a_reg_16_ ( clk, n1347_r, a8_k3a[16], a8_v3[16] );
not U_inv2509 ( n1347_r, n1347 );
dff a8_out_1_reg_16_ ( clk, n1347_r, k8[16], k7b[16] );
not U_inv2510 ( n1347_r, n1347 );
dff a8_k3a_reg_17_ ( clk, n1347_r, a8_k3a[17], a8_v3[17] );
not U_inv2511 ( n1347_r, n1347 );
dff a8_out_1_reg_17_ ( clk, n1347_r, k8[17], k7b[17] );
not U_inv2512 ( n1347_r, n1347 );
dff a8_k3a_reg_18_ ( clk, n1347_r, a8_k3a[18], a8_v3[18] );
not U_inv2513 ( n1347_r, n1347 );
dff a8_out_1_reg_18_ ( clk, n1347_r, k8[18], k7b[18] );
not U_inv2514 ( n1347_r, n1347 );
dff a8_k3a_reg_19_ ( clk, n1347_r, a8_k3a[19], a8_v3[19] );
not U_inv2515 ( n1347_r, n1347 );
dff a8_out_1_reg_19_ ( clk, n1347_r, k8[19], k7b[19] );
not U_inv2516 ( n1347_r, n1347 );
dff a8_k3a_reg_20_ ( clk, n1347_r, a8_k3a[20], a8_v3[20] );
not U_inv2517 ( n1347_r, n1347 );
dff a8_out_1_reg_20_ ( clk, n1346_r, k8[20], k7b[20] );
not U_inv2518 ( n1346_r, n1346 );
dff a8_k3a_reg_21_ ( clk, n1346_r, a8_k3a[21], a8_v3[21] );
not U_inv2519 ( n1346_r, n1346 );
dff a8_out_1_reg_21_ ( clk, n1346_r, k8[21], k7b[21] );
not U_inv2520 ( n1346_r, n1346 );
dff a8_k3a_reg_22_ ( clk, n1346_r, a8_k3a[22], a8_v3[22] );
not U_inv2521 ( n1346_r, n1346 );
dff a8_out_1_reg_22_ ( clk, n1346_r, k8[22], k7b[22] );
not U_inv2522 ( n1346_r, n1346 );
dff a8_k3a_reg_23_ ( clk, n1346_r, a8_k3a[23], a8_v3[23] );
not U_inv2523 ( n1346_r, n1346 );
dff a8_out_1_reg_23_ ( clk, n1346_r, k8[23], k7b[23] );
not U_inv2524 ( n1346_r, n1346 );
dff a8_k3a_reg_24_ ( clk, n1346_r, a8_k3a[24], a8_v3[24] );
not U_inv2525 ( n1346_r, n1346 );
dff a8_out_1_reg_24_ ( clk, n1346_r, k8[24], k7b[24] );
not U_inv2526 ( n1346_r, n1346 );
dff a8_k3a_reg_25_ ( clk, n1346_r, a8_k3a[25], a8_v3[25] );
not U_inv2527 ( n1346_r, n1346 );
dff a8_out_1_reg_25_ ( clk, n1346_r, k8[25], k7b[25] );
not U_inv2528 ( n1346_r, n1346 );
dff a8_k3a_reg_26_ ( clk, n1346_r, a8_k3a[26], a8_v3[26] );
not U_inv2529 ( n1346_r, n1346 );
dff a8_out_1_reg_26_ ( clk, n1345_r, k8[26], k7b[26] );
not U_inv2530 ( n1345_r, n1345 );
dff a8_k3a_reg_27_ ( clk, n1345_r, a8_k3a[27], a8_v3[27] );
not U_inv2531 ( n1345_r, n1345 );
dff a8_out_1_reg_27_ ( clk, n1345_r, k8[27], k7b[27] );
not U_inv2532 ( n1345_r, n1345 );
dff a8_k3a_reg_28_ ( clk, n1345_r, a8_k3a[28], a8_v3[28] );
not U_inv2533 ( n1345_r, n1345 );
dff a8_out_1_reg_28_ ( clk, n1345_r, k8[28], k7b[28] );
not U_inv2534 ( n1345_r, n1345 );
dff a8_k3a_reg_29_ ( clk, n1345_r, a8_k3a[29], a8_v3[29] );
not U_inv2535 ( n1345_r, n1345 );
dff a8_out_1_reg_29_ ( clk, n1345_r, k8[29], k7b[29] );
not U_inv2536 ( n1345_r, n1345 );
dff a8_k3a_reg_30_ ( clk, n1345_r, a8_k3a[30], a8_v3[30] );
not U_inv2537 ( n1345_r, n1345 );
dff a8_out_1_reg_30_ ( clk, n1345_r, k8[30], k7b[30] );
not U_inv2538 ( n1345_r, n1345 );
dff a8_k2a_reg_0_ ( clk, n1345_r, a8_k2a[0], a8_v2[0] );
not U_inv2539 ( n1345_r, n1345 );
dff a8_out_1_reg_32_ ( clk, n1345_r, k8[32], k7b[32] );
not U_inv2540 ( n1345_r, n1345 );
dff a8_k2a_reg_1_ ( clk, n1345_r, a8_k2a[1], a8_v2[1] );
not U_inv2541 ( n1345_r, n1345 );
dff a8_out_1_reg_33_ ( clk, n1344_r, k8[33], k7b[33] );
not U_inv2542 ( n1344_r, n1344 );
dff a8_k2a_reg_2_ ( clk, n1344_r, a8_k2a[2], a8_v2[2] );
not U_inv2543 ( n1344_r, n1344 );
dff a8_out_1_reg_34_ ( clk, n1344_r, k8[34], k7b[34] );
not U_inv2544 ( n1344_r, n1344 );
dff a8_k2a_reg_3_ ( clk, n1344_r, a8_k2a[3], a8_v2[3] );
not U_inv2545 ( n1344_r, n1344 );
dff a8_out_1_reg_35_ ( clk, n1344_r, k8[35], k7b[35] );
not U_inv2546 ( n1344_r, n1344 );
dff a8_k2a_reg_4_ ( clk, n1344_r, a8_k2a[4], a8_v2[4] );
not U_inv2547 ( n1344_r, n1344 );
dff a8_out_1_reg_36_ ( clk, n1344_r, k8[36], k7b[36] );
not U_inv2548 ( n1344_r, n1344 );
dff a8_k2a_reg_5_ ( clk, n1344_r, a8_k2a[5], a8_v2[5] );
not U_inv2549 ( n1344_r, n1344 );
dff a8_out_1_reg_37_ ( clk, n1344_r, k8[37], k7b[37] );
not U_inv2550 ( n1344_r, n1344 );
dff a8_k2a_reg_6_ ( clk, n1344_r, a8_k2a[6], a8_v2[6] );
not U_inv2551 ( n1344_r, n1344 );
dff a8_out_1_reg_38_ ( clk, n1344_r, k8[38], k7b[38] );
not U_inv2552 ( n1344_r, n1344 );
dff a8_k2a_reg_7_ ( clk, n1344_r, a8_k2a[7], a8_v2[7] );
not U_inv2553 ( n1344_r, n1344 );
dff a8_out_1_reg_39_ ( clk, n1343_r, k8[39], k7b[39] );
not U_inv2554 ( n1343_r, n1343 );
dff a8_k2a_reg_8_ ( clk, n1343_r, a8_k2a[8], a8_v2[8] );
not U_inv2555 ( n1343_r, n1343 );
dff a8_out_1_reg_40_ ( clk, n1343_r, k8[40], k7b[40] );
not U_inv2556 ( n1343_r, n1343 );
dff a8_k2a_reg_9_ ( clk, n1343_r, a8_k2a[9], a8_v2[9] );
not U_inv2557 ( n1343_r, n1343 );
dff a8_out_1_reg_41_ ( clk, n1343_r, k8[41], k7b[41] );
not U_inv2558 ( n1343_r, n1343 );
dff a8_k2a_reg_10_ ( clk, n1343_r, a8_k2a[10], a8_v2[10] );
not U_inv2559 ( n1343_r, n1343 );
dff a8_out_1_reg_42_ ( clk, n1343_r, k8[42], k7b[42] );
not U_inv2560 ( n1343_r, n1343 );
dff a8_k2a_reg_11_ ( clk, n1343_r, a8_k2a[11], a8_v2[11] );
not U_inv2561 ( n1343_r, n1343 );
dff a8_out_1_reg_43_ ( clk, n1343_r, k8[43], k7b[43] );
not U_inv2562 ( n1343_r, n1343 );
dff a8_k2a_reg_12_ ( clk, n1343_r, a8_k2a[12], a8_v2[12] );
not U_inv2563 ( n1343_r, n1343 );
dff a8_out_1_reg_44_ ( clk, n1343_r, k8[44], k7b[44] );
not U_inv2564 ( n1343_r, n1343 );
dff a8_k2a_reg_13_ ( clk, n1343_r, a8_k2a[13], a8_v2[13] );
not U_inv2565 ( n1343_r, n1343 );
dff a8_out_1_reg_45_ ( clk, n1342_r, k8[45], k7b[45] );
not U_inv2566 ( n1342_r, n1342 );
dff a8_k2a_reg_14_ ( clk, n1342_r, a8_k2a[14], a8_v2[14] );
not U_inv2567 ( n1342_r, n1342 );
dff a8_out_1_reg_46_ ( clk, n1342_r, k8[46], k7b[46] );
not U_inv2568 ( n1342_r, n1342 );
dff a8_k2a_reg_15_ ( clk, n1342_r, a8_k2a[15], a8_v2[15] );
not U_inv2569 ( n1342_r, n1342 );
dff a8_out_1_reg_47_ ( clk, n1342_r, k8[47], k7b[47] );
not U_inv2570 ( n1342_r, n1342 );
dff a8_k2a_reg_16_ ( clk, n1342_r, a8_k2a[16], a8_v2[16] );
not U_inv2571 ( n1342_r, n1342 );
dff a8_out_1_reg_48_ ( clk, n1342_r, k8[48], k7b[48] );
not U_inv2572 ( n1342_r, n1342 );
dff a8_k2a_reg_17_ ( clk, n1342_r, a8_k2a[17], a8_v2[17] );
not U_inv2573 ( n1342_r, n1342 );
dff a8_out_1_reg_49_ ( clk, n1342_r, k8[49], k7b[49] );
not U_inv2574 ( n1342_r, n1342 );
dff a8_k2a_reg_18_ ( clk, n1342_r, a8_k2a[18], a8_v2[18] );
not U_inv2575 ( n1342_r, n1342 );
dff a8_out_1_reg_50_ ( clk, n1342_r, k8[50], k7b[50] );
not U_inv2576 ( n1342_r, n1342 );
dff a8_k2a_reg_19_ ( clk, n1342_r, a8_k2a[19], a8_v2[19] );
not U_inv2577 ( n1342_r, n1342 );
dff a8_out_1_reg_51_ ( clk, n1341_r, k8[51], k7b[51] );
not U_inv2578 ( n1341_r, n1341 );
dff a8_k2a_reg_20_ ( clk, n1341_r, a8_k2a[20], a8_v2[20] );
not U_inv2579 ( n1341_r, n1341 );
dff a8_out_1_reg_52_ ( clk, n1341_r, k8[52], k7b[52] );
not U_inv2580 ( n1341_r, n1341 );
dff a8_k2a_reg_21_ ( clk, n1341_r, a8_k2a[21], a8_v2[21] );
not U_inv2581 ( n1341_r, n1341 );
dff a8_out_1_reg_53_ ( clk, n1341_r, k8[53], k7b[53] );
not U_inv2582 ( n1341_r, n1341 );
dff a8_k2a_reg_22_ ( clk, n1341_r, a8_k2a[22], a8_v2[22] );
not U_inv2583 ( n1341_r, n1341 );
dff a8_out_1_reg_54_ ( clk, n1341_r, k8[54], k7b[54] );
not U_inv2584 ( n1341_r, n1341 );
dff a8_k2a_reg_23_ ( clk, n1341_r, a8_k2a[23], a8_v2[23] );
not U_inv2585 ( n1341_r, n1341 );
dff a8_out_1_reg_55_ ( clk, n1341_r, k8[55], k7b[55] );
not U_inv2586 ( n1341_r, n1341 );
dff a8_k2a_reg_24_ ( clk, n1341_r, a8_k2a[24], a8_v2[24] );
not U_inv2587 ( n1341_r, n1341 );
dff a8_out_1_reg_56_ ( clk, n1341_r, k8[56], k7b[56] );
not U_inv2588 ( n1341_r, n1341 );
dff a8_k2a_reg_25_ ( clk, n1341_r, a8_k2a[25], a8_v2[25] );
not U_inv2589 ( n1341_r, n1341 );
dff a8_out_1_reg_57_ ( clk, n1340_r, k8[57], k7b[57] );
not U_inv2590 ( n1340_r, n1340 );
dff a8_k2a_reg_26_ ( clk, n1340_r, a8_k2a[26], a8_v2[26] );
not U_inv2591 ( n1340_r, n1340 );
dff a8_out_1_reg_58_ ( clk, n1340_r, k8[58], k7b[58] );
not U_inv2592 ( n1340_r, n1340 );
dff a8_k2a_reg_27_ ( clk, n1340_r, a8_k2a[27], a8_v2[27] );
not U_inv2593 ( n1340_r, n1340 );
dff a8_out_1_reg_59_ ( clk, n1340_r, k8[59], k7b[59] );
not U_inv2594 ( n1340_r, n1340 );
dff a8_k2a_reg_28_ ( clk, n1340_r, a8_k2a[28], a8_v2[28] );
not U_inv2595 ( n1340_r, n1340 );
dff a8_out_1_reg_60_ ( clk, n1340_r, k8[60], k7b[60] );
not U_inv2596 ( n1340_r, n1340 );
dff a8_k2a_reg_29_ ( clk, n1340_r, a8_k2a[29], a8_v2[29] );
not U_inv2597 ( n1340_r, n1340 );
dff a8_out_1_reg_61_ ( clk, n1340_r, k8[61], k7b[61] );
not U_inv2598 ( n1340_r, n1340 );
dff a8_k2a_reg_30_ ( clk, n1340_r, a8_k2a[30], a8_v2[30] );
not U_inv2599 ( n1340_r, n1340 );
dff a8_out_1_reg_62_ ( clk, n1340_r, k8[62], k7b[62] );
not U_inv2600 ( n1340_r, n1340 );
dff a8_k2a_reg_31_ ( clk, n1340_r, a8_k2a[31], a8_v2[31] );
not U_inv2601 ( n1340_r, n1340 );
dff a8_out_1_reg_63_ ( clk, n1339_r, k8[63], k7b[63] );
not U_inv2602 ( n1339_r, n1339 );
dff a8_k1a_reg_0_ ( clk, n1339_r, a8_k1a[0], a8_v1[0] );
not U_inv2603 ( n1339_r, n1339 );
dff a8_out_1_reg_64_ ( clk, n1339_r, ex_wire105, k7b[64] );
not U_inv2604 ( n896, ex_wire105 );
not U_inv2605 ( n1339_r, n1339 );
dff a8_k1a_reg_1_ ( clk, n1339_r, a8_k1a[1], a8_v1[1] );
not U_inv2606 ( n1339_r, n1339 );
dff a8_out_1_reg_65_ ( clk, n1339_r, ex_wire106, k7b[65] );
not U_inv2607 ( n907, ex_wire106 );
not U_inv2608 ( n1339_r, n1339 );
dff a8_k1a_reg_2_ ( clk, n1339_r, a8_k1a[2], a8_v1[2] );
not U_inv2609 ( n1339_r, n1339 );
dff a8_out_1_reg_66_ ( clk, n1339_r, ex_wire107, k7b[66] );
not U_inv2610 ( n914, ex_wire107 );
not U_inv2611 ( n1339_r, n1339 );
dff a8_k1a_reg_3_ ( clk, n1339_r, a8_k1a[3], a8_v1[3] );
not U_inv2612 ( n1339_r, n1339 );
dff a8_out_1_reg_67_ ( clk, n1339_r, ex_wire108, k7b[67] );
not U_inv2613 ( n917, ex_wire108 );
not U_inv2614 ( n1339_r, n1339 );
dff a8_k1a_reg_4_ ( clk, n1339_r, a8_k1a[4], a8_v1[4] );
not U_inv2615 ( n1339_r, n1339 );
dff a8_out_1_reg_68_ ( clk, n1339_r, k8[68], k7b[68] );
not U_inv2616 ( n1339_r, n1339 );
dff a8_k1a_reg_5_ ( clk, n1339_r, a8_k1a[5], a8_v1[5] );
not U_inv2617 ( n1339_r, n1339 );
dff a8_out_1_reg_69_ ( clk, n1338_r, k8[69], k7b[69] );
not U_inv2618 ( n1338_r, n1338 );
dff a8_k1a_reg_6_ ( clk, n1338_r, a8_k1a[6], a8_v1[6] );
not U_inv2619 ( n1338_r, n1338 );
dff a8_out_1_reg_70_ ( clk, n1338_r, k8[70], k7b[70] );
not U_inv2620 ( n1338_r, n1338 );
dff a8_k1a_reg_7_ ( clk, n1338_r, a8_k1a[7], a8_v1[7] );
not U_inv2621 ( n1338_r, n1338 );
dff a8_out_1_reg_71_ ( clk, n1338_r, k8[71], k7b[71] );
not U_inv2622 ( n1338_r, n1338 );
dff a8_k1a_reg_8_ ( clk, n1338_r, a8_k1a[8], a8_v1[8] );
not U_inv2623 ( n1338_r, n1338 );
dff a8_out_1_reg_72_ ( clk, n1338_r, k8[72], k7b[72] );
not U_inv2624 ( n1338_r, n1338 );
dff a8_k1a_reg_9_ ( clk, n1338_r, a8_k1a[9], a8_v1[9] );
not U_inv2625 ( n1338_r, n1338 );
dff a8_out_1_reg_73_ ( clk, n1338_r, k8[73], k7b[73] );
not U_inv2626 ( n1338_r, n1338 );
dff a8_k1a_reg_10_ ( clk, n1338_r, a8_k1a[10], a8_v1[10] );
not U_inv2627 ( n1338_r, n1338 );
dff a8_out_1_reg_74_ ( clk, n1338_r, k8[74], k7b[74] );
not U_inv2628 ( n1338_r, n1338 );
dff a8_k1a_reg_11_ ( clk, n1338_r, a8_k1a[11], a8_v1[11] );
not U_inv2629 ( n1338_r, n1338 );
dff a8_out_1_reg_75_ ( clk, n1337_r, k8[75], k7b[75] );
not U_inv2630 ( n1337_r, n1337 );
dff a8_k1a_reg_12_ ( clk, n1337_r, a8_k1a[12], a8_v1[12] );
not U_inv2631 ( n1337_r, n1337 );
dff a8_out_1_reg_76_ ( clk, n1337_r, k8[76], k7b[76] );
not U_inv2632 ( n1337_r, n1337 );
dff a8_k1a_reg_13_ ( clk, n1337_r, a8_k1a[13], a8_v1[13] );
not U_inv2633 ( n1337_r, n1337 );
dff a8_out_1_reg_77_ ( clk, n1337_r, k8[77], k7b[77] );
not U_inv2634 ( n1337_r, n1337 );
dff a8_k1a_reg_14_ ( clk, n1337_r, a8_k1a[14], a8_v1[14] );
not U_inv2635 ( n1337_r, n1337 );
dff a8_out_1_reg_78_ ( clk, n1337_r, k8[78], k7b[78] );
not U_inv2636 ( n1337_r, n1337 );
dff a8_k1a_reg_15_ ( clk, n1337_r, a8_k1a[15], a8_v1[15] );
not U_inv2637 ( n1337_r, n1337 );
dff a8_out_1_reg_79_ ( clk, n1337_r, k8[79], k7b[79] );
not U_inv2638 ( n1337_r, n1337 );
dff a8_k1a_reg_16_ ( clk, n1337_r, a8_k1a[16], a8_v1[16] );
not U_inv2639 ( n1337_r, n1337 );
dff a8_out_1_reg_80_ ( clk, n1337_r, k8[80], k7b[80] );
not U_inv2640 ( n1337_r, n1337 );
dff a8_k1a_reg_17_ ( clk, n1337_r, a8_k1a[17], a8_v1[17] );
not U_inv2641 ( n1337_r, n1337 );
dff a8_out_1_reg_81_ ( clk, n1336_r, k8[81], k7b[81] );
not U_inv2642 ( n1336_r, n1336 );
dff a8_k1a_reg_18_ ( clk, n1336_r, a8_k1a[18], a8_v1[18] );
not U_inv2643 ( n1336_r, n1336 );
dff a8_out_1_reg_82_ ( clk, n1336_r, k8[82], k7b[82] );
not U_inv2644 ( n1336_r, n1336 );
dff a8_k1a_reg_19_ ( clk, n1336_r, a8_k1a[19], a8_v1[19] );
not U_inv2645 ( n1336_r, n1336 );
dff a8_out_1_reg_83_ ( clk, n1336_r, k8[83], k7b[83] );
not U_inv2646 ( n1336_r, n1336 );
dff a8_k1a_reg_20_ ( clk, n1336_r, a8_k1a[20], a8_v1[20] );
not U_inv2647 ( n1336_r, n1336 );
dff a8_out_1_reg_84_ ( clk, n1336_r, k8[84], k7b[84] );
not U_inv2648 ( n1336_r, n1336 );
dff a8_k1a_reg_21_ ( clk, n1336_r, a8_k1a[21], a8_v1[21] );
not U_inv2649 ( n1336_r, n1336 );
dff a8_out_1_reg_85_ ( clk, n1336_r, k8[85], k7b[85] );
not U_inv2650 ( n1336_r, n1336 );
dff a8_k1a_reg_22_ ( clk, n1336_r, a8_k1a[22], a8_v1[22] );
not U_inv2651 ( n1336_r, n1336 );
dff a8_out_1_reg_86_ ( clk, n1336_r, k8[86], k7b[86] );
not U_inv2652 ( n1336_r, n1336 );
dff a8_k1a_reg_23_ ( clk, n1336_r, a8_k1a[23], a8_v1[23] );
not U_inv2653 ( n1336_r, n1336 );
dff a8_out_1_reg_87_ ( clk, n1335_r, k8[87], k7b[87] );
not U_inv2654 ( n1335_r, n1335 );
dff a8_k1a_reg_24_ ( clk, n1335_r, a8_k1a[24], a8_v1[24] );
not U_inv2655 ( n1335_r, n1335 );
dff a8_out_1_reg_88_ ( clk, n1335_r, k8[88], k7b[88] );
not U_inv2656 ( n1335_r, n1335 );
dff a8_k1a_reg_25_ ( clk, n1335_r, a8_k1a[25], a8_v1[25] );
not U_inv2657 ( n1335_r, n1335 );
dff a8_out_1_reg_89_ ( clk, n1335_r, k8[89], k7b[89] );
not U_inv2658 ( n1335_r, n1335 );
dff a8_k1a_reg_26_ ( clk, n1335_r, a8_k1a[26], a8_v1[26] );
not U_inv2659 ( n1335_r, n1335 );
dff a8_out_1_reg_90_ ( clk, n1335_r, k8[90], k7b[90] );
not U_inv2660 ( n1335_r, n1335 );
dff a8_k1a_reg_27_ ( clk, n1335_r, a8_k1a[27], a8_v1[27] );
not U_inv2661 ( n1335_r, n1335 );
dff a8_out_1_reg_91_ ( clk, n1335_r, k8[91], k7b[91] );
not U_inv2662 ( n1335_r, n1335 );
dff a8_k1a_reg_28_ ( clk, n1335_r, a8_k1a[28], a8_v1[28] );
not U_inv2663 ( n1335_r, n1335 );
dff a8_out_1_reg_92_ ( clk, n1335_r, k8[92], k7b[92] );
not U_inv2664 ( n1335_r, n1335 );
dff a8_k1a_reg_29_ ( clk, n1335_r, a8_k1a[29], a8_v1[29] );
not U_inv2665 ( n1335_r, n1335 );
dff a8_out_1_reg_93_ ( clk, n1334_r, k8[93], k7b[93] );
not U_inv2666 ( n1334_r, n1334 );
dff a8_k1a_reg_30_ ( clk, n1334_r, a8_k1a[30], a8_v1[30] );
not U_inv2667 ( n1334_r, n1334 );
dff a8_out_1_reg_94_ ( clk, n1334_r, k8[94], k7b[94] );
not U_inv2668 ( n1334_r, n1334 );
dff a8_out_1_reg_95_ ( clk, n1334_r, k8[95], k7b[95] );
not U_inv2669 ( n1334_r, n1334 );
dff a9_k0a_reg_0_ ( clk, n1334_r, a9_k0a[0], k8[96] );
not U_inv2670 ( n1334_r, n1334 );
dff a9_out_1_reg_96_ ( clk, n1334_r, k9[96], k8b[96] );
not U_inv2671 ( n1334_r, n1334 );
dff a9_k0a_reg_1_ ( clk, n1334_r, a9_k0a[1], k8[97] );
not U_inv2672 ( n1334_r, n1334 );
dff a9_out_1_reg_97_ ( clk, n1334_r, k9[97], k8b[97] );
not U_inv2673 ( n1334_r, n1334 );
dff a9_k0a_reg_2_ ( clk, n1334_r, a9_k0a[2], k8[98] );
not U_inv2674 ( n1334_r, n1334 );
dff a9_out_1_reg_98_ ( clk, n1334_r, k9[98], k8b[98] );
not U_inv2675 ( n1334_r, n1334 );
dff a9_k0a_reg_3_ ( clk, n1334_r, a9_k0a[3], k8[99] );
not U_inv2676 ( n1334_r, n1334 );
dff a9_out_1_reg_99_ ( clk, n1334_r, k9[99], k8b[99] );
not U_inv2677 ( n1334_r, n1334 );
dff a9_k0a_reg_4_ ( clk, n1333_r, a9_k0a[4], k8[100] );
not U_inv2678 ( n1333_r, n1333 );
dff a9_out_1_reg_100_ ( clk, n1333_r, k9[100], k8b[100] );
not U_inv2679 ( n673, k9[100] );
not U_inv2680 ( n1333_r, n1333 );
dff a9_k0a_reg_5_ ( clk, n1333_r, a9_k0a[5], k8[101] );
not U_inv2681 ( n1333_r, n1333 );
dff a9_out_1_reg_101_ ( clk, n1333_r, k9[101], k8b[101] );
not U_inv2682 ( n674, k9[101] );
not U_inv2683 ( n1333_r, n1333 );
dff a9_k0a_reg_6_ ( clk, n1333_r, a9_k0a[6], k8[102] );
not U_inv2684 ( n1333_r, n1333 );
dff a9_out_1_reg_102_ ( clk, n1333_r, k9[102], k8b[102] );
not U_inv2685 ( n675, k9[102] );
not U_inv2686 ( n1333_r, n1333 );
dff a9_k0a_reg_7_ ( clk, n1333_r, a9_k0a[7], k8[103] );
not U_inv2687 ( n1333_r, n1333 );
dff a9_out_1_reg_103_ ( clk, n1333_r, k9[103], k8b[103] );
not U_inv2688 ( n676, k9[103] );
not U_inv2689 ( n1333_r, n1333 );
dff a9_k0a_reg_8_ ( clk, n1333_r, a9_k0a[8], k8[104] );
not U_inv2690 ( n1333_r, n1333 );
dff a9_out_1_reg_104_ ( clk, n1333_r, k9[104], k8b[104] );
not U_inv2691 ( n677, k9[104] );
not U_inv2692 ( n1333_r, n1333 );
dff a9_k0a_reg_9_ ( clk, n1333_r, a9_k0a[9], k8[105] );
not U_inv2693 ( n1333_r, n1333 );
dff a9_out_1_reg_105_ ( clk, n1333_r, k9[105], k8b[105] );
not U_inv2694 ( n678, k9[105] );
not U_inv2695 ( n1333_r, n1333 );
dff a9_k0a_reg_10_ ( clk, n1332_r, a9_k0a[10], k8[106] );
not U_inv2696 ( n1332_r, n1332 );
dff a9_out_1_reg_106_ ( clk, n1332_r, k9[106], k8b[106] );
not U_inv2697 ( n652, k9[106] );
not U_inv2698 ( n1332_r, n1332 );
dff a9_k0a_reg_11_ ( clk, n1332_r, a9_k0a[11], k8[107] );
not U_inv2699 ( n1332_r, n1332 );
dff a9_out_1_reg_107_ ( clk, n1332_r, k9[107], k8b[107] );
not U_inv2700 ( n653, k9[107] );
not U_inv2701 ( n1332_r, n1332 );
dff a9_k0a_reg_12_ ( clk, n1332_r, a9_k0a[12], k8[108] );
not U_inv2702 ( n1332_r, n1332 );
dff a9_out_1_reg_108_ ( clk, n1332_r, k9[108], k8b[108] );
not U_inv2703 ( n654, k9[108] );
not U_inv2704 ( n1332_r, n1332 );
dff a9_k0a_reg_13_ ( clk, n1332_r, a9_k0a[13], k8[109] );
not U_inv2705 ( n1332_r, n1332 );
dff a9_out_1_reg_109_ ( clk, n1332_r, k9[109], k8b[109] );
not U_inv2706 ( n655, k9[109] );
not U_inv2707 ( n1332_r, n1332 );
dff a9_k0a_reg_14_ ( clk, n1332_r, a9_k0a[14], k8[110] );
not U_inv2708 ( n1332_r, n1332 );
dff a9_out_1_reg_110_ ( clk, n1332_r, k9[110], k8b[110] );
not U_inv2709 ( n656, k9[110] );
not U_inv2710 ( n1332_r, n1332 );
dff a9_k0a_reg_15_ ( clk, n1332_r, a9_k0a[15], k8[111] );
not U_inv2711 ( n1332_r, n1332 );
dff a9_out_1_reg_111_ ( clk, n1332_r, k9[111], k8b[111] );
not U_inv2712 ( n657, k9[111] );
not U_inv2713 ( n1332_r, n1332 );
dff a9_k0a_reg_16_ ( clk, n1331_r, a9_k0a[16], k8[112] );
not U_inv2714 ( n1331_r, n1331 );
dff a9_out_1_reg_112_ ( clk, n1331_r, k9[112], k8b[112] );
not U_inv2715 ( n658, k9[112] );
not U_inv2716 ( n1331_r, n1331 );
dff a9_k0a_reg_17_ ( clk, n1331_r, a9_k0a[17], k8[113] );
not U_inv2717 ( n1331_r, n1331 );
dff a9_out_1_reg_113_ ( clk, n1331_r, k9[113], k8b[113] );
not U_inv2718 ( n659, k9[113] );
not U_inv2719 ( n1331_r, n1331 );
dff a9_k0a_reg_18_ ( clk, n1331_r, a9_k0a[18], k8[114] );
not U_inv2720 ( n1331_r, n1331 );
dff a9_out_1_reg_114_ ( clk, n1331_r, k9[114], k8b[114] );
not U_inv2721 ( n660, k9[114] );
not U_inv2722 ( n1331_r, n1331 );
dff a9_k0a_reg_19_ ( clk, n1331_r, a9_k0a[19], k8[115] );
not U_inv2723 ( n1331_r, n1331 );
dff a9_out_1_reg_115_ ( clk, n1331_r, k9[115], k8b[115] );
not U_inv2724 ( n661, k9[115] );
not U_inv2725 ( n1331_r, n1331 );
dff a9_k0a_reg_20_ ( clk, n1331_r, a9_k0a[20], k8[116] );
not U_inv2726 ( n1331_r, n1331 );
dff a9_out_1_reg_116_ ( clk, n1331_r, k9[116], k8b[116] );
not U_inv2727 ( n663, k9[116] );
not U_inv2728 ( n1331_r, n1331 );
dff a9_k0a_reg_21_ ( clk, n1331_r, a9_k0a[21], k8[117] );
not U_inv2729 ( n1331_r, n1331 );
dff a9_out_1_reg_117_ ( clk, n1331_r, k9[117], k8b[117] );
not U_inv2730 ( n664, k9[117] );
not U_inv2731 ( n1331_r, n1331 );
dff a9_k0a_reg_22_ ( clk, n1330_r, a9_k0a[22], k8[118] );
not U_inv2732 ( n1330_r, n1330 );
dff a9_out_1_reg_118_ ( clk, n1330_r, k9[118], k8b[118] );
not U_inv2733 ( n665, k9[118] );
not U_inv2734 ( n1330_r, n1330 );
dff a9_k0a_reg_23_ ( clk, n1330_r, a9_k0a[23], k8[119] );
not U_inv2735 ( n1330_r, n1330 );
dff a9_out_1_reg_119_ ( clk, n1330_r, k9[119], k8b[119] );
not U_inv2736 ( n666, k9[119] );
not U_inv2737 ( n1330_r, n1330 );
dff a9_k0a_reg_24_ ( clk, n1330_r, a9_k0a[24], n1292 );
not U_inv2738 ( n1330_r, n1330 );
dff a9_out_1_reg_120_ ( clk, n1330_r, k9[120], k8b[120] );
not U_inv2739 ( n667, k9[120] );
not U_inv2740 ( n1330_r, n1330 );
dff a9_k0a_reg_25_ ( clk, n1330_r, a9_k0a[25], n1293 );
not U_inv2741 ( n1330_r, n1330 );
dff a9_out_1_reg_121_ ( clk, n1330_r, ex_wire109, k8b[121] );
not U_inv2742 ( n1296, ex_wire109 );
not U_inv2743 ( n1330_r, n1330 );
dff a9_k0a_reg_26_ ( clk, n1330_r, a9_k0a[26], k8[122] );
not U_inv2744 ( n1330_r, n1330 );
dff a9_out_1_reg_122_ ( clk, n1330_r, ex_wire110, k8b[122] );
not U_inv2745 ( n1297, ex_wire110 );
not U_inv2746 ( n1330_r, n1330 );
dff a9_k0a_reg_27_ ( clk, n1330_r, a9_k0a[27], n1294 );
not U_inv2747 ( n1330_r, n1330 );
dff a9_out_1_reg_123_ ( clk, n1330_r, k9[123], k8b[123] );
not U_inv2748 ( n668, k9[123] );
not U_inv2749 ( n1330_r, n1330 );
dff a9_k0a_reg_28_ ( clk, n1329_r, a9_k0a[28], n1295 );
not U_inv2750 ( n1329_r, n1329 );
dff a9_out_1_reg_124_ ( clk, n1329_r, ex_wire111, k8b[124] );
not U_inv2751 ( n1298, ex_wire111 );
not U_inv2752 ( n1329_r, n1329 );
dff a9_k0a_reg_29_ ( clk, n1329_r, a9_k0a[29], k8[125] );
not U_inv2753 ( n1329_r, n1329 );
dff a9_out_1_reg_125_ ( clk, n1329_r, ex_wire112, k8b[125] );
not U_inv2754 ( n1299, ex_wire112 );
not U_inv2755 ( n1329_r, n1329 );
dff a9_k0a_reg_30_ ( clk, n1329_r, a9_k0a[30], k8[126] );
not U_inv2756 ( n1329_r, n1329 );
dff a9_out_1_reg_126_ ( clk, n1329_r, k9[126], k8b[126] );
not U_inv2757 ( n670, k9[126] );
not U_inv2758 ( n1329_r, n1329 );
dff a9_k0a_reg_31_ ( clk, n1329_r, a9_k0a[31], k8[127] );
not U_inv2759 ( n1329_r, n1329 );
dff a9_out_1_reg_127_ ( clk, n1329_r, k9[127], k8b[127] );
not U_inv2760 ( n671, k9[127] );
not U_inv2761 ( n1329_r, n1329 );
dff a9_k3a_reg_0_ ( clk, n1329_r, a9_k3a[0], a9_v3[0] );
not U_inv2762 ( n1329_r, n1329 );
dff a9_out_1_reg_0_ ( clk, n1329_r, k9[0], k8b[0] );
not U_inv2763 ( n1329_r, n1329 );
dff a9_k3a_reg_1_ ( clk, n1329_r, a9_k3a[1], a9_v3[1] );
not U_inv2764 ( n1329_r, n1329 );
dff a9_out_1_reg_1_ ( clk, n1329_r, k9[1], k8b[1] );
not U_inv2765 ( n1329_r, n1329 );
dff a9_k3a_reg_2_ ( clk, n1328_r, a9_k3a[2], a9_v3[2] );
not U_inv2766 ( n1328_r, n1328 );
dff a9_out_1_reg_2_ ( clk, n1328_r, k9[2], k8b[2] );
not U_inv2767 ( n1328_r, n1328 );
dff a9_k3a_reg_3_ ( clk, n1328_r, a9_k3a[3], a9_v3[3] );
not U_inv2768 ( n1328_r, n1328 );
dff a9_out_1_reg_3_ ( clk, n1328_r, k9[3], k8b[3] );
not U_inv2769 ( n1328_r, n1328 );
dff a9_k3a_reg_4_ ( clk, n1328_r, a9_k3a[4], a9_v3[4] );
not U_inv2770 ( n1328_r, n1328 );
dff a9_out_1_reg_4_ ( clk, n1328_r, k9[4], k8b[4] );
not U_inv2771 ( n1328_r, n1328 );
dff a9_k3a_reg_5_ ( clk, n1328_r, a9_k3a[5], a9_v3[5] );
not U_inv2772 ( n1328_r, n1328 );
dff a9_out_1_reg_5_ ( clk, n1328_r, k9[5], k8b[5] );
not U_inv2773 ( n1328_r, n1328 );
dff a9_k3a_reg_6_ ( clk, n1328_r, a9_k3a[6], a9_v3[6] );
not U_inv2774 ( n1328_r, n1328 );
dff a9_out_1_reg_6_ ( clk, n1328_r, k9[6], k8b[6] );
not U_inv2775 ( n1328_r, n1328 );
dff a9_k3a_reg_7_ ( clk, n1328_r, a9_k3a[7], a9_v3[7] );
not U_inv2776 ( n1328_r, n1328 );
dff a9_out_1_reg_7_ ( clk, n1328_r, k9[7], k8b[7] );
not U_inv2777 ( n1328_r, n1328 );
dff a9_k3a_reg_8_ ( clk, n1327_r, a9_k3a[8], a9_v3[8] );
not U_inv2778 ( n1327_r, n1327 );
dff a9_out_1_reg_8_ ( clk, n1327_r, k9[8], k8b[8] );
not U_inv2779 ( n1327_r, n1327 );
dff a9_k3a_reg_9_ ( clk, n1327_r, a9_k3a[9], a9_v3[9] );
not U_inv2780 ( n1327_r, n1327 );
dff a9_out_1_reg_9_ ( clk, n1327_r, k9[9], k8b[9] );
not U_inv2781 ( n1327_r, n1327 );
dff a9_k3a_reg_10_ ( clk, n1327_r, a9_k3a[10], a9_v3[10] );
not U_inv2782 ( n1327_r, n1327 );
dff a9_out_1_reg_10_ ( clk, n1327_r, k9[10], k8b[10] );
not U_inv2783 ( n1327_r, n1327 );
dff a9_k3a_reg_11_ ( clk, n1327_r, a9_k3a[11], a9_v3[11] );
not U_inv2784 ( n1327_r, n1327 );
dff a9_out_1_reg_11_ ( clk, n1327_r, k9[11], k8b[11] );
not U_inv2785 ( n1327_r, n1327 );
dff a9_k3a_reg_12_ ( clk, n1327_r, a9_k3a[12], a9_v3[12] );
not U_inv2786 ( n1327_r, n1327 );
dff a9_out_1_reg_12_ ( clk, n1327_r, k9[12], k8b[12] );
not U_inv2787 ( n1327_r, n1327 );
dff a9_k3a_reg_13_ ( clk, n1327_r, a9_k3a[13], a9_v3[13] );
not U_inv2788 ( n1327_r, n1327 );
dff a9_out_1_reg_13_ ( clk, n1327_r, k9[13], k8b[13] );
not U_inv2789 ( n1327_r, n1327 );
dff a9_k3a_reg_14_ ( clk, n1326_r, a9_k3a[14], a9_v3[14] );
not U_inv2790 ( n1326_r, n1326 );
dff a9_out_1_reg_14_ ( clk, n1326_r, k9[14], k8b[14] );
not U_inv2791 ( n1326_r, n1326 );
dff a9_k3a_reg_15_ ( clk, n1326_r, a9_k3a[15], a9_v3[15] );
not U_inv2792 ( n1326_r, n1326 );
dff a9_out_1_reg_15_ ( clk, n1326_r, k9[15], k8b[15] );
not U_inv2793 ( n1326_r, n1326 );
dff a9_k3a_reg_16_ ( clk, n1326_r, a9_k3a[16], a9_v3[16] );
not U_inv2794 ( n1326_r, n1326 );
dff a9_out_1_reg_16_ ( clk, n1326_r, k9[16], k8b[16] );
not U_inv2795 ( n1326_r, n1326 );
dff a9_k3a_reg_17_ ( clk, n1326_r, a9_k3a[17], a9_v3[17] );
not U_inv2796 ( n1326_r, n1326 );
dff a9_out_1_reg_17_ ( clk, n1326_r, k9[17], k8b[17] );
not U_inv2797 ( n1326_r, n1326 );
dff a9_k3a_reg_18_ ( clk, n1326_r, a9_k3a[18], a9_v3[18] );
not U_inv2798 ( n1326_r, n1326 );
dff a9_out_1_reg_18_ ( clk, n1326_r, k9[18], k8b[18] );
not U_inv2799 ( n1326_r, n1326 );
dff a9_k3a_reg_19_ ( clk, n1326_r, a9_k3a[19], a9_v3[19] );
not U_inv2800 ( n1326_r, n1326 );
dff a9_out_1_reg_19_ ( clk, n1326_r, k9[19], k8b[19] );
not U_inv2801 ( n1326_r, n1326 );
dff a9_k3a_reg_20_ ( clk, n1325_r, a9_k3a[20], a9_v3[20] );
not U_inv2802 ( n1325_r, n1325 );
dff a9_out_1_reg_20_ ( clk, n1325_r, k9[20], k8b[20] );
not U_inv2803 ( n1325_r, n1325 );
dff a9_k3a_reg_21_ ( clk, n1325_r, a9_k3a[21], a9_v3[21] );
not U_inv2804 ( n1325_r, n1325 );
dff a9_out_1_reg_21_ ( clk, n1325_r, k9[21], k8b[21] );
not U_inv2805 ( n1325_r, n1325 );
dff a9_k3a_reg_22_ ( clk, n1325_r, a9_k3a[22], a9_v3[22] );
not U_inv2806 ( n1325_r, n1325 );
dff a9_out_1_reg_22_ ( clk, n1325_r, k9[22], k8b[22] );
not U_inv2807 ( n1325_r, n1325 );
dff a9_k3a_reg_23_ ( clk, n1325_r, a9_k3a[23], a9_v3[23] );
not U_inv2808 ( n1325_r, n1325 );
dff a9_out_1_reg_23_ ( clk, n1325_r, k9[23], k8b[23] );
not U_inv2809 ( n1325_r, n1325 );
dff a9_k3a_reg_24_ ( clk, n1325_r, a9_k3a[24], a9_v3[24] );
not U_inv2810 ( n1325_r, n1325 );
dff a9_out_1_reg_24_ ( clk, n1325_r, k9[24], k8b[24] );
not U_inv2811 ( n1325_r, n1325 );
dff a9_k3a_reg_25_ ( clk, n1325_r, a9_k3a[25], a9_v3[25] );
not U_inv2812 ( n1325_r, n1325 );
dff a9_out_1_reg_25_ ( clk, n1325_r, k9[25], k8b[25] );
not U_inv2813 ( n1325_r, n1325 );
dff a9_k3a_reg_26_ ( clk, n1324_r, a9_k3a[26], a9_v3[26] );
not U_inv2814 ( n1324_r, n1324 );
dff a9_out_1_reg_26_ ( clk, n1324_r, k9[26], k8b[26] );
not U_inv2815 ( n1324_r, n1324 );
dff a9_k3a_reg_27_ ( clk, n1324_r, a9_k3a[27], a9_v3[27] );
not U_inv2816 ( n1324_r, n1324 );
dff a9_out_1_reg_27_ ( clk, n1324_r, k9[27], k8b[27] );
not U_inv2817 ( n1324_r, n1324 );
dff a9_k3a_reg_28_ ( clk, n1324_r, a9_k3a[28], a9_v3[28] );
not U_inv2818 ( n1324_r, n1324 );
dff a9_out_1_reg_28_ ( clk, n1324_r, k9[28], k8b[28] );
not U_inv2819 ( n1324_r, n1324 );
dff a9_k3a_reg_29_ ( clk, n1324_r, a9_k3a[29], a9_v3[29] );
not U_inv2820 ( n1324_r, n1324 );
dff a9_out_1_reg_29_ ( clk, n1324_r, k9[29], k8b[29] );
not U_inv2821 ( n1324_r, n1324 );
dff a9_k3a_reg_30_ ( clk, n1324_r, a9_k3a[30], a9_v3[30] );
not U_inv2822 ( n1324_r, n1324 );
dff a9_out_1_reg_30_ ( clk, n1324_r, k9[30], k8b[30] );
not U_inv2823 ( n1324_r, n1324 );
dff a9_k2a_reg_0_ ( clk, n1324_r, a9_k2a[0], a9_v2[0] );
not U_inv2824 ( n1324_r, n1324 );
dff a9_out_1_reg_32_ ( clk, n1324_r, k9[32], k8b[32] );
not U_inv2825 ( n1324_r, n1324 );
dff a9_k2a_reg_1_ ( clk, n1323_r, a9_k2a[1], a9_v2[1] );
not U_inv2826 ( n1323_r, n1323 );
dff a9_out_1_reg_33_ ( clk, n1323_r, k9[33], k8b[33] );
not U_inv2827 ( n1323_r, n1323 );
dff a9_k2a_reg_2_ ( clk, n1323_r, a9_k2a[2], a9_v2[2] );
not U_inv2828 ( n1323_r, n1323 );
dff a9_out_1_reg_34_ ( clk, n1323_r, k9[34], k8b[34] );
not U_inv2829 ( n1323_r, n1323 );
dff a9_k2a_reg_3_ ( clk, n1323_r, a9_k2a[3], a9_v2[3] );
not U_inv2830 ( n1323_r, n1323 );
dff a9_out_1_reg_35_ ( clk, n1323_r, k9[35], k8b[35] );
not U_inv2831 ( n1323_r, n1323 );
dff a9_k2a_reg_4_ ( clk, n1323_r, a9_k2a[4], a9_v2[4] );
not U_inv2832 ( n1323_r, n1323 );
dff a9_out_1_reg_36_ ( clk, n1323_r, k9[36], k8b[36] );
not U_inv2833 ( n1323_r, n1323 );
dff a9_k2a_reg_5_ ( clk, n1323_r, a9_k2a[5], a9_v2[5] );
not U_inv2834 ( n1323_r, n1323 );
dff a9_out_1_reg_37_ ( clk, n1323_r, k9[37], k8b[37] );
not U_inv2835 ( n1323_r, n1323 );
dff a9_k2a_reg_6_ ( clk, n1323_r, a9_k2a[6], a9_v2[6] );
not U_inv2836 ( n1323_r, n1323 );
dff a9_out_1_reg_38_ ( clk, n1323_r, k9[38], k8b[38] );
not U_inv2837 ( n1323_r, n1323 );
dff a9_k2a_reg_7_ ( clk, n1322_r, a9_k2a[7], a9_v2[7] );
not U_inv2838 ( n1322_r, n1322 );
dff a9_out_1_reg_39_ ( clk, n1322_r, k9[39], k8b[39] );
not U_inv2839 ( n1322_r, n1322 );
dff a9_k2a_reg_8_ ( clk, n1322_r, a9_k2a[8], a9_v2[8] );
not U_inv2840 ( n1322_r, n1322 );
dff a9_out_1_reg_40_ ( clk, n1322_r, k9[40], k8b[40] );
not U_inv2841 ( n1322_r, n1322 );
dff a9_k2a_reg_9_ ( clk, n1322_r, a9_k2a[9], a9_v2[9] );
not U_inv2842 ( n1322_r, n1322 );
dff a9_out_1_reg_41_ ( clk, n1322_r, k9[41], k8b[41] );
not U_inv2843 ( n1322_r, n1322 );
dff a9_k2a_reg_10_ ( clk, n1322_r, a9_k2a[10], a9_v2[10] );
not U_inv2844 ( n1322_r, n1322 );
dff a9_out_1_reg_42_ ( clk, n1322_r, k9[42], k8b[42] );
not U_inv2845 ( n1322_r, n1322 );
dff a9_k2a_reg_11_ ( clk, n1322_r, a9_k2a[11], a9_v2[11] );
not U_inv2846 ( n1322_r, n1322 );
dff a9_out_1_reg_43_ ( clk, n1322_r, k9[43], k8b[43] );
not U_inv2847 ( n1322_r, n1322 );
dff a9_k2a_reg_12_ ( clk, n1322_r, a9_k2a[12], a9_v2[12] );
not U_inv2848 ( n1322_r, n1322 );
dff a9_out_1_reg_44_ ( clk, n1322_r, k9[44], k8b[44] );
not U_inv2849 ( n1322_r, n1322 );
dff a9_k2a_reg_13_ ( clk, n1321_r, a9_k2a[13], a9_v2[13] );
not U_inv2850 ( n1321_r, n1321 );
dff a9_out_1_reg_45_ ( clk, n1321_r, k9[45], k8b[45] );
not U_inv2851 ( n1321_r, n1321 );
dff a9_k2a_reg_14_ ( clk, n1321_r, a9_k2a[14], a9_v2[14] );
not U_inv2852 ( n1321_r, n1321 );
dff a9_out_1_reg_46_ ( clk, n1321_r, k9[46], k8b[46] );
not U_inv2853 ( n1321_r, n1321 );
dff a9_k2a_reg_15_ ( clk, n1321_r, a9_k2a[15], a9_v2[15] );
not U_inv2854 ( n1321_r, n1321 );
dff a9_out_1_reg_47_ ( clk, n1321_r, k9[47], k8b[47] );
not U_inv2855 ( n1321_r, n1321 );
dff a9_k2a_reg_16_ ( clk, n1321_r, a9_k2a[16], a9_v2[16] );
not U_inv2856 ( n1321_r, n1321 );
dff a9_out_1_reg_48_ ( clk, n1321_r, k9[48], k8b[48] );
not U_inv2857 ( n1321_r, n1321 );
dff a9_k2a_reg_17_ ( clk, n1321_r, a9_k2a[17], a9_v2[17] );
not U_inv2858 ( n1321_r, n1321 );
dff a9_out_1_reg_49_ ( clk, n1321_r, k9[49], k8b[49] );
not U_inv2859 ( n1321_r, n1321 );
dff a9_k2a_reg_18_ ( clk, n1321_r, a9_k2a[18], a9_v2[18] );
not U_inv2860 ( n1321_r, n1321 );
dff a9_out_1_reg_50_ ( clk, n1321_r, k9[50], k8b[50] );
not U_inv2861 ( n1321_r, n1321 );
dff a9_k2a_reg_19_ ( clk, n1320_r, a9_k2a[19], a9_v2[19] );
not U_inv2862 ( n1320_r, n1320 );
dff a9_out_1_reg_51_ ( clk, n1320_r, k9[51], k8b[51] );
not U_inv2863 ( n1320_r, n1320 );
dff a9_k2a_reg_20_ ( clk, n1320_r, a9_k2a[20], a9_v2[20] );
not U_inv2864 ( n1320_r, n1320 );
dff a9_out_1_reg_52_ ( clk, n1320_r, k9[52], k8b[52] );
not U_inv2865 ( n1320_r, n1320 );
dff a9_k2a_reg_21_ ( clk, n1320_r, a9_k2a[21], a9_v2[21] );
not U_inv2866 ( n1320_r, n1320 );
dff a9_out_1_reg_53_ ( clk, n1320_r, k9[53], k8b[53] );
not U_inv2867 ( n1320_r, n1320 );
dff a9_k2a_reg_22_ ( clk, n1320_r, a9_k2a[22], a9_v2[22] );
not U_inv2868 ( n1320_r, n1320 );
dff a9_out_1_reg_54_ ( clk, n1320_r, k9[54], k8b[54] );
not U_inv2869 ( n1320_r, n1320 );
dff a9_k2a_reg_23_ ( clk, n1320_r, a9_k2a[23], a9_v2[23] );
not U_inv2870 ( n1320_r, n1320 );
dff a9_out_1_reg_55_ ( clk, n1320_r, k9[55], k8b[55] );
not U_inv2871 ( n1320_r, n1320 );
dff a9_k2a_reg_24_ ( clk, n1320_r, a9_k2a[24], a9_v2[24] );
not U_inv2872 ( n1320_r, n1320 );
dff a9_out_1_reg_56_ ( clk, n1320_r, k9[56], k8b[56] );
not U_inv2873 ( n1320_r, n1320 );
dff a9_k2a_reg_25_ ( clk, n1319_r, a9_k2a[25], a9_v2[25] );
not U_inv2874 ( n1319_r, n1319 );
dff a9_out_1_reg_57_ ( clk, n1319_r, k9[57], k8b[57] );
not U_inv2875 ( n1319_r, n1319 );
dff a9_k2a_reg_26_ ( clk, n1319_r, a9_k2a[26], a9_v2[26] );
not U_inv2876 ( n1319_r, n1319 );
dff a9_out_1_reg_58_ ( clk, n1319_r, k9[58], k8b[58] );
not U_inv2877 ( n1319_r, n1319 );
dff a9_k2a_reg_27_ ( clk, n1319_r, a9_k2a[27], a9_v2[27] );
not U_inv2878 ( n1319_r, n1319 );
dff a9_out_1_reg_59_ ( clk, n1319_r, k9[59], k8b[59] );
not U_inv2879 ( n1319_r, n1319 );
dff a9_k2a_reg_28_ ( clk, n1319_r, a9_k2a[28], a9_v2[28] );
not U_inv2880 ( n1319_r, n1319 );
dff a9_out_1_reg_60_ ( clk, n1319_r, k9[60], k8b[60] );
not U_inv2881 ( n1319_r, n1319 );
dff a9_k2a_reg_29_ ( clk, n1319_r, a9_k2a[29], a9_v2[29] );
not U_inv2882 ( n1319_r, n1319 );
dff a9_out_1_reg_61_ ( clk, n1319_r, k9[61], k8b[61] );
not U_inv2883 ( n1319_r, n1319 );
dff a9_k2a_reg_30_ ( clk, n1319_r, a9_k2a[30], a9_v2[30] );
not U_inv2884 ( n1319_r, n1319 );
dff a9_out_1_reg_62_ ( clk, n1319_r, k9[62], k8b[62] );
not U_inv2885 ( n1319_r, n1319 );
dff a9_k2a_reg_31_ ( clk, n1318_r, a9_k2a[31], a9_v2[31] );
not U_inv2886 ( n1318_r, n1318 );
dff a9_out_1_reg_63_ ( clk, n1318_r, k9[63], k8b[63] );
not U_inv2887 ( n1318_r, n1318 );
dff a9_k1a_reg_0_ ( clk, n1318_r, a9_k1a[0], a9_v1[0] );
not U_inv2888 ( n1318_r, n1318 );
dff a9_out_1_reg_64_ ( clk, n1318_r, ex_wire113, k8b[64] );
not U_inv2889 ( n651, ex_wire113 );
not U_inv2890 ( n1318_r, n1318 );
dff a9_k1a_reg_1_ ( clk, n1318_r, a9_k1a[1], a9_v1[1] );
not U_inv2891 ( n1318_r, n1318 );
dff a9_out_1_reg_65_ ( clk, n1318_r, ex_wire114, k8b[65] );
not U_inv2892 ( n662, ex_wire114 );
not U_inv2893 ( n1318_r, n1318 );
dff a9_k1a_reg_2_ ( clk, n1318_r, a9_k1a[2], a9_v1[2] );
not U_inv2894 ( n1318_r, n1318 );
dff a9_out_1_reg_66_ ( clk, n1318_r, ex_wire115, k8b[66] );
not U_inv2895 ( n669, ex_wire115 );
not U_inv2896 ( n1318_r, n1318 );
dff a9_k1a_reg_3_ ( clk, n1318_r, a9_k1a[3], a9_v1[3] );
not U_inv2897 ( n1318_r, n1318 );
dff a9_out_1_reg_67_ ( clk, n1318_r, ex_wire116, k8b[67] );
not U_inv2898 ( n672, ex_wire116 );
not U_inv2899 ( n1318_r, n1318 );
dff a9_k1a_reg_4_ ( clk, n1318_r, a9_k1a[4], a9_v1[4] );
not U_inv2900 ( n1318_r, n1318 );
dff a9_out_1_reg_68_ ( clk, n1318_r, k9[68], k8b[68] );
not U_inv2901 ( n1318_r, n1318 );
dff a9_k1a_reg_5_ ( clk, n1317_r, a9_k1a[5], a9_v1[5] );
not U_inv2902 ( n1317_r, n1317 );
dff a9_out_1_reg_69_ ( clk, n1317_r, k9[69], k8b[69] );
not U_inv2903 ( n1317_r, n1317 );
dff a9_k1a_reg_6_ ( clk, n1317_r, a9_k1a[6], a9_v1[6] );
not U_inv2904 ( n1317_r, n1317 );
dff a9_out_1_reg_70_ ( clk, n1317_r, k9[70], k8b[70] );
not U_inv2905 ( n1317_r, n1317 );
dff a9_k1a_reg_7_ ( clk, n1317_r, a9_k1a[7], a9_v1[7] );
not U_inv2906 ( n1317_r, n1317 );
dff a9_out_1_reg_71_ ( clk, n1317_r, k9[71], k8b[71] );
not U_inv2907 ( n1317_r, n1317 );
dff a9_k1a_reg_8_ ( clk, n1317_r, a9_k1a[8], a9_v1[8] );
not U_inv2908 ( n1317_r, n1317 );
dff a9_out_1_reg_72_ ( clk, n1317_r, k9[72], k8b[72] );
not U_inv2909 ( n1317_r, n1317 );
dff a9_k1a_reg_9_ ( clk, n1317_r, a9_k1a[9], a9_v1[9] );
not U_inv2910 ( n1317_r, n1317 );
dff a9_out_1_reg_73_ ( clk, n1317_r, k9[73], k8b[73] );
not U_inv2911 ( n1317_r, n1317 );
dff a9_k1a_reg_10_ ( clk, n1317_r, a9_k1a[10], a9_v1[10] );
not U_inv2912 ( n1317_r, n1317 );
dff a9_out_1_reg_74_ ( clk, n1317_r, k9[74], k8b[74] );
not U_inv2913 ( n1317_r, n1317 );
dff a9_k1a_reg_11_ ( clk, n1316_r, a9_k1a[11], a9_v1[11] );
not U_inv2914 ( n1316_r, n1316 );
dff a9_out_1_reg_75_ ( clk, n1316_r, k9[75], k8b[75] );
not U_inv2915 ( n1316_r, n1316 );
dff a9_k1a_reg_12_ ( clk, n1316_r, a9_k1a[12], a9_v1[12] );
not U_inv2916 ( n1316_r, n1316 );
dff a9_out_1_reg_76_ ( clk, n1316_r, k9[76], k8b[76] );
not U_inv2917 ( n1316_r, n1316 );
dff a9_k1a_reg_13_ ( clk, n1316_r, a9_k1a[13], a9_v1[13] );
not U_inv2918 ( n1316_r, n1316 );
dff a9_out_1_reg_77_ ( clk, n1316_r, k9[77], k8b[77] );
not U_inv2919 ( n1316_r, n1316 );
dff a9_k1a_reg_14_ ( clk, n1316_r, a9_k1a[14], a9_v1[14] );
not U_inv2920 ( n1316_r, n1316 );
dff a9_out_1_reg_78_ ( clk, n1316_r, k9[78], k8b[78] );
not U_inv2921 ( n1316_r, n1316 );
dff a9_k1a_reg_15_ ( clk, n1316_r, a9_k1a[15], a9_v1[15] );
not U_inv2922 ( n1316_r, n1316 );
dff a9_out_1_reg_79_ ( clk, n1316_r, k9[79], k8b[79] );
not U_inv2923 ( n1316_r, n1316 );
dff a9_k1a_reg_16_ ( clk, n1316_r, a9_k1a[16], a9_v1[16] );
not U_inv2924 ( n1316_r, n1316 );
dff a9_out_1_reg_80_ ( clk, n1316_r, k9[80], k8b[80] );
not U_inv2925 ( n1316_r, n1316 );
dff a9_k1a_reg_17_ ( clk, n1315_r, a9_k1a[17], a9_v1[17] );
not U_inv2926 ( n1315_r, n1315 );
dff a9_out_1_reg_81_ ( clk, n1315_r, k9[81], k8b[81] );
not U_inv2927 ( n1315_r, n1315 );
dff a9_k1a_reg_18_ ( clk, n1315_r, a9_k1a[18], a9_v1[18] );
not U_inv2928 ( n1315_r, n1315 );
dff a9_out_1_reg_82_ ( clk, n1315_r, k9[82], k8b[82] );
not U_inv2929 ( n1315_r, n1315 );
dff a9_k1a_reg_19_ ( clk, n1315_r, a9_k1a[19], a9_v1[19] );
not U_inv2930 ( n1315_r, n1315 );
dff a9_out_1_reg_83_ ( clk, n1315_r, k9[83], k8b[83] );
not U_inv2931 ( n1315_r, n1315 );
dff a9_k1a_reg_20_ ( clk, n1315_r, a9_k1a[20], a9_v1[20] );
not U_inv2932 ( n1315_r, n1315 );
dff a9_out_1_reg_84_ ( clk, n1315_r, k9[84], k8b[84] );
not U_inv2933 ( n1315_r, n1315 );
dff a9_k1a_reg_21_ ( clk, n1315_r, a9_k1a[21], a9_v1[21] );
not U_inv2934 ( n1315_r, n1315 );
dff a9_out_1_reg_85_ ( clk, n1315_r, k9[85], k8b[85] );
not U_inv2935 ( n1315_r, n1315 );
dff a9_k1a_reg_22_ ( clk, n1315_r, a9_k1a[22], a9_v1[22] );
not U_inv2936 ( n1315_r, n1315 );
dff a9_out_1_reg_86_ ( clk, n1315_r, k9[86], k8b[86] );
not U_inv2937 ( n1315_r, n1315 );
dff a9_k1a_reg_23_ ( clk, n1314_r, a9_k1a[23], a9_v1[23] );
not U_inv2938 ( n1314_r, n1314 );
dff a9_out_1_reg_87_ ( clk, n1314_r, k9[87], k8b[87] );
not U_inv2939 ( n1314_r, n1314 );
dff a9_k1a_reg_24_ ( clk, n1314_r, a9_k1a[24], a9_v1[24] );
not U_inv2940 ( n1314_r, n1314 );
dff a9_out_1_reg_88_ ( clk, n1314_r, k9[88], k8b[88] );
not U_inv2941 ( n1314_r, n1314 );
dff a9_k1a_reg_25_ ( clk, n1314_r, a9_k1a[25], a9_v1[25] );
not U_inv2942 ( n1314_r, n1314 );
dff a9_out_1_reg_89_ ( clk, n1314_r, k9[89], k8b[89] );
not U_inv2943 ( n1314_r, n1314 );
dff a9_k1a_reg_26_ ( clk, n1314_r, a9_k1a[26], a9_v1[26] );
not U_inv2944 ( n1314_r, n1314 );
dff a9_out_1_reg_90_ ( clk, n1314_r, k9[90], k8b[90] );
not U_inv2945 ( n1314_r, n1314 );
dff a9_k1a_reg_27_ ( clk, n1314_r, a9_k1a[27], a9_v1[27] );
not U_inv2946 ( n1314_r, n1314 );
dff a9_out_1_reg_91_ ( clk, n1314_r, k9[91], k8b[91] );
not U_inv2947 ( n1314_r, n1314 );
dff a9_k1a_reg_28_ ( clk, n1314_r, a9_k1a[28], a9_v1[28] );
not U_inv2948 ( n1314_r, n1314 );
dff a9_out_1_reg_92_ ( clk, n1314_r, k9[92], k8b[92] );
not U_inv2949 ( n1314_r, n1314 );
dff a9_k1a_reg_29_ ( clk, n1313_r, a9_k1a[29], a9_v1[29] );
not U_inv2950 ( n1313_r, n1313 );
dff a9_out_1_reg_93_ ( clk, n1313_r, k9[93], k8b[93] );
not U_inv2951 ( n1313_r, n1313 );
dff a9_k1a_reg_30_ ( clk, n1313_r, a9_k1a[30], a9_v1[30] );
not U_inv2952 ( n1313_r, n1313 );
dff a9_out_1_reg_94_ ( clk, n1313_r, k9[94], k8b[94] );
not U_inv2953 ( n1313_r, n1313 );
dff a9_out_1_reg_95_ ( clk, n1313_r, k9[95], k8b[95] );
not U_inv2954 ( n1313_r, n1313 );
dff a10_k0a_reg_0_ ( clk, n1313_r, a10_k0a[0], k9[96] );
not U_inv2955 ( n1313_r, n1313 );
dff a10_k0a_reg_1_ ( clk, n1313_r, a10_k0a[1], k9[97] );
not U_inv2956 ( n1313_r, n1313 );
dff a10_k0a_reg_2_ ( clk, n1313_r, a10_k0a[2], k9[98] );
not U_inv2957 ( n1313_r, n1313 );
dff a10_k0a_reg_3_ ( clk, n1313_r, a10_k0a[3], k9[99] );
not U_inv2958 ( n1313_r, n1313 );
dff a10_k0a_reg_4_ ( clk, n1313_r, a10_k0a[4], k9[100] );
not U_inv2959 ( n1313_r, n1313 );
dff a10_k0a_reg_5_ ( clk, n1313_r, a10_k0a[5], k9[101] );
not U_inv2960 ( n1313_r, n1313 );
dff a10_k0a_reg_6_ ( clk, n1313_r, a10_k0a[6], k9[102] );
not U_inv2961 ( n1313_r, n1313 );
dff a10_k0a_reg_7_ ( clk, n1312_r, a10_k0a[7], k9[103] );
not U_inv2962 ( n1312_r, n1312 );
dff a10_k0a_reg_8_ ( clk, n1312_r, a10_k0a[8], k9[104] );
not U_inv2963 ( n1312_r, n1312 );
dff a10_k0a_reg_9_ ( clk, n1312_r, a10_k0a[9], k9[105] );
not U_inv2964 ( n1312_r, n1312 );
dff a10_k0a_reg_10_ ( clk, n1312_r, a10_k0a[10], k9[106] );
not U_inv2965 ( n1312_r, n1312 );
dff a10_k0a_reg_11_ ( clk, n1312_r, a10_k0a[11], k9[107] );
not U_inv2966 ( n1312_r, n1312 );
dff a10_k0a_reg_12_ ( clk, n1312_r, a10_k0a[12], k9[108] );
not U_inv2967 ( n1312_r, n1312 );
dff a10_k0a_reg_13_ ( clk, n1312_r, a10_k0a[13], k9[109] );
not U_inv2968 ( n1312_r, n1312 );
dff a10_k0a_reg_14_ ( clk, n1312_r, a10_k0a[14], k9[110] );
not U_inv2969 ( n1312_r, n1312 );
dff a10_k0a_reg_15_ ( clk, n1312_r, a10_k0a[15], k9[111] );
not U_inv2970 ( n1312_r, n1312 );
dff a10_k0a_reg_16_ ( clk, n1312_r, a10_k0a[16], k9[112] );
not U_inv2971 ( n1312_r, n1312 );
dff a10_k0a_reg_17_ ( clk, n1312_r, a10_k0a[17], k9[113] );
not U_inv2972 ( n1312_r, n1312 );
dff a10_k0a_reg_18_ ( clk, n1312_r, a10_k0a[18], k9[114] );
not U_inv2973 ( n1312_r, n1312 );
dff a10_k0a_reg_19_ ( clk, n1311_r, a10_k0a[19], k9[115] );
not U_inv2974 ( n1311_r, n1311 );
dff a10_k0a_reg_20_ ( clk, n1311_r, a10_k0a[20], k9[116] );
not U_inv2975 ( n1311_r, n1311 );
dff a10_k0a_reg_21_ ( clk, n1311_r, a10_k0a[21], k9[117] );
not U_inv2976 ( n1311_r, n1311 );
dff a10_k0a_reg_22_ ( clk, n1311_r, a10_k0a[22], k9[118] );
not U_inv2977 ( n1311_r, n1311 );
dff a10_k0a_reg_23_ ( clk, n1311_r, a10_k0a[23], k9[119] );
not U_inv2978 ( n1311_r, n1311 );
dff a10_k0a_reg_24_ ( clk, n1311_r, a10_k0a[24], k9[120] );
not U_inv2979 ( n1311_r, n1311 );
dff a10_k0a_reg_25_ ( clk, n1311_r, a10_k0a[25], n1296 );
not U_inv2980 ( n1311_r, n1311 );
dff a10_k0a_reg_26_ ( clk, n1311_r, a10_k0a[26], n1297 );
not U_inv2981 ( n1311_r, n1311 );
dff a10_k0a_reg_27_ ( clk, n1311_r, a10_k0a[27], k9[123] );
not U_inv2982 ( n1311_r, n1311 );
dff a10_k0a_reg_28_ ( clk, n1311_r, a10_k0a[28], n1298 );
not U_inv2983 ( n1311_r, n1311 );
dff a10_k0a_reg_29_ ( clk, n1311_r, a10_k0a[29], n1299 );
not U_inv2984 ( n1311_r, n1311 );
dff a10_k0a_reg_30_ ( clk, n1311_r, a10_k0a[30], k9[126] );
not U_inv2985 ( n1311_r, n1311 );
dff a10_k0a_reg_31_ ( clk, n1310_r, a10_k0a[31], k9[127] );
not U_inv2986 ( n1310_r, n1310 );
dff a10_k3a_reg_0_ ( clk, n1310_r, a10_k3a[0], a10_v3[0] );
not U_inv2987 ( n1310_r, n1310 );
dff a10_k3a_reg_1_ ( clk, n1310_r, a10_k3a[1], a10_v3[1] );
not U_inv2988 ( n1310_r, n1310 );
dff a10_k3a_reg_2_ ( clk, n1310_r, a10_k3a[2], a10_v3[2] );
not U_inv2989 ( n1310_r, n1310 );
dff a10_k3a_reg_3_ ( clk, n1310_r, a10_k3a[3], a10_v3[3] );
not U_inv2990 ( n1310_r, n1310 );
dff a10_k3a_reg_4_ ( clk, n1310_r, a10_k3a[4], a10_v3[4] );
not U_inv2991 ( n1310_r, n1310 );
dff a10_k3a_reg_5_ ( clk, n1310_r, a10_k3a[5], a10_v3[5] );
not U_inv2992 ( n1310_r, n1310 );
dff a10_k3a_reg_6_ ( clk, n1310_r, a10_k3a[6], a10_v3[6] );
not U_inv2993 ( n1310_r, n1310 );
dff a10_k3a_reg_7_ ( clk, n1310_r, a10_k3a[7], a10_v3[7] );
not U_inv2994 ( n1310_r, n1310 );
dff a10_k3a_reg_8_ ( clk, n1310_r, a10_k3a[8], a10_v3[8] );
not U_inv2995 ( n1310_r, n1310 );
dff a10_k3a_reg_9_ ( clk, n1310_r, a10_k3a[9], a10_v3[9] );
not U_inv2996 ( n1310_r, n1310 );
dff a10_k3a_reg_10_ ( clk, n1310_r, a10_k3a[10], a10_v3[10] );
not U_inv2997 ( n1310_r, n1310 );
dff a10_k3a_reg_11_ ( clk, n1309_r, a10_k3a[11], a10_v3[11] );
not U_inv2998 ( n1309_r, n1309 );
dff a10_k3a_reg_12_ ( clk, n1309_r, a10_k3a[12], a10_v3[12] );
not U_inv2999 ( n1309_r, n1309 );
dff a10_k3a_reg_13_ ( clk, n1309_r, a10_k3a[13], a10_v3[13] );
not U_inv3000 ( n1309_r, n1309 );
dff a10_k3a_reg_14_ ( clk, n1309_r, a10_k3a[14], a10_v3[14] );
not U_inv3001 ( n1309_r, n1309 );
dff a10_k3a_reg_15_ ( clk, n1309_r, a10_k3a[15], a10_v3[15] );
not U_inv3002 ( n1309_r, n1309 );
dff a10_k3a_reg_16_ ( clk, n1309_r, a10_k3a[16], a10_v3[16] );
not U_inv3003 ( n1309_r, n1309 );
dff a10_k3a_reg_17_ ( clk, n1309_r, a10_k3a[17], a10_v3[17] );
not U_inv3004 ( n1309_r, n1309 );
dff a10_k3a_reg_18_ ( clk, n1309_r, a10_k3a[18], a10_v3[18] );
not U_inv3005 ( n1309_r, n1309 );
dff a10_k3a_reg_19_ ( clk, n1309_r, a10_k3a[19], a10_v3[19] );
not U_inv3006 ( n1309_r, n1309 );
dff a10_k3a_reg_20_ ( clk, n1309_r, a10_k3a[20], a10_v3[20] );
not U_inv3007 ( n1309_r, n1309 );
dff a10_k3a_reg_21_ ( clk, n1309_r, a10_k3a[21], a10_v3[21] );
not U_inv3008 ( n1309_r, n1309 );
dff a10_k3a_reg_22_ ( clk, n1309_r, a10_k3a[22], a10_v3[22] );
not U_inv3009 ( n1309_r, n1309 );
dff a10_k3a_reg_23_ ( clk, n1308_r, a10_k3a[23], a10_v3[23] );
not U_inv3010 ( n1308_r, n1308 );
dff a10_k3a_reg_24_ ( clk, n1308_r, a10_k3a[24], a10_v3[24] );
not U_inv3011 ( n1308_r, n1308 );
dff a10_k3a_reg_25_ ( clk, n1308_r, a10_k3a[25], a10_v3[25] );
not U_inv3012 ( n1308_r, n1308 );
dff a10_k3a_reg_26_ ( clk, n1308_r, a10_k3a[26], a10_v3[26] );
not U_inv3013 ( n1308_r, n1308 );
dff a10_k3a_reg_27_ ( clk, n1308_r, a10_k3a[27], a10_v3[27] );
not U_inv3014 ( n1308_r, n1308 );
dff a10_k3a_reg_28_ ( clk, n1308_r, a10_k3a[28], a10_v3[28] );
not U_inv3015 ( n1308_r, n1308 );
dff a10_k3a_reg_29_ ( clk, n1308_r, a10_k3a[29], a10_v3[29] );
not U_inv3016 ( n1308_r, n1308 );
dff a10_k3a_reg_30_ ( clk, n1308_r, a10_k3a[30], a10_v3[30] );
not U_inv3017 ( n1308_r, n1308 );
dff a10_k3a_reg_31_ ( clk, n1308_r, a10_k3a[31], a10_v3[31] );
not U_inv3018 ( n1308_r, n1308 );
dff a10_k2a_reg_0_ ( clk, n1308_r, a10_k2a[0], a10_v2[0] );
not U_inv3019 ( n1308_r, n1308 );
dff a10_k2a_reg_1_ ( clk, n1308_r, a10_k2a[1], a10_v2[1] );
not U_inv3020 ( n1308_r, n1308 );
dff a10_k2a_reg_2_ ( clk, n1308_r, a10_k2a[2], a10_v2[2] );
not U_inv3021 ( n1308_r, n1308 );
dff a10_k2a_reg_3_ ( clk, n1307_r, a10_k2a[3], a10_v2[3] );
not U_inv3022 ( n1307_r, n1307 );
dff a10_k2a_reg_4_ ( clk, n1307_r, a10_k2a[4], a10_v2[4] );
not U_inv3023 ( n1307_r, n1307 );
dff a10_k2a_reg_5_ ( clk, n1307_r, a10_k2a[5], a10_v2[5] );
not U_inv3024 ( n1307_r, n1307 );
dff a10_k2a_reg_6_ ( clk, n1307_r, a10_k2a[6], a10_v2[6] );
not U_inv3025 ( n1307_r, n1307 );
dff a10_k2a_reg_7_ ( clk, n1307_r, a10_k2a[7], a10_v2[7] );
not U_inv3026 ( n1307_r, n1307 );
dff a10_k2a_reg_8_ ( clk, n1307_r, a10_k2a[8], a10_v2[8] );
not U_inv3027 ( n1307_r, n1307 );
dff a10_k2a_reg_9_ ( clk, n1307_r, a10_k2a[9], a10_v2[9] );
not U_inv3028 ( n1307_r, n1307 );
dff a10_k2a_reg_10_ ( clk, n1307_r, a10_k2a[10], a10_v2[10] );
not U_inv3029 ( n1307_r, n1307 );
dff a10_k2a_reg_11_ ( clk, n1307_r, a10_k2a[11], a10_v2[11] );
not U_inv3030 ( n1307_r, n1307 );
dff a10_k2a_reg_12_ ( clk, n1307_r, a10_k2a[12], a10_v2[12] );
not U_inv3031 ( n1307_r, n1307 );
dff a10_k2a_reg_13_ ( clk, n1307_r, a10_k2a[13], a10_v2[13] );
not U_inv3032 ( n1307_r, n1307 );
dff a10_k2a_reg_14_ ( clk, n1307_r, a10_k2a[14], a10_v2[14] );
not U_inv3033 ( n1307_r, n1307 );
dff a10_k2a_reg_15_ ( clk, n1306_r, a10_k2a[15], a10_v2[15] );
not U_inv3034 ( n1306_r, n1306 );
dff a10_k2a_reg_16_ ( clk, n1306_r, a10_k2a[16], a10_v2[16] );
not U_inv3035 ( n1306_r, n1306 );
dff a10_k2a_reg_17_ ( clk, n1306_r, a10_k2a[17], a10_v2[17] );
not U_inv3036 ( n1306_r, n1306 );
dff a10_k2a_reg_18_ ( clk, n1306_r, a10_k2a[18], a10_v2[18] );
not U_inv3037 ( n1306_r, n1306 );
dff a10_k2a_reg_19_ ( clk, n1306_r, a10_k2a[19], a10_v2[19] );
not U_inv3038 ( n1306_r, n1306 );
dff a10_k2a_reg_20_ ( clk, n1306_r, a10_k2a[20], a10_v2[20] );
not U_inv3039 ( n1306_r, n1306 );
dff a10_k2a_reg_21_ ( clk, n1306_r, a10_k2a[21], a10_v2[21] );
not U_inv3040 ( n1306_r, n1306 );
dff a10_k2a_reg_22_ ( clk, n1306_r, a10_k2a[22], a10_v2[22] );
not U_inv3041 ( n1306_r, n1306 );
dff a10_k2a_reg_23_ ( clk, n1306_r, a10_k2a[23], a10_v2[23] );
not U_inv3042 ( n1306_r, n1306 );
dff a10_k2a_reg_24_ ( clk, n1306_r, a10_k2a[24], a10_v2[24] );
not U_inv3043 ( n1306_r, n1306 );
dff a10_k2a_reg_25_ ( clk, n1306_r, a10_k2a[25], a10_v2[25] );
not U_inv3044 ( n1306_r, n1306 );
dff a10_k2a_reg_26_ ( clk, n1306_r, a10_k2a[26], a10_v2[26] );
not U_inv3045 ( n1306_r, n1306 );
dff a10_k2a_reg_27_ ( clk, n1305_r, a10_k2a[27], a10_v2[27] );
not U_inv3046 ( n1305_r, n1305 );
dff a10_k2a_reg_28_ ( clk, n1305_r, a10_k2a[28], a10_v2[28] );
not U_inv3047 ( n1305_r, n1305 );
dff a10_k2a_reg_29_ ( clk, n1305_r, a10_k2a[29], a10_v2[29] );
not U_inv3048 ( n1305_r, n1305 );
dff a10_k2a_reg_30_ ( clk, n1305_r, a10_k2a[30], a10_v2[30] );
not U_inv3049 ( n1305_r, n1305 );
dff a10_k2a_reg_31_ ( clk, n1305_r, a10_k2a[31], a10_v2[31] );
not U_inv3050 ( n1305_r, n1305 );
dff a10_k1a_reg_0_ ( clk, n1305_r, a10_k1a[0], a10_v1[0] );
not U_inv3051 ( n1305_r, n1305 );
dff a10_k1a_reg_1_ ( clk, n1305_r, a10_k1a[1], a10_v1[1] );
not U_inv3052 ( n1305_r, n1305 );
dff a10_k1a_reg_2_ ( clk, n1305_r, a10_k1a[2], a10_v1[2] );
not U_inv3053 ( n1305_r, n1305 );
dff a10_k1a_reg_3_ ( clk, n1305_r, a10_k1a[3], a10_v1[3] );
not U_inv3054 ( n1305_r, n1305 );
dff a10_k1a_reg_4_ ( clk, n1305_r, a10_k1a[4], a10_v1[4] );
not U_inv3055 ( n1305_r, n1305 );
dff a10_k1a_reg_5_ ( clk, n1305_r, a10_k1a[5], a10_v1[5] );
not U_inv3056 ( n1305_r, n1305 );
dff a10_k1a_reg_6_ ( clk, n1305_r, a10_k1a[6], a10_v1[6] );
not U_inv3057 ( n1305_r, n1305 );
dff a10_k1a_reg_7_ ( clk, n1304_r, a10_k1a[7], a10_v1[7] );
not U_inv3058 ( n1304_r, n1304 );
dff a10_k1a_reg_8_ ( clk, n1304_r, a10_k1a[8], a10_v1[8] );
not U_inv3059 ( n1304_r, n1304 );
dff a10_k1a_reg_9_ ( clk, n1304_r, a10_k1a[9], a10_v1[9] );
not U_inv3060 ( n1304_r, n1304 );
dff a10_k1a_reg_10_ ( clk, n1304_r, a10_k1a[10], a10_v1[10] );
not U_inv3061 ( n1304_r, n1304 );
dff a10_k1a_reg_11_ ( clk, n1304_r, a10_k1a[11], a10_v1[11] );
not U_inv3062 ( n1304_r, n1304 );
dff a10_k1a_reg_12_ ( clk, n1304_r, a10_k1a[12], a10_v1[12] );
not U_inv3063 ( n1304_r, n1304 );
dff a10_k1a_reg_13_ ( clk, n1304_r, a10_k1a[13], a10_v1[13] );
not U_inv3064 ( n1304_r, n1304 );
dff a10_k1a_reg_14_ ( clk, n1304_r, a10_k1a[14], a10_v1[14] );
not U_inv3065 ( n1304_r, n1304 );
dff a10_k1a_reg_15_ ( clk, n1304_r, a10_k1a[15], a10_v1[15] );
not U_inv3066 ( n1304_r, n1304 );
dff a10_k1a_reg_16_ ( clk, n1304_r, a10_k1a[16], a10_v1[16] );
not U_inv3067 ( n1304_r, n1304 );
dff a10_k1a_reg_17_ ( clk, n1304_r, a10_k1a[17], a10_v1[17] );
not U_inv3068 ( n1304_r, n1304 );
dff a10_k1a_reg_18_ ( clk, n1304_r, a10_k1a[18], a10_v1[18] );
not U_inv3069 ( n1304_r, n1304 );
dff a10_k1a_reg_19_ ( clk, n1303_r, a10_k1a[19], a10_v1[19] );
not U_inv3070 ( n1303_r, n1303 );
dff a10_k1a_reg_20_ ( clk, n1303_r, a10_k1a[20], a10_v1[20] );
not U_inv3071 ( n1303_r, n1303 );
dff a10_k1a_reg_21_ ( clk, n1303_r, a10_k1a[21], a10_v1[21] );
not U_inv3072 ( n1303_r, n1303 );
dff a10_k1a_reg_22_ ( clk, n1303_r, a10_k1a[22], a10_v1[22] );
not U_inv3073 ( n1303_r, n1303 );
dff a10_k1a_reg_23_ ( clk, n1303_r, a10_k1a[23], a10_v1[23] );
not U_inv3074 ( n1303_r, n1303 );
dff a10_k1a_reg_24_ ( clk, n1303_r, a10_k1a[24], a10_v1[24] );
not U_inv3075 ( n1303_r, n1303 );
dff a10_k1a_reg_25_ ( clk, n1303_r, a10_k1a[25], a10_v1[25] );
not U_inv3076 ( n1303_r, n1303 );
dff a10_k1a_reg_26_ ( clk, n1303_r, a10_k1a[26], a10_v1[26] );
not U_inv3077 ( n1303_r, n1303 );
dff a10_k1a_reg_27_ ( clk, n1303_r, a10_k1a[27], a10_v1[27] );
not U_inv3078 ( n1303_r, n1303 );
dff a10_k1a_reg_28_ ( clk, n1303_r, a10_k1a[28], a10_v1[28] );
not U_inv3079 ( n1303_r, n1303 );
dff a10_k1a_reg_29_ ( clk, n1303_r, a10_k1a[29], a10_v1[29] );
not U_inv3080 ( n1303_r, n1303 );
dff a10_k1a_reg_30_ ( clk, n1303_r, a10_k1a[30], a10_v1[30] );
not U_inv3081 ( n1303_r, n1303 );
one_round r1 ( .p1(clk), .p2(reset), .p3(s0), .p4(k0b), .p5({s1_127_, s1_126_,
s1_125_, s1_124_, s1_123_, s1_122_, s1_121_, s1_120_, s1_119_, s1_118_,
s1_117_, s1_116_, s1_115_, s1_114_, s1_113_, s1_112_, s1_111_, s1_110_,
s1_109_, s1_108_, s1_107_, s1_106_, s1_105_, s1_104_, s1_103_, s1_102_,
s1_101_, s1_100_, s1_99_, s1_98_, s1_97_, s1_96_, s1_95_, s1_94_,
s1_93_, s1_92_, s1_91_, s1_90_, s1_89_, s1_88_, s1_87_, s1_86_, s1_85_,
s1_84_, s1_83_, s1_82_, s1_81_, s1_80_, s1_79_, s1_78_, s1_77_, s1_76_,
s1_75_, s1_74_, s1_73_, s1_72_, s1_71_, s1_70_, s1_69_, s1_68_, s1_67_,
s1_66_, s1_65_, s1_64_, s1_63_, s1_62_, s1_61_, s1_60_, s1_59_, s1_58_,
s1_57_, s1_56_, s1_55_, s1_54_, s1_53_, s1_52_, s1_51_, s1_50_, s1_49_,
s1_48_, s1_47_, s1_46_, s1_45_, s1_44_, s1_43_, s1_42_, s1_41_, s1_40_,
s1_39_, s1_38_, s1_37_, s1_36_, s1_35_, s1_34_, s1_33_, s1_32_, s1_31_,
s1_30_, s1_29_, s1_28_, s1_27_, s1_26_, s1_25_, s1_24_, s1_23_, s1_22_,
s1_21_, s1_20_, s1_19_, s1_18_, s1_17_, s1_16_, s1_15_, s1_14_, s1_13_,
s1_12_, s1_11_, s1_10_, s1_9_, s1_8_, s1_7_, s1_6_, s1_5_, s1_4_,
s1_3_, s1_2_, s1_1_, s1_0_}) );
one_round r2 ( .p1(clk), .p2(reset), .p3({s1_127_, s1_126_, s1_125_, s1_124_,
s1_123_, s1_122_, s1_121_, s1_120_, s1_119_, s1_118_, s1_117_, s1_116_,
s1_115_, s1_114_, s1_113_, s1_112_, s1_111_, s1_110_, s1_109_, s1_108_,
s1_107_, s1_106_, s1_105_, s1_104_, s1_103_, s1_102_, s1_101_, s1_100_,
s1_99_, s1_98_, s1_97_, s1_96_, s1_95_, s1_94_, s1_93_, s1_92_, s1_91_,
s1_90_, s1_89_, s1_88_, s1_87_, s1_86_, s1_85_, s1_84_, s1_83_, s1_82_,
s1_81_, s1_80_, s1_79_, s1_78_, s1_77_, s1_76_, s1_75_, s1_74_, s1_73_,
s1_72_, s1_71_, s1_70_, s1_69_, s1_68_, s1_67_, s1_66_, s1_65_, s1_64_,
s1_63_, s1_62_, s1_61_, s1_60_, s1_59_, s1_58_, s1_57_, s1_56_, s1_55_,
s1_54_, s1_53_, s1_52_, s1_51_, s1_50_, s1_49_, s1_48_, s1_47_, s1_46_,
s1_45_, s1_44_, s1_43_, s1_42_, s1_41_, s1_40_, s1_39_, s1_38_, s1_37_,
s1_36_, s1_35_, s1_34_, s1_33_, s1_32_, s1_31_, s1_30_, s1_29_, s1_28_,
s1_27_, s1_26_, s1_25_, s1_24_, s1_23_, s1_22_, s1_21_, s1_20_, s1_19_,
s1_18_, s1_17_, s1_16_, s1_15_, s1_14_, s1_13_, s1_12_, s1_11_, s1_10_,
s1_9_, s1_8_, s1_7_, s1_6_, s1_5_, s1_4_, s1_3_, s1_2_, s1_1_, s1_0_}),
.p4(k1b), .p5({s2_127_, s2_126_, s2_125_, s2_124_, s2_123_, s2_122_,
s2_121_, s2_120_, s2_119_, s2_118_, s2_117_, s2_116_, s2_115_, s2_114_,
s2_113_, s2_112_, s2_111_, s2_110_, s2_109_, s2_108_, s2_107_, s2_106_,
s2_105_, s2_104_, s2_103_, s2_102_, s2_101_, s2_100_, s2_99_, s2_98_,
s2_97_, s2_96_, s2_95_, s2_94_, s2_93_, s2_92_, s2_91_, s2_90_, s2_89_,
s2_88_, s2_87_, s2_86_, s2_85_, s2_84_, s2_83_, s2_82_, s2_81_, s2_80_,
s2_79_, s2_78_, s2_77_, s2_76_, s2_75_, s2_74_, s2_73_, s2_72_, s2_71_,
s2_70_, s2_69_, s2_68_, s2_67_, s2_66_, s2_65_, s2_64_, s2_63_, s2_62_,
s2_61_, s2_60_, s2_59_, s2_58_, s2_57_, s2_56_, s2_55_, s2_54_, s2_53_,
s2_52_, s2_51_, s2_50_, s2_49_, s2_48_, s2_47_, s2_46_, s2_45_, s2_44_,
s2_43_, s2_42_, s2_41_, s2_40_, s2_39_, s2_38_, s2_37_, s2_36_, s2_35_,
s2_34_, s2_33_, s2_32_, s2_31_, s2_30_, s2_29_, s2_28_, s2_27_, s2_26_,
s2_25_, s2_24_, s2_23_, s2_22_, s2_21_, s2_20_, s2_19_, s2_18_, s2_17_,
s2_16_, s2_15_, s2_14_, s2_13_, s2_12_, s2_11_, s2_10_, s2_9_, s2_8_,
s2_7_, s2_6_, s2_5_, s2_4_, s2_3_, s2_2_, s2_1_, s2_0_}) );
one_round r3 ( .p1(clk), .p2(reset), .p3({s2_127_, s2_126_, s2_125_, s2_124_,
s2_123_, s2_122_, s2_121_, s2_120_, s2_119_, s2_118_, s2_117_, s2_116_,
s2_115_, s2_114_, s2_113_, s2_112_, s2_111_, s2_110_, s2_109_, s2_108_,
s2_107_, s2_106_, s2_105_, s2_104_, s2_103_, s2_102_, s2_101_, s2_100_,
s2_99_, s2_98_, s2_97_, s2_96_, s2_95_, s2_94_, s2_93_, s2_92_, s2_91_,
s2_90_, s2_89_, s2_88_, s2_87_, s2_86_, s2_85_, s2_84_, s2_83_, s2_82_,
s2_81_, s2_80_, s2_79_, s2_78_, s2_77_, s2_76_, s2_75_, s2_74_, s2_73_,
s2_72_, s2_71_, s2_70_, s2_69_, s2_68_, s2_67_, s2_66_, s2_65_, s2_64_,
s2_63_, s2_62_, s2_61_, s2_60_, s2_59_, s2_58_, s2_57_, s2_56_, s2_55_,
s2_54_, s2_53_, s2_52_, s2_51_, s2_50_, s2_49_, s2_48_, s2_47_, s2_46_,
s2_45_, s2_44_, s2_43_, s2_42_, s2_41_, s2_40_, s2_39_, s2_38_, s2_37_,
s2_36_, s2_35_, s2_34_, s2_33_, s2_32_, s2_31_, s2_30_, s2_29_, s2_28_,
s2_27_, s2_26_, s2_25_, s2_24_, s2_23_, s2_22_, s2_21_, s2_20_, s2_19_,
s2_18_, s2_17_, s2_16_, s2_15_, s2_14_, s2_13_, s2_12_, s2_11_, s2_10_,
s2_9_, s2_8_, s2_7_, s2_6_, s2_5_, s2_4_, s2_3_, s2_2_, s2_1_, s2_0_}),
.p4(k2b), .p5({s3_127_, s3_126_, s3_125_, s3_124_, s3_123_, s3_122_,
s3_121_, s3_120_, s3_119_, s3_118_, s3_117_, s3_116_, s3_115_, s3_114_,
s3_113_, s3_112_, s3_111_, s3_110_, s3_109_, s3_108_, s3_107_, s3_106_,
s3_105_, s3_104_, s3_103_, s3_102_, s3_101_, s3_100_, s3_99_, s3_98_,
s3_97_, s3_96_, s3_95_, s3_94_, s3_93_, s3_92_, s3_91_, s3_90_, s3_89_,
s3_88_, s3_87_, s3_86_, s3_85_, s3_84_, s3_83_, s3_82_, s3_81_, s3_80_,
s3_79_, s3_78_, s3_77_, s3_76_, s3_75_, s3_74_, s3_73_, s3_72_, s3_71_,
s3_70_, s3_69_, s3_68_, s3_67_, s3_66_, s3_65_, s3_64_, s3_63_, s3_62_,
s3_61_, s3_60_, s3_59_, s3_58_, s3_57_, s3_56_, s3_55_, s3_54_, s3_53_,
s3_52_, s3_51_, s3_50_, s3_49_, s3_48_, s3_47_, s3_46_, s3_45_, s3_44_,
s3_43_, s3_42_, s3_41_, s3_40_, s3_39_, s3_38_, s3_37_, s3_36_, s3_35_,
s3_34_, s3_33_, s3_32_, s3_31_, s3_30_, s3_29_, s3_28_, s3_27_, s3_26_,
s3_25_, s3_24_, s3_23_, s3_22_, s3_21_, s3_20_, s3_19_, s3_18_, s3_17_,
s3_16_, s3_15_, s3_14_, s3_13_, s3_12_, s3_11_, s3_10_, s3_9_, s3_8_,
s3_7_, s3_6_, s3_5_, s3_4_, s3_3_, s3_2_, s3_1_, s3_0_}) );
one_round r4 ( .p1(clk), .p2(reset), .p3({s3_127_, s3_126_, s3_125_, s3_124_,
s3_123_, s3_122_, s3_121_, s3_120_, s3_119_, s3_118_, s3_117_, s3_116_,
s3_115_, s3_114_, s3_113_, s3_112_, s3_111_, s3_110_, s3_109_, s3_108_,
s3_107_, s3_106_, s3_105_, s3_104_, s3_103_, s3_102_, s3_101_, s3_100_,
s3_99_, s3_98_, s3_97_, s3_96_, s3_95_, s3_94_, s3_93_, s3_92_, s3_91_,
s3_90_, s3_89_, s3_88_, s3_87_, s3_86_, s3_85_, s3_84_, s3_83_, s3_82_,
s3_81_, s3_80_, s3_79_, s3_78_, s3_77_, s3_76_, s3_75_, s3_74_, s3_73_,
s3_72_, s3_71_, s3_70_, s3_69_, s3_68_, s3_67_, s3_66_, s3_65_, s3_64_,
s3_63_, s3_62_, s3_61_, s3_60_, s3_59_, s3_58_, s3_57_, s3_56_, s3_55_,
s3_54_, s3_53_, s3_52_, s3_51_, s3_50_, s3_49_, s3_48_, s3_47_, s3_46_,
s3_45_, s3_44_, s3_43_, s3_42_, s3_41_, s3_40_, s3_39_, s3_38_, s3_37_,
s3_36_, s3_35_, s3_34_, s3_33_, s3_32_, s3_31_, s3_30_, s3_29_, s3_28_,
s3_27_, s3_26_, s3_25_, s3_24_, s3_23_, s3_22_, s3_21_, s3_20_, s3_19_,
s3_18_, s3_17_, s3_16_, s3_15_, s3_14_, s3_13_, s3_12_, s3_11_, s3_10_,
s3_9_, s3_8_, s3_7_, s3_6_, s3_5_, s3_4_, s3_3_, s3_2_, s3_1_, s3_0_}),
.p4(k3b), .p5({s4_127_, s4_126_, s4_125_, s4_124_, s4_123_, s4_122_,
s4_121_, s4_120_, s4_119_, s4_118_, s4_117_, s4_116_, s4_115_, s4_114_,
s4_113_, s4_112_, s4_111_, s4_110_, s4_109_, s4_108_, s4_107_, s4_106_,
s4_105_, s4_104_, s4_103_, s4_102_, s4_101_, s4_100_, s4_99_, s4_98_,
s4_97_, s4_96_, s4_95_, s4_94_, s4_93_, s4_92_, s4_91_, s4_90_, s4_89_,
s4_88_, s4_87_, s4_86_, s4_85_, s4_84_, s4_83_, s4_82_, s4_81_, s4_80_,
s4_79_, s4_78_, s4_77_, s4_76_, s4_75_, s4_74_, s4_73_, s4_72_, s4_71_,
s4_70_, s4_69_, s4_68_, s4_67_, s4_66_, s4_65_, s4_64_, s4_63_, s4_62_,
s4_61_, s4_60_, s4_59_, s4_58_, s4_57_, s4_56_, s4_55_, s4_54_, s4_53_,
s4_52_, s4_51_, s4_50_, s4_49_, s4_48_, s4_47_, s4_46_, s4_45_, s4_44_,
s4_43_, s4_42_, s4_41_, s4_40_, s4_39_, s4_38_, s4_37_, s4_36_, s4_35_,
s4_34_, s4_33_, s4_32_, s4_31_, s4_30_, s4_29_, s4_28_, s4_27_, s4_26_,
s4_25_, s4_24_, s4_23_, s4_22_, s4_21_, s4_20_, s4_19_, s4_18_, s4_17_,
s4_16_, s4_15_, s4_14_, s4_13_, s4_12_, s4_11_, s4_10_, s4_9_, s4_8_,
s4_7_, s4_6_, s4_5_, s4_4_, s4_3_, s4_2_, s4_1_, s4_0_}) );
one_round r5 ( .p1(clk), .p2(reset), .p3({s4_127_, s4_126_, s4_125_, s4_124_,
s4_123_, s4_122_, s4_121_, s4_120_, s4_119_, s4_118_, s4_117_, s4_116_,
s4_115_, s4_114_, s4_113_, s4_112_, s4_111_, s4_110_, s4_109_, s4_108_,
s4_107_, s4_106_, s4_105_, s4_104_, s4_103_, s4_102_, s4_101_, s4_100_,
s4_99_, s4_98_, s4_97_, s4_96_, s4_95_, s4_94_, s4_93_, s4_92_, s4_91_,
s4_90_, s4_89_, s4_88_, s4_87_, s4_86_, s4_85_, s4_84_, s4_83_, s4_82_,
s4_81_, s4_80_, s4_79_, s4_78_, s4_77_, s4_76_, s4_75_, s4_74_, s4_73_,
s4_72_, s4_71_, s4_70_, s4_69_, s4_68_, s4_67_, s4_66_, s4_65_, s4_64_,
s4_63_, s4_62_, s4_61_, s4_60_, s4_59_, s4_58_, s4_57_, s4_56_, s4_55_,
s4_54_, s4_53_, s4_52_, s4_51_, s4_50_, s4_49_, s4_48_, s4_47_, s4_46_,
s4_45_, s4_44_, s4_43_, s4_42_, s4_41_, s4_40_, s4_39_, s4_38_, s4_37_,
s4_36_, s4_35_, s4_34_, s4_33_, s4_32_, s4_31_, s4_30_, s4_29_, s4_28_,
s4_27_, s4_26_, s4_25_, s4_24_, s4_23_, s4_22_, s4_21_, s4_20_, s4_19_,
s4_18_, s4_17_, s4_16_, s4_15_, s4_14_, s4_13_, s4_12_, s4_11_, s4_10_,
s4_9_, s4_8_, s4_7_, s4_6_, s4_5_, s4_4_, s4_3_, s4_2_, s4_1_, s4_0_}),
.p4(k4b), .p5({s5_127_, s5_126_, s5_125_, s5_124_, s5_123_, s5_122_,
s5_121_, s5_120_, s5_119_, s5_118_, s5_117_, s5_116_, s5_115_, s5_114_,
s5_113_, s5_112_, s5_111_, s5_110_, s5_109_, s5_108_, s5_107_, s5_106_,
s5_105_, s5_104_, s5_103_, s5_102_, s5_101_, s5_100_, s5_99_, s5_98_,
s5_97_, s5_96_, s5_95_, s5_94_, s5_93_, s5_92_, s5_91_, s5_90_, s5_89_,
s5_88_, s5_87_, s5_86_, s5_85_, s5_84_, s5_83_, s5_82_, s5_81_, s5_80_,
s5_79_, s5_78_, s5_77_, s5_76_, s5_75_, s5_74_, s5_73_, s5_72_, s5_71_,
s5_70_, s5_69_, s5_68_, s5_67_, s5_66_, s5_65_, s5_64_, s5_63_, s5_62_,
s5_61_, s5_60_, s5_59_, s5_58_, s5_57_, s5_56_, s5_55_, s5_54_, s5_53_,
s5_52_, s5_51_, s5_50_, s5_49_, s5_48_, s5_47_, s5_46_, s5_45_, s5_44_,
s5_43_, s5_42_, s5_41_, s5_40_, s5_39_, s5_38_, s5_37_, s5_36_, s5_35_,
s5_34_, s5_33_, s5_32_, s5_31_, s5_30_, s5_29_, s5_28_, s5_27_, s5_26_,
s5_25_, s5_24_, s5_23_, s5_22_, s5_21_, s5_20_, s5_19_, s5_18_, s5_17_,
s5_16_, s5_15_, s5_14_, s5_13_, s5_12_, s5_11_, s5_10_, s5_9_, s5_8_,
s5_7_, s5_6_, s5_5_, s5_4_, s5_3_, s5_2_, s5_1_, s5_0_}) );
one_round r6 ( .p1(clk), .p2(reset), .p3({s5_127_, s5_126_, s5_125_, s5_124_,
s5_123_, s5_122_, s5_121_, s5_120_, s5_119_, s5_118_, s5_117_, s5_116_,
s5_115_, s5_114_, s5_113_, s5_112_, s5_111_, s5_110_, s5_109_, s5_108_,
s5_107_, s5_106_, s5_105_, s5_104_, s5_103_, s5_102_, s5_101_, s5_100_,
s5_99_, s5_98_, s5_97_, s5_96_, s5_95_, s5_94_, s5_93_, s5_92_, s5_91_,
s5_90_, s5_89_, s5_88_, s5_87_, s5_86_, s5_85_, s5_84_, s5_83_, s5_82_,
s5_81_, s5_80_, s5_79_, s5_78_, s5_77_, s5_76_, s5_75_, s5_74_, s5_73_,
s5_72_, s5_71_, s5_70_, s5_69_, s5_68_, s5_67_, s5_66_, s5_65_, s5_64_,
s5_63_, s5_62_, s5_61_, s5_60_, s5_59_, s5_58_, s5_57_, s5_56_, s5_55_,
s5_54_, s5_53_, s5_52_, s5_51_, s5_50_, s5_49_, s5_48_, s5_47_, s5_46_,
s5_45_, s5_44_, s5_43_, s5_42_, s5_41_, s5_40_, s5_39_, s5_38_, s5_37_,
s5_36_, s5_35_, s5_34_, s5_33_, s5_32_, s5_31_, s5_30_, s5_29_, s5_28_,
s5_27_, s5_26_, s5_25_, s5_24_, s5_23_, s5_22_, s5_21_, s5_20_, s5_19_,
s5_18_, s5_17_, s5_16_, s5_15_, s5_14_, s5_13_, s5_12_, s5_11_, s5_10_,
s5_9_, s5_8_, s5_7_, s5_6_, s5_5_, s5_4_, s5_3_, s5_2_, s5_1_, s5_0_}),
.p4(k5b), .p5({s6_127_, s6_126_, s6_125_, s6_124_, s6_123_, s6_122_,
s6_121_, s6_120_, s6_119_, s6_118_, s6_117_, s6_116_, s6_115_, s6_114_,
s6_113_, s6_112_, s6_111_, s6_110_, s6_109_, s6_108_, s6_107_, s6_106_,
s6_105_, s6_104_, s6_103_, s6_102_, s6_101_, s6_100_, s6_99_, s6_98_,
s6_97_, s6_96_, s6_95_, s6_94_, s6_93_, s6_92_, s6_91_, s6_90_, s6_89_,
s6_88_, s6_87_, s6_86_, s6_85_, s6_84_, s6_83_, s6_82_, s6_81_, s6_80_,
s6_79_, s6_78_, s6_77_, s6_76_, s6_75_, s6_74_, s6_73_, s6_72_, s6_71_,
s6_70_, s6_69_, s6_68_, s6_67_, s6_66_, s6_65_, s6_64_, s6_63_, s6_62_,
s6_61_, s6_60_, s6_59_, s6_58_, s6_57_, s6_56_, s6_55_, s6_54_, s6_53_,
s6_52_, s6_51_, s6_50_, s6_49_, s6_48_, s6_47_, s6_46_, s6_45_, s6_44_,
s6_43_, s6_42_, s6_41_, s6_40_, s6_39_, s6_38_, s6_37_, s6_36_, s6_35_,
s6_34_, s6_33_, s6_32_, s6_31_, s6_30_, s6_29_, s6_28_, s6_27_, s6_26_,
s6_25_, s6_24_, s6_23_, s6_22_, s6_21_, s6_20_, s6_19_, s6_18_, s6_17_,
s6_16_, s6_15_, s6_14_, s6_13_, s6_12_, s6_11_, s6_10_, s6_9_, s6_8_,
s6_7_, s6_6_, s6_5_, s6_4_, s6_3_, s6_2_, s6_1_, s6_0_}) );
one_round r7 ( .p1(clk), .p2(reset), .p3({s6_127_, s6_126_, s6_125_, s6_124_,
s6_123_, s6_122_, s6_121_, s6_120_, s6_119_, s6_118_, s6_117_, s6_116_,
s6_115_, s6_114_, s6_113_, s6_112_, s6_111_, s6_110_, s6_109_, s6_108_,
s6_107_, s6_106_, s6_105_, s6_104_, s6_103_, s6_102_, s6_101_, s6_100_,
s6_99_, s6_98_, s6_97_, s6_96_, s6_95_, s6_94_, s6_93_, s6_92_, s6_91_,
s6_90_, s6_89_, s6_88_, s6_87_, s6_86_, s6_85_, s6_84_, s6_83_, s6_82_,
s6_81_, s6_80_, s6_79_, s6_78_, s6_77_, s6_76_, s6_75_, s6_74_, s6_73_,
s6_72_, s6_71_, s6_70_, s6_69_, s6_68_, s6_67_, s6_66_, s6_65_, s6_64_,
s6_63_, s6_62_, s6_61_, s6_60_, s6_59_, s6_58_, s6_57_, s6_56_, s6_55_,
s6_54_, s6_53_, s6_52_, s6_51_, s6_50_, s6_49_, s6_48_, s6_47_, s6_46_,
s6_45_, s6_44_, s6_43_, s6_42_, s6_41_, s6_40_, s6_39_, s6_38_, s6_37_,
s6_36_, s6_35_, s6_34_, s6_33_, s6_32_, s6_31_, s6_30_, s6_29_, s6_28_,
s6_27_, s6_26_, s6_25_, s6_24_, s6_23_, s6_22_, s6_21_, s6_20_, s6_19_,
s6_18_, s6_17_, s6_16_, s6_15_, s6_14_, s6_13_, s6_12_, s6_11_, s6_10_,
s6_9_, s6_8_, s6_7_, s6_6_, s6_5_, s6_4_, s6_3_, s6_2_, s6_1_, s6_0_}),
.p4(k6b), .p5({s7_127_, s7_126_, s7_125_, s7_124_, s7_123_, s7_122_,
s7_121_, s7_120_, s7_119_, s7_118_, s7_117_, s7_116_, s7_115_, s7_114_,
s7_113_, s7_112_, s7_111_, s7_110_, s7_109_, s7_108_, s7_107_, s7_106_,
s7_105_, s7_104_, s7_103_, s7_102_, s7_101_, s7_100_, s7_99_, s7_98_,
s7_97_, s7_96_, s7_95_, s7_94_, s7_93_, s7_92_, s7_91_, s7_90_, s7_89_,
s7_88_, s7_87_, s7_86_, s7_85_, s7_84_, s7_83_, s7_82_, s7_81_, s7_80_,
s7_79_, s7_78_, s7_77_, s7_76_, s7_75_, s7_74_, s7_73_, s7_72_, s7_71_,
s7_70_, s7_69_, s7_68_, s7_67_, s7_66_, s7_65_, s7_64_, s7_63_, s7_62_,
s7_61_, s7_60_, s7_59_, s7_58_, s7_57_, s7_56_, s7_55_, s7_54_, s7_53_,
s7_52_, s7_51_, s7_50_, s7_49_, s7_48_, s7_47_, s7_46_, s7_45_, s7_44_,
s7_43_, s7_42_, s7_41_, s7_40_, s7_39_, s7_38_, s7_37_, s7_36_, s7_35_,
s7_34_, s7_33_, s7_32_, s7_31_, s7_30_, s7_29_, s7_28_, s7_27_, s7_26_,
s7_25_, s7_24_, s7_23_, s7_22_, s7_21_, s7_20_, s7_19_, s7_18_, s7_17_,
s7_16_, s7_15_, s7_14_, s7_13_, s7_12_, s7_11_, s7_10_, s7_9_, s7_8_,
s7_7_, s7_6_, s7_5_, s7_4_, s7_3_, s7_2_, s7_1_, s7_0_}) );
one_round r8 ( .p1(clk), .p2(reset), .p3({s7_127_, s7_126_, s7_125_, s7_124_,
s7_123_, s7_122_, s7_121_, s7_120_, s7_119_, s7_118_, s7_117_, s7_116_,
s7_115_, s7_114_, s7_113_, s7_112_, s7_111_, s7_110_, s7_109_, s7_108_,
s7_107_, s7_106_, s7_105_, s7_104_, s7_103_, s7_102_, s7_101_, s7_100_,
s7_99_, s7_98_, s7_97_, s7_96_, s7_95_, s7_94_, s7_93_, s7_92_, s7_91_,
s7_90_, s7_89_, s7_88_, s7_87_, s7_86_, s7_85_, s7_84_, s7_83_, s7_82_,
s7_81_, s7_80_, s7_79_, s7_78_, s7_77_, s7_76_, s7_75_, s7_74_, s7_73_,
s7_72_, s7_71_, s7_70_, s7_69_, s7_68_, s7_67_, s7_66_, s7_65_, s7_64_,
s7_63_, s7_62_, s7_61_, s7_60_, s7_59_, s7_58_, s7_57_, s7_56_, s7_55_,
s7_54_, s7_53_, s7_52_, s7_51_, s7_50_, s7_49_, s7_48_, s7_47_, s7_46_,
s7_45_, s7_44_, s7_43_, s7_42_, s7_41_, s7_40_, s7_39_, s7_38_, s7_37_,
s7_36_, s7_35_, s7_34_, s7_33_, s7_32_, s7_31_, s7_30_, s7_29_, s7_28_,
s7_27_, s7_26_, s7_25_, s7_24_, s7_23_, s7_22_, s7_21_, s7_20_, s7_19_,
s7_18_, s7_17_, s7_16_, s7_15_, s7_14_, s7_13_, s7_12_, s7_11_, s7_10_,
s7_9_, s7_8_, s7_7_, s7_6_, s7_5_, s7_4_, s7_3_, s7_2_, s7_1_, s7_0_}),
.p4(k7b), .p5({s8_127_, s8_126_, s8_125_, s8_124_, s8_123_, s8_122_,
s8_121_, s8_120_, s8_119_, s8_118_, s8_117_, s8_116_, s8_115_, s8_114_,
s8_113_, s8_112_, s8_111_, s8_110_, s8_109_, s8_108_, s8_107_, s8_106_,
s8_105_, s8_104_, s8_103_, s8_102_, s8_101_, s8_100_, s8_99_, s8_98_,
s8_97_, s8_96_, s8_95_, s8_94_, s8_93_, s8_92_, s8_91_, s8_90_, s8_89_,
s8_88_, s8_87_, s8_86_, s8_85_, s8_84_, s8_83_, s8_82_, s8_81_, s8_80_,
s8_79_, s8_78_, s8_77_, s8_76_, s8_75_, s8_74_, s8_73_, s8_72_, s8_71_,
s8_70_, s8_69_, s8_68_, s8_67_, s8_66_, s8_65_, s8_64_, s8_63_, s8_62_,
s8_61_, s8_60_, s8_59_, s8_58_, s8_57_, s8_56_, s8_55_, s8_54_, s8_53_,
s8_52_, s8_51_, s8_50_, s8_49_, s8_48_, s8_47_, s8_46_, s8_45_, s8_44_,
s8_43_, s8_42_, s8_41_, s8_40_, s8_39_, s8_38_, s8_37_, s8_36_, s8_35_,
s8_34_, s8_33_, s8_32_, s8_31_, s8_30_, s8_29_, s8_28_, s8_27_, s8_26_,
s8_25_, s8_24_, s8_23_, s8_22_, s8_21_, s8_20_, s8_19_, s8_18_, s8_17_,
s8_16_, s8_15_, s8_14_, s8_13_, s8_12_, s8_11_, s8_10_, s8_9_, s8_8_,
s8_7_, s8_6_, s8_5_, s8_4_, s8_3_, s8_2_, s8_1_, s8_0_}) );
one_round r9 ( .p1(clk), .p2(reset), .p3({s8_127_, s8_126_, s8_125_, s8_124_,
s8_123_, s8_122_, s8_121_, s8_120_, s8_119_, s8_118_, s8_117_, s8_116_,
s8_115_, s8_114_, s8_113_, s8_112_, s8_111_, s8_110_, s8_109_, s8_108_,
s8_107_, s8_106_, s8_105_, s8_104_, s8_103_, s8_102_, s8_101_, s8_100_,
s8_99_, s8_98_, s8_97_, s8_96_, s8_95_, s8_94_, s8_93_, s8_92_, s8_91_,
s8_90_, s8_89_, s8_88_, s8_87_, s8_86_, s8_85_, s8_84_, s8_83_, s8_82_,
s8_81_, s8_80_, s8_79_, s8_78_, s8_77_, s8_76_, s8_75_, s8_74_, s8_73_,
s8_72_, s8_71_, s8_70_, s8_69_, s8_68_, s8_67_, s8_66_, s8_65_, s8_64_,
s8_63_, s8_62_, s8_61_, s8_60_, s8_59_, s8_58_, s8_57_, s8_56_, s8_55_,
s8_54_, s8_53_, s8_52_, s8_51_, s8_50_, s8_49_, s8_48_, s8_47_, s8_46_,
s8_45_, s8_44_, s8_43_, s8_42_, s8_41_, s8_40_, s8_39_, s8_38_, s8_37_,
s8_36_, s8_35_, s8_34_, s8_33_, s8_32_, s8_31_, s8_30_, s8_29_, s8_28_,
s8_27_, s8_26_, s8_25_, s8_24_, s8_23_, s8_22_, s8_21_, s8_20_, s8_19_,
s8_18_, s8_17_, s8_16_, s8_15_, s8_14_, s8_13_, s8_12_, s8_11_, s8_10_,
s8_9_, s8_8_, s8_7_, s8_6_, s8_5_, s8_4_, s8_3_, s8_2_, s8_1_, s8_0_}),
.p4(k8b), .p5({s9_127_, s9_126_, s9_125_, s9_124_, s9_123_, s9_122_,
s9_121_, s9_120_, s9_119_, s9_118_, s9_117_, s9_116_, s9_115_, s9_114_,
s9_113_, s9_112_, s9_111_, s9_110_, s9_109_, s9_108_, s9_107_, s9_106_,
s9_105_, s9_104_, s9_103_, s9_102_, s9_101_, s9_100_, s9_99_, s9_98_,
s9_97_, s9_96_, s9_95_, s9_94_, s9_93_, s9_92_, s9_91_, s9_90_, s9_89_,
s9_88_, s9_87_, s9_86_, s9_85_, s9_84_, s9_83_, s9_82_, s9_81_, s9_80_,
s9_79_, s9_78_, s9_77_, s9_76_, s9_75_, s9_74_, s9_73_, s9_72_, s9_71_,
s9_70_, s9_69_, s9_68_, s9_67_, s9_66_, s9_65_, s9_64_, s9_63_, s9_62_,
s9_61_, s9_60_, s9_59_, s9_58_, s9_57_, s9_56_, s9_55_, s9_54_, s9_53_,
s9_52_, s9_51_, s9_50_, s9_49_, s9_48_, s9_47_, s9_46_, s9_45_, s9_44_,
s9_43_, s9_42_, s9_41_, s9_40_, s9_39_, s9_38_, s9_37_, s9_36_, s9_35_,
s9_34_, s9_33_, s9_32_, s9_31_, s9_30_, s9_29_, s9_28_, s9_27_, s9_26_,
s9_25_, s9_24_, s9_23_, s9_22_, s9_21_, s9_20_, s9_19_, s9_18_, s9_17_,
s9_16_, s9_15_, s9_14_, s9_13_, s9_12_, s9_11_, s9_10_, s9_9_, s9_8_,
s9_7_, s9_6_, s9_5_, s9_4_, s9_3_, s9_2_, s9_1_, s9_0_}) );
final_round rf ( .p1(clk), .p2(reset), .p3({s9_127_, s9_126_, s9_125_, s9_124_,
s9_123_, s9_122_, s9_121_, s9_120_, s9_119_, s9_118_, s9_117_, s9_116_,
s9_115_, s9_114_, s9_113_, s9_112_, s9_111_, s9_110_, s9_109_, s9_108_,
s9_107_, s9_106_, s9_105_, s9_104_, s9_103_, s9_102_, s9_101_, s9_100_,
s9_99_, s9_98_, s9_97_, s9_96_, s9_95_, s9_94_, s9_93_, s9_92_, s9_91_,
s9_90_, s9_89_, s9_88_, s9_87_, s9_86_, s9_85_, s9_84_, s9_83_, s9_82_,
s9_81_, s9_80_, s9_79_, s9_78_, s9_77_, s9_76_, s9_75_, s9_74_, s9_73_,
s9_72_, s9_71_, s9_70_, s9_69_, s9_68_, s9_67_, s9_66_, s9_65_, s9_64_,
s9_63_, s9_62_, s9_61_, s9_60_, s9_59_, s9_58_, s9_57_, s9_56_, s9_55_,
s9_54_, s9_53_, s9_52_, s9_51_, s9_50_, s9_49_, s9_48_, s9_47_, s9_46_,
s9_45_, s9_44_, s9_43_, s9_42_, s9_41_, s9_40_, s9_39_, s9_38_, s9_37_,
s9_36_, s9_35_, s9_34_, s9_33_, s9_32_, s9_31_, s9_30_, s9_29_, s9_28_,
s9_27_, s9_26_, s9_25_, s9_24_, s9_23_, s9_22_, s9_21_, s9_20_, s9_19_,
s9_18_, s9_17_, s9_16_, s9_15_, s9_14_, s9_13_, s9_12_, s9_11_, s9_10_,
s9_9_, s9_8_, s9_7_, s9_6_, s9_5_, s9_4_, s9_3_, s9_2_, s9_1_, s9_0_}),
.p4(k9b), .p5(out) );
S4 a1_S4_0 ( .p1(clk), .p2({k0[23:0], k0[31:24]}), .p3(a1_k4a) );
S4 a2_S4_0 ( .p1(clk), .p2({k1[23:0], k1[31:24]}), .p3(a2_k4a) );
S4 a3_S4_0 ( .p1(clk), .p2({k2[23:0], k2[31:24]}), .p3(a3_k4a) );
S4 a4_S4_0 ( .p1(clk), .p2({k3[23:0], k3[31:24]}), .p3(a4_k4a) );
S4 a5_S4_0 ( .p1(clk), .p2({k4[23:0], k4[31:24]}), .p3(a5_k4a) );
S4 a6_S4_0 ( .p1(clk), .p2({k5[23:0], k5[31:24]}), .p3(a6_k4a) );
S4 a7_S4_0 ( .p1(clk), .p2({k6[23:0], k6[31:24]}), .p3(a7_k4a) );
S4 a8_S4_0 ( .p1(clk), .p2({k7[23:0], k7[31:24]}), .p3(a8_k4a) );
S4 a9_S4_0 ( .p1(clk), .p2({k8[23:0], k8[31:24]}), .p3(a9_k4a) );
S4 a10_S4_0 ( .p1(clk), .p2({k9[23:0], k9[31:24]}), .p3(a10_k4a) );
xor a10_C865 ( k9b[127], a10_k0a[31], a10_k4a[31] );
xor a10_C866 ( k9b[126], a10_k0a[30], a10_k4a[30] );
xor a10_C867 ( k9b[125], a10_k0a[29], a10_k4a[29] );
xor a10_C868 ( k9b[124], a10_k0a[28], a10_k4a[28] );
xor a10_C869 ( k9b[123], a10_k0a[27], a10_k4a[27] );
xor a10_C870 ( k9b[122], a10_k0a[26], a10_k4a[26] );
xor a10_C871 ( k9b[121], a10_k0a[25], a10_k4a[25] );
xor a10_C872 ( k9b[120], a10_k0a[24], a10_k4a[24] );
xor a10_C873 ( k9b[119], a10_k0a[23], a10_k4a[23] );
xor a10_C874 ( k9b[118], a10_k0a[22], a10_k4a[22] );
xor a10_C875 ( k9b[117], a10_k0a[21], a10_k4a[21] );
xor a10_C876 ( k9b[116], a10_k0a[20], a10_k4a[20] );
xor a10_C877 ( k9b[115], a10_k0a[19], a10_k4a[19] );
xor a10_C878 ( k9b[114], a10_k0a[18], a10_k4a[18] );
xor a10_C879 ( k9b[113], a10_k0a[17], a10_k4a[17] );
xor a10_C880 ( k9b[112], a10_k0a[16], a10_k4a[16] );
xor a10_C881 ( k9b[111], a10_k0a[15], a10_k4a[15] );
xor a10_C882 ( k9b[110], a10_k0a[14], a10_k4a[14] );
xor a10_C883 ( k9b[109], a10_k0a[13], a10_k4a[13] );
xor a10_C884 ( k9b[108], a10_k0a[12], a10_k4a[12] );
xor a10_C885 ( k9b[107], a10_k0a[11], a10_k4a[11] );
xor a10_C886 ( k9b[106], a10_k0a[10], a10_k4a[10] );
xor a10_C887 ( k9b[105], a10_k0a[9], a10_k4a[9] );
xor a10_C888 ( k9b[104], a10_k0a[8], a10_k4a[8] );
xor a10_C889 ( k9b[103], a10_k0a[7], a10_k4a[7] );
xor a10_C890 ( k9b[102], a10_k0a[6], a10_k4a[6] );
xor a10_C891 ( k9b[101], a10_k0a[5], a10_k4a[5] );
xor a10_C892 ( k9b[100], a10_k0a[4], a10_k4a[4] );
xor a10_C893 ( k9b[99], a10_k0a[3], a10_k4a[3] );
xor a10_C894 ( k9b[98], a10_k0a[2], a10_k4a[2] );
xor a10_C895 ( k9b[97], a10_k0a[1], a10_k4a[1] );
xor a10_C896 ( k9b[96], a10_k0a[0], a10_k4a[0] );
xor a10_C897 ( k9b[95], a10_k1a[31], a10_k4a[31] );
xor a10_C898 ( k9b[94], a10_k1a[30], a10_k4a[30] );
xor a10_C899 ( k9b[93], a10_k1a[29], a10_k4a[29] );
xor a10_C900 ( k9b[92], a10_k1a[28], a10_k4a[28] );
xor a10_C901 ( k9b[91], a10_k1a[27], a10_k4a[27] );
xor a10_C902 ( k9b[90], a10_k1a[26], a10_k4a[26] );
xor a10_C903 ( k9b[89], a10_k1a[25], a10_k4a[25] );
xor a10_C904 ( k9b[88], a10_k1a[24], a10_k4a[24] );
xor a10_C905 ( k9b[87], a10_k1a[23], a10_k4a[23] );
xor a10_C906 ( k9b[86], a10_k1a[22], a10_k4a[22] );
xor a10_C907 ( k9b[85], a10_k1a[21], a10_k4a[21] );
xor a10_C908 ( k9b[84], a10_k1a[20], a10_k4a[20] );
xor a10_C909 ( k9b[83], a10_k1a[19], a10_k4a[19] );
xor a10_C910 ( k9b[82], a10_k1a[18], a10_k4a[18] );
xor a10_C911 ( k9b[81], a10_k1a[17], a10_k4a[17] );
xor a10_C912 ( k9b[80], a10_k1a[16], a10_k4a[16] );
xor a10_C913 ( k9b[79], a10_k1a[15], a10_k4a[15] );
xor a10_C914 ( k9b[78], a10_k1a[14], a10_k4a[14] );
xor a10_C915 ( k9b[77], a10_k1a[13], a10_k4a[13] );
xor a10_C916 ( k9b[76], a10_k1a[12], a10_k4a[12] );
xor a10_C917 ( k9b[75], a10_k1a[11], a10_k4a[11] );
xor a10_C918 ( k9b[74], a10_k1a[10], a10_k4a[10] );
xor a10_C919 ( k9b[73], a10_k1a[9], a10_k4a[9] );
xor a10_C920 ( k9b[72], a10_k1a[8], a10_k4a[8] );
xor a10_C921 ( k9b[71], a10_k1a[7], a10_k4a[7] );
xor a10_C922 ( k9b[70], a10_k1a[6], a10_k4a[6] );
xor a10_C923 ( k9b[69], a10_k1a[5], a10_k4a[5] );
xor a10_C924 ( k9b[68], a10_k1a[4], a10_k4a[4] );
xor a10_C925 ( k9b[67], a10_k1a[3], a10_k4a[3] );
xor a10_C926 ( k9b[66], a10_k1a[2], a10_k4a[2] );
xor a10_C927 ( k9b[65], a10_k1a[1], a10_k4a[1] );
xor a10_C928 ( k9b[64], a10_k1a[0], a10_k4a[0] );
xor a10_C929 ( k9b[63], a10_k2a[31], a10_k4a[31] );
xor a10_C930 ( k9b[62], a10_k2a[30], a10_k4a[30] );
xor a10_C931 ( k9b[61], a10_k2a[29], a10_k4a[29] );
xor a10_C932 ( k9b[60], a10_k2a[28], a10_k4a[28] );
xor a10_C933 ( k9b[59], a10_k2a[27], a10_k4a[27] );
xor a10_C934 ( k9b[58], a10_k2a[26], a10_k4a[26] );
xor a10_C935 ( k9b[57], a10_k2a[25], a10_k4a[25] );
xor a10_C936 ( k9b[56], a10_k2a[24], a10_k4a[24] );
xor a10_C937 ( k9b[55], a10_k2a[23], a10_k4a[23] );
xor a10_C938 ( k9b[54], a10_k2a[22], a10_k4a[22] );
xor a10_C939 ( k9b[53], a10_k2a[21], a10_k4a[21] );
xor a10_C940 ( k9b[52], a10_k2a[20], a10_k4a[20] );
xor a10_C941 ( k9b[51], a10_k2a[19], a10_k4a[19] );
xor a10_C942 ( k9b[50], a10_k2a[18], a10_k4a[18] );
xor a10_C943 ( k9b[49], a10_k2a[17], a10_k4a[17] );
xor a10_C944 ( k9b[48], a10_k2a[16], a10_k4a[16] );
xor a10_C945 ( k9b[47], a10_k2a[15], a10_k4a[15] );
xor a10_C946 ( k9b[46], a10_k2a[14], a10_k4a[14] );
xor a10_C947 ( k9b[45], a10_k2a[13], a10_k4a[13] );
xor a10_C948 ( k9b[44], a10_k2a[12], a10_k4a[12] );
xor a10_C949 ( k9b[43], a10_k2a[11], a10_k4a[11] );
xor a10_C950 ( k9b[42], a10_k2a[10], a10_k4a[10] );
xor a10_C951 ( k9b[41], a10_k2a[9], a10_k4a[9] );
xor a10_C952 ( k9b[40], a10_k2a[8], a10_k4a[8] );
xor a10_C953 ( k9b[39], a10_k2a[7], a10_k4a[7] );
xor a10_C954 ( k9b[38], a10_k2a[6], a10_k4a[6] );
xor a10_C955 ( k9b[37], a10_k2a[5], a10_k4a[5] );
xor a10_C956 ( k9b[36], a10_k2a[4], a10_k4a[4] );
xor a10_C957 ( k9b[35], a10_k2a[3], a10_k4a[3] );
xor a10_C958 ( k9b[34], a10_k2a[2], a10_k4a[2] );
xor a10_C959 ( k9b[33], a10_k2a[1], a10_k4a[1] );
xor a10_C960 ( k9b[32], a10_k2a[0], a10_k4a[0] );
xor a10_C961 ( k9b[31], a10_k3a[31], a10_k4a[31] );
xor a10_C962 ( k9b[30], a10_k3a[30], a10_k4a[30] );
xor a10_C963 ( k9b[29], a10_k3a[29], a10_k4a[29] );
xor a10_C964 ( k9b[28], a10_k3a[28], a10_k4a[28] );
xor a10_C965 ( k9b[27], a10_k3a[27], a10_k4a[27] );
xor a10_C966 ( k9b[26], a10_k3a[26], a10_k4a[26] );
xor a10_C967 ( k9b[25], a10_k3a[25], a10_k4a[25] );
xor a10_C968 ( k9b[24], a10_k3a[24], a10_k4a[24] );
xor a10_C969 ( k9b[23], a10_k3a[23], a10_k4a[23] );
xor a10_C970 ( k9b[22], a10_k3a[22], a10_k4a[22] );
xor a10_C971 ( k9b[21], a10_k3a[21], a10_k4a[21] );
xor a10_C972 ( k9b[20], a10_k3a[20], a10_k4a[20] );
xor a10_C973 ( k9b[19], a10_k3a[19], a10_k4a[19] );
xor a10_C974 ( k9b[18], a10_k3a[18], a10_k4a[18] );
xor a10_C975 ( k9b[17], a10_k3a[17], a10_k4a[17] );
xor a10_C976 ( k9b[16], a10_k3a[16], a10_k4a[16] );
xor a10_C977 ( k9b[15], a10_k3a[15], a10_k4a[15] );
xor a10_C978 ( k9b[14], a10_k3a[14], a10_k4a[14] );
xor a10_C979 ( k9b[13], a10_k3a[13], a10_k4a[13] );
xor a10_C980 ( k9b[12], a10_k3a[12], a10_k4a[12] );
xor a10_C981 ( k9b[11], a10_k3a[11], a10_k4a[11] );
xor a10_C982 ( k9b[10], a10_k3a[10], a10_k4a[10] );
xor a10_C983 ( k9b[9], a10_k3a[9], a10_k4a[9] );
xor a10_C984 ( k9b[8], a10_k3a[8], a10_k4a[8] );
xor a10_C985 ( k9b[7], a10_k3a[7], a10_k4a[7] );
xor a10_C986 ( k9b[6], a10_k3a[6], a10_k4a[6] );
xor a10_C987 ( k9b[5], a10_k3a[5], a10_k4a[5] );
xor a10_C988 ( k9b[4], a10_k3a[4], a10_k4a[4] );
xor a10_C989 ( k9b[3], a10_k3a[3], a10_k4a[3] );
xor a10_C990 ( k9b[2], a10_k3a[2], a10_k4a[2] );
xor a10_C991 ( k9b[1], a10_k3a[1], a10_k4a[1] );
xor a10_C992 ( k9b[0], a10_k3a[0], a10_k4a[0] );
xor a9_C961 ( k8b[31], a9_k3a[31], a9_k4a[31] );
xor a8_C961 ( k7b[31], a8_k3a[31], a8_k4a[31] );
xor a7_C961 ( k6b[31], a7_k3a[31], a7_k4a[31] );
xor a6_C961 ( k5b[31], a6_k3a[31], a6_k4a[31] );
xor a5_C961 ( k4b[31], a5_k3a[31], a5_k4a[31] );
xor a4_C961 ( k3b[31], a4_k3a[31], a4_k4a[31] );
xor a3_C961 ( k2b[31], a3_k3a[31], a3_k4a[31] );
xor a2_C961 ( k1b[31], a2_k3a[31], a2_k4a[31] );
xor a1_C961 ( k0b[31], a1_k3a[31], a1_k4a[31] );
xor a1_C896 ( k0b[96], a1_k0a[0], a1_k4a[0] );
xor a1_C895 ( k0b[97], a1_k0a[1], a1_k4a[1] );
xor a1_C894 ( k0b[98], a1_k0a[2], a1_k4a[2] );
xor a1_C893 ( k0b[99], a1_k0a[3], a1_k4a[3] );
xor a1_C892 ( k0b[100], a1_k0a[4], a1_k4a[4] );
xor a1_C891 ( k0b[101], a1_k0a[5], a1_k4a[5] );
xor a1_C890 ( k0b[102], a1_k0a[6], a1_k4a[6] );
xor a1_C889 ( k0b[103], a1_k0a[7], a1_k4a[7] );
xor a1_C888 ( k0b[104], a1_k0a[8], a1_k4a[8] );
xor a1_C887 ( k0b[105], a1_k0a[9], a1_k4a[9] );
xor a1_C886 ( k0b[106], a1_k0a[10], a1_k4a[10] );
xor a1_C885 ( k0b[107], a1_k0a[11], a1_k4a[11] );
xor a1_C884 ( k0b[108], a1_k0a[12], a1_k4a[12] );
xor a1_C883 ( k0b[109], a1_k0a[13], a1_k4a[13] );
xor a1_C882 ( k0b[110], a1_k0a[14], a1_k4a[14] );
xor a1_C881 ( k0b[111], a1_k0a[15], a1_k4a[15] );
xor a1_C880 ( k0b[112], a1_k0a[16], a1_k4a[16] );
xor a1_C879 ( k0b[113], a1_k0a[17], a1_k4a[17] );
xor a1_C878 ( k0b[114], a1_k0a[18], a1_k4a[18] );
xor a1_C877 ( k0b[115], a1_k0a[19], a1_k4a[19] );
xor a1_C876 ( k0b[116], a1_k0a[20], a1_k4a[20] );
xor a1_C875 ( k0b[117], a1_k0a[21], a1_k4a[21] );
xor a1_C874 ( k0b[118], a1_k0a[22], a1_k4a[22] );
xor a1_C873 ( k0b[119], a1_k0a[23], a1_k4a[23] );
xor a1_C872 ( k0b[120], a1_k0a[24], a1_k4a[24] );
xor a1_C871 ( k0b[121], a1_k0a[25], a1_k4a[25] );
xor a1_C870 ( k0b[122], a1_k0a[26], a1_k4a[26] );
xor a1_C869 ( k0b[123], a1_k0a[27], a1_k4a[27] );
xor a1_C868 ( k0b[124], a1_k0a[28], a1_k4a[28] );
xor a1_C867 ( k0b[125], a1_k0a[29], a1_k4a[29] );
xor a1_C866 ( k0b[126], a1_k0a[30], a1_k4a[30] );
xor a1_C865 ( k0b[127], a1_k0a[31], a1_k4a[31] );
xor a1_C992 ( k0b[0], a1_k3a[0], a1_k4a[0] );
xor a1_C991 ( k0b[1], a1_k3a[1], a1_k4a[1] );
xor a1_C990 ( k0b[2], a1_k3a[2], a1_k4a[2] );
xor a1_C989 ( k0b[3], a1_k3a[3], a1_k4a[3] );
xor a1_C988 ( k0b[4], a1_k3a[4], a1_k4a[4] );
xor a1_C987 ( k0b[5], a1_k3a[5], a1_k4a[5] );
xor a1_C986 ( k0b[6], a1_k3a[6], a1_k4a[6] );
xor a1_C985 ( k0b[7], a1_k3a[7], a1_k4a[7] );
xor a1_C984 ( k0b[8], a1_k3a[8], a1_k4a[8] );
xor a1_C983 ( k0b[9], a1_k3a[9], a1_k4a[9] );
xor a1_C982 ( k0b[10], a1_k3a[10], a1_k4a[10] );
xor a1_C981 ( k0b[11], a1_k3a[11], a1_k4a[11] );
xor a1_C980 ( k0b[12], a1_k3a[12], a1_k4a[12] );
xor a1_C979 ( k0b[13], a1_k3a[13], a1_k4a[13] );
xor a1_C978 ( k0b[14], a1_k3a[14], a1_k4a[14] );
xor a1_C977 ( k0b[15], a1_k3a[15], a1_k4a[15] );
xor a1_C976 ( k0b[16], a1_k3a[16], a1_k4a[16] );
xor a1_C975 ( k0b[17], a1_k3a[17], a1_k4a[17] );
xor a1_C974 ( k0b[18], a1_k3a[18], a1_k4a[18] );
xor a1_C973 ( k0b[19], a1_k3a[19], a1_k4a[19] );
xor a1_C972 ( k0b[20], a1_k3a[20], a1_k4a[20] );
xor a1_C971 ( k0b[21], a1_k3a[21], a1_k4a[21] );
xor a1_C970 ( k0b[22], a1_k3a[22], a1_k4a[22] );
xor a1_C969 ( k0b[23], a1_k3a[23], a1_k4a[23] );
xor a1_C968 ( k0b[24], a1_k3a[24], a1_k4a[24] );
xor a1_C967 ( k0b[25], a1_k3a[25], a1_k4a[25] );
xor a1_C966 ( k0b[26], a1_k3a[26], a1_k4a[26] );
xor a1_C965 ( k0b[27], a1_k3a[27], a1_k4a[27] );
xor a1_C964 ( k0b[28], a1_k3a[28], a1_k4a[28] );
xor a1_C963 ( k0b[29], a1_k3a[29], a1_k4a[29] );
xor a1_C962 ( k0b[30], a1_k3a[30], a1_k4a[30] );
xor a1_C960 ( k0b[32], a1_k2a[0], a1_k4a[0] );
xor a1_C959 ( k0b[33], a1_k2a[1], a1_k4a[1] );
xor a1_C958 ( k0b[34], a1_k2a[2], a1_k4a[2] );
xor a1_C957 ( k0b[35], a1_k2a[3], a1_k4a[3] );
xor a1_C956 ( k0b[36], a1_k2a[4], a1_k4a[4] );
xor a1_C955 ( k0b[37], a1_k2a[5], a1_k4a[5] );
xor a1_C954 ( k0b[38], a1_k2a[6], a1_k4a[6] );
xor a1_C953 ( k0b[39], a1_k2a[7], a1_k4a[7] );
xor a1_C952 ( k0b[40], a1_k2a[8], a1_k4a[8] );
xor a1_C951 ( k0b[41], a1_k2a[9], a1_k4a[9] );
xor a1_C950 ( k0b[42], a1_k2a[10], a1_k4a[10] );
xor a1_C949 ( k0b[43], a1_k2a[11], a1_k4a[11] );
xor a1_C948 ( k0b[44], a1_k2a[12], a1_k4a[12] );
xor a1_C947 ( k0b[45], a1_k2a[13], a1_k4a[13] );
xor a1_C946 ( k0b[46], a1_k2a[14], a1_k4a[14] );
xor a1_C945 ( k0b[47], a1_k2a[15], a1_k4a[15] );
xor a1_C944 ( k0b[48], a1_k2a[16], a1_k4a[16] );
xor a1_C943 ( k0b[49], a1_k2a[17], a1_k4a[17] );
xor a1_C942 ( k0b[50], a1_k2a[18], a1_k4a[18] );
xor a1_C941 ( k0b[51], a1_k2a[19], a1_k4a[19] );
xor a1_C940 ( k0b[52], a1_k2a[20], a1_k4a[20] );
xor a1_C939 ( k0b[53], a1_k2a[21], a1_k4a[21] );
xor a1_C938 ( k0b[54], a1_k2a[22], a1_k4a[22] );
xor a1_C937 ( k0b[55], a1_k2a[23], a1_k4a[23] );
xor a1_C936 ( k0b[56], a1_k2a[24], a1_k4a[24] );
xor a1_C935 ( k0b[57], a1_k2a[25], a1_k4a[25] );
xor a1_C934 ( k0b[58], a1_k2a[26], a1_k4a[26] );
xor a1_C933 ( k0b[59], a1_k2a[27], a1_k4a[27] );
xor a1_C932 ( k0b[60], a1_k2a[28], a1_k4a[28] );
xor a1_C931 ( k0b[61], a1_k2a[29], a1_k4a[29] );
xor a1_C930 ( k0b[62], a1_k2a[30], a1_k4a[30] );
xor a1_C929 ( k0b[63], a1_k2a[31], a1_k4a[31] );
xor a1_C928 ( k0b[64], a1_k1a[0], a1_k4a[0] );
xor a1_C927 ( k0b[65], a1_k1a[1], a1_k4a[1] );
xor a1_C926 ( k0b[66], a1_k1a[2], a1_k4a[2] );
xor a1_C925 ( k0b[67], a1_k1a[3], a1_k4a[3] );
xor a1_C924 ( k0b[68], a1_k1a[4], a1_k4a[4] );
xor a1_C923 ( k0b[69], a1_k1a[5], a1_k4a[5] );
xor a1_C922 ( k0b[70], a1_k1a[6], a1_k4a[6] );
xor a1_C921 ( k0b[71], a1_k1a[7], a1_k4a[7] );
xor a1_C920 ( k0b[72], a1_k1a[8], a1_k4a[8] );
xor a1_C919 ( k0b[73], a1_k1a[9], a1_k4a[9] );
xor a1_C918 ( k0b[74], a1_k1a[10], a1_k4a[10] );
xor a1_C917 ( k0b[75], a1_k1a[11], a1_k4a[11] );
xor a1_C916 ( k0b[76], a1_k1a[12], a1_k4a[12] );
xor a1_C915 ( k0b[77], a1_k1a[13], a1_k4a[13] );
xor a1_C914 ( k0b[78], a1_k1a[14], a1_k4a[14] );
xor a1_C913 ( k0b[79], a1_k1a[15], a1_k4a[15] );
xor a1_C912 ( k0b[80], a1_k1a[16], a1_k4a[16] );
xor a1_C911 ( k0b[81], a1_k1a[17], a1_k4a[17] );
xor a1_C910 ( k0b[82], a1_k1a[18], a1_k4a[18] );
xor a1_C909 ( k0b[83], a1_k1a[19], a1_k4a[19] );
xor a1_C908 ( k0b[84], a1_k1a[20], a1_k4a[20] );
xor a1_C907 ( k0b[85], a1_k1a[21], a1_k4a[21] );
xor a1_C906 ( k0b[86], a1_k1a[22], a1_k4a[22] );
xor a1_C905 ( k0b[87], a1_k1a[23], a1_k4a[23] );
xor a1_C904 ( k0b[88], a1_k1a[24], a1_k4a[24] );
xor a1_C903 ( k0b[89], a1_k1a[25], a1_k4a[25] );
xor a1_C902 ( k0b[90], a1_k1a[26], a1_k4a[26] );
xor a1_C901 ( k0b[91], a1_k1a[27], a1_k4a[27] );
xor a1_C900 ( k0b[92], a1_k1a[28], a1_k4a[28] );
xor a1_C899 ( k0b[93], a1_k1a[29], a1_k4a[29] );
xor a1_C898 ( k0b[94], a1_k1a[30], a1_k4a[30] );
xor a1_C897 ( k0b[95], a1_k1a[31], a1_k4a[31] );
xor a2_C896 ( k1b[96], a2_k0a[0], a2_k4a[0] );
xor a2_C895 ( k1b[97], a2_k0a[1], a2_k4a[1] );
xor a2_C894 ( k1b[98], a2_k0a[2], a2_k4a[2] );
xor a2_C893 ( k1b[99], a2_k0a[3], a2_k4a[3] );
xor a2_C892 ( k1b[100], a2_k0a[4], a2_k4a[4] );
xor a2_C891 ( k1b[101], a2_k0a[5], a2_k4a[5] );
xor a2_C890 ( k1b[102], a2_k0a[6], a2_k4a[6] );
xor a2_C889 ( k1b[103], a2_k0a[7], a2_k4a[7] );
xor a2_C888 ( k1b[104], a2_k0a[8], a2_k4a[8] );
xor a2_C887 ( k1b[105], a2_k0a[9], a2_k4a[9] );
xor a2_C886 ( k1b[106], a2_k0a[10], a2_k4a[10] );
xor a2_C885 ( k1b[107], a2_k0a[11], a2_k4a[11] );
xor a2_C884 ( k1b[108], a2_k0a[12], a2_k4a[12] );
xor a2_C883 ( k1b[109], a2_k0a[13], a2_k4a[13] );
xor a2_C882 ( k1b[110], a2_k0a[14], a2_k4a[14] );
xor a2_C881 ( k1b[111], a2_k0a[15], a2_k4a[15] );
xor a2_C880 ( k1b[112], a2_k0a[16], a2_k4a[16] );
xor a2_C879 ( k1b[113], a2_k0a[17], a2_k4a[17] );
xor a2_C878 ( k1b[114], a2_k0a[18], a2_k4a[18] );
xor a2_C877 ( k1b[115], a2_k0a[19], a2_k4a[19] );
xor a2_C876 ( k1b[116], a2_k0a[20], a2_k4a[20] );
xor a2_C875 ( k1b[117], a2_k0a[21], a2_k4a[21] );
xor a2_C874 ( k1b[118], a2_k0a[22], a2_k4a[22] );
xor a2_C873 ( k1b[119], a2_k0a[23], a2_k4a[23] );
xor a2_C872 ( k1b[120], a2_k0a[24], a2_k4a[24] );
xor a2_C871 ( k1b[121], a2_k0a[25], a2_k4a[25] );
xor a2_C870 ( k1b[122], a2_k0a[26], a2_k4a[26] );
xor a2_C869 ( k1b[123], a2_k0a[27], a2_k4a[27] );
xor a2_C868 ( k1b[124], a2_k0a[28], a2_k4a[28] );
xor a2_C867 ( k1b[125], a2_k0a[29], a2_k4a[29] );
xor a2_C866 ( k1b[126], a2_k0a[30], a2_k4a[30] );
xor a2_C865 ( k1b[127], a2_k0a[31], a2_k4a[31] );
xor a2_C992 ( k1b[0], a2_k3a[0], a2_k4a[0] );
xor a2_C991 ( k1b[1], a2_k3a[1], a2_k4a[1] );
xor a2_C990 ( k1b[2], a2_k3a[2], a2_k4a[2] );
xor a2_C989 ( k1b[3], a2_k3a[3], a2_k4a[3] );
xor a2_C988 ( k1b[4], a2_k3a[4], a2_k4a[4] );
xor a2_C987 ( k1b[5], a2_k3a[5], a2_k4a[5] );
xor a2_C986 ( k1b[6], a2_k3a[6], a2_k4a[6] );
xor a2_C985 ( k1b[7], a2_k3a[7], a2_k4a[7] );
xor a2_C984 ( k1b[8], a2_k3a[8], a2_k4a[8] );
xor a2_C983 ( k1b[9], a2_k3a[9], a2_k4a[9] );
xor a2_C982 ( k1b[10], a2_k3a[10], a2_k4a[10] );
xor a2_C981 ( k1b[11], a2_k3a[11], a2_k4a[11] );
xor a2_C980 ( k1b[12], a2_k3a[12], a2_k4a[12] );
xor a2_C979 ( k1b[13], a2_k3a[13], a2_k4a[13] );
xor a2_C978 ( k1b[14], a2_k3a[14], a2_k4a[14] );
xor a2_C977 ( k1b[15], a2_k3a[15], a2_k4a[15] );
xor a2_C976 ( k1b[16], a2_k3a[16], a2_k4a[16] );
xor a2_C975 ( k1b[17], a2_k3a[17], a2_k4a[17] );
xor a2_C974 ( k1b[18], a2_k3a[18], a2_k4a[18] );
xor a2_C973 ( k1b[19], a2_k3a[19], a2_k4a[19] );
xor a2_C972 ( k1b[20], a2_k3a[20], a2_k4a[20] );
xor a2_C971 ( k1b[21], a2_k3a[21], a2_k4a[21] );
xor a2_C970 ( k1b[22], a2_k3a[22], a2_k4a[22] );
xor a2_C969 ( k1b[23], a2_k3a[23], a2_k4a[23] );
xor a2_C968 ( k1b[24], a2_k3a[24], a2_k4a[24] );
xor a2_C967 ( k1b[25], a2_k3a[25], a2_k4a[25] );
xor a2_C966 ( k1b[26], a2_k3a[26], a2_k4a[26] );
xor a2_C965 ( k1b[27], a2_k3a[27], a2_k4a[27] );
xor a2_C964 ( k1b[28], a2_k3a[28], a2_k4a[28] );
xor a2_C963 ( k1b[29], a2_k3a[29], a2_k4a[29] );
xor a2_C962 ( k1b[30], a2_k3a[30], a2_k4a[30] );
xor a2_C960 ( k1b[32], a2_k2a[0], a2_k4a[0] );
xor a2_C959 ( k1b[33], a2_k2a[1], a2_k4a[1] );
xor a2_C958 ( k1b[34], a2_k2a[2], a2_k4a[2] );
xor a2_C957 ( k1b[35], a2_k2a[3], a2_k4a[3] );
xor a2_C956 ( k1b[36], a2_k2a[4], a2_k4a[4] );
xor a2_C955 ( k1b[37], a2_k2a[5], a2_k4a[5] );
xor a2_C954 ( k1b[38], a2_k2a[6], a2_k4a[6] );
xor a2_C953 ( k1b[39], a2_k2a[7], a2_k4a[7] );
xor a2_C952 ( k1b[40], a2_k2a[8], a2_k4a[8] );
xor a2_C951 ( k1b[41], a2_k2a[9], a2_k4a[9] );
xor a2_C950 ( k1b[42], a2_k2a[10], a2_k4a[10] );
xor a2_C949 ( k1b[43], a2_k2a[11], a2_k4a[11] );
xor a2_C948 ( k1b[44], a2_k2a[12], a2_k4a[12] );
xor a2_C947 ( k1b[45], a2_k2a[13], a2_k4a[13] );
xor a2_C946 ( k1b[46], a2_k2a[14], a2_k4a[14] );
xor a2_C945 ( k1b[47], a2_k2a[15], a2_k4a[15] );
xor a2_C944 ( k1b[48], a2_k2a[16], a2_k4a[16] );
xor a2_C943 ( k1b[49], a2_k2a[17], a2_k4a[17] );
xor a2_C942 ( k1b[50], a2_k2a[18], a2_k4a[18] );
xor a2_C941 ( k1b[51], a2_k2a[19], a2_k4a[19] );
xor a2_C940 ( k1b[52], a2_k2a[20], a2_k4a[20] );
xor a2_C939 ( k1b[53], a2_k2a[21], a2_k4a[21] );
xor a2_C938 ( k1b[54], a2_k2a[22], a2_k4a[22] );
xor a2_C937 ( k1b[55], a2_k2a[23], a2_k4a[23] );
xor a2_C936 ( k1b[56], a2_k2a[24], a2_k4a[24] );
xor a2_C935 ( k1b[57], a2_k2a[25], a2_k4a[25] );
xor a2_C934 ( k1b[58], a2_k2a[26], a2_k4a[26] );
xor a2_C933 ( k1b[59], a2_k2a[27], a2_k4a[27] );
xor a2_C932 ( k1b[60], a2_k2a[28], a2_k4a[28] );
xor a2_C931 ( k1b[61], a2_k2a[29], a2_k4a[29] );
xor a2_C930 ( k1b[62], a2_k2a[30], a2_k4a[30] );
xor a2_C929 ( k1b[63], a2_k2a[31], a2_k4a[31] );
xor a2_C928 ( k1b[64], a2_k1a[0], a2_k4a[0] );
xor a2_C927 ( k1b[65], a2_k1a[1], a2_k4a[1] );
xor a2_C926 ( k1b[66], a2_k1a[2], a2_k4a[2] );
xor a2_C925 ( k1b[67], a2_k1a[3], a2_k4a[3] );
xor a2_C924 ( k1b[68], a2_k1a[4], a2_k4a[4] );
xor a2_C923 ( k1b[69], a2_k1a[5], a2_k4a[5] );
xor a2_C922 ( k1b[70], a2_k1a[6], a2_k4a[6] );
xor a2_C921 ( k1b[71], a2_k1a[7], a2_k4a[7] );
xor a2_C920 ( k1b[72], a2_k1a[8], a2_k4a[8] );
xor a2_C919 ( k1b[73], a2_k1a[9], a2_k4a[9] );
xor a2_C918 ( k1b[74], a2_k1a[10], a2_k4a[10] );
xor a2_C917 ( k1b[75], a2_k1a[11], a2_k4a[11] );
xor a2_C916 ( k1b[76], a2_k1a[12], a2_k4a[12] );
xor a2_C915 ( k1b[77], a2_k1a[13], a2_k4a[13] );
xor a2_C914 ( k1b[78], a2_k1a[14], a2_k4a[14] );
xor a2_C913 ( k1b[79], a2_k1a[15], a2_k4a[15] );
xor a2_C912 ( k1b[80], a2_k1a[16], a2_k4a[16] );
xor a2_C911 ( k1b[81], a2_k1a[17], a2_k4a[17] );
xor a2_C910 ( k1b[82], a2_k1a[18], a2_k4a[18] );
xor a2_C909 ( k1b[83], a2_k1a[19], a2_k4a[19] );
xor a2_C908 ( k1b[84], a2_k1a[20], a2_k4a[20] );
xor a2_C907 ( k1b[85], a2_k1a[21], a2_k4a[21] );
xor a2_C906 ( k1b[86], a2_k1a[22], a2_k4a[22] );
xor a2_C905 ( k1b[87], a2_k1a[23], a2_k4a[23] );
xor a2_C904 ( k1b[88], a2_k1a[24], a2_k4a[24] );
xor a2_C903 ( k1b[89], a2_k1a[25], a2_k4a[25] );
xor a2_C902 ( k1b[90], a2_k1a[26], a2_k4a[26] );
xor a2_C901 ( k1b[91], a2_k1a[27], a2_k4a[27] );
xor a2_C900 ( k1b[92], a2_k1a[28], a2_k4a[28] );
xor a2_C899 ( k1b[93], a2_k1a[29], a2_k4a[29] );
xor a2_C898 ( k1b[94], a2_k1a[30], a2_k4a[30] );
xor a2_C897 ( k1b[95], a2_k1a[31], a2_k4a[31] );
xor a3_C896 ( k2b[96], a3_k0a[0], a3_k4a[0] );
xor a3_C895 ( k2b[97], a3_k0a[1], a3_k4a[1] );
xor a3_C894 ( k2b[98], a3_k0a[2], a3_k4a[2] );
xor a3_C893 ( k2b[99], a3_k0a[3], a3_k4a[3] );
xor a3_C892 ( k2b[100], a3_k0a[4], a3_k4a[4] );
xor a3_C891 ( k2b[101], a3_k0a[5], a3_k4a[5] );
xor a3_C890 ( k2b[102], a3_k0a[6], a3_k4a[6] );
xor a3_C889 ( k2b[103], a3_k0a[7], a3_k4a[7] );
xor a3_C888 ( k2b[104], a3_k0a[8], a3_k4a[8] );
xor a3_C887 ( k2b[105], a3_k0a[9], a3_k4a[9] );
xor a3_C886 ( k2b[106], a3_k0a[10], a3_k4a[10] );
xor a3_C885 ( k2b[107], a3_k0a[11], a3_k4a[11] );
xor a3_C884 ( k2b[108], a3_k0a[12], a3_k4a[12] );
xor a3_C883 ( k2b[109], a3_k0a[13], a3_k4a[13] );
xor a3_C882 ( k2b[110], a3_k0a[14], a3_k4a[14] );
xor a3_C881 ( k2b[111], a3_k0a[15], a3_k4a[15] );
xor a3_C880 ( k2b[112], a3_k0a[16], a3_k4a[16] );
xor a3_C879 ( k2b[113], a3_k0a[17], a3_k4a[17] );
xor a3_C878 ( k2b[114], a3_k0a[18], a3_k4a[18] );
xor a3_C877 ( k2b[115], a3_k0a[19], a3_k4a[19] );
xor a3_C876 ( k2b[116], a3_k0a[20], a3_k4a[20] );
xor a3_C875 ( k2b[117], a3_k0a[21], a3_k4a[21] );
xor a3_C874 ( k2b[118], a3_k0a[22], a3_k4a[22] );
xor a3_C873 ( k2b[119], a3_k0a[23], a3_k4a[23] );
xor a3_C872 ( k2b[120], a3_k0a[24], a3_k4a[24] );
xor a3_C871 ( k2b[121], a3_k0a[25], a3_k4a[25] );
xor a3_C870 ( k2b[122], a3_k0a[26], a3_k4a[26] );
xor a3_C869 ( k2b[123], a3_k0a[27], a3_k4a[27] );
xor a3_C868 ( k2b[124], a3_k0a[28], a3_k4a[28] );
xor a3_C867 ( k2b[125], a3_k0a[29], a3_k4a[29] );
xor a3_C866 ( k2b[126], a3_k0a[30], a3_k4a[30] );
xor a3_C865 ( k2b[127], a3_k0a[31], a3_k4a[31] );
xor a3_C992 ( k2b[0], a3_k3a[0], a3_k4a[0] );
xor a3_C991 ( k2b[1], a3_k3a[1], a3_k4a[1] );
xor a3_C990 ( k2b[2], a3_k3a[2], a3_k4a[2] );
xor a3_C989 ( k2b[3], a3_k3a[3], a3_k4a[3] );
xor a3_C988 ( k2b[4], a3_k3a[4], a3_k4a[4] );
xor a3_C987 ( k2b[5], a3_k3a[5], a3_k4a[5] );
xor a3_C986 ( k2b[6], a3_k3a[6], a3_k4a[6] );
xor a3_C985 ( k2b[7], a3_k3a[7], a3_k4a[7] );
xor a3_C984 ( k2b[8], a3_k3a[8], a3_k4a[8] );
xor a3_C983 ( k2b[9], a3_k3a[9], a3_k4a[9] );
xor a3_C982 ( k2b[10], a3_k3a[10], a3_k4a[10] );
xor a3_C981 ( k2b[11], a3_k3a[11], a3_k4a[11] );
xor a3_C980 ( k2b[12], a3_k3a[12], a3_k4a[12] );
xor a3_C979 ( k2b[13], a3_k3a[13], a3_k4a[13] );
xor a3_C978 ( k2b[14], a3_k3a[14], a3_k4a[14] );
xor a3_C977 ( k2b[15], a3_k3a[15], a3_k4a[15] );
xor a3_C976 ( k2b[16], a3_k3a[16], a3_k4a[16] );
xor a3_C975 ( k2b[17], a3_k3a[17], a3_k4a[17] );
xor a3_C974 ( k2b[18], a3_k3a[18], a3_k4a[18] );
xor a3_C973 ( k2b[19], a3_k3a[19], a3_k4a[19] );
xor a3_C972 ( k2b[20], a3_k3a[20], a3_k4a[20] );
xor a3_C971 ( k2b[21], a3_k3a[21], a3_k4a[21] );
xor a3_C970 ( k2b[22], a3_k3a[22], a3_k4a[22] );
xor a3_C969 ( k2b[23], a3_k3a[23], a3_k4a[23] );
xor a3_C968 ( k2b[24], a3_k3a[24], a3_k4a[24] );
xor a3_C967 ( k2b[25], a3_k3a[25], a3_k4a[25] );
xor a3_C966 ( k2b[26], a3_k3a[26], a3_k4a[26] );
xor a3_C965 ( k2b[27], a3_k3a[27], a3_k4a[27] );
xor a3_C964 ( k2b[28], a3_k3a[28], a3_k4a[28] );
xor a3_C963 ( k2b[29], a3_k3a[29], a3_k4a[29] );
xor a3_C962 ( k2b[30], a3_k3a[30], a3_k4a[30] );
xor a3_C960 ( k2b[32], a3_k2a[0], a3_k4a[0] );
xor a3_C959 ( k2b[33], a3_k2a[1], a3_k4a[1] );
xor a3_C958 ( k2b[34], a3_k2a[2], a3_k4a[2] );
xor a3_C957 ( k2b[35], a3_k2a[3], a3_k4a[3] );
xor a3_C956 ( k2b[36], a3_k2a[4], a3_k4a[4] );
xor a3_C955 ( k2b[37], a3_k2a[5], a3_k4a[5] );
xor a3_C954 ( k2b[38], a3_k2a[6], a3_k4a[6] );
xor a3_C953 ( k2b[39], a3_k2a[7], a3_k4a[7] );
xor a3_C952 ( k2b[40], a3_k2a[8], a3_k4a[8] );
xor a3_C951 ( k2b[41], a3_k2a[9], a3_k4a[9] );
xor a3_C950 ( k2b[42], a3_k2a[10], a3_k4a[10] );
xor a3_C949 ( k2b[43], a3_k2a[11], a3_k4a[11] );
xor a3_C948 ( k2b[44], a3_k2a[12], a3_k4a[12] );
xor a3_C947 ( k2b[45], a3_k2a[13], a3_k4a[13] );
xor a3_C946 ( k2b[46], a3_k2a[14], a3_k4a[14] );
xor a3_C945 ( k2b[47], a3_k2a[15], a3_k4a[15] );
xor a3_C944 ( k2b[48], a3_k2a[16], a3_k4a[16] );
xor a3_C943 ( k2b[49], a3_k2a[17], a3_k4a[17] );
xor a3_C942 ( k2b[50], a3_k2a[18], a3_k4a[18] );
xor a3_C941 ( k2b[51], a3_k2a[19], a3_k4a[19] );
xor a3_C940 ( k2b[52], a3_k2a[20], a3_k4a[20] );
xor a3_C939 ( k2b[53], a3_k2a[21], a3_k4a[21] );
xor a3_C938 ( k2b[54], a3_k2a[22], a3_k4a[22] );
xor a3_C937 ( k2b[55], a3_k2a[23], a3_k4a[23] );
xor a3_C936 ( k2b[56], a3_k2a[24], a3_k4a[24] );
xor a3_C935 ( k2b[57], a3_k2a[25], a3_k4a[25] );
xor a3_C934 ( k2b[58], a3_k2a[26], a3_k4a[26] );
xor a3_C933 ( k2b[59], a3_k2a[27], a3_k4a[27] );
xor a3_C932 ( k2b[60], a3_k2a[28], a3_k4a[28] );
xor a3_C931 ( k2b[61], a3_k2a[29], a3_k4a[29] );
xor a3_C930 ( k2b[62], a3_k2a[30], a3_k4a[30] );
xor a3_C929 ( k2b[63], a3_k2a[31], a3_k4a[31] );
xor a3_C928 ( k2b[64], a3_k1a[0], a3_k4a[0] );
xor a3_C927 ( k2b[65], a3_k1a[1], a3_k4a[1] );
xor a3_C926 ( k2b[66], a3_k1a[2], a3_k4a[2] );
xor a3_C925 ( k2b[67], a3_k1a[3], a3_k4a[3] );
xor a3_C924 ( k2b[68], a3_k1a[4], a3_k4a[4] );
xor a3_C923 ( k2b[69], a3_k1a[5], a3_k4a[5] );
xor a3_C922 ( k2b[70], a3_k1a[6], a3_k4a[6] );
xor a3_C921 ( k2b[71], a3_k1a[7], a3_k4a[7] );
xor a3_C920 ( k2b[72], a3_k1a[8], a3_k4a[8] );
xor a3_C919 ( k2b[73], a3_k1a[9], a3_k4a[9] );
xor a3_C918 ( k2b[74], a3_k1a[10], a3_k4a[10] );
xor a3_C917 ( k2b[75], a3_k1a[11], a3_k4a[11] );
xor a3_C916 ( k2b[76], a3_k1a[12], a3_k4a[12] );
xor a3_C915 ( k2b[77], a3_k1a[13], a3_k4a[13] );
xor a3_C914 ( k2b[78], a3_k1a[14], a3_k4a[14] );
xor a3_C913 ( k2b[79], a3_k1a[15], a3_k4a[15] );
xor a3_C912 ( k2b[80], a3_k1a[16], a3_k4a[16] );
xor a3_C911 ( k2b[81], a3_k1a[17], a3_k4a[17] );
xor a3_C910 ( k2b[82], a3_k1a[18], a3_k4a[18] );
xor a3_C909 ( k2b[83], a3_k1a[19], a3_k4a[19] );
xor a3_C908 ( k2b[84], a3_k1a[20], a3_k4a[20] );
xor a3_C907 ( k2b[85], a3_k1a[21], a3_k4a[21] );
xor a3_C906 ( k2b[86], a3_k1a[22], a3_k4a[22] );
xor a3_C905 ( k2b[87], a3_k1a[23], a3_k4a[23] );
xor a3_C904 ( k2b[88], a3_k1a[24], a3_k4a[24] );
xor a3_C903 ( k2b[89], a3_k1a[25], a3_k4a[25] );
xor a3_C902 ( k2b[90], a3_k1a[26], a3_k4a[26] );
xor a3_C901 ( k2b[91], a3_k1a[27], a3_k4a[27] );
xor a3_C900 ( k2b[92], a3_k1a[28], a3_k4a[28] );
xor a3_C899 ( k2b[93], a3_k1a[29], a3_k4a[29] );
xor a3_C898 ( k2b[94], a3_k1a[30], a3_k4a[30] );
xor a3_C897 ( k2b[95], a3_k1a[31], a3_k4a[31] );
xor a4_C896 ( k3b[96], a4_k0a[0], a4_k4a[0] );
xor a4_C895 ( k3b[97], a4_k0a[1], a4_k4a[1] );
xor a4_C894 ( k3b[98], a4_k0a[2], a4_k4a[2] );
xor a4_C893 ( k3b[99], a4_k0a[3], a4_k4a[3] );
xor a4_C892 ( k3b[100], a4_k0a[4], a4_k4a[4] );
xor a4_C891 ( k3b[101], a4_k0a[5], a4_k4a[5] );
xor a4_C890 ( k3b[102], a4_k0a[6], a4_k4a[6] );
xor a4_C889 ( k3b[103], a4_k0a[7], a4_k4a[7] );
xor a4_C888 ( k3b[104], a4_k0a[8], a4_k4a[8] );
xor a4_C887 ( k3b[105], a4_k0a[9], a4_k4a[9] );
xor a4_C886 ( k3b[106], a4_k0a[10], a4_k4a[10] );
xor a4_C885 ( k3b[107], a4_k0a[11], a4_k4a[11] );
xor a4_C884 ( k3b[108], a4_k0a[12], a4_k4a[12] );
xor a4_C883 ( k3b[109], a4_k0a[13], a4_k4a[13] );
xor a4_C882 ( k3b[110], a4_k0a[14], a4_k4a[14] );
xor a4_C881 ( k3b[111], a4_k0a[15], a4_k4a[15] );
xor a4_C880 ( k3b[112], a4_k0a[16], a4_k4a[16] );
xor a4_C879 ( k3b[113], a4_k0a[17], a4_k4a[17] );
xor a4_C878 ( k3b[114], a4_k0a[18], a4_k4a[18] );
xor a4_C877 ( k3b[115], a4_k0a[19], a4_k4a[19] );
xor a4_C876 ( k3b[116], a4_k0a[20], a4_k4a[20] );
xor a4_C875 ( k3b[117], a4_k0a[21], a4_k4a[21] );
xor a4_C874 ( k3b[118], a4_k0a[22], a4_k4a[22] );
xor a4_C873 ( k3b[119], a4_k0a[23], a4_k4a[23] );
xor a4_C872 ( k3b[120], a4_k0a[24], a4_k4a[24] );
xor a4_C871 ( k3b[121], a4_k0a[25], a4_k4a[25] );
xor a4_C870 ( k3b[122], a4_k0a[26], a4_k4a[26] );
xor a4_C869 ( k3b[123], a4_k0a[27], a4_k4a[27] );
xor a4_C868 ( k3b[124], a4_k0a[28], a4_k4a[28] );
xor a4_C867 ( k3b[125], a4_k0a[29], a4_k4a[29] );
xor a4_C866 ( k3b[126], a4_k0a[30], a4_k4a[30] );
xor a4_C865 ( k3b[127], a4_k0a[31], a4_k4a[31] );
xor a4_C992 ( k3b[0], a4_k3a[0], a4_k4a[0] );
xor a4_C991 ( k3b[1], a4_k3a[1], a4_k4a[1] );
xor a4_C990 ( k3b[2], a4_k3a[2], a4_k4a[2] );
xor a4_C989 ( k3b[3], a4_k3a[3], a4_k4a[3] );
xor a4_C988 ( k3b[4], a4_k3a[4], a4_k4a[4] );
xor a4_C987 ( k3b[5], a4_k3a[5], a4_k4a[5] );
xor a4_C986 ( k3b[6], a4_k3a[6], a4_k4a[6] );
xor a4_C985 ( k3b[7], a4_k3a[7], a4_k4a[7] );
xor a4_C984 ( k3b[8], a4_k3a[8], a4_k4a[8] );
xor a4_C983 ( k3b[9], a4_k3a[9], a4_k4a[9] );
xor a4_C982 ( k3b[10], a4_k3a[10], a4_k4a[10] );
xor a4_C981 ( k3b[11], a4_k3a[11], a4_k4a[11] );
xor a4_C980 ( k3b[12], a4_k3a[12], a4_k4a[12] );
xor a4_C979 ( k3b[13], a4_k3a[13], a4_k4a[13] );
xor a4_C978 ( k3b[14], a4_k3a[14], a4_k4a[14] );
xor a4_C977 ( k3b[15], a4_k3a[15], a4_k4a[15] );
xor a4_C976 ( k3b[16], a4_k3a[16], a4_k4a[16] );
xor a4_C975 ( k3b[17], a4_k3a[17], a4_k4a[17] );
xor a4_C974 ( k3b[18], a4_k3a[18], a4_k4a[18] );
xor a4_C973 ( k3b[19], a4_k3a[19], a4_k4a[19] );
xor a4_C972 ( k3b[20], a4_k3a[20], a4_k4a[20] );
xor a4_C971 ( k3b[21], a4_k3a[21], a4_k4a[21] );
xor a4_C970 ( k3b[22], a4_k3a[22], a4_k4a[22] );
xor a4_C969 ( k3b[23], a4_k3a[23], a4_k4a[23] );
xor a4_C968 ( k3b[24], a4_k3a[24], a4_k4a[24] );
xor a4_C967 ( k3b[25], a4_k3a[25], a4_k4a[25] );
xor a4_C966 ( k3b[26], a4_k3a[26], a4_k4a[26] );
xor a4_C965 ( k3b[27], a4_k3a[27], a4_k4a[27] );
xor a4_C964 ( k3b[28], a4_k3a[28], a4_k4a[28] );
xor a4_C963 ( k3b[29], a4_k3a[29], a4_k4a[29] );
xor a4_C962 ( k3b[30], a4_k3a[30], a4_k4a[30] );
xor a4_C960 ( k3b[32], a4_k2a[0], a4_k4a[0] );
xor a4_C959 ( k3b[33], a4_k2a[1], a4_k4a[1] );
xor a4_C958 ( k3b[34], a4_k2a[2], a4_k4a[2] );
xor a4_C957 ( k3b[35], a4_k2a[3], a4_k4a[3] );
xor a4_C956 ( k3b[36], a4_k2a[4], a4_k4a[4] );
xor a4_C955 ( k3b[37], a4_k2a[5], a4_k4a[5] );
xor a4_C954 ( k3b[38], a4_k2a[6], a4_k4a[6] );
xor a4_C953 ( k3b[39], a4_k2a[7], a4_k4a[7] );
xor a4_C952 ( k3b[40], a4_k2a[8], a4_k4a[8] );
xor a4_C951 ( k3b[41], a4_k2a[9], a4_k4a[9] );
xor a4_C950 ( k3b[42], a4_k2a[10], a4_k4a[10] );
xor a4_C949 ( k3b[43], a4_k2a[11], a4_k4a[11] );
xor a4_C948 ( k3b[44], a4_k2a[12], a4_k4a[12] );
xor a4_C947 ( k3b[45], a4_k2a[13], a4_k4a[13] );
xor a4_C946 ( k3b[46], a4_k2a[14], a4_k4a[14] );
xor a4_C945 ( k3b[47], a4_k2a[15], a4_k4a[15] );
xor a4_C944 ( k3b[48], a4_k2a[16], a4_k4a[16] );
xor a4_C943 ( k3b[49], a4_k2a[17], a4_k4a[17] );
xor a4_C942 ( k3b[50], a4_k2a[18], a4_k4a[18] );
xor a4_C941 ( k3b[51], a4_k2a[19], a4_k4a[19] );
xor a4_C940 ( k3b[52], a4_k2a[20], a4_k4a[20] );
xor a4_C939 ( k3b[53], a4_k2a[21], a4_k4a[21] );
xor a4_C938 ( k3b[54], a4_k2a[22], a4_k4a[22] );
xor a4_C937 ( k3b[55], a4_k2a[23], a4_k4a[23] );
xor a4_C936 ( k3b[56], a4_k2a[24], a4_k4a[24] );
xor a4_C935 ( k3b[57], a4_k2a[25], a4_k4a[25] );
xor a4_C934 ( k3b[58], a4_k2a[26], a4_k4a[26] );
xor a4_C933 ( k3b[59], a4_k2a[27], a4_k4a[27] );
xor a4_C932 ( k3b[60], a4_k2a[28], a4_k4a[28] );
xor a4_C931 ( k3b[61], a4_k2a[29], a4_k4a[29] );
xor a4_C930 ( k3b[62], a4_k2a[30], a4_k4a[30] );
xor a4_C929 ( k3b[63], a4_k2a[31], a4_k4a[31] );
xor a4_C928 ( k3b[64], a4_k1a[0], a4_k4a[0] );
xor a4_C927 ( k3b[65], a4_k1a[1], a4_k4a[1] );
xor a4_C926 ( k3b[66], a4_k1a[2], a4_k4a[2] );
xor a4_C925 ( k3b[67], a4_k1a[3], a4_k4a[3] );
xor a4_C924 ( k3b[68], a4_k1a[4], a4_k4a[4] );
xor a4_C923 ( k3b[69], a4_k1a[5], a4_k4a[5] );
xor a4_C922 ( k3b[70], a4_k1a[6], a4_k4a[6] );
xor a4_C921 ( k3b[71], a4_k1a[7], a4_k4a[7] );
xor a4_C920 ( k3b[72], a4_k1a[8], a4_k4a[8] );
xor a4_C919 ( k3b[73], a4_k1a[9], a4_k4a[9] );
xor a4_C918 ( k3b[74], a4_k1a[10], a4_k4a[10] );
xor a4_C917 ( k3b[75], a4_k1a[11], a4_k4a[11] );
xor a4_C916 ( k3b[76], a4_k1a[12], a4_k4a[12] );
xor a4_C915 ( k3b[77], a4_k1a[13], a4_k4a[13] );
xor a4_C914 ( k3b[78], a4_k1a[14], a4_k4a[14] );
xor a4_C913 ( k3b[79], a4_k1a[15], a4_k4a[15] );
xor a4_C912 ( k3b[80], a4_k1a[16], a4_k4a[16] );
xor a4_C911 ( k3b[81], a4_k1a[17], a4_k4a[17] );
xor a4_C910 ( k3b[82], a4_k1a[18], a4_k4a[18] );
xor a4_C909 ( k3b[83], a4_k1a[19], a4_k4a[19] );
xor a4_C908 ( k3b[84], a4_k1a[20], a4_k4a[20] );
xor a4_C907 ( k3b[85], a4_k1a[21], a4_k4a[21] );
xor a4_C906 ( k3b[86], a4_k1a[22], a4_k4a[22] );
xor a4_C905 ( k3b[87], a4_k1a[23], a4_k4a[23] );
xor a4_C904 ( k3b[88], a4_k1a[24], a4_k4a[24] );
xor a4_C903 ( k3b[89], a4_k1a[25], a4_k4a[25] );
xor a4_C902 ( k3b[90], a4_k1a[26], a4_k4a[26] );
xor a4_C901 ( k3b[91], a4_k1a[27], a4_k4a[27] );
xor a4_C900 ( k3b[92], a4_k1a[28], a4_k4a[28] );
xor a4_C899 ( k3b[93], a4_k1a[29], a4_k4a[29] );
xor a4_C898 ( k3b[94], a4_k1a[30], a4_k4a[30] );
xor a4_C897 ( k3b[95], a4_k1a[31], a4_k4a[31] );
xor a5_C896 ( k4b[96], a5_k0a[0], a5_k4a[0] );
xor a5_C895 ( k4b[97], a5_k0a[1], a5_k4a[1] );
xor a5_C894 ( k4b[98], a5_k0a[2], a5_k4a[2] );
xor a5_C893 ( k4b[99], a5_k0a[3], a5_k4a[3] );
xor a5_C892 ( k4b[100], a5_k0a[4], a5_k4a[4] );
xor a5_C891 ( k4b[101], a5_k0a[5], a5_k4a[5] );
xor a5_C890 ( k4b[102], a5_k0a[6], a5_k4a[6] );
xor a5_C889 ( k4b[103], a5_k0a[7], a5_k4a[7] );
xor a5_C888 ( k4b[104], a5_k0a[8], a5_k4a[8] );
xor a5_C887 ( k4b[105], a5_k0a[9], a5_k4a[9] );
xor a5_C886 ( k4b[106], a5_k0a[10], a5_k4a[10] );
xor a5_C885 ( k4b[107], a5_k0a[11], a5_k4a[11] );
xor a5_C884 ( k4b[108], a5_k0a[12], a5_k4a[12] );
xor a5_C883 ( k4b[109], a5_k0a[13], a5_k4a[13] );
xor a5_C882 ( k4b[110], a5_k0a[14], a5_k4a[14] );
xor a5_C881 ( k4b[111], a5_k0a[15], a5_k4a[15] );
xor a5_C880 ( k4b[112], a5_k0a[16], a5_k4a[16] );
xor a5_C879 ( k4b[113], a5_k0a[17], a5_k4a[17] );
xor a5_C878 ( k4b[114], a5_k0a[18], a5_k4a[18] );
xor a5_C877 ( k4b[115], a5_k0a[19], a5_k4a[19] );
xor a5_C876 ( k4b[116], a5_k0a[20], a5_k4a[20] );
xor a5_C875 ( k4b[117], a5_k0a[21], a5_k4a[21] );
xor a5_C874 ( k4b[118], a5_k0a[22], a5_k4a[22] );
xor a5_C873 ( k4b[119], a5_k0a[23], a5_k4a[23] );
xor a5_C872 ( k4b[120], a5_k0a[24], a5_k4a[24] );
xor a5_C871 ( k4b[121], a5_k0a[25], a5_k4a[25] );
xor a5_C870 ( k4b[122], a5_k0a[26], a5_k4a[26] );
xor a5_C869 ( k4b[123], a5_k0a[27], a5_k4a[27] );
xor a5_C868 ( k4b[124], a5_k0a[28], a5_k4a[28] );
xor a5_C867 ( k4b[125], a5_k0a[29], a5_k4a[29] );
xor a5_C866 ( k4b[126], a5_k0a[30], a5_k4a[30] );
xor a5_C865 ( k4b[127], a5_k0a[31], a5_k4a[31] );
xor a5_C992 ( k4b[0], a5_k3a[0], a5_k4a[0] );
xor a5_C991 ( k4b[1], a5_k3a[1], a5_k4a[1] );
xor a5_C990 ( k4b[2], a5_k3a[2], a5_k4a[2] );
xor a5_C989 ( k4b[3], a5_k3a[3], a5_k4a[3] );
xor a5_C988 ( k4b[4], a5_k3a[4], a5_k4a[4] );
xor a5_C987 ( k4b[5], a5_k3a[5], a5_k4a[5] );
xor a5_C986 ( k4b[6], a5_k3a[6], a5_k4a[6] );
xor a5_C985 ( k4b[7], a5_k3a[7], a5_k4a[7] );
xor a5_C984 ( k4b[8], a5_k3a[8], a5_k4a[8] );
xor a5_C983 ( k4b[9], a5_k3a[9], a5_k4a[9] );
xor a5_C982 ( k4b[10], a5_k3a[10], a5_k4a[10] );
xor a5_C981 ( k4b[11], a5_k3a[11], a5_k4a[11] );
xor a5_C980 ( k4b[12], a5_k3a[12], a5_k4a[12] );
xor a5_C979 ( k4b[13], a5_k3a[13], a5_k4a[13] );
xor a5_C978 ( k4b[14], a5_k3a[14], a5_k4a[14] );
xor a5_C977 ( k4b[15], a5_k3a[15], a5_k4a[15] );
xor a5_C976 ( k4b[16], a5_k3a[16], a5_k4a[16] );
xor a5_C975 ( k4b[17], a5_k3a[17], a5_k4a[17] );
xor a5_C974 ( k4b[18], a5_k3a[18], a5_k4a[18] );
xor a5_C973 ( k4b[19], a5_k3a[19], a5_k4a[19] );
xor a5_C972 ( k4b[20], a5_k3a[20], a5_k4a[20] );
xor a5_C971 ( k4b[21], a5_k3a[21], a5_k4a[21] );
xor a5_C970 ( k4b[22], a5_k3a[22], a5_k4a[22] );
xor a5_C969 ( k4b[23], a5_k3a[23], a5_k4a[23] );
xor a5_C968 ( k4b[24], a5_k3a[24], a5_k4a[24] );
xor a5_C967 ( k4b[25], a5_k3a[25], a5_k4a[25] );
xor a5_C966 ( k4b[26], a5_k3a[26], a5_k4a[26] );
xor a5_C965 ( k4b[27], a5_k3a[27], a5_k4a[27] );
xor a5_C964 ( k4b[28], a5_k3a[28], a5_k4a[28] );
xor a5_C963 ( k4b[29], a5_k3a[29], a5_k4a[29] );
xor a5_C962 ( k4b[30], a5_k3a[30], a5_k4a[30] );
xor a5_C960 ( k4b[32], a5_k2a[0], a5_k4a[0] );
xor a5_C959 ( k4b[33], a5_k2a[1], a5_k4a[1] );
xor a5_C958 ( k4b[34], a5_k2a[2], a5_k4a[2] );
xor a5_C957 ( k4b[35], a5_k2a[3], a5_k4a[3] );
xor a5_C956 ( k4b[36], a5_k2a[4], a5_k4a[4] );
xor a5_C955 ( k4b[37], a5_k2a[5], a5_k4a[5] );
xor a5_C954 ( k4b[38], a5_k2a[6], a5_k4a[6] );
xor a5_C953 ( k4b[39], a5_k2a[7], a5_k4a[7] );
xor a5_C952 ( k4b[40], a5_k2a[8], a5_k4a[8] );
xor a5_C951 ( k4b[41], a5_k2a[9], a5_k4a[9] );
xor a5_C950 ( k4b[42], a5_k2a[10], a5_k4a[10] );
xor a5_C949 ( k4b[43], a5_k2a[11], a5_k4a[11] );
xor a5_C948 ( k4b[44], a5_k2a[12], a5_k4a[12] );
xor a5_C947 ( k4b[45], a5_k2a[13], a5_k4a[13] );
xor a5_C946 ( k4b[46], a5_k2a[14], a5_k4a[14] );
xor a5_C945 ( k4b[47], a5_k2a[15], a5_k4a[15] );
xor a5_C944 ( k4b[48], a5_k2a[16], a5_k4a[16] );
xor a5_C943 ( k4b[49], a5_k2a[17], a5_k4a[17] );
xor a5_C942 ( k4b[50], a5_k2a[18], a5_k4a[18] );
xor a5_C941 ( k4b[51], a5_k2a[19], a5_k4a[19] );
xor a5_C940 ( k4b[52], a5_k2a[20], a5_k4a[20] );
xor a5_C939 ( k4b[53], a5_k2a[21], a5_k4a[21] );
xor a5_C938 ( k4b[54], a5_k2a[22], a5_k4a[22] );
xor a5_C937 ( k4b[55], a5_k2a[23], a5_k4a[23] );
xor a5_C936 ( k4b[56], a5_k2a[24], a5_k4a[24] );
xor a5_C935 ( k4b[57], a5_k2a[25], a5_k4a[25] );
xor a5_C934 ( k4b[58], a5_k2a[26], a5_k4a[26] );
xor a5_C933 ( k4b[59], a5_k2a[27], a5_k4a[27] );
xor a5_C932 ( k4b[60], a5_k2a[28], a5_k4a[28] );
xor a5_C931 ( k4b[61], a5_k2a[29], a5_k4a[29] );
xor a5_C930 ( k4b[62], a5_k2a[30], a5_k4a[30] );
xor a5_C929 ( k4b[63], a5_k2a[31], a5_k4a[31] );
xor a5_C928 ( k4b[64], a5_k1a[0], a5_k4a[0] );
xor a5_C927 ( k4b[65], a5_k1a[1], a5_k4a[1] );
xor a5_C926 ( k4b[66], a5_k1a[2], a5_k4a[2] );
xor a5_C925 ( k4b[67], a5_k1a[3], a5_k4a[3] );
xor a5_C924 ( k4b[68], a5_k1a[4], a5_k4a[4] );
xor a5_C923 ( k4b[69], a5_k1a[5], a5_k4a[5] );
xor a5_C922 ( k4b[70], a5_k1a[6], a5_k4a[6] );
xor a5_C921 ( k4b[71], a5_k1a[7], a5_k4a[7] );
xor a5_C920 ( k4b[72], a5_k1a[8], a5_k4a[8] );
xor a5_C919 ( k4b[73], a5_k1a[9], a5_k4a[9] );
xor a5_C918 ( k4b[74], a5_k1a[10], a5_k4a[10] );
xor a5_C917 ( k4b[75], a5_k1a[11], a5_k4a[11] );
xor a5_C916 ( k4b[76], a5_k1a[12], a5_k4a[12] );
xor a5_C915 ( k4b[77], a5_k1a[13], a5_k4a[13] );
xor a5_C914 ( k4b[78], a5_k1a[14], a5_k4a[14] );
xor a5_C913 ( k4b[79], a5_k1a[15], a5_k4a[15] );
xor a5_C912 ( k4b[80], a5_k1a[16], a5_k4a[16] );
xor a5_C911 ( k4b[81], a5_k1a[17], a5_k4a[17] );
xor a5_C910 ( k4b[82], a5_k1a[18], a5_k4a[18] );
xor a5_C909 ( k4b[83], a5_k1a[19], a5_k4a[19] );
xor a5_C908 ( k4b[84], a5_k1a[20], a5_k4a[20] );
xor a5_C907 ( k4b[85], a5_k1a[21], a5_k4a[21] );
xor a5_C906 ( k4b[86], a5_k1a[22], a5_k4a[22] );
xor a5_C905 ( k4b[87], a5_k1a[23], a5_k4a[23] );
xor a5_C904 ( k4b[88], a5_k1a[24], a5_k4a[24] );
xor a5_C903 ( k4b[89], a5_k1a[25], a5_k4a[25] );
xor a5_C902 ( k4b[90], a5_k1a[26], a5_k4a[26] );
xor a5_C901 ( k4b[91], a5_k1a[27], a5_k4a[27] );
xor a5_C900 ( k4b[92], a5_k1a[28], a5_k4a[28] );
xor a5_C899 ( k4b[93], a5_k1a[29], a5_k4a[29] );
xor a5_C898 ( k4b[94], a5_k1a[30], a5_k4a[30] );
xor a5_C897 ( k4b[95], a5_k1a[31], a5_k4a[31] );
xor a6_C896 ( k5b[96], a6_k0a[0], a6_k4a[0] );
xor a6_C895 ( k5b[97], a6_k0a[1], a6_k4a[1] );
xor a6_C894 ( k5b[98], a6_k0a[2], a6_k4a[2] );
xor a6_C893 ( k5b[99], a6_k0a[3], a6_k4a[3] );
xor a6_C892 ( k5b[100], a6_k0a[4], a6_k4a[4] );
xor a6_C891 ( k5b[101], a6_k0a[5], a6_k4a[5] );
xor a6_C890 ( k5b[102], a6_k0a[6], a6_k4a[6] );
xor a6_C889 ( k5b[103], a6_k0a[7], a6_k4a[7] );
xor a6_C888 ( k5b[104], a6_k0a[8], a6_k4a[8] );
xor a6_C887 ( k5b[105], a6_k0a[9], a6_k4a[9] );
xor a6_C886 ( k5b[106], a6_k0a[10], a6_k4a[10] );
xor a6_C885 ( k5b[107], a6_k0a[11], a6_k4a[11] );
xor a6_C884 ( k5b[108], a6_k0a[12], a6_k4a[12] );
xor a6_C883 ( k5b[109], a6_k0a[13], a6_k4a[13] );
xor a6_C882 ( k5b[110], a6_k0a[14], a6_k4a[14] );
xor a6_C881 ( k5b[111], a6_k0a[15], a6_k4a[15] );
xor a6_C880 ( k5b[112], a6_k0a[16], a6_k4a[16] );
xor a6_C879 ( k5b[113], a6_k0a[17], a6_k4a[17] );
xor a6_C878 ( k5b[114], a6_k0a[18], a6_k4a[18] );
xor a6_C877 ( k5b[115], a6_k0a[19], a6_k4a[19] );
xor a6_C876 ( k5b[116], a6_k0a[20], a6_k4a[20] );
xor a6_C875 ( k5b[117], a6_k0a[21], a6_k4a[21] );
xor a6_C874 ( k5b[118], a6_k0a[22], a6_k4a[22] );
xor a6_C873 ( k5b[119], a6_k0a[23], a6_k4a[23] );
xor a6_C872 ( k5b[120], a6_k0a[24], a6_k4a[24] );
xor a6_C871 ( k5b[121], a6_k0a[25], a6_k4a[25] );
xor a6_C870 ( k5b[122], a6_k0a[26], a6_k4a[26] );
xor a6_C869 ( k5b[123], a6_k0a[27], a6_k4a[27] );
xor a6_C868 ( k5b[124], a6_k0a[28], a6_k4a[28] );
xor a6_C867 ( k5b[125], a6_k0a[29], a6_k4a[29] );
xor a6_C866 ( k5b[126], a6_k0a[30], a6_k4a[30] );
xor a6_C865 ( k5b[127], a6_k0a[31], a6_k4a[31] );
xor a6_C992 ( k5b[0], a6_k3a[0], a6_k4a[0] );
xor a6_C991 ( k5b[1], a6_k3a[1], a6_k4a[1] );
xor a6_C990 ( k5b[2], a6_k3a[2], a6_k4a[2] );
xor a6_C989 ( k5b[3], a6_k3a[3], a6_k4a[3] );
xor a6_C988 ( k5b[4], a6_k3a[4], a6_k4a[4] );
xor a6_C987 ( k5b[5], a6_k3a[5], a6_k4a[5] );
xor a6_C986 ( k5b[6], a6_k3a[6], a6_k4a[6] );
xor a6_C985 ( k5b[7], a6_k3a[7], a6_k4a[7] );
xor a6_C984 ( k5b[8], a6_k3a[8], a6_k4a[8] );
xor a6_C983 ( k5b[9], a6_k3a[9], a6_k4a[9] );
xor a6_C982 ( k5b[10], a6_k3a[10], a6_k4a[10] );
xor a6_C981 ( k5b[11], a6_k3a[11], a6_k4a[11] );
xor a6_C980 ( k5b[12], a6_k3a[12], a6_k4a[12] );
xor a6_C979 ( k5b[13], a6_k3a[13], a6_k4a[13] );
xor a6_C978 ( k5b[14], a6_k3a[14], a6_k4a[14] );
xor a6_C977 ( k5b[15], a6_k3a[15], a6_k4a[15] );
xor a6_C976 ( k5b[16], a6_k3a[16], a6_k4a[16] );
xor a6_C975 ( k5b[17], a6_k3a[17], a6_k4a[17] );
xor a6_C974 ( k5b[18], a6_k3a[18], a6_k4a[18] );
xor a6_C973 ( k5b[19], a6_k3a[19], a6_k4a[19] );
xor a6_C972 ( k5b[20], a6_k3a[20], a6_k4a[20] );
xor a6_C971 ( k5b[21], a6_k3a[21], a6_k4a[21] );
xor a6_C970 ( k5b[22], a6_k3a[22], a6_k4a[22] );
xor a6_C969 ( k5b[23], a6_k3a[23], a6_k4a[23] );
xor a6_C968 ( k5b[24], a6_k3a[24], a6_k4a[24] );
xor a6_C967 ( k5b[25], a6_k3a[25], a6_k4a[25] );
xor a6_C966 ( k5b[26], a6_k3a[26], a6_k4a[26] );
xor a6_C965 ( k5b[27], a6_k3a[27], a6_k4a[27] );
xor a6_C964 ( k5b[28], a6_k3a[28], a6_k4a[28] );
xor a6_C963 ( k5b[29], a6_k3a[29], a6_k4a[29] );
xor a6_C962 ( k5b[30], a6_k3a[30], a6_k4a[30] );
xor a6_C960 ( k5b[32], a6_k2a[0], a6_k4a[0] );
xor a6_C959 ( k5b[33], a6_k2a[1], a6_k4a[1] );
xor a6_C958 ( k5b[34], a6_k2a[2], a6_k4a[2] );
xor a6_C957 ( k5b[35], a6_k2a[3], a6_k4a[3] );
xor a6_C956 ( k5b[36], a6_k2a[4], a6_k4a[4] );
xor a6_C955 ( k5b[37], a6_k2a[5], a6_k4a[5] );
xor a6_C954 ( k5b[38], a6_k2a[6], a6_k4a[6] );
xor a6_C953 ( k5b[39], a6_k2a[7], a6_k4a[7] );
xor a6_C952 ( k5b[40], a6_k2a[8], a6_k4a[8] );
xor a6_C951 ( k5b[41], a6_k2a[9], a6_k4a[9] );
xor a6_C950 ( k5b[42], a6_k2a[10], a6_k4a[10] );
xor a6_C949 ( k5b[43], a6_k2a[11], a6_k4a[11] );
xor a6_C948 ( k5b[44], a6_k2a[12], a6_k4a[12] );
xor a6_C947 ( k5b[45], a6_k2a[13], a6_k4a[13] );
xor a6_C946 ( k5b[46], a6_k2a[14], a6_k4a[14] );
xor a6_C945 ( k5b[47], a6_k2a[15], a6_k4a[15] );
xor a6_C944 ( k5b[48], a6_k2a[16], a6_k4a[16] );
xor a6_C943 ( k5b[49], a6_k2a[17], a6_k4a[17] );
xor a6_C942 ( k5b[50], a6_k2a[18], a6_k4a[18] );
xor a6_C941 ( k5b[51], a6_k2a[19], a6_k4a[19] );
xor a6_C940 ( k5b[52], a6_k2a[20], a6_k4a[20] );
xor a6_C939 ( k5b[53], a6_k2a[21], a6_k4a[21] );
xor a6_C938 ( k5b[54], a6_k2a[22], a6_k4a[22] );
xor a6_C937 ( k5b[55], a6_k2a[23], a6_k4a[23] );
xor a6_C936 ( k5b[56], a6_k2a[24], a6_k4a[24] );
xor a6_C935 ( k5b[57], a6_k2a[25], a6_k4a[25] );
xor a6_C934 ( k5b[58], a6_k2a[26], a6_k4a[26] );
xor a6_C933 ( k5b[59], a6_k2a[27], a6_k4a[27] );
xor a6_C932 ( k5b[60], a6_k2a[28], a6_k4a[28] );
xor a6_C931 ( k5b[61], a6_k2a[29], a6_k4a[29] );
xor a6_C930 ( k5b[62], a6_k2a[30], a6_k4a[30] );
xor a6_C929 ( k5b[63], a6_k2a[31], a6_k4a[31] );
xor a6_C928 ( k5b[64], a6_k1a[0], a6_k4a[0] );
xor a6_C927 ( k5b[65], a6_k1a[1], a6_k4a[1] );
xor a6_C926 ( k5b[66], a6_k1a[2], a6_k4a[2] );
xor a6_C925 ( k5b[67], a6_k1a[3], a6_k4a[3] );
xor a6_C924 ( k5b[68], a6_k1a[4], a6_k4a[4] );
xor a6_C923 ( k5b[69], a6_k1a[5], a6_k4a[5] );
xor a6_C922 ( k5b[70], a6_k1a[6], a6_k4a[6] );
xor a6_C921 ( k5b[71], a6_k1a[7], a6_k4a[7] );
xor a6_C920 ( k5b[72], a6_k1a[8], a6_k4a[8] );
xor a6_C919 ( k5b[73], a6_k1a[9], a6_k4a[9] );
xor a6_C918 ( k5b[74], a6_k1a[10], a6_k4a[10] );
xor a6_C917 ( k5b[75], a6_k1a[11], a6_k4a[11] );
xor a6_C916 ( k5b[76], a6_k1a[12], a6_k4a[12] );
xor a6_C915 ( k5b[77], a6_k1a[13], a6_k4a[13] );
xor a6_C914 ( k5b[78], a6_k1a[14], a6_k4a[14] );
xor a6_C913 ( k5b[79], a6_k1a[15], a6_k4a[15] );
xor a6_C912 ( k5b[80], a6_k1a[16], a6_k4a[16] );
xor a6_C911 ( k5b[81], a6_k1a[17], a6_k4a[17] );
xor a6_C910 ( k5b[82], a6_k1a[18], a6_k4a[18] );
xor a6_C909 ( k5b[83], a6_k1a[19], a6_k4a[19] );
xor a6_C908 ( k5b[84], a6_k1a[20], a6_k4a[20] );
xor a6_C907 ( k5b[85], a6_k1a[21], a6_k4a[21] );
xor a6_C906 ( k5b[86], a6_k1a[22], a6_k4a[22] );
xor a6_C905 ( k5b[87], a6_k1a[23], a6_k4a[23] );
xor a6_C904 ( k5b[88], a6_k1a[24], a6_k4a[24] );
xor a6_C903 ( k5b[89], a6_k1a[25], a6_k4a[25] );
xor a6_C902 ( k5b[90], a6_k1a[26], a6_k4a[26] );
xor a6_C901 ( k5b[91], a6_k1a[27], a6_k4a[27] );
xor a6_C900 ( k5b[92], a6_k1a[28], a6_k4a[28] );
xor a6_C899 ( k5b[93], a6_k1a[29], a6_k4a[29] );
xor a6_C898 ( k5b[94], a6_k1a[30], a6_k4a[30] );
xor a6_C897 ( k5b[95], a6_k1a[31], a6_k4a[31] );
xor a7_C896 ( k6b[96], a7_k0a[0], a7_k4a[0] );
xor a7_C895 ( k6b[97], a7_k0a[1], a7_k4a[1] );
xor a7_C894 ( k6b[98], a7_k0a[2], a7_k4a[2] );
xor a7_C893 ( k6b[99], a7_k0a[3], a7_k4a[3] );
xor a7_C892 ( k6b[100], a7_k0a[4], a7_k4a[4] );
xor a7_C891 ( k6b[101], a7_k0a[5], a7_k4a[5] );
xor a7_C890 ( k6b[102], a7_k0a[6], a7_k4a[6] );
xor a7_C889 ( k6b[103], a7_k0a[7], a7_k4a[7] );
xor a7_C888 ( k6b[104], a7_k0a[8], a7_k4a[8] );
xor a7_C887 ( k6b[105], a7_k0a[9], a7_k4a[9] );
xor a7_C886 ( k6b[106], a7_k0a[10], a7_k4a[10] );
xor a7_C885 ( k6b[107], a7_k0a[11], a7_k4a[11] );
xor a7_C884 ( k6b[108], a7_k0a[12], a7_k4a[12] );
xor a7_C883 ( k6b[109], a7_k0a[13], a7_k4a[13] );
xor a7_C882 ( k6b[110], a7_k0a[14], a7_k4a[14] );
xor a7_C881 ( k6b[111], a7_k0a[15], a7_k4a[15] );
xor a7_C880 ( k6b[112], a7_k0a[16], a7_k4a[16] );
xor a7_C879 ( k6b[113], a7_k0a[17], a7_k4a[17] );
xor a7_C878 ( k6b[114], a7_k0a[18], a7_k4a[18] );
xor a7_C877 ( k6b[115], a7_k0a[19], a7_k4a[19] );
xor a7_C876 ( k6b[116], a7_k0a[20], a7_k4a[20] );
xor a7_C875 ( k6b[117], a7_k0a[21], a7_k4a[21] );
xor a7_C874 ( k6b[118], a7_k0a[22], a7_k4a[22] );
xor a7_C873 ( k6b[119], a7_k0a[23], a7_k4a[23] );
xor a7_C872 ( k6b[120], a7_k0a[24], a7_k4a[24] );
xor a7_C871 ( k6b[121], a7_k0a[25], a7_k4a[25] );
xor a7_C870 ( k6b[122], a7_k0a[26], a7_k4a[26] );
xor a7_C869 ( k6b[123], a7_k0a[27], a7_k4a[27] );
xor a7_C868 ( k6b[124], a7_k0a[28], a7_k4a[28] );
xor a7_C867 ( k6b[125], a7_k0a[29], a7_k4a[29] );
xor a7_C866 ( k6b[126], a7_k0a[30], a7_k4a[30] );
xor a7_C865 ( k6b[127], a7_k0a[31], a7_k4a[31] );
xor a7_C992 ( k6b[0], a7_k3a[0], a7_k4a[0] );
xor a7_C991 ( k6b[1], a7_k3a[1], a7_k4a[1] );
xor a7_C990 ( k6b[2], a7_k3a[2], a7_k4a[2] );
xor a7_C989 ( k6b[3], a7_k3a[3], a7_k4a[3] );
xor a7_C988 ( k6b[4], a7_k3a[4], a7_k4a[4] );
xor a7_C987 ( k6b[5], a7_k3a[5], a7_k4a[5] );
xor a7_C986 ( k6b[6], a7_k3a[6], a7_k4a[6] );
xor a7_C985 ( k6b[7], a7_k3a[7], a7_k4a[7] );
xor a7_C984 ( k6b[8], a7_k3a[8], a7_k4a[8] );
xor a7_C983 ( k6b[9], a7_k3a[9], a7_k4a[9] );
xor a7_C982 ( k6b[10], a7_k3a[10], a7_k4a[10] );
xor a7_C981 ( k6b[11], a7_k3a[11], a7_k4a[11] );
xor a7_C980 ( k6b[12], a7_k3a[12], a7_k4a[12] );
xor a7_C979 ( k6b[13], a7_k3a[13], a7_k4a[13] );
xor a7_C978 ( k6b[14], a7_k3a[14], a7_k4a[14] );
xor a7_C977 ( k6b[15], a7_k3a[15], a7_k4a[15] );
xor a7_C976 ( k6b[16], a7_k3a[16], a7_k4a[16] );
xor a7_C975 ( k6b[17], a7_k3a[17], a7_k4a[17] );
xor a7_C974 ( k6b[18], a7_k3a[18], a7_k4a[18] );
xor a7_C973 ( k6b[19], a7_k3a[19], a7_k4a[19] );
xor a7_C972 ( k6b[20], a7_k3a[20], a7_k4a[20] );
xor a7_C971 ( k6b[21], a7_k3a[21], a7_k4a[21] );
xor a7_C970 ( k6b[22], a7_k3a[22], a7_k4a[22] );
xor a7_C969 ( k6b[23], a7_k3a[23], a7_k4a[23] );
xor a7_C968 ( k6b[24], a7_k3a[24], a7_k4a[24] );
xor a7_C967 ( k6b[25], a7_k3a[25], a7_k4a[25] );
xor a7_C966 ( k6b[26], a7_k3a[26], a7_k4a[26] );
xor a7_C965 ( k6b[27], a7_k3a[27], a7_k4a[27] );
xor a7_C964 ( k6b[28], a7_k3a[28], a7_k4a[28] );
xor a7_C963 ( k6b[29], a7_k3a[29], a7_k4a[29] );
xor a7_C962 ( k6b[30], a7_k3a[30], a7_k4a[30] );
xor a7_C960 ( k6b[32], a7_k2a[0], a7_k4a[0] );
xor a7_C959 ( k6b[33], a7_k2a[1], a7_k4a[1] );
xor a7_C958 ( k6b[34], a7_k2a[2], a7_k4a[2] );
xor a7_C957 ( k6b[35], a7_k2a[3], a7_k4a[3] );
xor a7_C956 ( k6b[36], a7_k2a[4], a7_k4a[4] );
xor a7_C955 ( k6b[37], a7_k2a[5], a7_k4a[5] );
xor a7_C954 ( k6b[38], a7_k2a[6], a7_k4a[6] );
xor a7_C953 ( k6b[39], a7_k2a[7], a7_k4a[7] );
xor a7_C952 ( k6b[40], a7_k2a[8], a7_k4a[8] );
xor a7_C951 ( k6b[41], a7_k2a[9], a7_k4a[9] );
xor a7_C950 ( k6b[42], a7_k2a[10], a7_k4a[10] );
xor a7_C949 ( k6b[43], a7_k2a[11], a7_k4a[11] );
xor a7_C948 ( k6b[44], a7_k2a[12], a7_k4a[12] );
xor a7_C947 ( k6b[45], a7_k2a[13], a7_k4a[13] );
xor a7_C946 ( k6b[46], a7_k2a[14], a7_k4a[14] );
xor a7_C945 ( k6b[47], a7_k2a[15], a7_k4a[15] );
xor a7_C944 ( k6b[48], a7_k2a[16], a7_k4a[16] );
xor a7_C943 ( k6b[49], a7_k2a[17], a7_k4a[17] );
xor a7_C942 ( k6b[50], a7_k2a[18], a7_k4a[18] );
xor a7_C941 ( k6b[51], a7_k2a[19], a7_k4a[19] );
xor a7_C940 ( k6b[52], a7_k2a[20], a7_k4a[20] );
xor a7_C939 ( k6b[53], a7_k2a[21], a7_k4a[21] );
xor a7_C938 ( k6b[54], a7_k2a[22], a7_k4a[22] );
xor a7_C937 ( k6b[55], a7_k2a[23], a7_k4a[23] );
xor a7_C936 ( k6b[56], a7_k2a[24], a7_k4a[24] );
xor a7_C935 ( k6b[57], a7_k2a[25], a7_k4a[25] );
xor a7_C934 ( k6b[58], a7_k2a[26], a7_k4a[26] );
xor a7_C933 ( k6b[59], a7_k2a[27], a7_k4a[27] );
xor a7_C932 ( k6b[60], a7_k2a[28], a7_k4a[28] );
xor a7_C931 ( k6b[61], a7_k2a[29], a7_k4a[29] );
xor a7_C930 ( k6b[62], a7_k2a[30], a7_k4a[30] );
xor a7_C929 ( k6b[63], a7_k2a[31], a7_k4a[31] );
xor a7_C928 ( k6b[64], a7_k1a[0], a7_k4a[0] );
xor a7_C927 ( k6b[65], a7_k1a[1], a7_k4a[1] );
xor a7_C926 ( k6b[66], a7_k1a[2], a7_k4a[2] );
xor a7_C925 ( k6b[67], a7_k1a[3], a7_k4a[3] );
xor a7_C924 ( k6b[68], a7_k1a[4], a7_k4a[4] );
xor a7_C923 ( k6b[69], a7_k1a[5], a7_k4a[5] );
xor a7_C922 ( k6b[70], a7_k1a[6], a7_k4a[6] );
xor a7_C921 ( k6b[71], a7_k1a[7], a7_k4a[7] );
xor a7_C920 ( k6b[72], a7_k1a[8], a7_k4a[8] );
xor a7_C919 ( k6b[73], a7_k1a[9], a7_k4a[9] );
xor a7_C918 ( k6b[74], a7_k1a[10], a7_k4a[10] );
xor a7_C917 ( k6b[75], a7_k1a[11], a7_k4a[11] );
xor a7_C916 ( k6b[76], a7_k1a[12], a7_k4a[12] );
xor a7_C915 ( k6b[77], a7_k1a[13], a7_k4a[13] );
xor a7_C914 ( k6b[78], a7_k1a[14], a7_k4a[14] );
xor a7_C913 ( k6b[79], a7_k1a[15], a7_k4a[15] );
xor a7_C912 ( k6b[80], a7_k1a[16], a7_k4a[16] );
xor a7_C911 ( k6b[81], a7_k1a[17], a7_k4a[17] );
xor a7_C910 ( k6b[82], a7_k1a[18], a7_k4a[18] );
xor a7_C909 ( k6b[83], a7_k1a[19], a7_k4a[19] );
xor a7_C908 ( k6b[84], a7_k1a[20], a7_k4a[20] );
xor a7_C907 ( k6b[85], a7_k1a[21], a7_k4a[21] );
xor a7_C906 ( k6b[86], a7_k1a[22], a7_k4a[22] );
xor a7_C905 ( k6b[87], a7_k1a[23], a7_k4a[23] );
xor a7_C904 ( k6b[88], a7_k1a[24], a7_k4a[24] );
xor a7_C903 ( k6b[89], a7_k1a[25], a7_k4a[25] );
xor a7_C902 ( k6b[90], a7_k1a[26], a7_k4a[26] );
xor a7_C901 ( k6b[91], a7_k1a[27], a7_k4a[27] );
xor a7_C900 ( k6b[92], a7_k1a[28], a7_k4a[28] );
xor a7_C899 ( k6b[93], a7_k1a[29], a7_k4a[29] );
xor a7_C898 ( k6b[94], a7_k1a[30], a7_k4a[30] );
xor a7_C897 ( k6b[95], a7_k1a[31], a7_k4a[31] );
xor a8_C896 ( k7b[96], a8_k0a[0], a8_k4a[0] );
xor a8_C895 ( k7b[97], a8_k0a[1], a8_k4a[1] );
xor a8_C894 ( k7b[98], a8_k0a[2], a8_k4a[2] );
xor a8_C893 ( k7b[99], a8_k0a[3], a8_k4a[3] );
xor a8_C892 ( k7b[100], a8_k0a[4], a8_k4a[4] );
xor a8_C891 ( k7b[101], a8_k0a[5], a8_k4a[5] );
xor a8_C890 ( k7b[102], a8_k0a[6], a8_k4a[6] );
xor a8_C889 ( k7b[103], a8_k0a[7], a8_k4a[7] );
xor a8_C888 ( k7b[104], a8_k0a[8], a8_k4a[8] );
xor a8_C887 ( k7b[105], a8_k0a[9], a8_k4a[9] );
xor a8_C886 ( k7b[106], a8_k0a[10], a8_k4a[10] );
xor a8_C885 ( k7b[107], a8_k0a[11], a8_k4a[11] );
xor a8_C884 ( k7b[108], a8_k0a[12], a8_k4a[12] );
xor a8_C883 ( k7b[109], a8_k0a[13], a8_k4a[13] );
xor a8_C882 ( k7b[110], a8_k0a[14], a8_k4a[14] );
xor a8_C881 ( k7b[111], a8_k0a[15], a8_k4a[15] );
xor a8_C880 ( k7b[112], a8_k0a[16], a8_k4a[16] );
xor a8_C879 ( k7b[113], a8_k0a[17], a8_k4a[17] );
xor a8_C878 ( k7b[114], a8_k0a[18], a8_k4a[18] );
xor a8_C877 ( k7b[115], a8_k0a[19], a8_k4a[19] );
xor a8_C876 ( k7b[116], a8_k0a[20], a8_k4a[20] );
xor a8_C875 ( k7b[117], a8_k0a[21], a8_k4a[21] );
xor a8_C874 ( k7b[118], a8_k0a[22], a8_k4a[22] );
xor a8_C873 ( k7b[119], a8_k0a[23], a8_k4a[23] );
xor a8_C872 ( k7b[120], a8_k0a[24], a8_k4a[24] );
xor a8_C871 ( k7b[121], a8_k0a[25], a8_k4a[25] );
xor a8_C870 ( k7b[122], a8_k0a[26], a8_k4a[26] );
xor a8_C869 ( k7b[123], a8_k0a[27], a8_k4a[27] );
xor a8_C868 ( k7b[124], a8_k0a[28], a8_k4a[28] );
xor a8_C867 ( k7b[125], a8_k0a[29], a8_k4a[29] );
xor a8_C866 ( k7b[126], a8_k0a[30], a8_k4a[30] );
xor a8_C865 ( k7b[127], a8_k0a[31], a8_k4a[31] );
xor a8_C992 ( k7b[0], a8_k3a[0], a8_k4a[0] );
xor a8_C991 ( k7b[1], a8_k3a[1], a8_k4a[1] );
xor a8_C990 ( k7b[2], a8_k3a[2], a8_k4a[2] );
xor a8_C989 ( k7b[3], a8_k3a[3], a8_k4a[3] );
xor a8_C988 ( k7b[4], a8_k3a[4], a8_k4a[4] );
xor a8_C987 ( k7b[5], a8_k3a[5], a8_k4a[5] );
xor a8_C986 ( k7b[6], a8_k3a[6], a8_k4a[6] );
xor a8_C985 ( k7b[7], a8_k3a[7], a8_k4a[7] );
xor a8_C984 ( k7b[8], a8_k3a[8], a8_k4a[8] );
xor a8_C983 ( k7b[9], a8_k3a[9], a8_k4a[9] );
xor a8_C982 ( k7b[10], a8_k3a[10], a8_k4a[10] );
xor a8_C981 ( k7b[11], a8_k3a[11], a8_k4a[11] );
xor a8_C980 ( k7b[12], a8_k3a[12], a8_k4a[12] );
xor a8_C979 ( k7b[13], a8_k3a[13], a8_k4a[13] );
xor a8_C978 ( k7b[14], a8_k3a[14], a8_k4a[14] );
xor a8_C977 ( k7b[15], a8_k3a[15], a8_k4a[15] );
xor a8_C976 ( k7b[16], a8_k3a[16], a8_k4a[16] );
xor a8_C975 ( k7b[17], a8_k3a[17], a8_k4a[17] );
xor a8_C974 ( k7b[18], a8_k3a[18], a8_k4a[18] );
xor a8_C973 ( k7b[19], a8_k3a[19], a8_k4a[19] );
xor a8_C972 ( k7b[20], a8_k3a[20], a8_k4a[20] );
xor a8_C971 ( k7b[21], a8_k3a[21], a8_k4a[21] );
xor a8_C970 ( k7b[22], a8_k3a[22], a8_k4a[22] );
xor a8_C969 ( k7b[23], a8_k3a[23], a8_k4a[23] );
xor a8_C968 ( k7b[24], a8_k3a[24], a8_k4a[24] );
xor a8_C967 ( k7b[25], a8_k3a[25], a8_k4a[25] );
xor a8_C966 ( k7b[26], a8_k3a[26], a8_k4a[26] );
xor a8_C965 ( k7b[27], a8_k3a[27], a8_k4a[27] );
xor a8_C964 ( k7b[28], a8_k3a[28], a8_k4a[28] );
xor a8_C963 ( k7b[29], a8_k3a[29], a8_k4a[29] );
xor a8_C962 ( k7b[30], a8_k3a[30], a8_k4a[30] );
xor a8_C960 ( k7b[32], a8_k2a[0], a8_k4a[0] );
xor a8_C959 ( k7b[33], a8_k2a[1], a8_k4a[1] );
xor a8_C958 ( k7b[34], a8_k2a[2], a8_k4a[2] );
xor a8_C957 ( k7b[35], a8_k2a[3], a8_k4a[3] );
xor a8_C956 ( k7b[36], a8_k2a[4], a8_k4a[4] );
xor a8_C955 ( k7b[37], a8_k2a[5], a8_k4a[5] );
xor a8_C954 ( k7b[38], a8_k2a[6], a8_k4a[6] );
xor a8_C953 ( k7b[39], a8_k2a[7], a8_k4a[7] );
xor a8_C952 ( k7b[40], a8_k2a[8], a8_k4a[8] );
xor a8_C951 ( k7b[41], a8_k2a[9], a8_k4a[9] );
xor a8_C950 ( k7b[42], a8_k2a[10], a8_k4a[10] );
xor a8_C949 ( k7b[43], a8_k2a[11], a8_k4a[11] );
xor a8_C948 ( k7b[44], a8_k2a[12], a8_k4a[12] );
xor a8_C947 ( k7b[45], a8_k2a[13], a8_k4a[13] );
xor a8_C946 ( k7b[46], a8_k2a[14], a8_k4a[14] );
xor a8_C945 ( k7b[47], a8_k2a[15], a8_k4a[15] );
xor a8_C944 ( k7b[48], a8_k2a[16], a8_k4a[16] );
xor a8_C943 ( k7b[49], a8_k2a[17], a8_k4a[17] );
xor a8_C942 ( k7b[50], a8_k2a[18], a8_k4a[18] );
xor a8_C941 ( k7b[51], a8_k2a[19], a8_k4a[19] );
xor a8_C940 ( k7b[52], a8_k2a[20], a8_k4a[20] );
xor a8_C939 ( k7b[53], a8_k2a[21], a8_k4a[21] );
xor a8_C938 ( k7b[54], a8_k2a[22], a8_k4a[22] );
xor a8_C937 ( k7b[55], a8_k2a[23], a8_k4a[23] );
xor a8_C936 ( k7b[56], a8_k2a[24], a8_k4a[24] );
xor a8_C935 ( k7b[57], a8_k2a[25], a8_k4a[25] );
xor a8_C934 ( k7b[58], a8_k2a[26], a8_k4a[26] );
xor a8_C933 ( k7b[59], a8_k2a[27], a8_k4a[27] );
xor a8_C932 ( k7b[60], a8_k2a[28], a8_k4a[28] );
xor a8_C931 ( k7b[61], a8_k2a[29], a8_k4a[29] );
xor a8_C930 ( k7b[62], a8_k2a[30], a8_k4a[30] );
xor a8_C929 ( k7b[63], a8_k2a[31], a8_k4a[31] );
xor a8_C928 ( k7b[64], a8_k1a[0], a8_k4a[0] );
xor a8_C927 ( k7b[65], a8_k1a[1], a8_k4a[1] );
xor a8_C926 ( k7b[66], a8_k1a[2], a8_k4a[2] );
xor a8_C925 ( k7b[67], a8_k1a[3], a8_k4a[3] );
xor a8_C924 ( k7b[68], a8_k1a[4], a8_k4a[4] );
xor a8_C923 ( k7b[69], a8_k1a[5], a8_k4a[5] );
xor a8_C922 ( k7b[70], a8_k1a[6], a8_k4a[6] );
xor a8_C921 ( k7b[71], a8_k1a[7], a8_k4a[7] );
xor a8_C920 ( k7b[72], a8_k1a[8], a8_k4a[8] );
xor a8_C919 ( k7b[73], a8_k1a[9], a8_k4a[9] );
xor a8_C918 ( k7b[74], a8_k1a[10], a8_k4a[10] );
xor a8_C917 ( k7b[75], a8_k1a[11], a8_k4a[11] );
xor a8_C916 ( k7b[76], a8_k1a[12], a8_k4a[12] );
xor a8_C915 ( k7b[77], a8_k1a[13], a8_k4a[13] );
xor a8_C914 ( k7b[78], a8_k1a[14], a8_k4a[14] );
xor a8_C913 ( k7b[79], a8_k1a[15], a8_k4a[15] );
xor a8_C912 ( k7b[80], a8_k1a[16], a8_k4a[16] );
xor a8_C911 ( k7b[81], a8_k1a[17], a8_k4a[17] );
xor a8_C910 ( k7b[82], a8_k1a[18], a8_k4a[18] );
xor a8_C909 ( k7b[83], a8_k1a[19], a8_k4a[19] );
xor a8_C908 ( k7b[84], a8_k1a[20], a8_k4a[20] );
xor a8_C907 ( k7b[85], a8_k1a[21], a8_k4a[21] );
xor a8_C906 ( k7b[86], a8_k1a[22], a8_k4a[22] );
xor a8_C905 ( k7b[87], a8_k1a[23], a8_k4a[23] );
xor a8_C904 ( k7b[88], a8_k1a[24], a8_k4a[24] );
xor a8_C903 ( k7b[89], a8_k1a[25], a8_k4a[25] );
xor a8_C902 ( k7b[90], a8_k1a[26], a8_k4a[26] );
xor a8_C901 ( k7b[91], a8_k1a[27], a8_k4a[27] );
xor a8_C900 ( k7b[92], a8_k1a[28], a8_k4a[28] );
xor a8_C899 ( k7b[93], a8_k1a[29], a8_k4a[29] );
xor a8_C898 ( k7b[94], a8_k1a[30], a8_k4a[30] );
xor a8_C897 ( k7b[95], a8_k1a[31], a8_k4a[31] );
xor a9_C896 ( k8b[96], a9_k0a[0], a9_k4a[0] );
xor a9_C895 ( k8b[97], a9_k0a[1], a9_k4a[1] );
xor a9_C894 ( k8b[98], a9_k0a[2], a9_k4a[2] );
xor a9_C893 ( k8b[99], a9_k0a[3], a9_k4a[3] );
xor a9_C892 ( k8b[100], a9_k0a[4], a9_k4a[4] );
xor a9_C891 ( k8b[101], a9_k0a[5], a9_k4a[5] );
xor a9_C890 ( k8b[102], a9_k0a[6], a9_k4a[6] );
xor a9_C889 ( k8b[103], a9_k0a[7], a9_k4a[7] );
xor a9_C888 ( k8b[104], a9_k0a[8], a9_k4a[8] );
xor a9_C887 ( k8b[105], a9_k0a[9], a9_k4a[9] );
xor a9_C886 ( k8b[106], a9_k0a[10], a9_k4a[10] );
xor a9_C885 ( k8b[107], a9_k0a[11], a9_k4a[11] );
xor a9_C884 ( k8b[108], a9_k0a[12], a9_k4a[12] );
xor a9_C883 ( k8b[109], a9_k0a[13], a9_k4a[13] );
xor a9_C882 ( k8b[110], a9_k0a[14], a9_k4a[14] );
xor a9_C881 ( k8b[111], a9_k0a[15], a9_k4a[15] );
xor a9_C880 ( k8b[112], a9_k0a[16], a9_k4a[16] );
xor a9_C879 ( k8b[113], a9_k0a[17], a9_k4a[17] );
xor a9_C878 ( k8b[114], a9_k0a[18], a9_k4a[18] );
xor a9_C877 ( k8b[115], a9_k0a[19], a9_k4a[19] );
xor a9_C876 ( k8b[116], a9_k0a[20], a9_k4a[20] );
xor a9_C875 ( k8b[117], a9_k0a[21], a9_k4a[21] );
xor a9_C874 ( k8b[118], a9_k0a[22], a9_k4a[22] );
xor a9_C873 ( k8b[119], a9_k0a[23], a9_k4a[23] );
xor a9_C872 ( k8b[120], a9_k0a[24], a9_k4a[24] );
xor a9_C871 ( k8b[121], a9_k0a[25], a9_k4a[25] );
xor a9_C870 ( k8b[122], a9_k0a[26], a9_k4a[26] );
xor a9_C869 ( k8b[123], a9_k0a[27], a9_k4a[27] );
xor a9_C868 ( k8b[124], a9_k0a[28], a9_k4a[28] );
xor a9_C867 ( k8b[125], a9_k0a[29], a9_k4a[29] );
xor a9_C866 ( k8b[126], a9_k0a[30], a9_k4a[30] );
xor a9_C865 ( k8b[127], a9_k0a[31], a9_k4a[31] );
xor a9_C992 ( k8b[0], a9_k3a[0], a9_k4a[0] );
xor a9_C991 ( k8b[1], a9_k3a[1], a9_k4a[1] );
xor a9_C990 ( k8b[2], a9_k3a[2], a9_k4a[2] );
xor a9_C989 ( k8b[3], a9_k3a[3], a9_k4a[3] );
xor a9_C988 ( k8b[4], a9_k3a[4], a9_k4a[4] );
xor a9_C987 ( k8b[5], a9_k3a[5], a9_k4a[5] );
xor a9_C986 ( k8b[6], a9_k3a[6], a9_k4a[6] );
xor a9_C985 ( k8b[7], a9_k3a[7], a9_k4a[7] );
xor a9_C984 ( k8b[8], a9_k3a[8], a9_k4a[8] );
xor a9_C983 ( k8b[9], a9_k3a[9], a9_k4a[9] );
xor a9_C982 ( k8b[10], a9_k3a[10], a9_k4a[10] );
xor a9_C981 ( k8b[11], a9_k3a[11], a9_k4a[11] );
xor a9_C980 ( k8b[12], a9_k3a[12], a9_k4a[12] );
xor a9_C979 ( k8b[13], a9_k3a[13], a9_k4a[13] );
xor a9_C978 ( k8b[14], a9_k3a[14], a9_k4a[14] );
xor a9_C977 ( k8b[15], a9_k3a[15], a9_k4a[15] );
xor a9_C976 ( k8b[16], a9_k3a[16], a9_k4a[16] );
xor a9_C975 ( k8b[17], a9_k3a[17], a9_k4a[17] );
xor a9_C974 ( k8b[18], a9_k3a[18], a9_k4a[18] );
xor a9_C973 ( k8b[19], a9_k3a[19], a9_k4a[19] );
xor a9_C972 ( k8b[20], a9_k3a[20], a9_k4a[20] );
xor a9_C971 ( k8b[21], a9_k3a[21], a9_k4a[21] );
xor a9_C970 ( k8b[22], a9_k3a[22], a9_k4a[22] );
xor a9_C969 ( k8b[23], a9_k3a[23], a9_k4a[23] );
xor a9_C968 ( k8b[24], a9_k3a[24], a9_k4a[24] );
xor a9_C967 ( k8b[25], a9_k3a[25], a9_k4a[25] );
xor a9_C966 ( k8b[26], a9_k3a[26], a9_k4a[26] );
xor a9_C965 ( k8b[27], a9_k3a[27], a9_k4a[27] );
xor a9_C964 ( k8b[28], a9_k3a[28], a9_k4a[28] );
xor a9_C963 ( k8b[29], a9_k3a[29], a9_k4a[29] );
xor a9_C962 ( k8b[30], a9_k3a[30], a9_k4a[30] );
xor a9_C960 ( k8b[32], a9_k2a[0], a9_k4a[0] );
xor a9_C959 ( k8b[33], a9_k2a[1], a9_k4a[1] );
xor a9_C958 ( k8b[34], a9_k2a[2], a9_k4a[2] );
xor a9_C957 ( k8b[35], a9_k2a[3], a9_k4a[3] );
xor a9_C956 ( k8b[36], a9_k2a[4], a9_k4a[4] );
xor a9_C955 ( k8b[37], a9_k2a[5], a9_k4a[5] );
xor a9_C954 ( k8b[38], a9_k2a[6], a9_k4a[6] );
xor a9_C953 ( k8b[39], a9_k2a[7], a9_k4a[7] );
xor a9_C952 ( k8b[40], a9_k2a[8], a9_k4a[8] );
xor a9_C951 ( k8b[41], a9_k2a[9], a9_k4a[9] );
xor a9_C950 ( k8b[42], a9_k2a[10], a9_k4a[10] );
xor a9_C949 ( k8b[43], a9_k2a[11], a9_k4a[11] );
xor a9_C948 ( k8b[44], a9_k2a[12], a9_k4a[12] );
xor a9_C947 ( k8b[45], a9_k2a[13], a9_k4a[13] );
xor a9_C946 ( k8b[46], a9_k2a[14], a9_k4a[14] );
xor a9_C945 ( k8b[47], a9_k2a[15], a9_k4a[15] );
xor a9_C944 ( k8b[48], a9_k2a[16], a9_k4a[16] );
xor a9_C943 ( k8b[49], a9_k2a[17], a9_k4a[17] );
xor a9_C942 ( k8b[50], a9_k2a[18], a9_k4a[18] );
xor a9_C941 ( k8b[51], a9_k2a[19], a9_k4a[19] );
xor a9_C940 ( k8b[52], a9_k2a[20], a9_k4a[20] );
xor a9_C939 ( k8b[53], a9_k2a[21], a9_k4a[21] );
xor a9_C938 ( k8b[54], a9_k2a[22], a9_k4a[22] );
xor a9_C937 ( k8b[55], a9_k2a[23], a9_k4a[23] );
xor a9_C936 ( k8b[56], a9_k2a[24], a9_k4a[24] );
xor a9_C935 ( k8b[57], a9_k2a[25], a9_k4a[25] );
xor a9_C934 ( k8b[58], a9_k2a[26], a9_k4a[26] );
xor a9_C933 ( k8b[59], a9_k2a[27], a9_k4a[27] );
xor a9_C932 ( k8b[60], a9_k2a[28], a9_k4a[28] );
xor a9_C931 ( k8b[61], a9_k2a[29], a9_k4a[29] );
xor a9_C930 ( k8b[62], a9_k2a[30], a9_k4a[30] );
xor a9_C929 ( k8b[63], a9_k2a[31], a9_k4a[31] );
xor a9_C928 ( k8b[64], a9_k1a[0], a9_k4a[0] );
xor a9_C927 ( k8b[65], a9_k1a[1], a9_k4a[1] );
xor a9_C926 ( k8b[66], a9_k1a[2], a9_k4a[2] );
xor a9_C925 ( k8b[67], a9_k1a[3], a9_k4a[3] );
xor a9_C924 ( k8b[68], a9_k1a[4], a9_k4a[4] );
xor a9_C923 ( k8b[69], a9_k1a[5], a9_k4a[5] );
xor a9_C922 ( k8b[70], a9_k1a[6], a9_k4a[6] );
xor a9_C921 ( k8b[71], a9_k1a[7], a9_k4a[7] );
xor a9_C920 ( k8b[72], a9_k1a[8], a9_k4a[8] );
xor a9_C919 ( k8b[73], a9_k1a[9], a9_k4a[9] );
xor a9_C918 ( k8b[74], a9_k1a[10], a9_k4a[10] );
xor a9_C917 ( k8b[75], a9_k1a[11], a9_k4a[11] );
xor a9_C916 ( k8b[76], a9_k1a[12], a9_k4a[12] );
xor a9_C915 ( k8b[77], a9_k1a[13], a9_k4a[13] );
xor a9_C914 ( k8b[78], a9_k1a[14], a9_k4a[14] );
xor a9_C913 ( k8b[79], a9_k1a[15], a9_k4a[15] );
xor a9_C912 ( k8b[80], a9_k1a[16], a9_k4a[16] );
xor a9_C911 ( k8b[81], a9_k1a[17], a9_k4a[17] );
xor a9_C910 ( k8b[82], a9_k1a[18], a9_k4a[18] );
xor a9_C909 ( k8b[83], a9_k1a[19], a9_k4a[19] );
xor a9_C908 ( k8b[84], a9_k1a[20], a9_k4a[20] );
xor a9_C907 ( k8b[85], a9_k1a[21], a9_k4a[21] );
xor a9_C906 ( k8b[86], a9_k1a[22], a9_k4a[22] );
xor a9_C905 ( k8b[87], a9_k1a[23], a9_k4a[23] );
xor a9_C904 ( k8b[88], a9_k1a[24], a9_k4a[24] );
xor a9_C903 ( k8b[89], a9_k1a[25], a9_k4a[25] );
xor a9_C902 ( k8b[90], a9_k1a[26], a9_k4a[26] );
xor a9_C901 ( k8b[91], a9_k1a[27], a9_k4a[27] );
xor a9_C900 ( k8b[92], a9_k1a[28], a9_k4a[28] );
xor a9_C899 ( k8b[93], a9_k1a[29], a9_k4a[29] );
xor a9_C898 ( k8b[94], a9_k1a[30], a9_k4a[30] );
xor a9_C897 ( k8b[95], a9_k1a[31], a9_k4a[31] );
buf U1876 ( n1548, n1555 );
buf U1877 ( n1549, n1555 );
buf U1878 ( n1550, n1555 );
buf U1879 ( n1551, n1554 );
buf U1880 ( n1552, n1554 );
buf U1881 ( n1555, n1283 );
buf U1882 ( n1554, n1283 );
buf U1883 ( n1547, n1556 );
not U1884 ( n1560, n1578 );
not U1885 ( n1561, n1578 );
not U1886 ( n1568, n1575 );
not U1887 ( n1572, n1573 );
not U1888 ( n1571, n1574 );
not U1889 ( n1569, n1575 );
not U1890 ( n1570, n1575 );
not U1891 ( n1565, n1576 );
not U1892 ( n1563, n1577 );
not U1893 ( n1567, n1576 );
not U1894 ( n1564, n1577 );
not U1895 ( n1566, n1576 );
not U1896 ( n1562, n1577 );
buf U1897 ( n1578, n1585 );
buf U1898 ( n1575, n1586 );
buf U1899 ( n1573, n1587 );
buf U1900 ( n1574, n1587 );
buf U1901 ( n1577, n1586 );
buf U1902 ( n1576, n1586 );
buf U1903 ( n1336, n1543 );
buf U1904 ( n1337, n1543 );
buf U1905 ( n1338, n1543 );
buf U1906 ( n1339, n1543 );
buf U1907 ( n1340, n1543 );
buf U1908 ( n1341, n1543 );
buf U1909 ( n1342, n1543 );
buf U1910 ( n1343, n1543 );
buf U1911 ( n1344, n1543 );
buf U1912 ( n1345, n1543 );
buf U1913 ( n1346, n1543 );
buf U1914 ( n1347, n1543 );
buf U1915 ( n1348, n1542 );
buf U1916 ( n1349, n1542 );
buf U1917 ( n1350, n1542 );
buf U1918 ( n1351, n1542 );
buf U1919 ( n1352, n1542 );
buf U1920 ( n1353, n1542 );
buf U1921 ( n1354, n1542 );
buf U1922 ( n1355, n1542 );
buf U1923 ( n1356, n1542 );
buf U1924 ( n1357, n1542 );
buf U1925 ( n1358, n1542 );
buf U1926 ( n1359, n1542 );
buf U1927 ( n1360, n1541 );
buf U1928 ( n1361, n1541 );
buf U1929 ( n1362, n1541 );
buf U1930 ( n1363, n1541 );
buf U1931 ( n1364, n1541 );
buf U1932 ( n1365, n1541 );
buf U1933 ( n1366, n1541 );
buf U1934 ( n1367, n1541 );
buf U1935 ( n1368, n1541 );
buf U1936 ( n1369, n1541 );
buf U1937 ( n1370, n1541 );
buf U1938 ( n1371, n1541 );
buf U1939 ( n1372, n1540 );
buf U1940 ( n1373, n1540 );
buf U1941 ( n1374, n1540 );
buf U1942 ( n1375, n1540 );
buf U1943 ( n1376, n1540 );
buf U1944 ( n1377, n1540 );
buf U1945 ( n1378, n1540 );
buf U1946 ( n1379, n1540 );
buf U1947 ( n1380, n1540 );
buf U1948 ( n1381, n1540 );
buf U1949 ( n1382, n1540 );
buf U1950 ( n1383, n1540 );
buf U1951 ( n1384, n1539 );
buf U1952 ( n1385, n1539 );
buf U1953 ( n1386, n1539 );
buf U1954 ( n1387, n1539 );
buf U1955 ( n1388, n1539 );
buf U1956 ( n1389, n1539 );
buf U1957 ( n1390, n1539 );
buf U1958 ( n1391, n1539 );
buf U1959 ( n1392, n1539 );
buf U1960 ( n1393, n1539 );
buf U1961 ( n1394, n1539 );
buf U1962 ( n1395, n1539 );
buf U1963 ( n1396, n1538 );
buf U1964 ( n1397, n1538 );
buf U1965 ( n1398, n1538 );
buf U1966 ( n1399, n1538 );
buf U1967 ( n1400, n1538 );
buf U1968 ( n1401, n1538 );
buf U1969 ( n1402, n1538 );
buf U1970 ( n1403, n1538 );
buf U1971 ( n1404, n1538 );
buf U1972 ( n1405, n1538 );
buf U1973 ( n1406, n1538 );
buf U1974 ( n1407, n1538 );
buf U1975 ( n1408, n1537 );
buf U1976 ( n1409, n1537 );
buf U1977 ( n1410, n1537 );
buf U1978 ( n1411, n1537 );
buf U1979 ( n1412, n1537 );
buf U1980 ( n1413, n1537 );
buf U1981 ( n1414, n1537 );
buf U1982 ( n1415, n1537 );
buf U1983 ( n1416, n1537 );
buf U1984 ( n1417, n1537 );
buf U1985 ( n1418, n1537 );
buf U1986 ( n1419, n1537 );
buf U1987 ( n1420, n1536 );
buf U1988 ( n1421, n1536 );
buf U1989 ( n1422, n1536 );
buf U1990 ( n1423, n1536 );
buf U1991 ( n1424, n1536 );
buf U1992 ( n1425, n1536 );
buf U1993 ( n1426, n1536 );
buf U1994 ( n1427, n1536 );
buf U1995 ( n1428, n1536 );
buf U1996 ( n1429, n1536 );
buf U1997 ( n1430, n1536 );
buf U1998 ( n1431, n1536 );
buf U1999 ( n1432, n1535 );
buf U2000 ( n1433, n1535 );
buf U2001 ( n1434, n1535 );
buf U2002 ( n1435, n1535 );
buf U2003 ( n1436, n1535 );
buf U2004 ( n1437, n1535 );
buf U2005 ( n1438, n1535 );
buf U2006 ( n1439, n1535 );
buf U2007 ( n1440, n1535 );
buf U2008 ( n1441, n1535 );
buf U2009 ( n1442, n1535 );
buf U2010 ( n1443, n1535 );
buf U2011 ( n1444, n1534 );
buf U2012 ( n1445, n1534 );
buf U2013 ( n1446, n1534 );
buf U2014 ( n1447, n1534 );
buf U2015 ( n1448, n1534 );
buf U2016 ( n1449, n1534 );
buf U2017 ( n1450, n1534 );
buf U2018 ( n1451, n1534 );
buf U2019 ( n1452, n1534 );
buf U2020 ( n1453, n1534 );
buf U2021 ( n1454, n1534 );
buf U2022 ( n1455, n1534 );
buf U2023 ( n1456, n1533 );
buf U2024 ( n1457, n1533 );
buf U2025 ( n1458, n1533 );
buf U2026 ( n1459, n1533 );
buf U2027 ( n1460, n1533 );
buf U2028 ( n1461, n1533 );
buf U2029 ( n1462, n1533 );
buf U2030 ( n1463, n1533 );
buf U2031 ( n1464, n1533 );
buf U2032 ( n1465, n1533 );
buf U2033 ( n1466, n1533 );
buf U2034 ( n1467, n1533 );
buf U2035 ( n1468, n1532 );
buf U2036 ( n1469, n1532 );
buf U2037 ( n1470, n1532 );
buf U2038 ( n1471, n1532 );
buf U2039 ( n1472, n1532 );
buf U2040 ( n1473, n1532 );
buf U2041 ( n1474, n1532 );
buf U2042 ( n1475, n1532 );
buf U2043 ( n1476, n1532 );
buf U2044 ( n1477, n1532 );
buf U2045 ( n1478, n1532 );
buf U2046 ( n1479, n1532 );
buf U2047 ( n1480, n1531 );
buf U2048 ( n1481, n1531 );
buf U2049 ( n1482, n1531 );
buf U2050 ( n1483, n1531 );
buf U2051 ( n1484, n1531 );
buf U2052 ( n1485, n1531 );
buf U2053 ( n1486, n1531 );
buf U2054 ( n1487, n1531 );
buf U2055 ( n1488, n1531 );
buf U2056 ( n1489, n1531 );
buf U2057 ( n1490, n1531 );
buf U2058 ( n1491, n1531 );
buf U2059 ( n1492, n1530 );
buf U2060 ( n1493, n1530 );
buf U2061 ( n1494, n1530 );
buf U2062 ( n1495, n1530 );
buf U2063 ( n1496, n1530 );
buf U2064 ( n1497, n1530 );
buf U2065 ( n1498, n1530 );
buf U2066 ( n1499, n1530 );
buf U2067 ( n1500, n1530 );
buf U2068 ( n1501, n1530 );
buf U2069 ( n1502, n1530 );
buf U2070 ( n1503, n1530 );
buf U2071 ( n1504, n1529 );
buf U2072 ( n1505, n1529 );
buf U2073 ( n1506, n1529 );
buf U2074 ( n1507, n1529 );
buf U2075 ( n1508, n1529 );
buf U2076 ( n1509, n1529 );
buf U2077 ( n1510, n1529 );
buf U2078 ( n1511, n1529 );
buf U2079 ( n1512, n1529 );
buf U2080 ( n1513, n1529 );
buf U2081 ( n1514, n1529 );
buf U2082 ( n1515, n1529 );
buf U2083 ( n1586, n1557 );
buf U2084 ( n1587, n1558 );
buf U2085 ( n1303, n1546 );
buf U2086 ( n1304, n1546 );
buf U2087 ( n1305, n1546 );
buf U2088 ( n1306, n1546 );
buf U2089 ( n1307, n1546 );
buf U2090 ( n1308, n1546 );
buf U2091 ( n1309, n1546 );
buf U2092 ( n1310, n1546 );
buf U2093 ( n1311, n1546 );
buf U2094 ( n1312, n1545 );
buf U2095 ( n1313, n1545 );
buf U2096 ( n1314, n1545 );
buf U2097 ( n1315, n1545 );
buf U2098 ( n1316, n1545 );
buf U2099 ( n1317, n1545 );
buf U2100 ( n1318, n1545 );
buf U2101 ( n1319, n1545 );
buf U2102 ( n1320, n1545 );
buf U2103 ( n1321, n1545 );
buf U2104 ( n1322, n1545 );
buf U2105 ( n1323, n1545 );
buf U2106 ( n1324, n1544 );
buf U2107 ( n1325, n1544 );
buf U2108 ( n1326, n1544 );
buf U2109 ( n1327, n1544 );
buf U2110 ( n1328, n1544 );
buf U2111 ( n1329, n1544 );
buf U2112 ( n1330, n1544 );
buf U2113 ( n1331, n1544 );
buf U2114 ( n1332, n1544 );
buf U2115 ( n1333, n1544 );
buf U2116 ( n1334, n1544 );
buf U2117 ( n1335, n1544 );
buf U2118 ( n1516, n1528 );
buf U2119 ( n1517, n1528 );
buf U2120 ( n1518, n1528 );
buf U2121 ( n1519, n1528 );
buf U2122 ( n1520, n1528 );
buf U2123 ( n1521, n1528 );
buf U2124 ( n1522, n1528 );
buf U2125 ( n1523, n1528 );
buf U2126 ( n1524, n1528 );
buf U2127 ( n1525, n1528 );
buf U2128 ( n1526, n1528 );
buf U2129 ( n1527, n1528 );
buf U2130 ( n1543, n1548 );
buf U2131 ( n1542, n1548 );
buf U2132 ( n1541, n1548 );
buf U2133 ( n1540, n1549 );
buf U2134 ( n1539, n1549 );
buf U2135 ( n1538, n1549 );
buf U2136 ( n1537, n1550 );
buf U2137 ( n1536, n1550 );
buf U2138 ( n1535, n1550 );
buf U2139 ( n1534, n1551 );
buf U2140 ( n1533, n1551 );
buf U2141 ( n1532, n1551 );
buf U2142 ( n1531, n1552 );
buf U2143 ( n1530, n1552 );
buf U2144 ( n1529, n1552 );
buf U2145 ( n1557, n1559 );
nor U2146 ( n4, out_valid, n1568 );
buf U2147 ( n1558, n1559 );
buf U2148 ( n1545, n1547 );
buf U2149 ( n1544, n1547 );
buf U2150 ( n1528, n1553 );
buf U2151 ( n1553, n1554 );
buf U2152 ( n1546, n1547 );
buf U2153 ( n1559, n2 );
not U2154 ( out_valid, n3 );
buf U2155 ( n1556, n1283 );
nand U2156 ( n2, start, n1019 );
nand U2157 ( n1059, n72, n73 );
nand U2158 ( n72, key[33], n1561 );
or U2159 ( n73, n1560, n925 );
nand U2160 ( n1083, n120, n121 );
nand U2161 ( n120, key[57], n1564 );
or U2162 ( n121, n1561, n949 );
nand U2163 ( n1087, n128, n129 );
nand U2164 ( n128, key[61], n1560 );
or U2165 ( n129, n1560, n953 );
nand U2166 ( n1088, n130, n131 );
nand U2167 ( n130, key[62], n1565 );
or U2168 ( n131, n1561, n954 );
nand U2169 ( n1097, n148, n149 );
nand U2170 ( n148, key[71], n1563 );
or U2171 ( n149, n1561, n963 );
nand U2172 ( n1144, n242, n243 );
nand U2173 ( n242, key[118], n1570 );
or U2174 ( n243, n1560, n1010 );
nand U2175 ( n1091, n136, n137 );
nand U2176 ( n136, key[65], n1562 );
or U2177 ( n137, n1560, n957 );
nand U2178 ( n1060, n74, n75 );
nand U2179 ( n74, key[34], n1570 );
or U2180 ( n75, n1561, n926 );
nand U2181 ( n1092, n138, n139 );
nand U2182 ( n138, key[66], n1566 );
or U2183 ( n139, n1561, n958 );
nand U2184 ( n1096, n146, n147 );
nand U2185 ( n146, key[70], n1562 );
or U2186 ( n147, n1560, n962 );
and U2187 ( n1023, n4, N137 );
xnor U2188 ( N137, validCounter[3], n1592 );
and U2189 ( n1025, n4, N135 );
nand U2190 ( N135, n1590, n1589 );
nand U2191 ( n1589, validCounter[1], validCounter[0] );
nand U2192 ( n1068, n90, n91 );
or U2193 ( n91, n1571, n934 );
nand U2194 ( n90, key[42], n1560 );
nand U2195 ( n1078, n110, n111 );
or U2196 ( n111, n1565, n944 );
nand U2197 ( n110, key[52], n1560 );
nand U2198 ( n1079, n112, n113 );
or U2199 ( n113, n1562, n945 );
nand U2200 ( n112, key[53], n1560 );
nand U2201 ( n1080, n114, n115 );
or U2202 ( n115, n1567, n946 );
nand U2203 ( n114, key[54], n1561 );
nand U2204 ( n1089, n132, n133 );
or U2205 ( n133, n1571, n955 );
nand U2206 ( n132, key[63], n1561 );
nand U2207 ( n1094, n142, n143 );
or U2208 ( n143, n1564, n960 );
nand U2209 ( n142, key[68], n1561 );
nand U2210 ( n1102, n158, n159 );
or U2211 ( n159, n1572, n968 );
nand U2212 ( n158, key[76], n1561 );
nand U2213 ( n1107, n168, n169 );
or U2214 ( n169, n1572, n973 );
nand U2215 ( n168, key[81], n1560 );
nand U2216 ( n1129, n212, n213 );
or U2217 ( n213, n1562, n995 );
nand U2218 ( n212, key[103], n1561 );
nand U2219 ( n1132, n218, n219 );
or U2220 ( n219, n1566, n998 );
nand U2221 ( n218, key[106], n1560 );
nand U2222 ( n1136, n226, n227 );
or U2223 ( n227, n1563, n1002 );
nand U2224 ( n226, key[110], n1560 );
nand U2225 ( n1139, n232, n233 );
or U2226 ( n233, n1564, n1005 );
nand U2227 ( n232, key[113], n1561 );
nand U2228 ( n1145, n244, n245 );
or U2229 ( n245, n1568, n1011 );
nand U2230 ( n244, key[119], n1561 );
nand U2231 ( n1153, n260, n261 );
or U2232 ( n261, n1563, n1018 );
nand U2233 ( n260, key[127], n1560 );
nand U2234 ( n1197, n391, n392 );
nand U2235 ( n391, s0[43], n1585 );
nand U2236 ( n392, n1560, n393 );
xor U2237 ( n393, state[43], key[43] );
nand U2238 ( n1208, n424, n425 );
nand U2239 ( n424, s0[54], n1584 );
nand U2240 ( n425, n1560, n426 );
xor U2241 ( n426, state[54], key[54] );
nand U2242 ( n1173, n319, n320 );
nand U2243 ( n319, s0[19], n1581 );
nand U2244 ( n320, n1561, n321 );
xor U2245 ( n321, state[19], key[19] );
nand U2246 ( n1253, n559, n560 );
nand U2247 ( n559, s0[99], n1581 );
nand U2248 ( n560, n1561, n561 );
xor U2249 ( n561, state[99], key[99] );
nand U2250 ( n1258, n574, n575 );
nand U2251 ( n574, s0[104], n1582 );
nand U2252 ( n575, n1560, n576 );
xor U2253 ( n576, state[104], key[104] );
nand U2254 ( n1268, n604, n605 );
nand U2255 ( n604, s0[114], n1580 );
nand U2256 ( n605, n1560, n606 );
xor U2257 ( n606, state[114], key[114] );
nand U2258 ( n1193, n379, n380 );
nand U2259 ( n379, s0[39], n1558 );
nand U2260 ( n380, n1560, n381 );
xor U2261 ( n381, state[39], key[39] );
nand U2262 ( n1224, n472, n473 );
nand U2263 ( n472, s0[70], n2 );
nand U2264 ( n473, n1561, n474 );
xor U2265 ( n474, state[70], key[70] );
nand U2266 ( n1158, n274, n275 );
nand U2267 ( n274, s0[4], n1577 );
nand U2268 ( n275, n1560, n276 );
xor U2269 ( n276, state[4], key[4] );
nand U2270 ( n1159, n277, n278 );
nand U2271 ( n277, s0[5], n1578 );
nand U2272 ( n278, n1561, n279 );
xor U2273 ( n279, state[5], key[5] );
nand U2274 ( n1172, n316, n317 );
nand U2275 ( n316, s0[18], n1587 );
nand U2276 ( n317, n1560, n318 );
xor U2277 ( n318, state[18], key[18] );
nand U2278 ( n1198, n394, n395 );
nand U2279 ( n394, s0[44], n1557 );
nand U2280 ( n395, n1561, n396 );
xor U2281 ( n396, state[44], key[44] );
nand U2282 ( n1257, n571, n572 );
nand U2283 ( n571, s0[103], n1574 );
nand U2284 ( n572, n1561, n573 );
xor U2285 ( n573, state[103], key[103] );
nand U2286 ( n1266, n598, n599 );
nand U2287 ( n598, s0[112], n1578 );
nand U2288 ( n599, n1561, n600 );
xor U2289 ( n600, state[112], key[112] );
nand U2290 ( n1267, n601, n602 );
nand U2291 ( n601, s0[113], n1578 );
nand U2292 ( n602, n1560, n603 );
xor U2293 ( n603, state[113], key[113] );
nand U2294 ( n1276, n628, n629 );
nand U2295 ( n628, s0[122], n1576 );
nand U2296 ( n629, n1561, n630 );
xor U2297 ( n630, state[122], key[122] );
nand U2298 ( n1072, n98, n99 );
nand U2299 ( n98, key[46], n1565 );
or U2300 ( n99, n1572, n938 );
nand U2301 ( n1112, n178, n179 );
nand U2302 ( n178, key[86], n1563 );
or U2303 ( n179, n1568, n978 );
nand U2304 ( n1122, n198, n199 );
nand U2305 ( n198, key[96], n1564 );
or U2306 ( n199, n1571, n988 );
nand U2307 ( n1146, n246, n247 );
nand U2308 ( n246, key[120], n1564 );
or U2309 ( n247, n1571, n1284 );
nand U2310 ( n1104, n162, n163 );
nand U2311 ( n162, key[78], n1565 );
or U2312 ( n163, n1572, n970 );
nand U2313 ( n1109, n172, n173 );
nand U2314 ( n172, key[83], n1565 );
or U2315 ( n173, n1564, n975 );
nand U2316 ( n1061, n76, n77 );
nand U2317 ( n76, key[35], n1569 );
or U2318 ( n77, n1572, n927 );
nand U2319 ( n1110, n174, n175 );
nand U2320 ( n174, key[84], n1569 );
or U2321 ( n175, n1572, n976 );
nand U2322 ( n1121, n196, n197 );
nand U2323 ( n196, key[95], n1569 );
or U2324 ( n197, n1572, n987 );
nand U2325 ( n1149, n252, n253 );
nand U2326 ( n252, key[123], n1563 );
or U2327 ( n253, n1568, n1014 );
nand U2328 ( n1101, n156, n157 );
nand U2329 ( n156, key[75], n1568 );
or U2330 ( n157, n1572, n967 );
nand U2331 ( n1106, n166, n167 );
nand U2332 ( n166, key[80], n1565 );
or U2333 ( n167, n1566, n972 );
nand U2334 ( n1135, n224, n225 );
nand U2335 ( n224, key[109], n1565 );
or U2336 ( n225, n1571, n1001 );
nand U2337 ( n1123, n200, n201 );
nand U2338 ( n200, key[97], n1563 );
or U2339 ( n201, n1571, n989 );
nand U2340 ( n1140, n234, n235 );
nand U2341 ( n234, key[114], n1564 );
or U2342 ( n235, n1571, n1006 );
nand U2343 ( n1071, n96, n97 );
nand U2344 ( n96, key[45], n1566 );
or U2345 ( n97, n1568, n937 );
nand U2346 ( n1103, n160, n161 );
nand U2347 ( n160, key[77], n1572 );
or U2348 ( n161, n1572, n969 );
nand U2349 ( n1108, n170, n171 );
nand U2350 ( n170, key[82], n1572 );
or U2351 ( n171, n1571, n974 );
nand U2352 ( n1111, n176, n177 );
nand U2353 ( n176, key[85], n1566 );
or U2354 ( n177, n1568, n977 );
nand U2355 ( n1074, n102, n103 );
nand U2356 ( n102, key[48], n1567 );
or U2357 ( n103, n1571, n940 );
nand U2358 ( n1058, n70, n71 );
nand U2359 ( n70, key[32], n1572 );
or U2360 ( n71, n1571, n924 );
nand U2361 ( n1114, n182, n183 );
nand U2362 ( n182, key[88], n1571 );
or U2363 ( n183, n1571, n980 );
nand U2364 ( n1131, n216, n217 );
nand U2365 ( n216, key[105], n1563 );
or U2366 ( n217, n1571, n997 );
nand U2367 ( n1151, n256, n257 );
nand U2368 ( n256, key[125], n1569 );
or U2369 ( n257, n1561, n1016 );
nand U2370 ( n1067, n88, n89 );
nand U2371 ( n88, key[41], n1564 );
or U2372 ( n89, n1564, n933 );
nand U2373 ( n1113, n180, n181 );
nand U2374 ( n180, key[87], n1570 );
or U2375 ( n181, n1571, n979 );
nand U2376 ( n1073, n100, n101 );
nand U2377 ( n100, key[47], n1567 );
or U2378 ( n101, n1560, n939 );
nand U2379 ( n1086, n126, n127 );
nand U2380 ( n126, key[60], n1566 );
or U2381 ( n127, n1561, n952 );
nand U2382 ( n1105, n164, n165 );
nand U2383 ( n164, key[79], n1566 );
or U2384 ( n165, n1560, n971 );
nand U2385 ( n1033, n20, n21 );
nand U2386 ( n21, k0[7], n1579 );
nand U2387 ( n20, key[7], n1561 );
nand U2388 ( n1028, n10, n11 );
nand U2389 ( n11, k0[2], n1559 );
nand U2390 ( n10, key[2], n1560 );
nand U2391 ( n1029, n12, n13 );
nand U2392 ( n13, k0[3], n1558 );
nand U2393 ( n12, key[3], n1571 );
nand U2394 ( n1090, n134, n135 );
or U2395 ( n135, n1570, n956 );
nand U2396 ( n134, key[64], n1567 );
nand U2397 ( n1116, n186, n187 );
or U2398 ( n187, n1570, n982 );
nand U2399 ( n186, key[90], n1562 );
nand U2400 ( n1128, n210, n211 );
or U2401 ( n211, n1564, n994 );
nand U2402 ( n210, key[102], n1572 );
nand U2403 ( n1040, n34, n35 );
nand U2404 ( n35, k0[14], n1302 );
nand U2405 ( n34, key[14], n1569 );
nand U2406 ( n1037, n28, n29 );
nand U2407 ( n29, k0[11], n1579 );
nand U2408 ( n28, key[11], n1572 );
nand U2409 ( n1043, n40, n41 );
nand U2410 ( n41, k0[17], n1580 );
nand U2411 ( n40, key[17], n1572 );
nand U2412 ( n1049, n52, n53 );
nand U2413 ( n53, k0[23], n1558 );
nand U2414 ( n52, key[23], n1572 );
nand U2415 ( n1030, n14, n15 );
nand U2416 ( n15, k0[4], n1575 );
nand U2417 ( n14, key[4], n1572 );
nand U2418 ( n1075, n104, n105 );
or U2419 ( n105, n1569, n941 );
nand U2420 ( n104, key[49], n1572 );
nand U2421 ( n1142, n238, n239 );
or U2422 ( n239, n1565, n1008 );
nand U2423 ( n238, key[116], n1572 );
nand U2424 ( n1045, n44, n45 );
nand U2425 ( n45, k0[19], n1582 );
nand U2426 ( n44, key[19], n1564 );
nand U2427 ( n1032, n18, n19 );
nand U2428 ( n19, k0[6], n1587 );
nand U2429 ( n18, key[6], n1566 );
nand U2430 ( n1138, n230, n231 );
or U2431 ( n231, n1566, n1004 );
nand U2432 ( n230, key[112], n1560 );
nand U2433 ( n1063, n80, n81 );
nand U2434 ( n80, key[37], n1567 );
or U2435 ( n81, n1569, n929 );
nand U2436 ( n1069, n92, n93 );
nand U2437 ( n92, key[43], n1563 );
or U2438 ( n93, n1569, n935 );
nand U2439 ( n1147, n248, n249 );
nand U2440 ( n248, key[121], n1565 );
or U2441 ( n249, n1569, n1012 );
nand U2442 ( n1124, n202, n203 );
nand U2443 ( n202, key[98], n1571 );
or U2444 ( n203, n1569, n990 );
nand U2445 ( n1259, n577, n578 );
nand U2446 ( n577, s0[105], n1302 );
nand U2447 ( n578, n1572, n579 );
xor U2448 ( n579, state[105], key[105] );
nand U2449 ( n1095, n144, n145 );
nand U2450 ( n144, key[69], n1567 );
or U2451 ( n145, n1570, n961 );
nand U2452 ( n1143, n240, n241 );
nand U2453 ( n240, key[117], n1570 );
or U2454 ( n241, n1570, n1009 );
nand U2455 ( n1150, n254, n255 );
nand U2456 ( n254, key[124], n1568 );
or U2457 ( n255, n1569, n1015 );
nand U2458 ( n1082, n118, n119 );
nand U2459 ( n118, key[56], n1562 );
or U2460 ( n119, n1570, n948 );
nand U2461 ( n1085, n124, n125 );
nand U2462 ( n124, key[59], n1568 );
or U2463 ( n125, n1570, n951 );
nand U2464 ( n1160, n280, n281 );
nand U2465 ( n280, s0[6], n1579 );
nand U2466 ( n281, n1572, n282 );
xor U2467 ( n282, state[6], key[6] );
nand U2468 ( n1174, n322, n323 );
nand U2469 ( n322, s0[20], n1579 );
nand U2470 ( n323, n1572, n324 );
xor U2471 ( n324, state[20], key[20] );
nand U2472 ( n1220, n460, n461 );
nand U2473 ( n460, s0[66], n1583 );
nand U2474 ( n461, n1572, n462 );
xor U2475 ( n462, state[66], key[66] );
nand U2476 ( n1161, n283, n284 );
nand U2477 ( n283, s0[7], n1580 );
nand U2478 ( n284, n1563, n285 );
xor U2479 ( n285, state[7], key[7] );
nand U2480 ( n1187, n361, n362 );
nand U2481 ( n361, s0[33], n1583 );
nand U2482 ( n362, n1567, n363 );
xor U2483 ( n363, state[33], key[33] );
nand U2484 ( n1243, n529, n530 );
nand U2485 ( n529, s0[89], n1583 );
nand U2486 ( n530, n1569, n531 );
xor U2487 ( n531, state[89], key[89] );
nand U2488 ( n1053, n60, n61 );
nand U2489 ( n61, k0[27], n1580 );
nand U2490 ( n60, key[27], n1566 );
nand U2491 ( n1050, n54, n55 );
nand U2492 ( n55, k0[24], n1557 );
nand U2493 ( n54, key[24], n1569 );
nand U2494 ( n1052, n58, n59 );
nand U2495 ( n59, k0[26], n1586 );
nand U2496 ( n58, key[26], n1563 );
nand U2497 ( n1099, n152, n153 );
or U2498 ( n153, n1563, n965 );
nand U2499 ( n152, key[73], n1567 );
nand U2500 ( n1115, n184, n185 );
or U2501 ( n185, n1564, n981 );
nand U2502 ( n184, key[89], n1564 );
nand U2503 ( n1127, n208, n209 );
or U2504 ( n209, n1566, n993 );
nand U2505 ( n208, key[101], n1566 );
nand U2506 ( n1242, n526, n527 );
nand U2507 ( n526, s0[88], n1582 );
nand U2508 ( n527, n1565, n528 );
xor U2509 ( n528, state[88], key[88] );
nand U2510 ( n1264, n592, n593 );
nand U2511 ( n592, s0[110], n1558 );
nand U2512 ( n593, n1565, n594 );
xor U2513 ( n594, state[110], key[110] );
nand U2514 ( n1199, n397, n398 );
nand U2515 ( n397, s0[45], n1587 );
nand U2516 ( n398, n1572, n399 );
xor U2517 ( n399, state[45], key[45] );
nand U2518 ( n1252, n556, n557 );
nand U2519 ( n556, s0[98], n1576 );
nand U2520 ( n557, n1572, n558 );
xor U2521 ( n558, state[98], key[98] );
nand U2522 ( n1084, n122, n123 );
or U2523 ( n123, n1564, n950 );
nand U2524 ( n122, key[58], n1571 );
nand U2525 ( n1100, n154, n155 );
or U2526 ( n155, n1562, n966 );
nand U2527 ( n154, key[74], n1571 );
nand U2528 ( n1119, n192, n193 );
or U2529 ( n193, n1567, n985 );
nand U2530 ( n192, key[93], n1571 );
nand U2531 ( n1125, n204, n205 );
or U2532 ( n205, n1567, n991 );
nand U2533 ( n204, key[99], n1571 );
nand U2534 ( n1137, n228, n229 );
or U2535 ( n229, n1568, n1003 );
nand U2536 ( n228, key[111], n1571 );
nand U2537 ( n1265, n595, n596 );
nand U2538 ( n595, s0[111], n1573 );
nand U2539 ( n596, n1572, n597 );
xor U2540 ( n597, state[111], key[111] );
nand U2541 ( n1256, n568, n569 );
nand U2542 ( n568, s0[102], n1574 );
nand U2543 ( n569, n1572, n570 );
xor U2544 ( n570, state[102], key[102] );
nand U2545 ( n1154, n262, n263 );
nand U2546 ( n262, s0[0], n1576 );
nand U2547 ( n263, n1561, n264 );
xor U2548 ( n264, state[0], key[0] );
nand U2549 ( n1255, n565, n566 );
nand U2550 ( n565, s0[101], n1573 );
nand U2551 ( n566, n1570, n567 );
xor U2552 ( n567, state[101], key[101] );
nand U2553 ( n1251, n553, n554 );
nand U2554 ( n553, s0[97], n1575 );
nand U2555 ( n554, n1562, n555 );
xor U2556 ( n555, state[97], key[97] );
nand U2557 ( n1031, n16, n17 );
nand U2558 ( n17, k0[5], n1576 );
nand U2559 ( n16, key[5], n1563 );
nand U2560 ( n1076, n106, n107 );
or U2561 ( n107, n1566, n942 );
nand U2562 ( n106, key[50], n1567 );
nand U2563 ( n1117, n188, n189 );
or U2564 ( n189, n1563, n983 );
nand U2565 ( n188, key[91], n1569 );
nand U2566 ( n1118, n190, n191 );
or U2567 ( n191, n1566, n984 );
nand U2568 ( n190, key[92], n1566 );
nand U2569 ( n1126, n206, n207 );
or U2570 ( n207, n1562, n992 );
nand U2571 ( n206, key[100], n1568 );
nand U2572 ( n1155, n265, n266 );
nand U2573 ( n265, s0[1], n1577 );
nand U2574 ( n266, n1570, n267 );
xor U2575 ( n267, state[1], key[1] );
nand U2576 ( n1188, n364, n365 );
nand U2577 ( n364, s0[34], n1587 );
nand U2578 ( n365, n1562, n366 );
xor U2579 ( n366, state[34], key[34] );
nand U2580 ( n1223, n469, n470 );
nand U2581 ( n469, s0[69], n1574 );
nand U2582 ( n470, n1560, n471 );
xor U2583 ( n471, state[69], key[69] );
nand U2584 ( n1237, n511, n512 );
nand U2585 ( n511, s0[83], n1573 );
nand U2586 ( n512, n1570, n513 );
xor U2587 ( n513, state[83], key[83] );
nand U2588 ( n1263, n589, n590 );
nand U2589 ( n589, s0[109], n1575 );
nand U2590 ( n590, n1561, n591 );
xor U2591 ( n591, state[109], key[109] );
nand U2592 ( n1195, n385, n386 );
nand U2593 ( n385, s0[41], n1302 );
nand U2594 ( n386, n1571, n387 );
xor U2595 ( n387, state[41], key[41] );
nand U2596 ( n1254, n562, n563 );
nand U2597 ( n562, s0[100], n1584 );
nand U2598 ( n563, n1565, n564 );
xor U2599 ( n564, state[100], key[100] );
nand U2600 ( n1222, n466, n467 );
nand U2601 ( n466, s0[68], n1581 );
nand U2602 ( n467, n1561, n468 );
xor U2603 ( n468, state[68], key[68] );
nand U2604 ( n1190, n370, n371 );
nand U2605 ( n370, s0[36], n1585 );
nand U2606 ( n371, n1571, n372 );
xor U2607 ( n372, state[36], key[36] );
nand U2608 ( n1236, n508, n509 );
nand U2609 ( n508, s0[82], n1585 );
nand U2610 ( n509, n1563, n510 );
xor U2611 ( n510, state[82], key[82] );
nand U2612 ( n1240, n520, n521 );
nand U2613 ( n520, s0[86], n1579 );
nand U2614 ( n521, n1571, n522 );
xor U2615 ( n522, state[86], key[86] );
nand U2616 ( n1250, n550, n551 );
nand U2617 ( n550, s0[96], n1579 );
nand U2618 ( n551, n1571, n552 );
xor U2619 ( n552, state[96], key[96] );
nand U2620 ( n1213, n439, n440 );
nand U2621 ( n439, s0[59], n1584 );
nand U2622 ( n440, n1567, n441 );
xor U2623 ( n441, state[59], key[59] );
nand U2624 ( n1178, n334, n335 );
nand U2625 ( n334, s0[24], n1582 );
nand U2626 ( n335, n1561, n336 );
xor U2627 ( n336, state[24], key[24] );
nand U2628 ( n1241, n523, n524 );
nand U2629 ( n523, s0[87], n1580 );
nand U2630 ( n524, n1564, n525 );
xor U2631 ( n525, state[87], key[87] );
nand U2632 ( n1191, n373, n374 );
nand U2633 ( n373, s0[37], n1586 );
nand U2634 ( n374, n1560, n375 );
xor U2635 ( n375, state[37], key[37] );
nand U2636 ( n1167, n301, n302 );
nand U2637 ( n301, s0[13], n1574 );
nand U2638 ( n302, n1569, n303 );
xor U2639 ( n303, state[13], key[13] );
nand U2640 ( n1239, n517, n518 );
nand U2641 ( n517, s0[85], n1578 );
nand U2642 ( n518, n1572, n519 );
xor U2643 ( n519, state[85], key[85] );
nand U2644 ( n1249, n547, n548 );
nand U2645 ( n547, s0[95], n1578 );
nand U2646 ( n548, n1562, n549 );
xor U2647 ( n549, state[95], key[95] );
nand U2648 ( n1278, n634, n635 );
nand U2649 ( n634, s0[124], n1557 );
nand U2650 ( n635, n1570, n636 );
xor U2651 ( n636, state[124], key[124] );
nand U2652 ( n1157, n271, n272 );
nand U2653 ( n271, s0[3], n1587 );
nand U2654 ( n272, n1571, n273 );
xor U2655 ( n273, state[3], key[3] );
nand U2656 ( n1235, n505, n506 );
nand U2657 ( n505, s0[81], n1586 );
nand U2658 ( n506, n1571, n507 );
xor U2659 ( n507, state[81], key[81] );
nand U2660 ( n1271, n613, n614 );
nand U2661 ( n613, s0[117], n1577 );
nand U2662 ( n614, n1571, n615 );
xor U2663 ( n615, state[117], key[117] );
nand U2664 ( n1279, n637, n638 );
nand U2665 ( n637, s0[125], n1587 );
nand U2666 ( n638, n1571, n639 );
xor U2667 ( n639, state[125], key[125] );
nand U2668 ( n1189, n367, n368 );
nand U2669 ( n367, s0[35], n1586 );
nand U2670 ( n368, n1569, n369 );
xor U2671 ( n369, state[35], key[35] );
nand U2672 ( n1156, n268, n269 );
nand U2673 ( n268, s0[2], n1578 );
nand U2674 ( n269, n1562, n270 );
xor U2675 ( n270, state[2], key[2] );
nand U2676 ( n1219, n457, n458 );
nand U2677 ( n457, s0[65], n1574 );
nand U2678 ( n458, n1565, n459 );
xor U2679 ( n459, state[65], key[65] );
nand U2680 ( n1141, n236, n237 );
nand U2681 ( n236, key[115], n1563 );
or U2682 ( n237, n1568, n1007 );
nand U2683 ( n1152, n258, n259 );
nand U2684 ( n258, key[126], n1563 );
or U2685 ( n259, n1568, n1017 );
nand U2686 ( n1062, n78, n79 );
nand U2687 ( n78, key[36], n1568 );
or U2688 ( n79, n1568, n928 );
nand U2689 ( n1081, n116, n117 );
nand U2690 ( n116, key[55], n1569 );
or U2691 ( n117, n1565, n947 );
nand U2692 ( n1070, n94, n95 );
nand U2693 ( n94, key[44], n1570 );
or U2694 ( n95, n1567, n936 );
nand U2695 ( n1077, n108, n109 );
nand U2696 ( n108, key[51], n1567 );
or U2697 ( n109, n1567, n943 );
nand U2698 ( n1093, n140, n141 );
nand U2699 ( n140, key[67], n1570 );
or U2700 ( n141, n1563, n959 );
nand U2701 ( n1130, n214, n215 );
nand U2702 ( n214, key[104], n1567 );
or U2703 ( n215, n1565, n996 );
nand U2704 ( n1134, n222, n223 );
nand U2705 ( n222, key[108], n1564 );
or U2706 ( n223, n1564, n1000 );
nand U2707 ( n1065, n84, n85 );
nand U2708 ( n84, key[39], n1562 );
or U2709 ( n85, n1567, n931 );
nand U2710 ( n1066, n86, n87 );
nand U2711 ( n86, key[40], n1566 );
or U2712 ( n87, n1565, n932 );
nand U2713 ( n1120, n194, n195 );
nand U2714 ( n194, key[94], n1568 );
or U2715 ( n195, n1565, n986 );
nand U2716 ( n1148, n250, n251 );
nand U2717 ( n250, key[122], n1562 );
or U2718 ( n251, n1563, n1013 );
nand U2719 ( n1034, n22, n23 );
nand U2720 ( n23, k0[8], n1302 );
nand U2721 ( n22, key[8], n1569 );
nand U2722 ( n1282, n646, n647 );
nand U2723 ( n647, k0[0], n1302 );
nand U2724 ( n646, key[0], n1569 );
nand U2725 ( n1057, n68, n69 );
nand U2726 ( n69, k0[31], n1582 );
nand U2727 ( n68, key[31], n1569 );
nand U2728 ( n1064, n82, n83 );
nand U2729 ( n82, key[38], n1570 );
or U2730 ( n83, n1566, n930 );
nand U2731 ( n1035, n24, n25 );
nand U2732 ( n25, k0[9], n1559 );
nand U2733 ( n24, key[9], n1570 );
nand U2734 ( n1098, n150, n151 );
or U2735 ( n151, n1562, n964 );
nand U2736 ( n150, key[72], n1570 );
nand U2737 ( n1133, n220, n221 );
nand U2738 ( n220, key[107], n1568 );
or U2739 ( n221, n1562, n999 );
nand U2740 ( n1163, n289, n290 );
nand U2741 ( n289, s0[9], n1585 );
nand U2742 ( n290, n1569, n291 );
xor U2743 ( n291, state[9], key[9] );
nand U2744 ( n1166, n298, n299 );
nand U2745 ( n298, s0[12], n1574 );
nand U2746 ( n299, n1569, n300 );
xor U2747 ( n300, state[12], key[12] );
nand U2748 ( n1169, n307, n308 );
nand U2749 ( n307, s0[15], n1558 );
nand U2750 ( n308, n1569, n309 );
xor U2751 ( n309, state[15], key[15] );
nand U2752 ( n1205, n415, n416 );
nand U2753 ( n415, s0[51], n1586 );
nand U2754 ( n416, n1569, n417 );
xor U2755 ( n417, state[51], key[51] );
nand U2756 ( n1209, n427, n428 );
nand U2757 ( n427, s0[55], n1573 );
nand U2758 ( n428, n1569, n429 );
xor U2759 ( n429, state[55], key[55] );
nand U2760 ( n1247, n541, n542 );
nand U2761 ( n541, s0[93], n1577 );
nand U2762 ( n542, n1569, n543 );
xor U2763 ( n543, state[93], key[93] );
nand U2764 ( n1261, n583, n584 );
nand U2765 ( n583, s0[107], n1559 );
nand U2766 ( n584, n1569, n585 );
xor U2767 ( n585, state[107], key[107] );
nand U2768 ( n1171, n313, n314 );
nand U2769 ( n313, s0[17], n1557 );
nand U2770 ( n314, n1570, n315 );
xor U2771 ( n315, state[17], key[17] );
nand U2772 ( n1192, n376, n377 );
nand U2773 ( n376, s0[38], n1585 );
nand U2774 ( n377, n1570, n378 );
xor U2775 ( n378, state[38], key[38] );
nand U2776 ( n1194, n382, n383 );
nand U2777 ( n382, s0[40], n1582 );
nand U2778 ( n383, n1570, n384 );
xor U2779 ( n384, state[40], key[40] );
nand U2780 ( n1196, n388, n389 );
nand U2781 ( n388, s0[42], n2 );
nand U2782 ( n389, n1570, n390 );
xor U2783 ( n390, state[42], key[42] );
nand U2784 ( n1225, n475, n476 );
nand U2785 ( n475, s0[71], n1585 );
nand U2786 ( n476, n1570, n477 );
xor U2787 ( n477, state[71], key[71] );
nand U2788 ( n1269, n607, n608 );
nand U2789 ( n607, s0[115], n1581 );
nand U2790 ( n608, n1570, n609 );
xor U2791 ( n609, state[115], key[115] );
nand U2792 ( n1272, n616, n617 );
nand U2793 ( n616, s0[118], n1578 );
nand U2794 ( n617, n1570, n618 );
xor U2795 ( n618, state[118], key[118] );
nand U2796 ( n1280, n640, n641 );
nand U2797 ( n640, s0[126], n1586 );
nand U2798 ( n641, n1570, n642 );
xor U2799 ( n642, state[126], key[126] );
nand U2800 ( n1055, n64, n65 );
nand U2801 ( n65, k0[29], n1558 );
nand U2802 ( n64, key[29], n1568 );
nand U2803 ( n1051, n56, n57 );
nand U2804 ( n57, k0[25], n1577 );
nand U2805 ( n56, key[25], n1568 );
nand U2806 ( n1204, n412, n413 );
nand U2807 ( n412, s0[50], n1302 );
nand U2808 ( n413, n1568, n414 );
xor U2809 ( n414, state[50], key[50] );
nand U2810 ( n1262, n586, n587 );
nand U2811 ( n586, s0[108], n1302 );
nand U2812 ( n587, n1568, n588 );
xor U2813 ( n588, state[108], key[108] );
nand U2814 ( n1238, n514, n515 );
nand U2815 ( n514, s0[84], n1577 );
nand U2816 ( n515, n1568, n516 );
xor U2817 ( n516, state[84], key[84] );
nand U2818 ( n1248, n544, n545 );
nand U2819 ( n544, s0[94], n1577 );
nand U2820 ( n545, n1568, n546 );
xor U2821 ( n546, state[94], key[94] );
nand U2822 ( n1168, n304, n305 );
nand U2823 ( n304, s0[14], n1559 );
nand U2824 ( n305, n1568, n306 );
xor U2825 ( n306, state[14], key[14] );
nand U2826 ( n1162, n286, n287 );
nand U2827 ( n286, s0[8], n1578 );
nand U2828 ( n287, n1568, n288 );
xor U2829 ( n288, state[8], key[8] );
nand U2830 ( n1221, n463, n464 );
nand U2831 ( n463, s0[67], n1575 );
nand U2832 ( n464, n1568, n465 );
xor U2833 ( n465, state[67], key[67] );
nand U2834 ( n1042, n38, n39 );
nand U2835 ( n39, k0[16], n1302 );
nand U2836 ( n38, key[16], n1564 );
nand U2837 ( n1036, n26, n27 );
nand U2838 ( n27, k0[10], n1584 );
nand U2839 ( n26, key[10], n1565 );
nand U2840 ( n1039, n32, n33 );
nand U2841 ( n33, k0[13], n1581 );
nand U2842 ( n32, key[13], n1565 );
nand U2843 ( n1044, n42, n43 );
nand U2844 ( n43, k0[18], n1581 );
nand U2845 ( n42, key[18], n1564 );
nand U2846 ( n1027, n8, n9 );
nand U2847 ( n9, k0[1], n2 );
nand U2848 ( n8, key[1], n1567 );
nand U2849 ( n1041, n36, n37 );
nand U2850 ( n37, k0[15], n2 );
nand U2851 ( n36, key[15], n1563 );
nand U2852 ( n1056, n66, n67 );
nand U2853 ( n67, k0[30], n1573 );
nand U2854 ( n66, key[30], n1567 );
nand U2855 ( n1179, n337, n338 );
nand U2856 ( n337, s0[25], n1302 );
nand U2857 ( n338, n1565, n339 );
xor U2858 ( n339, state[25], key[25] );
nand U2859 ( n1281, n643, n644 );
nand U2860 ( n643, s0[127], n1585 );
nand U2861 ( n644, n1564, n645 );
xor U2862 ( n645, state[127], key[127] );
nand U2863 ( n1211, n433, n434 );
nand U2864 ( n433, s0[57], n1584 );
nand U2865 ( n434, n1567, n435 );
xor U2866 ( n435, state[57], key[57] );
nand U2867 ( n1217, n451, n452 );
nand U2868 ( n451, s0[63], n1584 );
nand U2869 ( n452, n1565, n453 );
xor U2870 ( n453, state[63], key[63] );
nand U2871 ( n1245, n535, n536 );
nand U2872 ( n535, s0[91], n1584 );
nand U2873 ( n536, n1567, n537 );
xor U2874 ( n537, state[91], key[91] );
nand U2875 ( n1175, n325, n326 );
nand U2876 ( n325, s0[21], n1580 );
nand U2877 ( n326, n1563, n327 );
xor U2878 ( n327, state[21], key[21] );
nand U2879 ( n1176, n328, n329 );
nand U2880 ( n328, s0[22], n1581 );
nand U2881 ( n329, n1564, n330 );
xor U2882 ( n330, state[22], key[22] );
nand U2883 ( n1182, n346, n347 );
nand U2884 ( n346, s0[28], n1579 );
nand U2885 ( n347, n1564, n348 );
xor U2886 ( n348, state[28], key[28] );
nand U2887 ( n1186, n358, n359 );
nand U2888 ( n358, s0[32], n1583 );
nand U2889 ( n359, n1565, n360 );
xor U2890 ( n360, state[32], key[32] );
nand U2891 ( n1202, n406, n407 );
nand U2892 ( n406, s0[48], n1580 );
nand U2893 ( n407, n1563, n408 );
xor U2894 ( n408, state[48], key[48] );
nand U2895 ( n1232, n496, n497 );
nand U2896 ( n496, s0[78], n1583 );
nand U2897 ( n497, n1565, n498 );
xor U2898 ( n498, state[78], key[78] );
nand U2899 ( n1270, n610, n611 );
nand U2900 ( n610, s0[116], n1582 );
nand U2901 ( n611, n1564, n612 );
xor U2902 ( n612, state[116], key[116] );
nand U2903 ( n1274, n622, n623 );
nand U2904 ( n622, s0[120], n1583 );
nand U2905 ( n623, n1563, n624 );
xor U2906 ( n624, state[120], key[120] );
nand U2907 ( n1277, n631, n632 );
nand U2908 ( n631, s0[123], n1583 );
nand U2909 ( n632, n1567, n633 );
xor U2910 ( n633, state[123], key[123] );
nand U2911 ( n1260, n580, n581 );
nand U2912 ( n580, s0[106], n2 );
nand U2913 ( n581, n1565, n582 );
xor U2914 ( n582, state[106], key[106] );
nand U2915 ( n1273, n619, n620 );
nand U2916 ( n619, s0[119], n1558 );
nand U2917 ( n620, n1564, n621 );
xor U2918 ( n621, state[119], key[119] );
nand U2919 ( n1165, n295, n296 );
nand U2920 ( n295, s0[11], n1557 );
nand U2921 ( n296, n1567, n297 );
xor U2922 ( n297, state[11], key[11] );
nand U2923 ( n1170, n310, n311 );
nand U2924 ( n310, s0[16], n1557 );
nand U2925 ( n311, n1564, n312 );
xor U2926 ( n312, state[16], key[16] );
nand U2927 ( n1177, n331, n332 );
nand U2928 ( n331, s0[23], n1586 );
nand U2929 ( n332, n1564, n333 );
xor U2930 ( n333, state[23], key[23] );
nand U2931 ( n1181, n343, n344 );
nand U2932 ( n343, s0[27], n1559 );
nand U2933 ( n344, n1563, n345 );
xor U2934 ( n345, state[27], key[27] );
nand U2935 ( n1185, n355, n356 );
nand U2936 ( n355, s0[31], n1587 );
nand U2937 ( n356, n1567, n357 );
xor U2938 ( n357, state[31], key[31] );
nand U2939 ( n1200, n400, n401 );
nand U2940 ( n400, s0[46], n1586 );
nand U2941 ( n401, n1567, n402 );
xor U2942 ( n402, state[46], key[46] );
nand U2943 ( n1203, n409, n410 );
nand U2944 ( n409, s0[49], n1573 );
nand U2945 ( n410, n1564, n411 );
xor U2946 ( n411, state[49], key[49] );
nand U2947 ( n1207, n421, n422 );
nand U2948 ( n421, s0[53], n1575 );
nand U2949 ( n422, n1567, n423 );
xor U2950 ( n423, state[53], key[53] );
nand U2951 ( n1212, n436, n437 );
nand U2952 ( n436, s0[58], n1573 );
nand U2953 ( n437, n1565, n438 );
xor U2954 ( n438, state[58], key[58] );
nand U2955 ( n1214, n442, n443 );
nand U2956 ( n442, s0[60], n1559 );
nand U2957 ( n443, n1565, n444 );
xor U2958 ( n444, state[60], key[60] );
nand U2959 ( n1216, n448, n449 );
nand U2960 ( n448, s0[62], n1557 );
nand U2961 ( n449, n1563, n450 );
xor U2962 ( n450, state[62], key[62] );
nand U2963 ( n1227, n481, n482 );
nand U2964 ( n481, s0[73], n1576 );
nand U2965 ( n482, n1563, n483 );
xor U2966 ( n483, state[73], key[73] );
nand U2967 ( n1229, n487, n488 );
nand U2968 ( n487, s0[75], n1575 );
nand U2969 ( n488, n1565, n489 );
xor U2970 ( n489, state[75], key[75] );
nand U2971 ( n1230, n490, n491 );
nand U2972 ( n490, s0[76], n1576 );
nand U2973 ( n491, n1563, n492 );
xor U2974 ( n492, state[76], key[76] );
nand U2975 ( n1233, n499, n500 );
nand U2976 ( n499, s0[79], n1576 );
nand U2977 ( n500, n1567, n501 );
xor U2978 ( n501, state[79], key[79] );
nand U2979 ( n1234, n502, n503 );
nand U2980 ( n502, s0[80], n1587 );
nand U2981 ( n503, n1563, n504 );
xor U2982 ( n504, state[80], key[80] );
nand U2983 ( n1048, n50, n51 );
nand U2984 ( n51, k0[22], n1559 );
nand U2985 ( n50, key[22], n1566 );
nand U2986 ( n1054, n62, n63 );
nand U2987 ( n63, k0[28], n2 );
nand U2988 ( n62, key[28], n1566 );
nand U2989 ( n1038, n30, n31 );
nand U2990 ( n31, k0[12], n1580 );
nand U2991 ( n30, key[12], n1562 );
nand U2992 ( n1046, n46, n47 );
nand U2993 ( n47, k0[20], n1579 );
nand U2994 ( n46, key[20], n1562 );
nand U2995 ( n1047, n48, n49 );
nand U2996 ( n49, k0[21], n2 );
nand U2997 ( n48, key[21], n1562 );
nand U2998 ( n1201, n403, n404 );
nand U2999 ( n403, s0[47], n1585 );
nand U3000 ( n404, n1562, n405 );
xor U3001 ( n405, state[47], key[47] );
nand U3002 ( n1183, n349, n350 );
nand U3003 ( n349, s0[29], n1584 );
nand U3004 ( n350, n1566, n351 );
xor U3005 ( n351, state[29], key[29] );
nand U3006 ( n1164, n292, n293 );
nand U3007 ( n292, s0[10], n1581 );
nand U3008 ( n293, n1566, n294 );
xor U3009 ( n294, state[10], key[10] );
nand U3010 ( n1184, n352, n353 );
nand U3011 ( n352, s0[30], n1582 );
nand U3012 ( n353, n1566, n354 );
xor U3013 ( n354, state[30], key[30] );
nand U3014 ( n1228, n484, n485 );
nand U3015 ( n484, s0[74], n1583 );
nand U3016 ( n485, n1562, n486 );
xor U3017 ( n486, state[74], key[74] );
nand U3018 ( n1226, n478, n479 );
nand U3019 ( n478, s0[72], n1576 );
nand U3020 ( n479, n1566, n480 );
xor U3021 ( n480, state[72], key[72] );
nand U3022 ( n1246, n538, n539 );
nand U3023 ( n538, s0[92], n1577 );
nand U3024 ( n539, n1566, n540 );
xor U3025 ( n540, state[92], key[92] );
nand U3026 ( n1180, n340, n341 );
nand U3027 ( n340, s0[26], n2 );
nand U3028 ( n341, n1562, n342 );
xor U3029 ( n342, state[26], key[26] );
nand U3030 ( n1215, n445, n446 );
nand U3031 ( n445, s0[61], n1558 );
nand U3032 ( n446, n1562, n447 );
xor U3033 ( n447, state[61], key[61] );
nand U3034 ( n1206, n418, n419 );
nand U3035 ( n418, s0[52], n1575 );
nand U3036 ( n419, n1566, n420 );
xor U3037 ( n420, state[52], key[52] );
nand U3038 ( n1210, n430, n431 );
nand U3039 ( n430, s0[56], n1574 );
nand U3040 ( n431, n1566, n432 );
xor U3041 ( n432, state[56], key[56] );
nand U3042 ( n1244, n532, n533 );
nand U3043 ( n532, s0[90], n1559 );
nand U3044 ( n533, n1562, n534 );
xor U3045 ( n534, state[90], key[90] );
nand U3046 ( n1218, n454, n455 );
nand U3047 ( n454, s0[64], n1573 );
nand U3048 ( n455, n1562, n456 );
xor U3049 ( n456, state[64], key[64] );
nand U3050 ( n1275, n625, n626 );
nand U3051 ( n625, s0[121], n1575 );
nand U3052 ( n626, n1562, n627 );
xor U3053 ( n627, state[121], key[121] );
nand U3054 ( n1231, n493, n494 );
nand U3055 ( n493, s0[77], n1574 );
nand U3056 ( n494, n1562, n495 );
xor U3057 ( n495, state[77], key[77] );
nand U3058 ( n1026, n1557, n7 );
nand U3059 ( n7, n1301, n3 );
nand U3060 ( n3, n648, n649 );
nor U3061 ( n649, validCounter[2], n650 );
nor U3062 ( n648, validCounter[1], validCounter[0] );
nand U3063 ( n650, n1020, n1021 );
nand U3064 ( n1022, n1, n1559 );
nand U3065 ( n1, N138, n3 );
xor U3066 ( N138, validCounter[4], n1593 );
nor U3067 ( n1593, validCounter[3], n1592 );
nand U3068 ( n1024, n2, n5 );
nand U3069 ( n5, N136, n3 );
nand U3070 ( N136, n1592, n1591 );
nand U3071 ( n1591, validCounter[2], n1590 );
or U3072 ( n1592, n1590, validCounter[2] );
or U3073 ( n1590, validCounter[1], validCounter[0] );
xor U3074 ( a10_v1[29], k9[93], n1299 );
xor U3075 ( a10_v1[28], k9[92], n1298 );
xor U3076 ( a10_v1[26], k9[90], n1297 );
xor U3077 ( a10_v1[25], k9[89], n1296 );
xor U3078 ( a10_v2[29], k9[61], a10_v1[29] );
xor U3079 ( a10_v2[28], k9[60], a10_v1[28] );
xor U3080 ( a10_v2[26], k9[58], a10_v1[26] );
xor U3081 ( a10_v2[25], k9[57], a10_v1[25] );
xor U3082 ( a9_v1[28], k8[92], n1295 );
xor U3083 ( a9_v1[27], k8[91], n1294 );
xor U3084 ( a9_v1[25], k8[89], n1293 );
xor U3085 ( a9_v1[24], k8[88], n1292 );
xor U3086 ( a9_v2[28], k8[60], a9_v1[28] );
xor U3087 ( a9_v2[27], k8[59], a9_v1[27] );
xor U3088 ( a9_v2[25], k8[57], a9_v1[25] );
xor U3089 ( a9_v2[24], k8[56], a9_v1[24] );
xor U3090 ( a8_v2[31], k7[63], a8_v1[31] );
xor U3091 ( a7_v1[30], k6[94], n1290 );
xor U3092 ( a7_v2[30], k6[62], a7_v1[30] );
xor U3093 ( a6_v1[29], k5[93], n1289 );
xor U3094 ( a6_v2[29], k5[61], a6_v1[29] );
xor U3095 ( a5_v1[28], k4[92], n1288 );
xor U3096 ( a5_v2[28], k4[60], a5_v1[28] );
xor U3097 ( a4_v1[27], k3[91], n1287 );
xor U3098 ( a4_v2[27], k3[59], a4_v1[27] );
xor U3099 ( a3_v1[26], k2[90], n1286 );
xor U3100 ( a3_v2[26], k2[58], a3_v1[26] );
xor U3101 ( a2_v1[25], k1[89], n1285 );
xor U3102 ( a2_v2[25], k1[57], a2_v1[25] );
xor U3103 ( a8_v1[31], k7[95], n1291 );
xor U3104 ( a10_v3[29], k9[29], a10_v2[29] );
xor U3105 ( a10_v3[28], k9[28], a10_v2[28] );
xor U3106 ( a10_v3[26], k9[26], a10_v2[26] );
xor U3107 ( a10_v3[25], k9[25], a10_v2[25] );
xor U3108 ( a9_v3[28], k8[28], a9_v2[28] );
xor U3109 ( a9_v3[27], k8[27], a9_v2[27] );
xor U3110 ( a9_v3[25], k8[25], a9_v2[25] );
xor U3111 ( a9_v3[24], k8[24], a9_v2[24] );
xor U3112 ( a7_v3[30], k6[30], a7_v2[30] );
xor U3113 ( a6_v3[29], k5[29], a6_v2[29] );
xor U3114 ( a5_v3[28], k4[28], a5_v2[28] );
xor U3115 ( a4_v3[27], k3[27], a4_v2[27] );
xor U3116 ( a3_v3[26], k2[26], a3_v2[26] );
xor U3117 ( a2_v3[25], k1[25], a2_v2[25] );
xor U3118 ( a8_v3[31], k7[31], a8_v2[31] );
xor U3119 ( a10_v2[3], k9[35], a10_v1[3] );
xor U3120 ( a10_v2[2], k9[34], a10_v1[2] );
xor U3121 ( a10_v2[1], k9[33], a10_v1[1] );
xor U3122 ( a10_v2[0], k9[32], a10_v1[0] );
xor U3123 ( a9_v2[3], k8[35], a9_v1[3] );
xor U3124 ( a9_v2[2], k8[34], a9_v1[2] );
xor U3125 ( a9_v2[1], k8[33], a9_v1[1] );
xor U3126 ( a9_v2[0], k8[32], a9_v1[0] );
xor U3127 ( a8_v2[3], k7[35], a8_v1[3] );
xor U3128 ( a8_v2[2], k7[34], a8_v1[2] );
xor U3129 ( a8_v2[1], k7[33], a8_v1[1] );
xor U3130 ( a8_v2[0], k7[32], a8_v1[0] );
xor U3131 ( a7_v2[3], k6[35], a7_v1[3] );
xor U3132 ( a7_v2[2], k6[34], a7_v1[2] );
xor U3133 ( a7_v2[1], k6[33], a7_v1[1] );
xor U3134 ( a7_v2[0], k6[32], a7_v1[0] );
xor U3135 ( a6_v2[3], k5[35], a6_v1[3] );
xor U3136 ( a6_v2[2], k5[34], a6_v1[2] );
xor U3137 ( a6_v2[1], k5[33], a6_v1[1] );
xor U3138 ( a6_v2[0], k5[32], a6_v1[0] );
xor U3139 ( a5_v2[3], k4[35], a5_v1[3] );
xor U3140 ( a5_v2[2], k4[34], a5_v1[2] );
xor U3141 ( a5_v2[1], k4[33], a5_v1[1] );
xor U3142 ( a5_v2[0], k4[32], a5_v1[0] );
xor U3143 ( a4_v2[3], k3[35], a4_v1[3] );
xor U3144 ( a4_v2[2], k3[34], a4_v1[2] );
xor U3145 ( a4_v2[1], k3[33], a4_v1[1] );
xor U3146 ( a4_v2[0], k3[32], a4_v1[0] );
xor U3147 ( a3_v2[3], k2[35], a3_v1[3] );
xor U3148 ( a3_v2[2], k2[34], a3_v1[2] );
xor U3149 ( a3_v2[1], k2[33], a3_v1[1] );
xor U3150 ( a3_v2[0], k2[32], a3_v1[0] );
xor U3151 ( a2_v2[3], k1[35], a2_v1[3] );
xor U3152 ( a2_v2[2], k1[34], a2_v1[2] );
xor U3153 ( a2_v2[1], k1[33], a2_v1[1] );
xor U3154 ( a2_v2[0], k1[32], a2_v1[0] );
xnor U3155 ( a10_v1[3], k9[99], n672 );
xnor U3156 ( a10_v1[2], k9[98], n669 );
xnor U3157 ( a10_v1[1], k9[97], n662 );
xnor U3158 ( a10_v1[0], k9[96], n651 );
xnor U3159 ( a9_v1[3], k8[99], n917 );
xnor U3160 ( a9_v1[2], k8[98], n914 );
xnor U3161 ( a9_v1[1], k8[97], n907 );
xnor U3162 ( a9_v1[0], k8[96], n896 );
xnor U3163 ( a8_v1[3], k7[99], n889 );
xnor U3164 ( a8_v1[2], k7[98], n887 );
xnor U3165 ( a8_v1[1], k7[97], n876 );
xnor U3166 ( a8_v1[0], k7[96], n865 );
xnor U3167 ( a7_v1[3], k6[99], n858 );
xnor U3168 ( a7_v1[2], k6[98], n856 );
xnor U3169 ( a7_v1[1], k6[97], n845 );
xnor U3170 ( a7_v1[0], k6[96], n834 );
xnor U3171 ( a6_v1[3], k5[99], n827 );
xnor U3172 ( a6_v1[2], k5[98], n824 );
xnor U3173 ( a6_v1[1], k5[97], n814 );
xnor U3174 ( a6_v1[0], k5[96], n803 );
xnor U3175 ( a5_v1[3], k4[99], n796 );
xnor U3176 ( a5_v1[2], k4[98], n793 );
xnor U3177 ( a5_v1[1], k4[97], n783 );
xnor U3178 ( a5_v1[0], k4[96], n772 );
xnor U3179 ( a4_v1[3], k3[99], n765 );
xnor U3180 ( a4_v1[2], k3[98], n762 );
xnor U3181 ( a4_v1[1], k3[97], n752 );
xnor U3182 ( a4_v1[0], k3[96], n741 );
xnor U3183 ( a3_v1[3], k2[99], n734 );
xnor U3184 ( a3_v1[2], k2[98], n731 );
xnor U3185 ( a3_v1[1], k2[97], n721 );
xnor U3186 ( a3_v1[0], k2[96], n710 );
xnor U3187 ( a2_v1[3], k1[99], n703 );
xnor U3188 ( a2_v1[2], k1[98], n700 );
xnor U3189 ( a2_v1[1], k1[97], n690 );
xnor U3190 ( a2_v1[0], k1[96], n679 );
xor U3191 ( a10_v3[3], a10_v2[3], k9[3] );
xor U3192 ( a10_v3[2], a10_v2[2], k9[2] );
xor U3193 ( a10_v3[1], a10_v2[1], k9[1] );
xor U3194 ( a10_v3[0], a10_v2[0], k9[0] );
xor U3195 ( a9_v3[3], a9_v2[3], k8[3] );
xor U3196 ( a9_v3[2], a9_v2[2], k8[2] );
xor U3197 ( a9_v3[1], a9_v2[1], k8[1] );
xor U3198 ( a9_v3[0], a9_v2[0], k8[0] );
xor U3199 ( a8_v3[3], a8_v2[3], k7[3] );
xor U3200 ( a8_v3[2], a8_v2[2], k7[2] );
xor U3201 ( a8_v3[1], a8_v2[1], k7[1] );
xor U3202 ( a8_v3[0], a8_v2[0], k7[0] );
xor U3203 ( a7_v3[3], a7_v2[3], k6[3] );
xor U3204 ( a7_v3[2], a7_v2[2], k6[2] );
xor U3205 ( a7_v3[1], a7_v2[1], k6[1] );
xor U3206 ( a7_v3[0], a7_v2[0], k6[0] );
xor U3207 ( a6_v3[3], a6_v2[3], k5[3] );
xor U3208 ( a6_v3[2], a6_v2[2], k5[2] );
xor U3209 ( a6_v3[1], a6_v2[1], k5[1] );
xor U3210 ( a6_v3[0], a6_v2[0], k5[0] );
xor U3211 ( a5_v3[3], a5_v2[3], k4[3] );
xor U3212 ( a5_v3[2], a5_v2[2], k4[2] );
xor U3213 ( a5_v3[1], a5_v2[1], k4[1] );
xor U3214 ( a5_v3[0], a5_v2[0], k4[0] );
xor U3215 ( a4_v3[3], a4_v2[3], k3[3] );
xor U3216 ( a4_v3[2], a4_v2[2], k3[2] );
xor U3217 ( a4_v3[1], a4_v2[1], k3[1] );
xor U3218 ( a4_v3[0], a4_v2[0], k3[0] );
xor U3219 ( a3_v3[3], a3_v2[3], k2[3] );
xor U3220 ( a3_v3[2], a3_v2[2], k2[2] );
xor U3221 ( a3_v3[1], a3_v2[1], k2[1] );
xor U3222 ( a3_v3[0], a3_v2[0], k2[0] );
xor U3223 ( a2_v3[3], a2_v2[3], k1[3] );
xor U3224 ( a2_v3[2], a2_v2[2], k1[2] );
xor U3225 ( a2_v3[1], a2_v2[1], k1[1] );
xor U3226 ( a2_v3[0], a2_v2[0], k1[0] );
xor U3227 ( a10_v2[31], k9[63], a10_v1[31] );
xor U3228 ( a10_v2[30], k9[62], a10_v1[30] );
xor U3229 ( a10_v2[27], k9[59], a10_v1[27] );
xor U3230 ( a10_v2[24], k9[56], a10_v1[24] );
xor U3231 ( a10_v2[23], k9[55], a10_v1[23] );
xor U3232 ( a10_v2[22], k9[54], a10_v1[22] );
xor U3233 ( a10_v2[21], k9[53], a10_v1[21] );
xor U3234 ( a10_v2[20], k9[52], a10_v1[20] );
xor U3235 ( a10_v2[19], k9[51], a10_v1[19] );
xor U3236 ( a10_v2[18], k9[50], a10_v1[18] );
xor U3237 ( a10_v2[17], k9[49], a10_v1[17] );
xor U3238 ( a10_v2[16], k9[48], a10_v1[16] );
xor U3239 ( a10_v2[15], k9[47], a10_v1[15] );
xor U3240 ( a10_v2[14], k9[46], a10_v1[14] );
xor U3241 ( a10_v2[13], k9[45], a10_v1[13] );
xor U3242 ( a10_v2[12], k9[44], a10_v1[12] );
xor U3243 ( a10_v2[11], k9[43], a10_v1[11] );
xor U3244 ( a10_v2[10], k9[42], a10_v1[10] );
xor U3245 ( a10_v2[9], k9[41], a10_v1[9] );
xor U3246 ( a10_v2[8], k9[40], a10_v1[8] );
xor U3247 ( a10_v2[7], k9[39], a10_v1[7] );
xor U3248 ( a10_v2[6], k9[38], a10_v1[6] );
xor U3249 ( a10_v2[5], k9[37], a10_v1[5] );
xor U3250 ( a10_v2[4], k9[36], a10_v1[4] );
xor U3251 ( a9_v2[31], k8[63], a9_v1[31] );
xor U3252 ( a9_v2[30], k8[62], a9_v1[30] );
xor U3253 ( a9_v2[29], k8[61], a9_v1[29] );
xor U3254 ( a9_v2[26], k8[58], a9_v1[26] );
xor U3255 ( a9_v2[23], k8[55], a9_v1[23] );
xor U3256 ( a9_v2[22], k8[54], a9_v1[22] );
xor U3257 ( a9_v2[21], k8[53], a9_v1[21] );
xor U3258 ( a9_v2[20], k8[52], a9_v1[20] );
xor U3259 ( a9_v2[19], k8[51], a9_v1[19] );
xor U3260 ( a9_v2[18], k8[50], a9_v1[18] );
xor U3261 ( a9_v2[17], k8[49], a9_v1[17] );
xor U3262 ( a9_v2[16], k8[48], a9_v1[16] );
xor U3263 ( a9_v2[15], k8[47], a9_v1[15] );
xor U3264 ( a9_v2[14], k8[46], a9_v1[14] );
xor U3265 ( a9_v2[13], k8[45], a9_v1[13] );
xor U3266 ( a9_v2[12], k8[44], a9_v1[12] );
xor U3267 ( a9_v2[11], k8[43], a9_v1[11] );
xor U3268 ( a9_v2[10], k8[42], a9_v1[10] );
xor U3269 ( a9_v2[9], k8[41], a9_v1[9] );
xor U3270 ( a9_v2[8], k8[40], a9_v1[8] );
xor U3271 ( a9_v2[7], k8[39], a9_v1[7] );
xor U3272 ( a9_v2[6], k8[38], a9_v1[6] );
xor U3273 ( a9_v2[5], k8[37], a9_v1[5] );
xor U3274 ( a9_v2[4], k8[36], a9_v1[4] );
xor U3275 ( a8_v2[30], k7[62], a8_v1[30] );
xor U3276 ( a8_v2[29], k7[61], a8_v1[29] );
xor U3277 ( a8_v2[28], k7[60], a8_v1[28] );
xor U3278 ( a8_v2[27], k7[59], a8_v1[27] );
xor U3279 ( a8_v2[26], k7[58], a8_v1[26] );
xor U3280 ( a8_v2[25], k7[57], a8_v1[25] );
xor U3281 ( a8_v2[24], k7[56], a8_v1[24] );
xor U3282 ( a8_v2[23], k7[55], a8_v1[23] );
xor U3283 ( a8_v2[22], k7[54], a8_v1[22] );
xor U3284 ( a8_v2[21], k7[53], a8_v1[21] );
xor U3285 ( a8_v2[20], k7[52], a8_v1[20] );
xor U3286 ( a8_v2[19], k7[51], a8_v1[19] );
xor U3287 ( a8_v2[18], k7[50], a8_v1[18] );
xor U3288 ( a8_v2[17], k7[49], a8_v1[17] );
xor U3289 ( a8_v2[16], k7[48], a8_v1[16] );
xor U3290 ( a8_v2[15], k7[47], a8_v1[15] );
xor U3291 ( a8_v2[14], k7[46], a8_v1[14] );
xor U3292 ( a8_v2[13], k7[45], a8_v1[13] );
xor U3293 ( a8_v2[12], k7[44], a8_v1[12] );
xor U3294 ( a8_v2[11], k7[43], a8_v1[11] );
xor U3295 ( a8_v2[10], k7[42], a8_v1[10] );
xor U3296 ( a8_v2[9], k7[41], a8_v1[9] );
xor U3297 ( a8_v2[8], k7[40], a8_v1[8] );
xor U3298 ( a8_v2[7], k7[39], a8_v1[7] );
xor U3299 ( a8_v2[6], k7[38], a8_v1[6] );
xor U3300 ( a8_v2[5], k7[37], a8_v1[5] );
xor U3301 ( a8_v2[4], k7[36], a8_v1[4] );
xor U3302 ( a7_v2[31], k6[63], a7_v1[31] );
xor U3303 ( a7_v2[29], k6[61], a7_v1[29] );
xor U3304 ( a7_v2[28], k6[60], a7_v1[28] );
xor U3305 ( a7_v2[27], k6[59], a7_v1[27] );
xor U3306 ( a7_v2[26], k6[58], a7_v1[26] );
xor U3307 ( a7_v2[25], k6[57], a7_v1[25] );
xor U3308 ( a7_v2[24], k6[56], a7_v1[24] );
xor U3309 ( a7_v2[23], k6[55], a7_v1[23] );
xor U3310 ( a7_v2[22], k6[54], a7_v1[22] );
xor U3311 ( a7_v2[21], k6[53], a7_v1[21] );
xor U3312 ( a7_v2[20], k6[52], a7_v1[20] );
xor U3313 ( a7_v2[19], k6[51], a7_v1[19] );
xor U3314 ( a7_v2[18], k6[50], a7_v1[18] );
xor U3315 ( a7_v2[17], k6[49], a7_v1[17] );
xor U3316 ( a7_v2[16], k6[48], a7_v1[16] );
xor U3317 ( a7_v2[15], k6[47], a7_v1[15] );
xor U3318 ( a7_v2[14], k6[46], a7_v1[14] );
xor U3319 ( a7_v2[13], k6[45], a7_v1[13] );
xor U3320 ( a7_v2[12], k6[44], a7_v1[12] );
xor U3321 ( a7_v2[11], k6[43], a7_v1[11] );
xor U3322 ( a7_v2[10], k6[42], a7_v1[10] );
xor U3323 ( a7_v2[9], k6[41], a7_v1[9] );
xor U3324 ( a7_v2[8], k6[40], a7_v1[8] );
xor U3325 ( a7_v2[7], k6[39], a7_v1[7] );
xor U3326 ( a7_v2[6], k6[38], a7_v1[6] );
xor U3327 ( a7_v2[5], k6[37], a7_v1[5] );
xor U3328 ( a7_v2[4], k6[36], a7_v1[4] );
xor U3329 ( a6_v2[31], k5[63], a6_v1[31] );
xor U3330 ( a6_v2[30], k5[62], a6_v1[30] );
xor U3331 ( a6_v2[28], k5[60], a6_v1[28] );
xor U3332 ( a6_v2[27], k5[59], a6_v1[27] );
xor U3333 ( a6_v2[26], k5[58], a6_v1[26] );
xor U3334 ( a6_v2[25], k5[57], a6_v1[25] );
xor U3335 ( a6_v2[24], k5[56], a6_v1[24] );
xor U3336 ( a6_v2[23], k5[55], a6_v1[23] );
xor U3337 ( a6_v2[22], k5[54], a6_v1[22] );
xor U3338 ( a6_v2[21], k5[53], a6_v1[21] );
xor U3339 ( a6_v2[20], k5[52], a6_v1[20] );
xor U3340 ( a6_v2[19], k5[51], a6_v1[19] );
xor U3341 ( a6_v2[18], k5[50], a6_v1[18] );
xor U3342 ( a6_v2[17], k5[49], a6_v1[17] );
xor U3343 ( a6_v2[16], k5[48], a6_v1[16] );
xor U3344 ( a6_v2[15], k5[47], a6_v1[15] );
xor U3345 ( a6_v2[14], k5[46], a6_v1[14] );
xor U3346 ( a6_v2[13], k5[45], a6_v1[13] );
xor U3347 ( a6_v2[12], k5[44], a6_v1[12] );
xor U3348 ( a6_v2[11], k5[43], a6_v1[11] );
xor U3349 ( a6_v2[10], k5[42], a6_v1[10] );
xor U3350 ( a6_v2[9], k5[41], a6_v1[9] );
xor U3351 ( a6_v2[8], k5[40], a6_v1[8] );
xor U3352 ( a6_v2[7], k5[39], a6_v1[7] );
xor U3353 ( a6_v2[6], k5[38], a6_v1[6] );
xor U3354 ( a6_v2[5], k5[37], a6_v1[5] );
xor U3355 ( a6_v2[4], k5[36], a6_v1[4] );
xor U3356 ( a5_v2[31], k4[63], a5_v1[31] );
xor U3357 ( a5_v2[30], k4[62], a5_v1[30] );
xor U3358 ( a5_v2[29], k4[61], a5_v1[29] );
xor U3359 ( a5_v2[27], k4[59], a5_v1[27] );
xor U3360 ( a5_v2[26], k4[58], a5_v1[26] );
xor U3361 ( a5_v2[25], k4[57], a5_v1[25] );
xor U3362 ( a5_v2[24], k4[56], a5_v1[24] );
xor U3363 ( a5_v2[23], k4[55], a5_v1[23] );
xor U3364 ( a5_v2[22], k4[54], a5_v1[22] );
xor U3365 ( a5_v2[21], k4[53], a5_v1[21] );
xor U3366 ( a5_v2[20], k4[52], a5_v1[20] );
xor U3367 ( a5_v2[19], k4[51], a5_v1[19] );
xor U3368 ( a5_v2[18], k4[50], a5_v1[18] );
xor U3369 ( a5_v2[17], k4[49], a5_v1[17] );
xor U3370 ( a5_v2[16], k4[48], a5_v1[16] );
xor U3371 ( a5_v2[15], k4[47], a5_v1[15] );
xor U3372 ( a5_v2[14], k4[46], a5_v1[14] );
xor U3373 ( a5_v2[13], k4[45], a5_v1[13] );
xor U3374 ( a5_v2[12], k4[44], a5_v1[12] );
xor U3375 ( a5_v2[11], k4[43], a5_v1[11] );
xor U3376 ( a5_v2[10], k4[42], a5_v1[10] );
xor U3377 ( a5_v2[9], k4[41], a5_v1[9] );
xor U3378 ( a5_v2[8], k4[40], a5_v1[8] );
xor U3379 ( a5_v2[7], k4[39], a5_v1[7] );
xor U3380 ( a5_v2[6], k4[38], a5_v1[6] );
xor U3381 ( a5_v2[5], k4[37], a5_v1[5] );
xor U3382 ( a5_v2[4], k4[36], a5_v1[4] );
xor U3383 ( a4_v2[31], k3[63], a4_v1[31] );
xor U3384 ( a4_v2[30], k3[62], a4_v1[30] );
xor U3385 ( a4_v2[29], k3[61], a4_v1[29] );
xor U3386 ( a4_v2[28], k3[60], a4_v1[28] );
xor U3387 ( a4_v2[26], k3[58], a4_v1[26] );
xor U3388 ( a4_v2[25], k3[57], a4_v1[25] );
xor U3389 ( a4_v2[24], k3[56], a4_v1[24] );
xor U3390 ( a4_v2[23], k3[55], a4_v1[23] );
xor U3391 ( a4_v2[22], k3[54], a4_v1[22] );
xor U3392 ( a4_v2[21], k3[53], a4_v1[21] );
xor U3393 ( a4_v2[20], k3[52], a4_v1[20] );
xor U3394 ( a4_v2[19], k3[51], a4_v1[19] );
xor U3395 ( a4_v2[18], k3[50], a4_v1[18] );
xor U3396 ( a4_v2[17], k3[49], a4_v1[17] );
xor U3397 ( a4_v2[16], k3[48], a4_v1[16] );
xor U3398 ( a4_v2[15], k3[47], a4_v1[15] );
xor U3399 ( a4_v2[14], k3[46], a4_v1[14] );
xor U3400 ( a4_v2[13], k3[45], a4_v1[13] );
xor U3401 ( a4_v2[12], k3[44], a4_v1[12] );
xor U3402 ( a4_v2[11], k3[43], a4_v1[11] );
xor U3403 ( a4_v2[10], k3[42], a4_v1[10] );
xor U3404 ( a4_v2[9], k3[41], a4_v1[9] );
xor U3405 ( a4_v2[8], k3[40], a4_v1[8] );
xor U3406 ( a4_v2[7], k3[39], a4_v1[7] );
xor U3407 ( a4_v2[6], k3[38], a4_v1[6] );
xor U3408 ( a4_v2[5], k3[37], a4_v1[5] );
xor U3409 ( a4_v2[4], k3[36], a4_v1[4] );
xor U3410 ( a3_v2[31], k2[63], a3_v1[31] );
xor U3411 ( a3_v2[30], k2[62], a3_v1[30] );
xor U3412 ( a3_v2[29], k2[61], a3_v1[29] );
xor U3413 ( a3_v2[28], k2[60], a3_v1[28] );
xor U3414 ( a3_v2[27], k2[59], a3_v1[27] );
xor U3415 ( a3_v2[25], k2[57], a3_v1[25] );
xor U3416 ( a3_v2[24], k2[56], a3_v1[24] );
xor U3417 ( a3_v2[23], k2[55], a3_v1[23] );
xor U3418 ( a3_v2[22], k2[54], a3_v1[22] );
xor U3419 ( a3_v2[21], k2[53], a3_v1[21] );
xor U3420 ( a3_v2[20], k2[52], a3_v1[20] );
xor U3421 ( a3_v2[19], k2[51], a3_v1[19] );
xor U3422 ( a3_v2[18], k2[50], a3_v1[18] );
xor U3423 ( a3_v2[17], k2[49], a3_v1[17] );
xor U3424 ( a3_v2[16], k2[48], a3_v1[16] );
xor U3425 ( a3_v2[15], k2[47], a3_v1[15] );
xor U3426 ( a3_v2[14], k2[46], a3_v1[14] );
xor U3427 ( a3_v2[13], k2[45], a3_v1[13] );
xor U3428 ( a3_v2[12], k2[44], a3_v1[12] );
xor U3429 ( a3_v2[11], k2[43], a3_v1[11] );
xor U3430 ( a3_v2[10], k2[42], a3_v1[10] );
xor U3431 ( a3_v2[9], k2[41], a3_v1[9] );
xor U3432 ( a3_v2[8], k2[40], a3_v1[8] );
xor U3433 ( a3_v2[7], k2[39], a3_v1[7] );
xor U3434 ( a3_v2[6], k2[38], a3_v1[6] );
xor U3435 ( a3_v2[5], k2[37], a3_v1[5] );
xor U3436 ( a3_v2[4], k2[36], a3_v1[4] );
xor U3437 ( a2_v2[31], k1[63], a2_v1[31] );
xor U3438 ( a2_v2[30], k1[62], a2_v1[30] );
xor U3439 ( a2_v2[29], k1[61], a2_v1[29] );
xor U3440 ( a2_v2[28], k1[60], a2_v1[28] );
xor U3441 ( a2_v2[27], k1[59], a2_v1[27] );
xor U3442 ( a2_v2[26], k1[58], a2_v1[26] );
xor U3443 ( a2_v2[24], k1[56], a2_v1[24] );
xor U3444 ( a2_v2[23], k1[55], a2_v1[23] );
xor U3445 ( a2_v2[22], k1[54], a2_v1[22] );
xor U3446 ( a2_v2[21], k1[53], a2_v1[21] );
xor U3447 ( a2_v2[20], k1[52], a2_v1[20] );
xor U3448 ( a2_v2[19], k1[51], a2_v1[19] );
xor U3449 ( a2_v2[18], k1[50], a2_v1[18] );
xor U3450 ( a2_v2[17], k1[49], a2_v1[17] );
xor U3451 ( a2_v2[16], k1[48], a2_v1[16] );
xor U3452 ( a2_v2[15], k1[47], a2_v1[15] );
xor U3453 ( a2_v2[14], k1[46], a2_v1[14] );
xor U3454 ( a2_v2[13], k1[45], a2_v1[13] );
xor U3455 ( a2_v2[12], k1[44], a2_v1[12] );
xor U3456 ( a2_v2[11], k1[43], a2_v1[11] );
xor U3457 ( a2_v2[10], k1[42], a2_v1[10] );
xor U3458 ( a2_v2[9], k1[41], a2_v1[9] );
xor U3459 ( a2_v2[8], k1[40], a2_v1[8] );
xor U3460 ( a2_v2[7], k1[39], a2_v1[7] );
xor U3461 ( a2_v2[6], k1[38], a2_v1[6] );
xor U3462 ( a2_v2[5], k1[37], a2_v1[5] );
xor U3463 ( a2_v2[4], k1[36], a2_v1[4] );
xnor U3464 ( a10_v1[30], k9[94], n670 );
xnor U3465 ( a10_v1[27], k9[91], n668 );
xnor U3466 ( a10_v1[24], k9[88], n667 );
xnor U3467 ( a10_v1[23], k9[87], n666 );
xnor U3468 ( a10_v1[22], k9[86], n665 );
xnor U3469 ( a10_v1[21], k9[85], n664 );
xnor U3470 ( a10_v1[20], k9[84], n663 );
xnor U3471 ( a10_v1[19], k9[83], n661 );
xnor U3472 ( a10_v1[18], k9[82], n660 );
xnor U3473 ( a10_v1[17], k9[81], n659 );
xnor U3474 ( a10_v1[16], k9[80], n658 );
xnor U3475 ( a10_v1[15], k9[79], n657 );
xnor U3476 ( a10_v1[14], k9[78], n656 );
xnor U3477 ( a10_v1[13], k9[77], n655 );
xnor U3478 ( a10_v1[12], k9[76], n654 );
xnor U3479 ( a10_v1[11], k9[75], n653 );
xnor U3480 ( a10_v1[10], k9[74], n652 );
xnor U3481 ( a10_v1[9], k9[73], n678 );
xnor U3482 ( a10_v1[8], k9[72], n677 );
xnor U3483 ( a10_v1[7], k9[71], n676 );
xnor U3484 ( a10_v1[6], k9[70], n675 );
xnor U3485 ( a10_v1[5], k9[69], n674 );
xnor U3486 ( a10_v1[4], k9[68], n673 );
xnor U3487 ( a9_v1[30], k8[94], n915 );
xnor U3488 ( a9_v1[29], k8[93], n913 );
xnor U3489 ( a9_v1[26], k8[90], n912 );
xnor U3490 ( a9_v1[23], k8[87], n911 );
xnor U3491 ( a9_v1[22], k8[86], n910 );
xnor U3492 ( a9_v1[21], k8[85], n909 );
xnor U3493 ( a9_v1[20], k8[84], n908 );
xnor U3494 ( a9_v1[19], k8[83], n906 );
xnor U3495 ( a9_v1[18], k8[82], n905 );
xnor U3496 ( a9_v1[17], k8[81], n904 );
xnor U3497 ( a9_v1[16], k8[80], n903 );
xnor U3498 ( a9_v1[15], k8[79], n902 );
xnor U3499 ( a9_v1[14], k8[78], n901 );
xnor U3500 ( a9_v1[13], k8[77], n900 );
xnor U3501 ( a9_v1[12], k8[76], n899 );
xnor U3502 ( a9_v1[11], k8[75], n898 );
xnor U3503 ( a9_v1[10], k8[74], n897 );
xnor U3504 ( a9_v1[9], k8[73], n923 );
xnor U3505 ( a9_v1[8], k8[72], n922 );
xnor U3506 ( a9_v1[7], k8[71], n921 );
xnor U3507 ( a9_v1[6], k8[70], n920 );
xnor U3508 ( a9_v1[5], k8[69], n919 );
xnor U3509 ( a9_v1[4], k8[68], n918 );
xnor U3510 ( a8_v1[30], k7[94], n888 );
xnor U3511 ( a8_v1[29], k7[93], n886 );
xnor U3512 ( a8_v1[28], k7[92], n885 );
xnor U3513 ( a8_v1[27], k7[91], n884 );
xnor U3514 ( a8_v1[26], k7[90], n883 );
xnor U3515 ( a8_v1[25], k7[89], n882 );
xnor U3516 ( a8_v1[24], k7[88], n881 );
xnor U3517 ( a8_v1[23], k7[87], n880 );
xnor U3518 ( a8_v1[22], k7[86], n879 );
xnor U3519 ( a8_v1[21], k7[85], n878 );
xnor U3520 ( a8_v1[20], k7[84], n877 );
xnor U3521 ( a8_v1[19], k7[83], n875 );
xnor U3522 ( a8_v1[18], k7[82], n874 );
xnor U3523 ( a8_v1[17], k7[81], n873 );
xnor U3524 ( a8_v1[16], k7[80], n872 );
xnor U3525 ( a8_v1[15], k7[79], n871 );
xnor U3526 ( a8_v1[14], k7[78], n870 );
xnor U3527 ( a8_v1[13], k7[77], n869 );
xnor U3528 ( a8_v1[12], k7[76], n868 );
xnor U3529 ( a8_v1[11], k7[75], n867 );
xnor U3530 ( a8_v1[10], k7[74], n866 );
xnor U3531 ( a8_v1[9], k7[73], n895 );
xnor U3532 ( a8_v1[8], k7[72], n894 );
xnor U3533 ( a8_v1[7], k7[71], n893 );
xnor U3534 ( a8_v1[6], k7[70], n892 );
xnor U3535 ( a8_v1[5], k7[69], n891 );
xnor U3536 ( a8_v1[4], k7[68], n890 );
xnor U3537 ( a7_v1[29], k6[93], n855 );
xnor U3538 ( a7_v1[28], k6[92], n854 );
xnor U3539 ( a7_v1[27], k6[91], n853 );
xnor U3540 ( a7_v1[26], k6[90], n852 );
xnor U3541 ( a7_v1[25], k6[89], n851 );
xnor U3542 ( a7_v1[24], k6[88], n850 );
xnor U3543 ( a7_v1[23], k6[87], n849 );
xnor U3544 ( a7_v1[22], k6[86], n848 );
xnor U3545 ( a7_v1[21], k6[85], n847 );
xnor U3546 ( a7_v1[20], k6[84], n846 );
xnor U3547 ( a7_v1[19], k6[83], n844 );
xnor U3548 ( a7_v1[18], k6[82], n843 );
xnor U3549 ( a7_v1[17], k6[81], n842 );
xnor U3550 ( a7_v1[16], k6[80], n841 );
xnor U3551 ( a7_v1[15], k6[79], n840 );
xnor U3552 ( a7_v1[14], k6[78], n839 );
xnor U3553 ( a7_v1[13], k6[77], n838 );
xnor U3554 ( a7_v1[12], k6[76], n837 );
xnor U3555 ( a7_v1[11], k6[75], n836 );
xnor U3556 ( a7_v1[10], k6[74], n835 );
xnor U3557 ( a7_v1[9], k6[73], n864 );
xnor U3558 ( a7_v1[8], k6[72], n863 );
xnor U3559 ( a7_v1[7], k6[71], n862 );
xnor U3560 ( a7_v1[6], k6[70], n861 );
xnor U3561 ( a7_v1[5], k6[69], n860 );
xnor U3562 ( a7_v1[4], k6[68], n859 );
xnor U3563 ( a6_v1[30], k5[94], n825 );
xnor U3564 ( a6_v1[28], k5[92], n823 );
xnor U3565 ( a6_v1[27], k5[91], n822 );
xnor U3566 ( a6_v1[26], k5[90], n821 );
xnor U3567 ( a6_v1[25], k5[89], n820 );
xnor U3568 ( a6_v1[24], k5[88], n819 );
xnor U3569 ( a6_v1[23], k5[87], n818 );
xnor U3570 ( a6_v1[22], k5[86], n817 );
xnor U3571 ( a6_v1[21], k5[85], n816 );
xnor U3572 ( a6_v1[20], k5[84], n815 );
xnor U3573 ( a6_v1[19], k5[83], n813 );
xnor U3574 ( a6_v1[18], k5[82], n812 );
xnor U3575 ( a6_v1[17], k5[81], n811 );
xnor U3576 ( a6_v1[16], k5[80], n810 );
xnor U3577 ( a6_v1[15], k5[79], n809 );
xnor U3578 ( a6_v1[14], k5[78], n808 );
xnor U3579 ( a6_v1[13], k5[77], n807 );
xnor U3580 ( a6_v1[12], k5[76], n806 );
xnor U3581 ( a6_v1[11], k5[75], n805 );
xnor U3582 ( a6_v1[10], k5[74], n804 );
xnor U3583 ( a6_v1[9], k5[73], n833 );
xnor U3584 ( a6_v1[8], k5[72], n832 );
xnor U3585 ( a6_v1[7], k5[71], n831 );
xnor U3586 ( a6_v1[6], k5[70], n830 );
xnor U3587 ( a6_v1[5], k5[69], n829 );
xnor U3588 ( a6_v1[4], k5[68], n828 );
xnor U3589 ( a5_v1[30], k4[94], n794 );
xnor U3590 ( a5_v1[29], k4[93], n792 );
xnor U3591 ( a5_v1[27], k4[91], n791 );
xnor U3592 ( a5_v1[26], k4[90], n790 );
xnor U3593 ( a5_v1[25], k4[89], n789 );
xnor U3594 ( a5_v1[24], k4[88], n788 );
xnor U3595 ( a5_v1[23], k4[87], n787 );
xnor U3596 ( a5_v1[22], k4[86], n786 );
xnor U3597 ( a5_v1[21], k4[85], n785 );
xnor U3598 ( a5_v1[20], k4[84], n784 );
xnor U3599 ( a5_v1[19], k4[83], n782 );
xnor U3600 ( a5_v1[18], k4[82], n781 );
xnor U3601 ( a5_v1[17], k4[81], n780 );
xnor U3602 ( a5_v1[16], k4[80], n779 );
xnor U3603 ( a5_v1[15], k4[79], n778 );
xnor U3604 ( a5_v1[14], k4[78], n777 );
xnor U3605 ( a5_v1[13], k4[77], n776 );
xnor U3606 ( a5_v1[12], k4[76], n775 );
xnor U3607 ( a5_v1[11], k4[75], n774 );
xnor U3608 ( a5_v1[10], k4[74], n773 );
xnor U3609 ( a5_v1[9], k4[73], n802 );
xnor U3610 ( a5_v1[8], k4[72], n801 );
xnor U3611 ( a5_v1[7], k4[71], n800 );
xnor U3612 ( a5_v1[6], k4[70], n799 );
xnor U3613 ( a5_v1[5], k4[69], n798 );
xnor U3614 ( a5_v1[4], k4[68], n797 );
xnor U3615 ( a4_v1[30], k3[94], n763 );
xnor U3616 ( a4_v1[29], k3[93], n761 );
xnor U3617 ( a4_v1[28], k3[92], n760 );
xnor U3618 ( a4_v1[26], k3[90], n759 );
xnor U3619 ( a4_v1[25], k3[89], n758 );
xnor U3620 ( a4_v1[24], k3[88], n757 );
xnor U3621 ( a4_v1[23], k3[87], n756 );
xnor U3622 ( a4_v1[22], k3[86], n755 );
xnor U3623 ( a4_v1[21], k3[85], n754 );
xnor U3624 ( a4_v1[20], k3[84], n753 );
xnor U3625 ( a4_v1[19], k3[83], n751 );
xnor U3626 ( a4_v1[18], k3[82], n750 );
xnor U3627 ( a4_v1[17], k3[81], n749 );
xnor U3628 ( a4_v1[16], k3[80], n748 );
xnor U3629 ( a4_v1[15], k3[79], n747 );
xnor U3630 ( a4_v1[14], k3[78], n746 );
xnor U3631 ( a4_v1[13], k3[77], n745 );
xnor U3632 ( a4_v1[12], k3[76], n744 );
xnor U3633 ( a4_v1[11], k3[75], n743 );
xnor U3634 ( a4_v1[10], k3[74], n742 );
xnor U3635 ( a4_v1[9], k3[73], n771 );
xnor U3636 ( a4_v1[8], k3[72], n770 );
xnor U3637 ( a4_v1[7], k3[71], n769 );
xnor U3638 ( a4_v1[6], k3[70], n768 );
xnor U3639 ( a4_v1[5], k3[69], n767 );
xnor U3640 ( a4_v1[4], k3[68], n766 );
xnor U3641 ( a3_v1[30], k2[94], n732 );
xnor U3642 ( a3_v1[29], k2[93], n730 );
xnor U3643 ( a3_v1[28], k2[92], n729 );
xnor U3644 ( a3_v1[27], k2[91], n728 );
xnor U3645 ( a3_v1[25], k2[89], n727 );
xnor U3646 ( a3_v1[24], k2[88], n726 );
xnor U3647 ( a3_v1[23], k2[87], n725 );
xnor U3648 ( a3_v1[22], k2[86], n724 );
xnor U3649 ( a3_v1[21], k2[85], n723 );
xnor U3650 ( a3_v1[20], k2[84], n722 );
xnor U3651 ( a3_v1[19], k2[83], n720 );
xnor U3652 ( a3_v1[18], k2[82], n719 );
xnor U3653 ( a3_v1[17], k2[81], n718 );
xnor U3654 ( a3_v1[16], k2[80], n717 );
xnor U3655 ( a3_v1[15], k2[79], n716 );
xnor U3656 ( a3_v1[14], k2[78], n715 );
xnor U3657 ( a3_v1[13], k2[77], n714 );
xnor U3658 ( a3_v1[12], k2[76], n713 );
xnor U3659 ( a3_v1[11], k2[75], n712 );
xnor U3660 ( a3_v1[10], k2[74], n711 );
xnor U3661 ( a3_v1[9], k2[73], n740 );
xnor U3662 ( a3_v1[8], k2[72], n739 );
xnor U3663 ( a3_v1[7], k2[71], n738 );
xnor U3664 ( a3_v1[6], k2[70], n737 );
xnor U3665 ( a3_v1[5], k2[69], n736 );
xnor U3666 ( a3_v1[4], k2[68], n735 );
xnor U3667 ( a2_v1[30], k1[94], n701 );
xnor U3668 ( a2_v1[29], k1[93], n699 );
xnor U3669 ( a2_v1[28], k1[92], n698 );
xnor U3670 ( a2_v1[27], k1[91], n697 );
xnor U3671 ( a2_v1[26], k1[90], n696 );
xnor U3672 ( a2_v1[24], k1[88], n695 );
xnor U3673 ( a2_v1[23], k1[87], n694 );
xnor U3674 ( a2_v1[22], k1[86], n693 );
xnor U3675 ( a2_v1[21], k1[85], n692 );
xnor U3676 ( a2_v1[20], k1[84], n691 );
xnor U3677 ( a2_v1[19], k1[83], n689 );
xnor U3678 ( a2_v1[18], k1[82], n688 );
xnor U3679 ( a2_v1[17], k1[81], n687 );
xnor U3680 ( a2_v1[16], k1[80], n686 );
xnor U3681 ( a2_v1[15], k1[79], n685 );
xnor U3682 ( a2_v1[14], k1[78], n684 );
xnor U3683 ( a2_v1[13], k1[77], n683 );
xnor U3684 ( a2_v1[12], k1[76], n682 );
xnor U3685 ( a2_v1[11], k1[75], n681 );
xnor U3686 ( a2_v1[10], k1[74], n680 );
xnor U3687 ( a2_v1[9], k1[73], n709 );
xnor U3688 ( a2_v1[8], k1[72], n708 );
xnor U3689 ( a2_v1[7], k1[71], n707 );
xnor U3690 ( a2_v1[6], k1[70], n706 );
xnor U3691 ( a2_v1[5], k1[69], n705 );
xnor U3692 ( a2_v1[4], k1[68], n704 );
xnor U3693 ( a2_v1[31], k1[95], n702 );
xnor U3694 ( a3_v1[31], k2[95], n733 );
xnor U3695 ( a4_v1[31], k3[95], n764 );
xnor U3696 ( a5_v1[31], k4[95], n795 );
xnor U3697 ( a6_v1[31], k5[95], n826 );
xnor U3698 ( a7_v1[31], k6[95], n857 );
xnor U3699 ( a9_v1[31], k8[95], n916 );
xnor U3700 ( a10_v1[31], k9[95], n671 );
xor U3701 ( a10_v3[31], a10_v2[31], k9[31] );
xor U3702 ( a10_v3[30], a10_v2[30], k9[30] );
xor U3703 ( a10_v3[27], a10_v2[27], k9[27] );
xor U3704 ( a10_v3[24], a10_v2[24], k9[24] );
xor U3705 ( a10_v3[23], a10_v2[23], k9[23] );
xor U3706 ( a10_v3[22], a10_v2[22], k9[22] );
xor U3707 ( a10_v3[21], a10_v2[21], k9[21] );
xor U3708 ( a10_v3[20], a10_v2[20], k9[20] );
xor U3709 ( a10_v3[19], a10_v2[19], k9[19] );
xor U3710 ( a10_v3[18], a10_v2[18], k9[18] );
xor U3711 ( a10_v3[17], a10_v2[17], k9[17] );
xor U3712 ( a10_v3[16], a10_v2[16], k9[16] );
xor U3713 ( a10_v3[15], a10_v2[15], k9[15] );
xor U3714 ( a10_v3[14], a10_v2[14], k9[14] );
xor U3715 ( a10_v3[13], a10_v2[13], k9[13] );
xor U3716 ( a10_v3[12], a10_v2[12], k9[12] );
xor U3717 ( a10_v3[11], a10_v2[11], k9[11] );
xor U3718 ( a10_v3[10], a10_v2[10], k9[10] );
xor U3719 ( a10_v3[9], a10_v2[9], k9[9] );
xor U3720 ( a10_v3[8], a10_v2[8], k9[8] );
xor U3721 ( a10_v3[7], a10_v2[7], k9[7] );
xor U3722 ( a10_v3[6], a10_v2[6], k9[6] );
xor U3723 ( a10_v3[5], a10_v2[5], k9[5] );
xor U3724 ( a10_v3[4], a10_v2[4], k9[4] );
xor U3725 ( a9_v3[30], a9_v2[30], k8[30] );
xor U3726 ( a9_v3[29], a9_v2[29], k8[29] );
xor U3727 ( a9_v3[26], a9_v2[26], k8[26] );
xor U3728 ( a9_v3[23], a9_v2[23], k8[23] );
xor U3729 ( a9_v3[22], a9_v2[22], k8[22] );
xor U3730 ( a9_v3[21], a9_v2[21], k8[21] );
xor U3731 ( a9_v3[20], a9_v2[20], k8[20] );
xor U3732 ( a9_v3[19], a9_v2[19], k8[19] );
xor U3733 ( a9_v3[18], a9_v2[18], k8[18] );
xor U3734 ( a9_v3[17], a9_v2[17], k8[17] );
xor U3735 ( a9_v3[16], a9_v2[16], k8[16] );
xor U3736 ( a9_v3[15], a9_v2[15], k8[15] );
xor U3737 ( a9_v3[14], a9_v2[14], k8[14] );
xor U3738 ( a9_v3[13], a9_v2[13], k8[13] );
xor U3739 ( a9_v3[12], a9_v2[12], k8[12] );
xor U3740 ( a9_v3[11], a9_v2[11], k8[11] );
xor U3741 ( a9_v3[10], a9_v2[10], k8[10] );
xor U3742 ( a9_v3[9], a9_v2[9], k8[9] );
xor U3743 ( a9_v3[8], a9_v2[8], k8[8] );
xor U3744 ( a9_v3[7], a9_v2[7], k8[7] );
xor U3745 ( a9_v3[6], a9_v2[6], k8[6] );
xor U3746 ( a9_v3[5], a9_v2[5], k8[5] );
xor U3747 ( a9_v3[4], a9_v2[4], k8[4] );
xor U3748 ( a8_v3[30], a8_v2[30], k7[30] );
xor U3749 ( a8_v3[29], a8_v2[29], k7[29] );
xor U3750 ( a8_v3[28], a8_v2[28], k7[28] );
xor U3751 ( a8_v3[27], a8_v2[27], k7[27] );
xor U3752 ( a8_v3[26], a8_v2[26], k7[26] );
xor U3753 ( a8_v3[25], a8_v2[25], k7[25] );
xor U3754 ( a8_v3[24], a8_v2[24], k7[24] );
xor U3755 ( a8_v3[23], a8_v2[23], k7[23] );
xor U3756 ( a8_v3[22], a8_v2[22], k7[22] );
xor U3757 ( a8_v3[21], a8_v2[21], k7[21] );
xor U3758 ( a8_v3[20], a8_v2[20], k7[20] );
xor U3759 ( a8_v3[19], a8_v2[19], k7[19] );
xor U3760 ( a8_v3[18], a8_v2[18], k7[18] );
xor U3761 ( a8_v3[17], a8_v2[17], k7[17] );
xor U3762 ( a8_v3[16], a8_v2[16], k7[16] );
xor U3763 ( a8_v3[15], a8_v2[15], k7[15] );
xor U3764 ( a8_v3[14], a8_v2[14], k7[14] );
xor U3765 ( a8_v3[13], a8_v2[13], k7[13] );
xor U3766 ( a8_v3[12], a8_v2[12], k7[12] );
xor U3767 ( a8_v3[11], a8_v2[11], k7[11] );
xor U3768 ( a8_v3[10], a8_v2[10], k7[10] );
xor U3769 ( a8_v3[9], a8_v2[9], k7[9] );
xor U3770 ( a8_v3[8], a8_v2[8], k7[8] );
xor U3771 ( a8_v3[7], a8_v2[7], k7[7] );
xor U3772 ( a8_v3[6], a8_v2[6], k7[6] );
xor U3773 ( a8_v3[5], a8_v2[5], k7[5] );
xor U3774 ( a8_v3[4], a8_v2[4], k7[4] );
xor U3775 ( a7_v3[29], a7_v2[29], k6[29] );
xor U3776 ( a7_v3[28], a7_v2[28], k6[28] );
xor U3777 ( a7_v3[27], a7_v2[27], k6[27] );
xor U3778 ( a7_v3[26], a7_v2[26], k6[26] );
xor U3779 ( a7_v3[25], a7_v2[25], k6[25] );
xor U3780 ( a7_v3[24], a7_v2[24], k6[24] );
xor U3781 ( a7_v3[23], a7_v2[23], k6[23] );
xor U3782 ( a7_v3[22], a7_v2[22], k6[22] );
xor U3783 ( a7_v3[21], a7_v2[21], k6[21] );
xor U3784 ( a7_v3[20], a7_v2[20], k6[20] );
xor U3785 ( a7_v3[19], a7_v2[19], k6[19] );
xor U3786 ( a7_v3[18], a7_v2[18], k6[18] );
xor U3787 ( a7_v3[17], a7_v2[17], k6[17] );
xor U3788 ( a7_v3[16], a7_v2[16], k6[16] );
xor U3789 ( a7_v3[15], a7_v2[15], k6[15] );
xor U3790 ( a7_v3[14], a7_v2[14], k6[14] );
xor U3791 ( a7_v3[13], a7_v2[13], k6[13] );
xor U3792 ( a7_v3[12], a7_v2[12], k6[12] );
xor U3793 ( a7_v3[11], a7_v2[11], k6[11] );
xor U3794 ( a7_v3[10], a7_v2[10], k6[10] );
xor U3795 ( a7_v3[9], a7_v2[9], k6[9] );
xor U3796 ( a7_v3[8], a7_v2[8], k6[8] );
xor U3797 ( a7_v3[7], a7_v2[7], k6[7] );
xor U3798 ( a7_v3[6], a7_v2[6], k6[6] );
xor U3799 ( a7_v3[5], a7_v2[5], k6[5] );
xor U3800 ( a7_v3[4], a7_v2[4], k6[4] );
xor U3801 ( a6_v3[30], a6_v2[30], k5[30] );
xor U3802 ( a6_v3[28], a6_v2[28], k5[28] );
xor U3803 ( a6_v3[27], a6_v2[27], k5[27] );
xor U3804 ( a6_v3[26], a6_v2[26], k5[26] );
xor U3805 ( a6_v3[25], a6_v2[25], k5[25] );
xor U3806 ( a6_v3[24], a6_v2[24], k5[24] );
xor U3807 ( a6_v3[23], a6_v2[23], k5[23] );
xor U3808 ( a6_v3[22], a6_v2[22], k5[22] );
xor U3809 ( a6_v3[21], a6_v2[21], k5[21] );
xor U3810 ( a6_v3[20], a6_v2[20], k5[20] );
xor U3811 ( a6_v3[19], a6_v2[19], k5[19] );
xor U3812 ( a6_v3[18], a6_v2[18], k5[18] );
xor U3813 ( a6_v3[17], a6_v2[17], k5[17] );
xor U3814 ( a6_v3[16], a6_v2[16], k5[16] );
xor U3815 ( a6_v3[15], a6_v2[15], k5[15] );
xor U3816 ( a6_v3[14], a6_v2[14], k5[14] );
xor U3817 ( a6_v3[13], a6_v2[13], k5[13] );
xor U3818 ( a6_v3[12], a6_v2[12], k5[12] );
xor U3819 ( a6_v3[11], a6_v2[11], k5[11] );
xor U3820 ( a6_v3[10], a6_v2[10], k5[10] );
xor U3821 ( a6_v3[9], a6_v2[9], k5[9] );
xor U3822 ( a6_v3[8], a6_v2[8], k5[8] );
xor U3823 ( a6_v3[7], a6_v2[7], k5[7] );
xor U3824 ( a6_v3[6], a6_v2[6], k5[6] );
xor U3825 ( a6_v3[5], a6_v2[5], k5[5] );
xor U3826 ( a6_v3[4], a6_v2[4], k5[4] );
xor U3827 ( a5_v3[30], a5_v2[30], k4[30] );
xor U3828 ( a5_v3[29], a5_v2[29], k4[29] );
xor U3829 ( a5_v3[27], a5_v2[27], k4[27] );
xor U3830 ( a5_v3[26], a5_v2[26], k4[26] );
xor U3831 ( a5_v3[25], a5_v2[25], k4[25] );
xor U3832 ( a5_v3[24], a5_v2[24], k4[24] );
xor U3833 ( a5_v3[23], a5_v2[23], k4[23] );
xor U3834 ( a5_v3[22], a5_v2[22], k4[22] );
xor U3835 ( a5_v3[21], a5_v2[21], k4[21] );
xor U3836 ( a5_v3[20], a5_v2[20], k4[20] );
xor U3837 ( a5_v3[19], a5_v2[19], k4[19] );
xor U3838 ( a5_v3[18], a5_v2[18], k4[18] );
xor U3839 ( a5_v3[17], a5_v2[17], k4[17] );
xor U3840 ( a5_v3[16], a5_v2[16], k4[16] );
xor U3841 ( a5_v3[15], a5_v2[15], k4[15] );
xor U3842 ( a5_v3[14], a5_v2[14], k4[14] );
xor U3843 ( a5_v3[13], a5_v2[13], k4[13] );
xor U3844 ( a5_v3[12], a5_v2[12], k4[12] );
xor U3845 ( a5_v3[11], a5_v2[11], k4[11] );
xor U3846 ( a5_v3[10], a5_v2[10], k4[10] );
xor U3847 ( a5_v3[9], a5_v2[9], k4[9] );
xor U3848 ( a5_v3[8], a5_v2[8], k4[8] );
xor U3849 ( a5_v3[7], a5_v2[7], k4[7] );
xor U3850 ( a5_v3[6], a5_v2[6], k4[6] );
xor U3851 ( a5_v3[5], a5_v2[5], k4[5] );
xor U3852 ( a5_v3[4], a5_v2[4], k4[4] );
xor U3853 ( a4_v3[30], a4_v2[30], k3[30] );
xor U3854 ( a4_v3[29], a4_v2[29], k3[29] );
xor U3855 ( a4_v3[28], a4_v2[28], k3[28] );
xor U3856 ( a4_v3[26], a4_v2[26], k3[26] );
xor U3857 ( a4_v3[25], a4_v2[25], k3[25] );
xor U3858 ( a4_v3[24], a4_v2[24], k3[24] );
xor U3859 ( a4_v3[23], a4_v2[23], k3[23] );
xor U3860 ( a4_v3[22], a4_v2[22], k3[22] );
xor U3861 ( a4_v3[21], a4_v2[21], k3[21] );
xor U3862 ( a4_v3[20], a4_v2[20], k3[20] );
xor U3863 ( a4_v3[19], a4_v2[19], k3[19] );
xor U3864 ( a4_v3[18], a4_v2[18], k3[18] );
xor U3865 ( a4_v3[17], a4_v2[17], k3[17] );
xor U3866 ( a4_v3[16], a4_v2[16], k3[16] );
xor U3867 ( a4_v3[15], a4_v2[15], k3[15] );
xor U3868 ( a4_v3[14], a4_v2[14], k3[14] );
xor U3869 ( a4_v3[13], a4_v2[13], k3[13] );
xor U3870 ( a4_v3[12], a4_v2[12], k3[12] );
xor U3871 ( a4_v3[11], a4_v2[11], k3[11] );
xor U3872 ( a4_v3[10], a4_v2[10], k3[10] );
xor U3873 ( a4_v3[9], a4_v2[9], k3[9] );
xor U3874 ( a4_v3[8], a4_v2[8], k3[8] );
xor U3875 ( a4_v3[7], a4_v2[7], k3[7] );
xor U3876 ( a4_v3[6], a4_v2[6], k3[6] );
xor U3877 ( a4_v3[5], a4_v2[5], k3[5] );
xor U3878 ( a4_v3[4], a4_v2[4], k3[4] );
xor U3879 ( a3_v3[30], a3_v2[30], k2[30] );
xor U3880 ( a3_v3[29], a3_v2[29], k2[29] );
xor U3881 ( a3_v3[28], a3_v2[28], k2[28] );
xor U3882 ( a3_v3[27], a3_v2[27], k2[27] );
xor U3883 ( a3_v3[25], a3_v2[25], k2[25] );
xor U3884 ( a3_v3[24], a3_v2[24], k2[24] );
xor U3885 ( a3_v3[23], a3_v2[23], k2[23] );
xor U3886 ( a3_v3[22], a3_v2[22], k2[22] );
xor U3887 ( a3_v3[21], a3_v2[21], k2[21] );
xor U3888 ( a3_v3[20], a3_v2[20], k2[20] );
xor U3889 ( a3_v3[19], a3_v2[19], k2[19] );
xor U3890 ( a3_v3[18], a3_v2[18], k2[18] );
xor U3891 ( a3_v3[17], a3_v2[17], k2[17] );
xor U3892 ( a3_v3[16], a3_v2[16], k2[16] );
xor U3893 ( a3_v3[15], a3_v2[15], k2[15] );
xor U3894 ( a3_v3[14], a3_v2[14], k2[14] );
xor U3895 ( a3_v3[13], a3_v2[13], k2[13] );
xor U3896 ( a3_v3[12], a3_v2[12], k2[12] );
xor U3897 ( a3_v3[11], a3_v2[11], k2[11] );
xor U3898 ( a3_v3[10], a3_v2[10], k2[10] );
xor U3899 ( a3_v3[9], a3_v2[9], k2[9] );
xor U3900 ( a3_v3[8], a3_v2[8], k2[8] );
xor U3901 ( a3_v3[7], a3_v2[7], k2[7] );
xor U3902 ( a3_v3[6], a3_v2[6], k2[6] );
xor U3903 ( a3_v3[5], a3_v2[5], k2[5] );
xor U3904 ( a3_v3[4], a3_v2[4], k2[4] );
xor U3905 ( a2_v3[30], a2_v2[30], k1[30] );
xor U3906 ( a2_v3[29], a2_v2[29], k1[29] );
xor U3907 ( a2_v3[28], a2_v2[28], k1[28] );
xor U3908 ( a2_v3[27], a2_v2[27], k1[27] );
xor U3909 ( a2_v3[26], a2_v2[26], k1[26] );
xor U3910 ( a2_v3[24], a2_v2[24], k1[24] );
xor U3911 ( a2_v3[23], a2_v2[23], k1[23] );
xor U3912 ( a2_v3[22], a2_v2[22], k1[22] );
xor U3913 ( a2_v3[21], a2_v2[21], k1[21] );
xor U3914 ( a2_v3[20], a2_v2[20], k1[20] );
xor U3915 ( a2_v3[19], a2_v2[19], k1[19] );
xor U3916 ( a2_v3[18], a2_v2[18], k1[18] );
xor U3917 ( a2_v3[17], a2_v2[17], k1[17] );
xor U3918 ( a2_v3[16], a2_v2[16], k1[16] );
xor U3919 ( a2_v3[15], a2_v2[15], k1[15] );
xor U3920 ( a2_v3[14], a2_v2[14], k1[14] );
xor U3921 ( a2_v3[13], a2_v2[13], k1[13] );
xor U3922 ( a2_v3[12], a2_v2[12], k1[12] );
xor U3923 ( a2_v3[11], a2_v2[11], k1[11] );
xor U3924 ( a2_v3[10], a2_v2[10], k1[10] );
xor U3925 ( a2_v3[9], a2_v2[9], k1[9] );
xor U3926 ( a2_v3[8], a2_v2[8], k1[8] );
xor U3927 ( a2_v3[7], a2_v2[7], k1[7] );
xor U3928 ( a2_v3[6], a2_v2[6], k1[6] );
xor U3929 ( a2_v3[5], a2_v2[5], k1[5] );
xor U3930 ( a2_v3[4], a2_v2[4], k1[4] );
xor U3931 ( a2_v3[31], a2_v2[31], k1[31] );
xor U3932 ( a3_v3[31], a3_v2[31], k2[31] );
xor U3933 ( a4_v3[31], a4_v2[31], k3[31] );
xor U3934 ( a5_v3[31], a5_v2[31], k4[31] );
xor U3935 ( a6_v3[31], a6_v2[31], k5[31] );
xor U3936 ( a7_v3[31], a7_v2[31], k6[31] );
xor U3937 ( a9_v3[31], a9_v2[31], k8[31] );
xor U3938 ( a1_v1[30], n1017, n986 );
xor U3939 ( a1_v1[29], n1016, n985 );
xor U3940 ( a1_v1[28], n1015, n984 );
xor U3941 ( a1_v1[27], n1014, n983 );
xor U3942 ( a1_v1[26], n1013, n982 );
xor U3943 ( a1_v1[25], n1012, n981 );
xor U3944 ( a1_v1[23], n1011, n979 );
xor U3945 ( a1_v1[22], n1010, n978 );
xor U3946 ( a1_v1[21], n1009, n977 );
xor U3947 ( a1_v1[20], n1008, n976 );
xor U3948 ( a1_v1[19], n1007, n975 );
xor U3949 ( a1_v1[18], n1006, n974 );
xor U3950 ( a1_v1[17], n1005, n973 );
xor U3951 ( a1_v1[16], n1004, n972 );
xor U3952 ( a1_v1[15], n1003, n971 );
xor U3953 ( a1_v1[14], n1002, n970 );
xor U3954 ( a1_v1[13], n1001, n969 );
xor U3955 ( a1_v1[12], n1000, n968 );
xor U3956 ( a1_v1[11], n999, n967 );
xor U3957 ( a1_v1[10], n998, n966 );
xor U3958 ( a1_v1[9], n997, n965 );
xor U3959 ( a1_v1[8], n996, n964 );
xor U3960 ( a1_v1[7], n995, n963 );
xor U3961 ( a1_v1[6], n994, n962 );
xor U3962 ( a1_v1[5], n993, n961 );
xor U3963 ( a1_v1[4], n992, n960 );
xor U3964 ( a1_v1[3], n991, n959 );
xor U3965 ( a1_v1[2], n990, n958 );
xor U3966 ( a1_v1[1], n989, n957 );
xor U3967 ( a1_v1[0], n988, n956 );
xor U3968 ( a1_v1[31], n1018, n987 );
xnor U3969 ( a1_v2[31], n955, a1_v1[31] );
xnor U3970 ( a1_v2[30], n954, a1_v1[30] );
xnor U3971 ( a1_v2[29], n953, a1_v1[29] );
xnor U3972 ( a1_v2[28], n952, a1_v1[28] );
xnor U3973 ( a1_v2[27], n951, a1_v1[27] );
xnor U3974 ( a1_v2[26], n950, a1_v1[26] );
xnor U3975 ( a1_v2[25], n949, a1_v1[25] );
xnor U3976 ( a1_v2[23], n947, a1_v1[23] );
xnor U3977 ( a1_v2[22], n946, a1_v1[22] );
xnor U3978 ( a1_v2[21], n945, a1_v1[21] );
xnor U3979 ( a1_v2[20], n944, a1_v1[20] );
xnor U3980 ( a1_v2[19], n943, a1_v1[19] );
xnor U3981 ( a1_v2[18], n942, a1_v1[18] );
xnor U3982 ( a1_v2[17], n941, a1_v1[17] );
xnor U3983 ( a1_v2[16], n940, a1_v1[16] );
xnor U3984 ( a1_v2[15], n939, a1_v1[15] );
xnor U3985 ( a1_v2[14], n938, a1_v1[14] );
xnor U3986 ( a1_v2[13], n937, a1_v1[13] );
xnor U3987 ( a1_v2[12], n936, a1_v1[12] );
xnor U3988 ( a1_v2[11], n935, a1_v1[11] );
xnor U3989 ( a1_v2[10], n934, a1_v1[10] );
xnor U3990 ( a1_v2[9], n933, a1_v1[9] );
xnor U3991 ( a1_v2[8], n932, a1_v1[8] );
xnor U3992 ( a1_v2[7], n931, a1_v1[7] );
xnor U3993 ( a1_v2[6], n930, a1_v1[6] );
xnor U3994 ( a1_v2[5], n929, a1_v1[5] );
xnor U3995 ( a1_v2[4], n928, a1_v1[4] );
xnor U3996 ( a1_v2[3], n927, a1_v1[3] );
xnor U3997 ( a1_v2[2], n926, a1_v1[2] );
xnor U3998 ( a1_v2[1], n925, a1_v1[1] );
xnor U3999 ( a1_v2[0], n924, a1_v1[0] );
xor U4000 ( a1_v3[30], a1_v2[30], k0[30] );
xor U4001 ( a1_v3[29], a1_v2[29], k0[29] );
xor U4002 ( a1_v3[28], a1_v2[28], k0[28] );
xor U4003 ( a1_v3[27], a1_v2[27], k0[27] );
xor U4004 ( a1_v3[26], a1_v2[26], k0[26] );
xor U4005 ( a1_v3[25], a1_v2[25], k0[25] );
xor U4006 ( a1_v3[23], a1_v2[23], k0[23] );
xor U4007 ( a1_v3[22], a1_v2[22], k0[22] );
xor U4008 ( a1_v3[21], a1_v2[21], k0[21] );
xor U4009 ( a1_v3[20], a1_v2[20], k0[20] );
xor U4010 ( a1_v3[19], a1_v2[19], k0[19] );
xor U4011 ( a1_v3[18], a1_v2[18], k0[18] );
xor U4012 ( a1_v3[17], a1_v2[17], k0[17] );
xor U4013 ( a1_v3[16], a1_v2[16], k0[16] );
xor U4014 ( a1_v3[15], a1_v2[15], k0[15] );
xor U4015 ( a1_v3[14], a1_v2[14], k0[14] );
xor U4016 ( a1_v3[13], a1_v2[13], k0[13] );
xor U4017 ( a1_v3[12], a1_v2[12], k0[12] );
xor U4018 ( a1_v3[11], a1_v2[11], k0[11] );
xor U4019 ( a1_v3[10], a1_v2[10], k0[10] );
xor U4020 ( a1_v3[9], a1_v2[9], k0[9] );
xor U4021 ( a1_v3[8], a1_v2[8], k0[8] );
xor U4022 ( a1_v3[7], a1_v2[7], k0[7] );
xor U4023 ( a1_v3[6], a1_v2[6], k0[6] );
xor U4024 ( a1_v3[5], a1_v2[5], k0[5] );
xor U4025 ( a1_v3[4], a1_v2[4], k0[4] );
xor U4026 ( a1_v3[3], a1_v2[3], k0[3] );
xor U4027 ( a1_v3[2], a1_v2[2], k0[2] );
xor U4028 ( a1_v3[1], a1_v2[1], k0[1] );
xor U4029 ( a1_v3[0], a1_v2[0], k0[0] );
xor U4030 ( a1_v3[31], a1_v2[31], k0[31] );
xnor U4031 ( a1_v1[24], n1284, n980 );
xnor U4032 ( a1_v2[24], n948, a1_v1[24] );
xor U4033 ( a1_v3[24], k0[24], a1_v2[24] );
not U4034 ( n1283, reset );
nand U4035 ( n1302, start, n1019 );
buf U4036 ( n1585, n1557 );
buf U4037 ( n1584, n1557 );
buf U4038 ( n1583, n1584 );
buf U4039 ( n1579, n1585 );
buf U4040 ( n1580, n1585 );
buf U4041 ( n1581, n1584 );
buf U4042 ( n1582, n1584 );
endmodule

