
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule


module s38584_ori ( clk, reset, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6753, g7243, g7245, g7257, g7260, g7540, g7916,
g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342,
g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784,
g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917,
g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615,
g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500,
g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238,
g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039,
g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895,
g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694,
g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656,
g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874,
g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519,
g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678,
g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764,
g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095,
g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245,
g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683,
g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584,
g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876,
g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212,
g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221,
g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946,
g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233,
g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425,
g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917,
g34919, g34921, g34923, g34925, g34927, g34956, g34972 );
input clk, reset, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750,
g6751, g6753;
output g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215,
g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398,
g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019,
g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741,
g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418,
g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368,
g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068,
g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259,
g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589,
g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041,
g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215,
g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329,
g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860,
g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945,
g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221,
g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239,
g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788,
g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925,
g34927, g34956, g34972;
wire ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, ex_wire30, ex_wire31, ex_wire32, ex_wire33, ex_wire34, ex_wire35, ex_wire36, ex_wire37, ex_wire38, ex_wire39, ex_wire40, ex_wire41, ex_wire42, ex_wire43, ex_wire44, ex_wire45, ex_wire46, ex_wire47, ex_wire48, ex_wire49, ex_wire50, ex_wire51, ex_wire52, ex_wire53, ex_wire54, ex_wire55, ex_wire56, ex_wire57, ex_wire58, ex_wire59, ex_wire60, ex_wire61, ex_wire62, ex_wire63, ex_wire64, ex_wire65, ex_wire66, ex_wire67, ex_wire68, ex_wire69, ex_wire70, ex_wire71, ex_wire72, ex_wire73, ex_wire74, ex_wire75, ex_wire76, ex_wire77, ex_wire78, ex_wire79, ex_wire80, ex_wire81, ex_wire82, ex_wire83, ex_wire84, ex_wire85, ex_wire86, ex_wire87, ex_wire88, ex_wire89, ex_wire90, ex_wire91, ex_wire92, ex_wire93, ex_wire94, ex_wire95, ex_wire96, ex_wire97, ex_wire98, ex_wire99, ex_wire100, ex_wire101, ex_wire102, ex_wire103, ex_wire104, ex_wire105, ex_wire106, ex_wire107, ex_wire108, ex_wire109, ex_wire110, ex_wire111, ex_wire112, ex_wire113, ex_wire114, ex_wire115, ex_wire116, ex_wire117, ex_wire118, ex_wire119, ex_wire120, ex_wire121, ex_wire122, ex_wire123, ex_wire124, ex_wire125, ex_wire126, ex_wire127, ex_wire128, ex_wire129, ex_wire130, ex_wire131, ex_wire132, ex_wire133, ex_wire134, ex_wire135, ex_wire136, ex_wire137, ex_wire138, ex_wire139, ex_wire140, ex_wire141, ex_wire142, ex_wire143, ex_wire144, ex_wire145, ex_wire146, ex_wire147, ex_wire148, ex_wire149, ex_wire150, ex_wire151, ex_wire152, ex_wire153, ex_wire154, ex_wire155, ex_wire156, ex_wire157, ex_wire158, ex_wire159, ex_wire160, ex_wire161, ex_wire162, ex_wire163, ex_wire164, ex_wire165, ex_wire166, ex_wire167, ex_wire168, ex_wire169, ex_wire170, ex_wire171, ex_wire172, ex_wire173, ex_wire174, ex_wire175, ex_wire176, ex_wire177, ex_wire178, ex_wire179, ex_wire180, ex_wire181, ex_wire182, ex_wire183, ex_wire184, ex_wire185, ex_wire186, ex_wire187, ex_wire188, ex_wire189, ex_wire190, ex_wire191, ex_wire192, ex_wire193, ex_wire194, ex_wire195, ex_wire196, ex_wire197, ex_wire198, ex_wire199, ex_wire200, ex_wire201, ex_wire202, ex_wire203, ex_wire204, ex_wire205, ex_wire206, ex_wire207, ex_wire208, ex_wire209, ex_wire210, ex_wire211, ex_wire212, ex_wire213, ex_wire214, ex_wire215, ex_wire216, ex_wire217, ex_wire218, ex_wire219, ex_wire220, ex_wire221, ex_wire222, ex_wire223, ex_wire224, ex_wire225, ex_wire226, ex_wire227, ex_wire228, ex_wire229, ex_wire230, ex_wire231, ex_wire232, ex_wire233, ex_wire234, ex_wire235, ex_wire236, ex_wire237, ex_wire238, ex_wire239, ex_wire240, ex_wire241, ex_wire242, ex_wire243, ex_wire244, ex_wire245, ex_wire246, ex_wire247, ex_wire248, ex_wire249, ex_wire250, ex_wire251, ex_wire252, ex_wire253, ex_wire254, ex_wire255, ex_wire256, ex_wire257, ex_wire258, ex_wire259, ex_wire260, ex_wire261, ex_wire262, ex_wire263, ex_wire264, ex_wire265, ex_wire266, ex_wire267, ex_wire268, ex_wire269, ex_wire270, ex_wire271, ex_wire272, ex_wire273, ex_wire274, ex_wire275, ex_wire276, ex_wire277, ex_wire278, ex_wire279, ex_wire280, ex_wire281, ex_wire282, ex_wire283, ex_wire284, ex_wire285, ex_wire286, ex_wire287, ex_wire288, ex_wire289, ex_wire290, ex_wire291, ex_wire292, ex_wire293, ex_wire294, ex_wire295, ex_wire296, ex_wire297, ex_wire298, ex_wire299, ex_wire300, ex_wire301, ex_wire302, ex_wire303, ex_wire304, ex_wire305, ex_wire306, ex_wire307, ex_wire308, ex_wire309, ex_wire310, ex_wire311, ex_wire312, ex_wire313, ex_wire314, ex_wire315, ex_wire316, ex_wire317, ex_wire318, ex_wire319, ex_wire320, ex_wire321, ex_wire322, ex_wire323, ex_wire324, ex_wire325, ex_wire326, ex_wire327, ex_wire328, ex_wire329, ex_wire330, ex_wire331, ex_wire332, ex_wire333, ex_wire334, ex_wire335, ex_wire336, ex_wire337, ex_wire338, ex_wire339, ex_wire340, ex_wire341, ex_wire342, ex_wire343, ex_wire344, ex_wire345, ex_wire346, ex_wire347, ex_wire348, ex_wire349, ex_wire350, ex_wire351, ex_wire352, ex_wire353, ex_wire354, ex_wire355, ex_wire356, ex_wire357, ex_wire358, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6753,
g496, g341, g21270, g4467, g4519, g4564, g4570, g4531, g4578, g20557,
g21245, g20763, g45, g46, g47, g48, g55, g53, g23683, g54, g56, g57,
g20049, g20899, g65, g64, g90, g91, g72, g73, g113, g124, g114,
g25219, g92, g99, g115, g125, g84, g100, g126, g127, g20652, g116,
g20654, g134, g120, g135, g21292, g20901, g44, g21176, g26801,
new_g10520_, g25167, g25259, g27831, new_g18597_, new_g24265_,
new_g24266_, new_g24298_, g31521, g31656, g31665, new_g25688_,
new_g25689_, new_g25690_, g33894, g29218, new_g34649_, new_g34657_,
new_g34663_, new_g34781_, new_g34783_, new_g34843_, new_g34809_,
new_g34970_, new_g34971_, new_g34974_, new_g34975_, new_g34976_,
new_g34977_, new_g34978_, new_g34979_, g4480, g4495, g4567, g4498,
g4501, g4540, g4543, g4546, g4455, n4694, n4595, n4575, n4580, n4585,
n4629, n4638, n4643, n4652, n4600, n4657, n5240, n5245, n5205, n5235,
n5230, n5225, n5220, n5215, n5210, n5195, n5295, n5413, n5320, n5040,
n5045, n5035, n5862, n6053, n6103, n6108, n6113, n6013, n6023, n5912,
n5963, n5977, n5990, n5949, n5972, n5929, n5958, n5934, n5536, n5727,
n5777, n5782, n5787, n5687, n5697, n5586, n5637, n5651, n5664, n5623,
n5646, n5603, n5632, n5608, n7293, n3353, n3394, n3399, n3404, n3712,
n3753, n3758, n3763, n4071, n4112, n4117, n4122, n4731, n4590, n1110,
n1119, n1164, n1169, n1558, n1599, n1604, n1609, n1917, n1958, n1963,
n1968, n2276, n2317, n2322, n2327, n2635, n2676, n2681, n2686, n2994,
n3035, n3040, n3045, n5527, n5513, n5522, n5438, n5001, n5015, n5010,
n5020, n5025, n5260, n5255, n5250, n5270, n5265, n5160, n5165, n5170,
n5175, n4823, n5135, n5140, n5310, n5060, n5065, n5050, n5867, n6058,
n6063, n6093, n6043, n6153, n6018, n5944, n5939, n5541, n5732, n5737,
n5767, n5717, n5827, n5692, n5618, n5613, n7298, n3419, n3433, n3428,
n3677, n3697, n3702, n3662, n3778, n3792, n3787, n4036, n4056, n4061,
n4021, n4137, n4151, n4146, n4395, n4415, n4420, n4380, n4450, n4455,
n4460, n4445, n1476, n1707, n1712, n1717, n1722, n1727, n1624, n1638,
n1633, n1647, n1702, n1882, n1902, n1907, n1867, n1983, n1997, n1992,
n2241, n2261, n2266, n2226, n2342, n2356, n2351, n2600, n2620, n2625,
n2585, n2701, n2715, n2710, n2959, n2979, n2984, n2944, n3060, n3074,
n3069, n3318, n3338, n3343, n3303, n4736, n4741, n4761, n4756, n4771,
n4766, n4746, n4751, n4805, n4800, n4776, n4785, n4790, n4795, n5180,
n4828, n5125, n5315, n5055, n5070, n4903, n4936, n4941, n4946, n4951,
n4956, n4961, n4966, n4971, n4981, n4986, n5872, n6098, n6048, n6133,
n6143, n6123, n6028, n5546, n5772, n5722, n5807, n5817, n5797, n5702,
n7303, n7343, n7348, n7353, n7358, n7393, n7398, n7403, n7408, n4465,
n4500, n4530, n1214, n1061, n1052, n1080, n1070, n1075, n1090, n1047,
n1042, n1023, n1014, n1032, n1037, n1105, n1100, n852, n916, n921,
n926, n897, n1004, n984, n994, n989, n837, n822, n887, n5443, n5185,
n4833, n5085, n5090, n5130, n5100, n5105, n5110, n5115, n5095, n5120,
n5075, n5877, n6068, n5551, n5742, n7308, n3652, n4011, n4370, n4470,
n4505, n4510, n4515, n4520, n892, n1518, n1528, n1538, n1548, n1351,
n1361, n1371, n1381, n1697, n1692, n1857, n2216, n2575, n2934, n3293,
n5200, n5190, n4838, n5145, n5150, n5155, n5333, n5080, n5882, n6118,
n6138, n6148, n6128, n5556, n5792, n5812, n5822, n5802, n6273, n6278,
n6403, n6408, n6533, n6538, n6663, n6668, n6818, n6823, n6948, n6953,
n7078, n7083, n7208, n7213, n7313, n3667, n3672, n3682, n3687, n3692,
n3657, n4026, n4031, n4041, n4046, n4051, n4016, n4385, n4390, n4400,
n4405, n4410, n4375, n4475, n1471, n1304, n1872, n1877, n1887, n1892,
n1897, n1862, n2231, n2236, n2246, n2251, n2256, n2221, n2590, n2595,
n2605, n2610, n2615, n2580, n2949, n2954, n2964, n2969, n2974, n2939,
n3308, n3313, n3323, n3328, n3333, n3298, n5473, n4843, n5338, n5887,
n6073, n6003, n6008, n6033, n6038, n5561, n5747, n5677, n5682, n5707,
n5712, n6248, n6283, n6288, n6308, n6313, n6378, n6413, n6418, n6438,
n6443, n6508, n6543, n6548, n6568, n6573, n6638, n6673, n6678, n6698,
n6703, n6793, n6828, n6833, n6853, n6858, n6923, n6958, n6963, n6983,
n6988, n7053, n7088, n7093, n7113, n7118, n7183, n7218, n7223, n7243,
n7248, n7318, n7388, n7438, n7383, n7433, n3527, n3552, n3577, n3602,
n3627, n3557, n3582, n3607, n3632, n3562, n3587, n3612, n3637, n3567,
n3592, n3617, n3642, n3572, n3597, n3622, n3647, n3886, n3911, n3936,
n3961, n3986, n3916, n3941, n3966, n3991, n3921, n3946, n3971, n3996,
n3926, n3951, n3976, n4001, n3931, n3956, n3981, n4006, n4245, n4270,
n4295, n4320, n4345, n4275, n4300, n4325, n4350, n4280, n4305, n4330,
n4355, n4285, n4310, n4335, n4360, n4290, n4315, n4340, n4365, n4480,
n4525, n812, n1732, n1757, n1782, n1807, n1832, n1762, n1787, n1812,
n1837, n1767, n1792, n1817, n1842, n1772, n1797, n1822, n1847, n1777,
n1802, n1827, n1852, n2091, n2116, n2141, n2166, n2191, n2121, n2146,
n2171, n2196, n2126, n2151, n2176, n2201, n2131, n2156, n2181, n2206,
n2136, n2161, n2186, n2211, n2450, n2475, n2500, n2525, n2550, n2480,
n2505, n2530, n2555, n2485, n2510, n2535, n2560, n2490, n2515, n2540,
n2565, n2495, n2520, n2545, n2570, n2809, n2834, n2859, n2884, n2909,
n2839, n2864, n2889, n2914, n2844, n2869, n2894, n2919, n2849, n2874,
n2899, n2924, n2854, n2879, n2904, n2929, n3168, n3193, n3218, n3243,
n3268, n3198, n3223, n3248, n3273, n3203, n3228, n3253, n3278, n3208,
n3233, n3258, n3283, n3213, n3238, n3263, n3288, n5478, n5448, n4848,
n5343, n5892, n6078, n5566, n5752, n7323, n4485, n1085, n857, n940,
n1652, n1667, n1672, n1677, n1657, n1682, n1662, n5483, n5453, n4853,
n5348, n5030, n5897, n5907, n6083, n5571, n5581, n5757, n6253, n6258,
n6268, n6263, n6383, n6388, n6398, n6393, n6513, n6518, n6528, n6523,
n6643, n6648, n6658, n6653, n6798, n6803, n6813, n6808, n6928, n6933,
n6943, n6938, n7058, n7063, n7073, n7068, n7188, n7193, n7203, n7198,
n7328, n3532, n3537, n3542, n3547, n3891, n3896, n3901, n3906, n4250,
n4255, n4260, n4265, n4490, n862, n867, n872, n877, n882, n960, n945,
n950, n965, n955, n1687, n1737, n1742, n1747, n1752, n2096, n2101,
n2106, n2111, n2455, n2460, n2465, n2470, n2814, n2819, n2824, n2829,
n3173, n3178, n3183, n3188, n5488, n5458, n5503, n5508, n4858, n5353,
n5902, n6088, n5576, n5762, n6188, n6198, n6203, n6213, n6293, n6298,
n6303, n6193, n6318, n6328, n6333, n6343, n6423, n6428, n6433, n6323,
n6448, n6458, n6463, n6473, n6553, n6558, n6563, n6453, n6578, n6588,
n6593, n6603, n6683, n6688, n6693, n6583, n6733, n6743, n6748, n6758,
n6838, n6843, n6848, n6738, n6863, n6873, n6878, n6888, n6968, n6973,
n6978, n6868, n6993, n7003, n7008, n7018, n7098, n7103, n7108, n6998,
n7123, n7133, n7138, n7148, n7228, n7233, n7238, n7128, n7333, n3409,
n3414, n3768, n3773, n4127, n4132, n4495, n902, n970, n1614, n1619,
n1973, n1978, n2332, n2337, n2691, n2696, n3050, n3055, n5493, n5463,
n5300, n5305, n4863, n5358, n6223, n6228, n6243, n6238, n6233, n6208,
n6218, n6353, n6358, n6373, n6368, n6363, n6338, n6348, n6483, n6488,
n6503, n6498, n6493, n6468, n6478, n6613, n6618, n6633, n6628, n6623,
n6598, n6608, n6768, n6773, n6788, n6783, n6778, n6753, n6763, n6898,
n6903, n6918, n6913, n6908, n6883, n6893, n7028, n7033, n7048, n7043,
n7038, n7013, n7023, n7158, n7163, n7178, n7173, n7168, n7143, n7153,
n7338, n999, n931, n1396, n1401, n1406, n1508, n1498, n1503, n1513,
n1493, n1229, n1234, n1239, n1341, n1331, n1336, n1346, n1326, n5498,
n5468, n4868, n5363, n817, n832, n842, n827, n1154, n1159, n1144,
n1391, n1523, n1533, n1543, n1553, n1224, n1356, n1366, n1376, n1386,
n4873, n5368, n4976, n7378, n7368, n7373, n7363, n7428, n7418, n7423,
n7413, n1174, n1179, n1189, n1194, n1199, n1204, n1184, n1209, n1134,
n1139, n1149, n1129, n1416, n1411, n1421, n1426, n1249, n1244, n1254,
n1259, n5428, n4878, n5373, n6158, n5832, n6708, n6713, n6718, n7253,
n7258, n7263, n7473, n7478, n7483, n7488, n7493, n7498, n7463, n7458,
n7548, n7553, n7558, n7563, n7568, n7573, n7578, n7453, n3707, n4066,
n4425, n4565, n4570, n4614, n4619, n4624, n1431, n1436, n1441, n1446,
n1451, n1264, n1269, n1274, n1279, n1284, n1912, n2271, n2630, n2989,
n3348, n5403, n5423, n5433, n5408, n5418, n4883, n5378, n6163, n6168,
n6173, n5837, n5842, n5847, n7448, n4555, n4560, n4609, n4888, n5383,
n7503, n7508, n7513, n7518, n7523, n7528, n7533, n7468, n7538, n7583,
n7588, n7593, n7613, n7443, n7598, n7603, n7608, n4893, n5388, n4898,
n5393, n1219, n5398, n7543, n911, n979, n40, n51, n137, n139, n145,
n177, g33959, n210, g31860, g30329, g30331, g30330, g30327, g34839,
n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
n20238;
assign g21698 = g36;
assign g18098 = g6744;
assign g18099 = g6745;
assign g18101 = g6746;
assign g18097 = g6747;
assign g18094 = g6748;
assign g18095 = g6749;
assign g18096 = g6750;
assign g18100 = g6751;
assign g18092 = g6753;
assign g29217 = g21270;
assign g29213 = g20557;
assign g29220 = g21245;
assign g29211 = g20763;
assign g30332 = g23683;
assign g29210 = g20049;
assign g29212 = g20899;
assign g31861 = g25219;
assign g29214 = g20652;
assign g29219 = g20654;
assign g29221 = g21292;
assign g29215 = g20901;
assign g29216 = g21176;
assign g32975 = g26801;
assign g31863 = g25167;
assign g31862 = g25259;
assign g33533 = g27831;
assign g34435 = g31521;
assign g34436 = g31656;
assign g34437 = g31665;
assign g34788 = g33894;
assign g18881 = g29218;
assign g28753 = g33959;
assign g25114 = g31860;
assign g23612 = g30329;
assign g23759 = g30331;
assign g23652 = g30330;
assign g23002 = g30327;
assign g34240 = 1'b1;
assign g34239 = 1'b1;
assign g34238 = 1'b1;
assign g34237 = 1'b1;
assign g34236 = 1'b1;
assign g34235 = 1'b1;
assign g34234 = 1'b1;
assign g34233 = 1'b1;
assign g34956 = g34839;
assign g33945 = 1'b1;
assign g32429 = 1'b1;
assign g33947 = 1'b1;
assign g33950 = 1'b1;
assign g34232 = 1'b1;
assign g33948 = 1'b1;
assign g33946 = 1'b1;
assign g33949 = 1'b1;
assign g32454 = 1'b1;
assign g24151 = 1'b1;
assign g25590 = 1'b1;
assign g25589 = 1'b1;
assign g25588 = 1'b1;
assign g25587 = 1'b1;
assign g25586 = 1'b1;
assign g25585 = 1'b1;
assign g25584 = 1'b1;
assign g25583 = 1'b1;
assign g25582 = 1'b1;
assign g34597 = 1'b0;

dff g72_reg ( clk, reset, g72, g72 );
not U_inv0 ( n19562, g72 );
dff g73_reg ( clk, reset, g73, g73 );
not U_inv1 ( n19563, g73 );
dff g84_reg ( clk, reset, g84, g84 );
not U_inv2 ( n19564, g84 );
dff g90_reg ( clk, reset, g90, g90 );
not U_inv3 ( n19502, g90 );
dff g91_reg ( clk, reset, g91, g91 );
dff g92_reg ( clk, reset, g92, g92 );
not U_inv4 ( n19330, g92 );
dff g99_reg ( clk, reset, g99, g99 );
dff g100_reg ( clk, reset, g100, g100 );
dff g113_reg ( clk, reset, g113, g113 );
not U_inv5 ( n19566, g113 );
dff g114_reg ( clk, reset, g114, g114 );
dff g115_reg ( clk, reset, g115, g115 );
not U_inv6 ( n19342, g115 );
dff g116_reg ( clk, reset, g116, g116 );
dff g120_reg ( clk, reset, g120, g120 );
dff g124_reg ( clk, reset, g124, g124 );
dff g125_reg ( clk, reset, g125, g125 );
not U_inv7 ( n19109, g125 );
dff g126_reg ( clk, reset, g126, g126 );
not U_inv8 ( n19343, g126 );
dff g127_reg ( clk, reset, g127, g127 );
dff g134_reg ( clk, reset, g134, g134 );
not U_inv9 ( n19567, g134 );
dff g135_reg ( clk, reset, g135, g135 );
not U_inv10 ( n19503, g135 );
dff g44_reg ( clk, reset, g44, g44 );
not U_inv11 ( n19568, g44 );
dff g53_reg ( clk, reset, g53, g53 );
not U_inv12 ( n19492, g53 );
dff g54_reg ( clk, reset, g54, g54 );
dff g56_reg ( clk, reset, g56, g56 );
not U_inv13 ( n19569, g56 );
dff g57_reg ( clk, reset, g57, g57 );
dff g64_reg ( clk, reset, g64, g64 );
dff g4308_reg ( clk, reset, ex_wire0, g9251 );
not U_inv14 ( n19506, ex_wire0 );
dff g4304_reg ( clk, reset, g9251, n1110 );
not U_inv15 ( n19505, g9251 );
dff g2932_reg ( clk, reset, ex_wire1, n1119 );
not U_inv16 ( n19581, ex_wire1 );
dff g4999_reg ( clk, reset, g8178, n1476 );
not U_inv17 ( n19451, g8178 );
dff g5002_reg ( clk, reset, g8283, g8178 );
not U_inv18 ( n19103, g8283 );
dff g5005_reg ( clk, reset, g8403, g8283 );
not U_inv19 ( n19104, g8403 );
dff g5008_reg ( clk, reset, n10893, g8403 );
dff g4809_reg ( clk, reset, g8132, n1476 );
not U_inv20 ( n19440, g8132 );
dff g4812_reg ( clk, reset, g8235, g8132 );
not U_inv21 ( n19105, g8235 );
dff g4815_reg ( clk, reset, g8353, g8235 );
not U_inv22 ( n19106, g8353 );
dff g4818_reg ( clk, reset, n10891, g8353 );
dff g5308_reg ( clk, reset, g13039, g17577 );
not U_inv23 ( n19435, g13039 );
dff g5313_reg ( clk, reset, g12238, n1558 );
not U_inv24 ( n19433, g12238 );
dff g5290_reg ( clk, reset, g14662, g12238 );
not U_inv25 ( n19627, g14662 );
dff g5320_reg ( clk, reset, g17674, g14662 );
not U_inv26 ( n19432, g17674 );
dff g5276_reg ( clk, reset, g17519, g17674 );
not U_inv27 ( n19628, g17519 );
dff g5283_reg ( clk, reset, g17577, g17519 );
not U_inv28 ( n19434, g17577 );
dff g5327_reg ( clk, reset, g17787, g13039 );
not U_inv29 ( n19422, g17787 );
dff g5331_reg ( clk, reset, g14597, g17787 );
not U_inv30 ( n19423, g14597 );
dff g5335_reg ( clk, reset, g17639, g14597 );
not U_inv31 ( n19421, g17639 );
dff g5339_reg ( clk, reset, ex_wire2, g17639 );
not U_inv32 ( n19431, ex_wire2 );
dff g5343_reg ( clk, reset, g25219, n1599 );
not U_inv33 ( n19629, g25219 );
dff g5352_reg ( clk, reset, n10691, n1609 );
not U_inv34 ( n19631, n10691 );
dff g5348_reg ( clk, reset, ex_wire3, n1604 );
not U_inv35 ( n19630, ex_wire3 );
dff g5654_reg ( clk, reset, g13049, g17604 );
not U_inv36 ( n19417, g13049 );
dff g5659_reg ( clk, reset, g12300, n1917 );
not U_inv37 ( n19415, g12300 );
dff g5637_reg ( clk, reset, g14694, g12300 );
not U_inv38 ( n19677, g14694 );
dff g5666_reg ( clk, reset, g17711, g14694 );
not U_inv39 ( n19678, g17711 );
dff g5623_reg ( clk, reset, g17580, g17711 );
not U_inv40 ( n19679, g17580 );
dff g5630_reg ( clk, reset, g17604, g17580 );
not U_inv41 ( n19416, g17604 );
dff g5673_reg ( clk, reset, g17813, g13049 );
not U_inv42 ( n19411, g17813 );
dff g5677_reg ( clk, reset, g14635, g17813 );
not U_inv43 ( n19413, g14635 );
dff g5681_reg ( clk, reset, g17678, g14635 );
not U_inv44 ( n19412, g17678 );
dff g5685_reg ( clk, reset, ex_wire4, g17678 );
not U_inv45 ( n19414, ex_wire4 );
dff g5689_reg ( clk, reset, n10330, n1958 );
not U_inv46 ( n19680, n10330 );
dff g5698_reg ( clk, reset, n10739, n1968 );
not U_inv47 ( n19682, n10739 );
dff g5694_reg ( clk, reset, ex_wire5, n1963 );
not U_inv48 ( n19681, ex_wire5 );
dff g6000_reg ( clk, reset, g13068, g17646 );
not U_inv49 ( n19407, g13068 );
dff g6005_reg ( clk, reset, g12350, n2276 );
not U_inv50 ( n19405, g12350 );
dff g5983_reg ( clk, reset, g14738, g12350 );
not U_inv51 ( n19713, g14738 );
dff g6012_reg ( clk, reset, g17739, g14738 );
not U_inv52 ( n19714, g17739 );
dff g5969_reg ( clk, reset, g17607, g17739 );
not U_inv53 ( n19715, g17607 );
dff g5976_reg ( clk, reset, g17646, g17607 );
not U_inv54 ( n19406, g17646 );
dff g6019_reg ( clk, reset, g17819, g13068 );
not U_inv55 ( n19401, g17819 );
dff g6023_reg ( clk, reset, g14673, g17819 );
not U_inv56 ( n19403, g14673 );
dff g6027_reg ( clk, reset, g17715, g14673 );
not U_inv57 ( n19402, g17715 );
dff g6031_reg ( clk, reset, ex_wire6, g17715 );
not U_inv58 ( n19404, ex_wire6 );
dff g6035_reg ( clk, reset, n10329, n2317 );
not U_inv59 ( n19716, n10329 );
dff g6044_reg ( clk, reset, n10690, n2327 );
not U_inv60 ( n19718, n10690 );
dff g6040_reg ( clk, reset, ex_wire7, n2322 );
not U_inv61 ( n19717, ex_wire7 );
dff g6346_reg ( clk, reset, g13085, g17685 );
not U_inv62 ( n19397, g13085 );
dff g6351_reg ( clk, reset, g12422, n2635 );
not U_inv63 ( n19395, g12422 );
dff g6329_reg ( clk, reset, g14779, g12422 );
not U_inv64 ( n19750, g14779 );
dff g6358_reg ( clk, reset, g17760, g14779 );
not U_inv65 ( n19751, g17760 );
dff g6315_reg ( clk, reset, g17649, g17760 );
not U_inv66 ( n19752, g17649 );
dff g6322_reg ( clk, reset, g17685, g17649 );
not U_inv67 ( n19396, g17685 );
dff g6365_reg ( clk, reset, g17845, g13085 );
not U_inv68 ( n19391, g17845 );
dff g6369_reg ( clk, reset, g14705, g17845 );
not U_inv69 ( n19393, g14705 );
dff g6373_reg ( clk, reset, g17743, g14705 );
not U_inv70 ( n19392, g17743 );
dff g6377_reg ( clk, reset, ex_wire8, g17743 );
not U_inv71 ( n19394, ex_wire8 );
dff g6381_reg ( clk, reset, n10328, n2676 );
not U_inv72 ( n19753, n10328 );
dff g6390_reg ( clk, reset, n10689, n2686 );
not U_inv73 ( n19755, n10689 );
dff g6386_reg ( clk, reset, ex_wire9, n2681 );
not U_inv74 ( n19754, ex_wire9 );
dff g6692_reg ( clk, reset, g13099, g17722 );
not U_inv75 ( n19387, g13099 );
dff g6697_reg ( clk, reset, g12470, n2994 );
not U_inv76 ( n19385, g12470 );
dff g6675_reg ( clk, reset, g14828, g12470 );
not U_inv77 ( n19786, g14828 );
dff g6704_reg ( clk, reset, g17778, g14828 );
not U_inv78 ( n19787, g17778 );
dff g6661_reg ( clk, reset, g17688, g17778 );
not U_inv79 ( n19788, g17688 );
dff g6668_reg ( clk, reset, g17722, g17688 );
not U_inv80 ( n19386, g17722 );
dff g6711_reg ( clk, reset, g17871, g13099 );
not U_inv81 ( n19381, g17871 );
dff g6715_reg ( clk, reset, g14749, g17871 );
not U_inv82 ( n19383, g14749 );
dff g6719_reg ( clk, reset, g17764, g14749 );
not U_inv83 ( n19382, g17764 );
dff g6723_reg ( clk, reset, ex_wire10, g17764 );
not U_inv84 ( n19384, ex_wire10 );
dff g6727_reg ( clk, reset, n10327, n3035 );
not U_inv85 ( n19789, n10327 );
dff g6736_reg ( clk, reset, n10694, n3045 );
not U_inv86 ( n19791, n10694 );
dff g6732_reg ( clk, reset, ex_wire11, n3040 );
not U_inv87 ( n19790, ex_wire11 );
dff g3298_reg ( clk, reset, g14421, g16624 );
not U_inv88 ( n19377, g14421 );
dff g3303_reg ( clk, reset, g11349, n3353 );
not U_inv89 ( n19375, g11349 );
dff g3281_reg ( clk, reset, g13895, g11349 );
not U_inv90 ( n19823, g13895 );
dff g3310_reg ( clk, reset, g16718, g13895 );
not U_inv91 ( n19824, g16718 );
dff g3267_reg ( clk, reset, g16603, g16718 );
not U_inv92 ( n19825, g16603 );
dff g3274_reg ( clk, reset, g16624, g16603 );
not U_inv93 ( n19376, g16624 );
dff g3317_reg ( clk, reset, g16874, g14421 );
not U_inv94 ( n19371, g16874 );
dff g3321_reg ( clk, reset, g13865, g16874 );
not U_inv95 ( n19373, g13865 );
dff g3325_reg ( clk, reset, g16686, g13865 );
not U_inv96 ( n19372, g16686 );
dff g3329_reg ( clk, reset, ex_wire12, g16686 );
not U_inv97 ( n19374, ex_wire12 );
dff g3338_reg ( clk, reset, n10326, n3394 );
not U_inv98 ( n19826, n10326 );
dff g3347_reg ( clk, reset, n10740, n3404 );
not U_inv99 ( n19828, n10740 );
dff g3343_reg ( clk, reset, ex_wire13, n3399 );
not U_inv100 ( n19827, ex_wire13 );
dff g3649_reg ( clk, reset, g14451, g16656 );
not U_inv101 ( n19367, g14451 );
dff g3654_reg ( clk, reset, g11388, n3712 );
not U_inv102 ( n19365, g11388 );
dff g3632_reg ( clk, reset, g13926, g11388 );
not U_inv103 ( n19860, g13926 );
dff g3661_reg ( clk, reset, g16744, g13926 );
not U_inv104 ( n19861, g16744 );
dff g3618_reg ( clk, reset, g16627, g16744 );
not U_inv105 ( n19862, g16627 );
dff g3625_reg ( clk, reset, g16656, g16627 );
not U_inv106 ( n19366, g16656 );
dff g3668_reg ( clk, reset, g16924, g14451 );
not U_inv107 ( n19361, g16924 );
dff g3672_reg ( clk, reset, g13881, g16924 );
not U_inv108 ( n19363, g13881 );
dff g3676_reg ( clk, reset, g16722, g13881 );
not U_inv109 ( n19362, g16722 );
dff g3680_reg ( clk, reset, ex_wire14, g16722 );
not U_inv110 ( n19364, ex_wire14 );
dff g3689_reg ( clk, reset, n10325, n3753 );
not U_inv111 ( n19863, n10325 );
dff g3698_reg ( clk, reset, n10693, n3763 );
not U_inv112 ( n19865, n10693 );
dff g3694_reg ( clk, reset, ex_wire15, n3758 );
not U_inv113 ( n19864, ex_wire15 );
dff g4000_reg ( clk, reset, g14518, g16693 );
not U_inv114 ( n19357, g14518 );
dff g4005_reg ( clk, reset, g11418, n4071 );
not U_inv115 ( n19355, g11418 );
dff g3983_reg ( clk, reset, g13966, g11418 );
not U_inv116 ( n19896, g13966 );
dff g4012_reg ( clk, reset, g16775, g13966 );
not U_inv117 ( n19897, g16775 );
dff g3969_reg ( clk, reset, g16659, g16775 );
not U_inv118 ( n19898, g16659 );
dff g3976_reg ( clk, reset, g16693, g16659 );
not U_inv119 ( n19356, g16693 );
dff g4019_reg ( clk, reset, g16955, g14518 );
not U_inv120 ( n19351, g16955 );
dff g4023_reg ( clk, reset, g13906, g16955 );
not U_inv121 ( n19353, g13906 );
dff g4027_reg ( clk, reset, g16748, g13906 );
not U_inv122 ( n19352, g16748 );
dff g4031_reg ( clk, reset, ex_wire16, g16748 );
not U_inv123 ( n19354, ex_wire16 );
dff g4040_reg ( clk, reset, n10324, n4112 );
not U_inv124 ( n19899, n10324 );
dff g4049_reg ( clk, reset, n10692, n4122 );
not U_inv125 ( n19901, n10692 );
dff g4045_reg ( clk, reset, ex_wire17, n4117 );
not U_inv126 ( n19900, ex_wire17 );
dff g4165_reg ( clk, reset, new_g25689_, new_g25688_ );
not U_inv127 ( n19107, new_g25689_ );
dff g4169_reg ( clk, reset, n10311, new_g25689_ );
not U_inv128 ( n19346, n10311 );
dff g4125_reg ( clk, reset, n10701, new_g25690_ );
not U_inv129 ( n19347, n10701 );
dff g4098_reg ( clk, reset, n10293, n4485 );
not U_inv130 ( n19939, n10293 );
dff g4072_reg ( clk, reset, ex_wire18, n4445 );
not U_inv131 ( n19345, ex_wire18 );
dff g4064_reg ( clk, reset, n10344, n4450 );
not U_inv132 ( n19932, n10344 );
dff g4057_reg ( clk, reset, n10446, n4455 );
not U_inv133 ( n19933, n10446 );
dff g4141_reg ( clk, reset, n10611, n4460 );
not U_inv134 ( n19934, n10611 );
dff g4082_reg ( clk, reset, ex_wire19, n4465 );
not U_inv135 ( n19935, ex_wire19 );
dff g4076_reg ( clk, reset, n10226, n4470 );
not U_inv136 ( n19936, n10226 );
dff g4087_reg ( clk, reset, n10232, n4475 );
not U_inv137 ( n19937, n10232 );
dff g4093_reg ( clk, reset, n10421, n4480 );
not U_inv138 ( n19938, n10421 );
dff g4108_reg ( clk, reset, n10462, n4490 );
not U_inv139 ( n19940, n10462 );
dff g4104_reg ( clk, reset, n10475, n4495 );
not U_inv140 ( n19426, n10475 );
dff g4258_reg ( clk, reset, n10477, n4575 );
not U_inv141 ( n19947, n10477 );
dff g4264_reg ( clk, reset, n10359, n4580 );
not U_inv142 ( n19318, n10359 );
dff g4269_reg ( clk, reset, n10903, n4585 );
not U_inv143 ( n19948, n10903 );
dff g4273_reg ( clk, reset, n10788, n4590 );
not U_inv144 ( n19317, n10788 );
dff g4239_reg ( clk, reset, ex_wire20, n4595 );
not U_inv145 ( n19316, ex_wire20 );
dff g4297_reg ( clk, reset, n10874, g10122 );
dff g4294_reg ( clk, reset, g10122, n4600 );
dff g305_reg ( clk, reset, n10255, n4736 );
not U_inv146 ( n19954, n10255 );
dff g311_reg ( clk, reset, ex_wire21, n4741 );
not U_inv147 ( n19955, ex_wire21 );
dff g324_reg ( clk, reset, n10395, n4751 );
dff g336_reg ( clk, reset, n10682, n4746 );
not U_inv148 ( n19956, n10682 );
dff g316_reg ( clk, reset, ex_wire22, n4756 );
not U_inv149 ( n19297, ex_wire22 );
dff g319_reg ( clk, reset, n4766, n4761 );
not U_inv150 ( n19957, n4766 );
dff g329_reg ( clk, reset, n10549, n4766 );
dff g333_reg ( clk, reset, n10280, n4771 );
dff g347_reg ( clk, reset, ex_wire23, g7540 );
not U_inv151 ( n19296, ex_wire23 );
dff g344_reg ( clk, reset, g7540, n4776 );
not U_inv152 ( n19295, g7540 );
dff g351_reg ( clk, reset, n10697, n4785 );
not U_inv153 ( n19294, n10697 );
dff g355_reg ( clk, reset, n10873, n4790 );
dff g74_reg ( clk, reset, g20763, n4795 );
dff g341_reg ( clk, reset, g341, n4805 );
dff g106_reg ( clk, reset, g21176, n4800 );
not U_inv154 ( n19293, g21176 );
dff g637_reg ( clk, reset, g12368, n139 );
dff g640_reg ( clk, reset, g9048, g12368 );
not U_inv155 ( n19958, g9048 );
dff g559_reg ( clk, reset, n10834, g9048 );
dff g632_reg ( clk, reset, n10657, n4898 );
not U_inv156 ( n19967, n10657 );
dff g562_reg ( clk, reset, n10403, n4823 );
not U_inv157 ( n19959, n10403 );
dff g568_reg ( clk, reset, n10653, n4828 );
not U_inv158 ( n19328, n10653 );
dff g572_reg ( clk, reset, n10652, n4833 );
not U_inv159 ( n19960, n10652 );
dff g586_reg ( clk, reset, n10505, n4838 );
not U_inv160 ( n19464, n10505 );
dff g577_reg ( clk, reset, n10504, n4843 );
not U_inv161 ( n19961, n10504 );
dff g582_reg ( clk, reset, n10651, n4848 );
not U_inv162 ( n19473, n10651 );
dff g590_reg ( clk, reset, n10650, n4853 );
not U_inv163 ( n19962, n10650 );
dff g595_reg ( clk, reset, n10503, n4858 );
not U_inv164 ( n19487, n10503 );
dff g599_reg ( clk, reset, n10502, n4863 );
not U_inv165 ( n19963, n10502 );
dff g604_reg ( clk, reset, n10649, n4868 );
not U_inv166 ( n19327, n10649 );
dff g608_reg ( clk, reset, n10648, n4873 );
not U_inv167 ( n19964, n10648 );
dff g613_reg ( clk, reset, n10647, n4878 );
not U_inv168 ( n19463, n10647 );
dff g617_reg ( clk, reset, n10646, n4883 );
not U_inv169 ( n19965, n10646 );
dff g622_reg ( clk, reset, n10639, n4888 );
not U_inv170 ( n19474, n10639 );
dff g626_reg ( clk, reset, n10372, n4893 );
not U_inv171 ( n19966, n10372 );
dff g859_reg ( clk, reset, g14189, n4903 );
not U_inv172 ( n19292, g14189 );
dff g869_reg ( clk, reset, g14201, g14189 );
not U_inv173 ( n19290, g14201 );
dff g875_reg ( clk, reset, g14217, g14201 );
not U_inv174 ( n19289, g14217 );
dff g878_reg ( clk, reset, g14096, g14217 );
not U_inv175 ( n19288, g14096 );
dff g881_reg ( clk, reset, g14125, g14096 );
not U_inv176 ( n19287, g14125 );
dff g884_reg ( clk, reset, g14147, g14125 );
not U_inv177 ( n19286, g14147 );
dff g887_reg ( clk, reset, g14167, g14147 );
not U_inv178 ( n19285, g14167 );
dff g872_reg ( clk, reset, ex_wire24, g14167 );
not U_inv179 ( n19291, ex_wire24 );
dff g358_reg ( clk, reset, ex_wire25, g8719 );
not U_inv180 ( n19278, ex_wire25 );
dff g365_reg ( clk, reset, g8719, n5001 );
not U_inv181 ( n19279, g8719 );
dff g385_reg ( clk, reset, n10347, n5020 );
not U_inv182 ( n19979, n10347 );
dff g370_reg ( clk, reset, ex_wire26, n5010 );
not U_inv183 ( n19280, ex_wire26 );
dff g376_reg ( clk, reset, ex_wire27, n5015 );
not U_inv184 ( n19978, ex_wire27 );
dff g203_reg ( clk, reset, ex_wire28, n5025 );
not U_inv185 ( n19264, ex_wire28 );
dff g452_reg ( clk, reset, ex_wire29, n5270 );
not U_inv186 ( n19283, ex_wire29 );
dff g854_reg ( clk, reset, n10773, n5030 );
not U_inv187 ( n19980, n10773 );
dff g847_reg ( clk, reset, n10433, n5035 );
not U_inv188 ( n19981, n10433 );
dff g703_reg ( clk, reset, n10300, n5040 );
not U_inv189 ( n19982, n10300 );
dff g837_reg ( clk, reset, n10256, n5045 );
not U_inv190 ( n19983, n10256 );
dff g843_reg ( clk, reset, n10899, n5050 );
not U_inv191 ( n19275, n10899 );
dff g812_reg ( clk, reset, n10456, n5055 );
not U_inv192 ( n19984, n10456 );
dff g817_reg ( clk, reset, n10599, n5060 );
not U_inv193 ( n19985, n10599 );
dff g832_reg ( clk, reset, ex_wire30, n5065 );
not U_inv194 ( n19276, ex_wire30 );
dff g822_reg ( clk, reset, n10664, n5070 );
not U_inv195 ( n19277, n10664 );
dff g827_reg ( clk, reset, n10605, n5075 );
not U_inv196 ( n19986, n10605 );
dff g723_reg ( clk, reset, n10904, n5080 );
not U_inv197 ( n19987, n10904 );
dff g890_reg ( clk, reset, n10600, n4976 );
not U_inv198 ( n19976, n10600 );
dff g862_reg ( clk, reset, n10331, n4981 );
dff g896_reg ( clk, reset, n10283, n4986 );
not U_inv199 ( n19977, n10283 );
dff g225_reg ( clk, reset, n10230, n4936 );
not U_inv200 ( n19968, n10230 );
dff g255_reg ( clk, reset, n10253, n4941 );
not U_inv201 ( n19969, n10253 );
dff g232_reg ( clk, reset, n10335, n4946 );
not U_inv202 ( n19970, n10335 );
dff g262_reg ( clk, reset, n10458, n4951 );
not U_inv203 ( n19971, n10458 );
dff g239_reg ( clk, reset, n10241, n4956 );
not U_inv204 ( n19972, n10241 );
dff g269_reg ( clk, reset, n10431, n4961 );
not U_inv205 ( n19973, n10431 );
dff g246_reg ( clk, reset, n10349, n4966 );
not U_inv206 ( n19974, n10349 );
dff g446_reg ( clk, reset, n10365, n4971 );
not U_inv207 ( n19975, n10365 );
dff g417_reg ( clk, reset, n10229, n5195 );
not U_inv208 ( n20000, n10229 );
dff g411_reg ( clk, reset, n10352, n5200 );
dff g424_reg ( clk, reset, n10506, n5205 );
not U_inv209 ( n20001, n10506 );
dff g475_reg ( clk, reset, ex_wire31, n5210 );
not U_inv210 ( n19267, ex_wire31 );
dff g441_reg ( clk, reset, n10548, n5215 );
dff g437_reg ( clk, reset, n10543, n5220 );
dff g433_reg ( clk, reset, ex_wire32, n5225 );
not U_inv211 ( n19266, ex_wire32 );
dff g429_reg ( clk, reset, n10871, n5230 );
dff g401_reg ( clk, reset, n10544, n5235 );
dff g392_reg ( clk, reset, n10271, n5240 );
not U_inv212 ( n20002, n10271 );
dff g405_reg ( clk, reset, n10415, n5245 );
not U_inv213 ( n19284, n10415 );
dff g182_reg ( clk, reset, n10278, n5250 );
not U_inv214 ( n19281, n10278 );
dff g174_reg ( clk, reset, n10561, n5255 );
not U_inv215 ( n19282, n10561 );
dff g168_reg ( clk, reset, n10578, n5260 );
not U_inv216 ( n19265, n10578 );
dff g460_reg ( clk, reset, n10870, n5265 );
dff g645_reg ( clk, reset, n10786, n5085 );
not U_inv217 ( n19988, n10786 );
dff g681_reg ( clk, reset, n10260, n5090 );
dff g699_reg ( clk, reset, n10836, n5095 );
not U_inv218 ( n19989, n10836 );
dff g650_reg ( clk, reset, n10722, n5100 );
not U_inv219 ( n19990, n10722 );
dff g655_reg ( clk, reset, n10277, n5105 );
not U_inv220 ( n19274, n10277 );
dff g718_reg ( clk, reset, n10333, n5110 );
not U_inv221 ( n19273, n10333 );
dff g661_reg ( clk, reset, n10662, n5115 );
not U_inv222 ( n19272, n10662 );
dff g728_reg ( clk, reset, ex_wire33, n5120 );
not U_inv223 ( n19271, ex_wire33 );
dff g79_reg ( clk, reset, g20899, n5125 );
dff g691_reg ( clk, reset, n10307, n5130 );
not U_inv224 ( n19991, n10307 );
dff g686_reg ( clk, reset, ex_wire34, n5135 );
not U_inv225 ( n19992, ex_wire34 );
dff g667_reg ( clk, reset, n10538, n5140 );
dff g504_reg ( clk, reset, n10404, n5165 );
not U_inv226 ( n19996, n10404 );
dff g513_reg ( clk, reset, n10384, n5170 );
not U_inv227 ( n19268, n10384 );
dff g518_reg ( clk, reset, n10224, n5175 );
not U_inv228 ( n19997, n10224 );
dff g528_reg ( clk, reset, n10345, n5180 );
not U_inv229 ( n19998, n10345 );
dff g482_reg ( clk, reset, ex_wire35, n5185 );
not U_inv230 ( n19999, ex_wire35 );
dff g490_reg ( clk, reset, ex_wire36, n5190 );
not U_inv231 ( n19270, ex_wire36 );
dff g499_reg ( clk, reset, n10661, n5160 );
not U_inv232 ( n19995, n10661 );
dff g671_reg ( clk, reset, ex_wire37, n5145 );
not U_inv233 ( n19269, ex_wire37 );
dff g676_reg ( clk, reset, n10656, n5150 );
not U_inv234 ( n19993, n10656 );
dff g714_reg ( clk, reset, n10663, n5155 );
not U_inv235 ( n19994, n10663 );
dff g479_reg ( clk, reset, ex_wire38, n5295 );
not U_inv236 ( n19263, ex_wire38 );
dff g102_reg ( clk, reset, g20901, n5300 );
dff g496_reg ( clk, reset, g496, n5305 );
dff g732_reg ( clk, reset, n10898, n5310 );
dff g753_reg ( clk, reset, n10814, n5315 );
not U_inv237 ( n20003, n10814 );
dff g799_reg ( clk, reset, g12184, n5320 );
dff g802_reg ( clk, reset, g11678, g12184 );
not U_inv238 ( n20004, g11678 );
dff g736_reg ( clk, reset, n10581, g11678 );
dff g554_reg ( clk, reset, n10794, n5398 );
not U_inv239 ( n20009, n10794 );
dff g739_reg ( clk, reset, ex_wire39, n5333 );
not U_inv240 ( n20005, ex_wire39 );
dff g744_reg ( clk, reset, n10501, n5338 );
not U_inv241 ( n20006, n10501 );
dff g749_reg ( clk, reset, n10500, n5343 );
not U_inv242 ( n19335, n10500 );
dff g758_reg ( clk, reset, n10645, n5348 );
not U_inv243 ( n20007, n10645 );
dff g763_reg ( clk, reset, n10644, n5353 );
not U_inv244 ( n19467, n10644 );
dff g767_reg ( clk, reset, n10499, n5358 );
not U_inv245 ( n19476, n10499 );
dff g772_reg ( clk, reset, n10498, n5363 );
not U_inv246 ( n19482, n10498 );
dff g776_reg ( clk, reset, n10496, n5368 );
not U_inv247 ( n19488, n10496 );
dff g781_reg ( clk, reset, n10497, n5373 );
not U_inv248 ( n19320, n10497 );
dff g785_reg ( clk, reset, n10643, n5378 );
not U_inv249 ( n19326, n10643 );
dff g790_reg ( clk, reset, n10494, n5383 );
not U_inv250 ( n19337, n10494 );
dff g794_reg ( clk, reset, n10495, n5388 );
not U_inv251 ( n19462, n10495 );
dff g807_reg ( clk, reset, n10608, n5393 );
not U_inv252 ( n20008, n10608 );
dff g278_reg ( clk, reset, n10900, n5438 );
not U_inv253 ( n20010, n10900 );
dff g283_reg ( clk, reset, n10902, n5443 );
not U_inv254 ( n20011, n10902 );
dff g287_reg ( clk, reset, ex_wire40, n5448 );
not U_inv255 ( n19260, ex_wire40 );
dff g291_reg ( clk, reset, n10750, n5453 );
not U_inv256 ( n20012, n10750 );
dff g294_reg ( clk, reset, n10681, n5458 );
not U_inv257 ( n19259, n10681 );
dff g298_reg ( clk, reset, n10522, n5463 );
not U_inv258 ( n19258, n10522 );
dff g142_reg ( clk, reset, n10699, n5468 );
not U_inv259 ( n19257, n10699 );
dff g146_reg ( clk, reset, ex_wire41, n5473 );
not U_inv260 ( n19256, ex_wire41 );
dff g164_reg ( clk, reset, n10749, n5478 );
not U_inv261 ( n20013, n10749 );
dff g150_reg ( clk, reset, n10748, n5483 );
not U_inv262 ( n19255, n10748 );
dff g153_reg ( clk, reset, n10747, n5488 );
not U_inv263 ( n20014, n10747 );
dff g157_reg ( clk, reset, n10680, n5493 );
not U_inv264 ( n19254, n10680 );
dff g160_reg ( clk, reset, ex_wire42, n5498 );
not U_inv265 ( n20015, ex_wire42 );
dff g301_reg ( clk, reset, ex_wire43, n5503 );
not U_inv266 ( n19262, ex_wire43 );
dff g222_reg ( clk, reset, ex_wire44, n5508 );
not U_inv267 ( n19261, ex_wire44 );
dff g218_reg ( clk, reset, ex_wire45, g8291 );
not U_inv268 ( n19253, ex_wire45 );
dff g194_reg ( clk, reset, g8358, n5513 );
not U_inv269 ( n19251, g8358 );
dff g191_reg ( clk, reset, ex_wire46, g8358 );
not U_inv270 ( n19252, ex_wire46 );
dff g209_reg ( clk, reset, n10252, n5522 );
dff g215_reg ( clk, reset, g8291, n5527 );
not U_inv271 ( n10941, g8291 );
dff g1389_reg ( clk, reset, n10618, n5772 );
not U_inv272 ( n20043, n10618 );
dff g1312_reg ( clk, reset, n10607, n5732 );
not U_inv273 ( n20036, n10607 );
dff g1418_reg ( clk, reset, g17320, n5586 );
not U_inv274 ( n20023, g17320 );
dff g1422_reg ( clk, reset, g17404, g17320 );
not U_inv275 ( n19247, g17404 );
dff g1426_reg ( clk, reset, g17423, g17404 );
not U_inv276 ( n19248, g17423 );
dff g1430_reg ( clk, reset, n10590, g17423 );
not U_inv277 ( n19246, n10590 );
dff g1548_reg ( clk, reset, n10660, n5603 );
not U_inv278 ( n19245, n10660 );
dff g1564_reg ( clk, reset, n10620, n5608 );
not U_inv279 ( n19244, n10620 );
dff g1559_reg ( clk, reset, n10480, n5613 );
not U_inv280 ( n19242, n10480 );
dff g1554_reg ( clk, reset, n10449, n5618 );
not U_inv281 ( n19243, n10449 );
dff g1570_reg ( clk, reset, g12923, n5623 );
not U_inv282 ( n20024, g12923 );
dff g1585_reg ( clk, reset, n10473, g12923 );
not U_inv283 ( n20025, n10473 );
dff g1589_reg ( clk, reset, n10337, n5632 );
not U_inv284 ( n20026, n10337 );
dff g1249_reg ( clk, reset, n10483, n5536 );
not U_inv285 ( n19250, n10483 );
dff g1266_reg ( clk, reset, n10670, n5541 );
not U_inv286 ( n19249, n10670 );
dff g1280_reg ( clk, reset, n10655, n5546 );
not U_inv287 ( n20016, n10655 );
dff g1252_reg ( clk, reset, n10746, n5551 );
not U_inv288 ( n20017, n10746 );
dff g1256_reg ( clk, reset, n10745, n5556 );
not U_inv289 ( n20018, n10745 );
dff g1259_reg ( clk, reset, n10744, n5561 );
not U_inv290 ( n20019, n10744 );
dff g1263_reg ( clk, reset, n10679, n5566 );
not U_inv291 ( n20020, n10679 );
dff g1270_reg ( clk, reset, n10521, n5571 );
not U_inv292 ( n20021, n10521 );
dff g1274_reg ( clk, reset, n10911, n5576 );
not U_inv293 ( n20022, n10911 );
dff g1576_reg ( clk, reset, g10527, n5637 );
dff g1579_reg ( clk, reset, ex_wire47, g10527 );
not U_inv294 ( n19241, ex_wire47 );
dff g1339_reg ( clk, reset, n10240, n5646 );
not U_inv295 ( n20027, n10240 );
dff g1500_reg ( clk, reset, g7946, n5651 );
not U_inv296 ( n20028, g7946 );
dff g1582_reg ( clk, reset, g8475, g7946 );
dff g1333_reg ( clk, reset, n10401, g8475 );
not U_inv297 ( n20029, n10401 );
dff g1399_reg ( clk, reset, g19357, n5664 );
not U_inv298 ( n19240, g19357 );
dff g1459_reg ( clk, reset, g13272, g19357 );
not U_inv299 ( n19239, g13272 );
dff g1322_reg ( clk, reset, n10286, g13272 );
not U_inv300 ( n20030, n10286 );
dff g1395_reg ( clk, reset, n10417, n5717 );
not U_inv301 ( n20034, n10417 );
dff g1404_reg ( clk, reset, n10642, n5722 );
not U_inv302 ( n20035, n10642 );
dff g1319_reg ( clk, reset, ex_wire48, n5727 );
not U_inv303 ( n19235, ex_wire48 );
dff g1351_reg ( clk, reset, ex_wire49, n5737 );
not U_inv304 ( n20037, ex_wire49 );
dff g1345_reg ( clk, reset, n10258, n5742 );
not U_inv305 ( n20038, n10258 );
dff g1361_reg ( clk, reset, ex_wire50, n5747 );
not U_inv306 ( n20039, ex_wire50 );
dff g1367_reg ( clk, reset, n10394, n5752 );
not U_inv307 ( n20040, n10394 );
dff g1373_reg ( clk, reset, n10318, n5757 );
not U_inv308 ( n20041, n10318 );
dff g1379_reg ( clk, reset, n10638, n5762 );
not U_inv309 ( n19238, n10638 );
dff g1384_reg ( clk, reset, n10519, n5767 );
not U_inv310 ( n20042, n10519 );
dff g1514_reg ( clk, reset, n10582, n5677 );
not U_inv311 ( n20031, n10582 );
dff g1526_reg ( clk, reset, n10303, n5682 );
not U_inv312 ( n20032, n10303 );
dff g1521_reg ( clk, reset, n10363, n5687 );
dff g1306_reg ( clk, reset, n10492, n5692 );
not U_inv313 ( n19523, n10492 );
dff g1532_reg ( clk, reset, n10361, n5697 );
dff g1536_reg ( clk, reset, n10676, n5702 );
not U_inv314 ( n20033, n10676 );
dff g1542_reg ( clk, reset, n10419, n5707 );
dff g1413_reg ( clk, reset, ex_wire51, n5712 );
not U_inv315 ( n19237, ex_wire51 );
dff g1277_reg ( clk, reset, ex_wire52, n5581 );
not U_inv316 ( n19230, ex_wire52 );
dff g1442_reg ( clk, reset, n10371, n5787 );
not U_inv317 ( n19236, n10371 );
dff g1489_reg ( clk, reset, ex_wire53, n5777 );
not U_inv318 ( n20044, ex_wire53 );
dff g1495_reg ( clk, reset, n10669, n5782 );
not U_inv319 ( n20045, n10669 );
dff g1478_reg ( clk, reset, n10455, n5797 );
not U_inv320 ( n20046, n10455 );
dff g1437_reg ( clk, reset, n10918, n5792 );
not U_inv321 ( n19234, n10918 );
dff g1448_reg ( clk, reset, n10323, n5807 );
not U_inv322 ( n20047, n10323 );
dff g1454_reg ( clk, reset, n10910, n5802 );
not U_inv323 ( n19233, n10910 );
dff g1472_reg ( clk, reset, n10453, n5817 );
not U_inv324 ( n20048, n10453 );
dff g1467_reg ( clk, reset, n10917, n5812 );
not U_inv325 ( n19232, n10917 );
dff g1300_reg ( clk, reset, n10622, n5827 );
not U_inv326 ( n20049, n10622 );
dff g1484_reg ( clk, reset, n10916, n5822 );
not U_inv327 ( n19231, n10916 );
dff g1046_reg ( clk, reset, n10617, n6098 );
not U_inv328 ( n20081, n10617 );
dff g969_reg ( clk, reset, n10606, n6058 );
not U_inv329 ( n20074, n10606 );
dff g1075_reg ( clk, reset, g17291, n5912 );
not U_inv330 ( n20059, g17291 );
dff g1079_reg ( clk, reset, g17316, g17291 );
not U_inv331 ( n19226, g17316 );
dff g1083_reg ( clk, reset, g17400, g17316 );
not U_inv332 ( n19227, g17400 );
dff g1087_reg ( clk, reset, n10589, g17400 );
not U_inv333 ( n19225, n10589 );
dff g1205_reg ( clk, reset, n10659, n5929 );
not U_inv334 ( n19224, n10659 );
dff g1221_reg ( clk, reset, n10619, n5934 );
not U_inv335 ( n19223, n10619 );
dff g1216_reg ( clk, reset, n10479, n5939 );
not U_inv336 ( n19221, n10479 );
dff g1211_reg ( clk, reset, n10448, n5944 );
not U_inv337 ( n19222, n10448 );
dff g1227_reg ( clk, reset, g12919, n5949 );
not U_inv338 ( n20060, g12919 );
dff g1242_reg ( clk, reset, g23683, g12919 );
not U_inv339 ( n20061, g23683 );
dff g1246_reg ( clk, reset, n10338, n5958 );
not U_inv340 ( n20062, n10338 );
dff g904_reg ( clk, reset, n10482, n5862 );
not U_inv341 ( n19229, n10482 );
dff g921_reg ( clk, reset, n10668, n5867 );
not U_inv342 ( n19228, n10668 );
dff g936_reg ( clk, reset, n10654, n5872 );
not U_inv343 ( n20052, n10654 );
dff g907_reg ( clk, reset, n10743, n5877 );
not U_inv344 ( n20053, n10743 );
dff g911_reg ( clk, reset, n10742, n5882 );
not U_inv345 ( n20054, n10742 );
dff g914_reg ( clk, reset, n10741, n5887 );
not U_inv346 ( n20055, n10741 );
dff g918_reg ( clk, reset, n10678, n5892 );
not U_inv347 ( n20056, n10678 );
dff g925_reg ( clk, reset, n10520, n5897 );
not U_inv348 ( n20057, n10520 );
dff g930_reg ( clk, reset, n10909, n5902 );
not U_inv349 ( n20058, n10909 );
dff g1233_reg ( clk, reset, g10500, n5963 );
dff g1236_reg ( clk, reset, ex_wire54, g10500 );
not U_inv350 ( n19220, ex_wire54 );
dff g996_reg ( clk, reset, n10239, n5972 );
not U_inv351 ( n20063, n10239 );
dff g1157_reg ( clk, reset, g7916, n5977 );
not U_inv352 ( n20064, g7916 );
dff g1239_reg ( clk, reset, g8416, g7916 );
dff g990_reg ( clk, reset, n10400, g8416 );
not U_inv353 ( n20065, n10400 );
dff g1056_reg ( clk, reset, g19334, n5990 );
not U_inv354 ( n19219, g19334 );
dff g1116_reg ( clk, reset, g13259, g19334 );
not U_inv355 ( n19218, g13259 );
dff g979_reg ( clk, reset, n10285, g13259 );
not U_inv356 ( n20066, n10285 );
dff g1052_reg ( clk, reset, n10416, n6043 );
not U_inv357 ( n20072, n10416 );
dff g1061_reg ( clk, reset, n10641, n6048 );
not U_inv358 ( n20073, n10641 );
dff g976_reg ( clk, reset, ex_wire55, n6053 );
not U_inv359 ( n19214, ex_wire55 );
dff g1008_reg ( clk, reset, ex_wire56, n6063 );
not U_inv360 ( n20075, ex_wire56 );
dff g1002_reg ( clk, reset, n10257, n6068 );
not U_inv361 ( n20076, n10257 );
dff g1018_reg ( clk, reset, ex_wire57, n6073 );
not U_inv362 ( n20077, ex_wire57 );
dff g1024_reg ( clk, reset, n10393, n6078 );
not U_inv363 ( n20078, n10393 );
dff g1030_reg ( clk, reset, n10317, n6083 );
not U_inv364 ( n20079, n10317 );
dff g1036_reg ( clk, reset, n10637, n6088 );
not U_inv365 ( n19217, n10637 );
dff g1041_reg ( clk, reset, n10518, n6093 );
not U_inv366 ( n20080, n10518 );
dff g1171_reg ( clk, reset, n10580, n6003 );
not U_inv367 ( n20067, n10580 );
dff g1183_reg ( clk, reset, n10294, n6008 );
not U_inv368 ( n20068, n10294 );
dff g1178_reg ( clk, reset, n10387, n6013 );
not U_inv369 ( n20069, n10387 );
dff g962_reg ( clk, reset, n10381, n6018 );
not U_inv370 ( n20070, n10381 );
dff g1189_reg ( clk, reset, n10360, n6023 );
dff g1193_reg ( clk, reset, n10675, n6028 );
not U_inv371 ( n20071, n10675 );
dff g1199_reg ( clk, reset, n10418, n6033 );
dff g1070_reg ( clk, reset, ex_wire58, n6038 );
not U_inv372 ( n19216, ex_wire58 );
dff g933_reg ( clk, reset, ex_wire59, n5907 );
not U_inv373 ( n19209, ex_wire59 );
dff g1099_reg ( clk, reset, n10370, n6113 );
not U_inv374 ( n19215, n10370 );
dff g1146_reg ( clk, reset, ex_wire60, n6103 );
not U_inv375 ( n20082, ex_wire60 );
dff g1152_reg ( clk, reset, n10667, n6108 );
not U_inv376 ( n20083, n10667 );
dff g1135_reg ( clk, reset, n10454, n6123 );
not U_inv377 ( n20084, n10454 );
dff g1094_reg ( clk, reset, n10915, n6118 );
not U_inv378 ( n19213, n10915 );
dff g1105_reg ( clk, reset, n10322, n6133 );
not U_inv379 ( n20085, n10322 );
dff g1111_reg ( clk, reset, n10908, n6128 );
not U_inv380 ( n19212, n10908 );
dff g1129_reg ( clk, reset, n10452, n6143 );
not U_inv381 ( n20086, n10452 );
dff g1124_reg ( clk, reset, n10914, n6138 );
not U_inv382 ( n19211, n10914 );
dff g956_reg ( clk, reset, n10621, n6153 );
not U_inv383 ( n20087, n10621 );
dff g1141_reg ( clk, reset, n10913, n6148 );
not U_inv384 ( n19210, n10913 );
dff g2837_reg ( clk, reset, new_g24265_, new_g25688_ );
not U_inv385 ( n19108, new_g24265_ );
dff g2841_reg ( clk, reset, n10476, new_g24265_ );
not U_inv386 ( n19141, n10476 );
dff g2712_reg ( clk, reset, n10922, new_g24266_ );
not U_inv387 ( n19140, n10922 );
dff g2715_reg ( clk, reset, n10225, n7293 );
not U_inv388 ( n20198, n10225 );
dff g2719_reg ( clk, reset, n10420, n7298 );
not U_inv389 ( n20199, n10420 );
dff g2724_reg ( clk, reset, n10228, n7303 );
not U_inv390 ( n20200, n10228 );
dff g2729_reg ( clk, reset, n10332, n7308 );
not U_inv391 ( n20201, n10332 );
dff g2735_reg ( clk, reset, n10437, n7313 );
not U_inv392 ( n20202, n10437 );
dff g2741_reg ( clk, reset, n10231, n7318 );
not U_inv393 ( n20203, n10231 );
dff g2748_reg ( clk, reset, n10222, n7323 );
not U_inv394 ( n20204, n10222 );
dff g2756_reg ( clk, reset, n10405, n7328 );
not U_inv395 ( n20205, n10405 );
dff g2759_reg ( clk, reset, n10461, n7333 );
not U_inv396 ( n20206, n10461 );
dff g2763_reg ( clk, reset, n10474, n7338 );
not U_inv397 ( n19201, n10474 );
dff g4927_reg ( clk, reset, n10703, n1284 );
not U_inv398 ( n19604, n10703 );
dff g49_reg ( clk, reset, ex_wire61, new_g34977_ );
not U_inv399 ( n19459, ex_wire61 );
dff g16_reg ( clk, reset, n10343, new_g34977_ );
not U_inv400 ( n20234, n10343 );
dff g4737_reg ( clk, reset, n10702, n1451 );
not U_inv401 ( n19619, n10702 );
dff g59_reg ( clk, reset, g20049, n210 );
not U_inv402 ( n19442, g20049 );
dff g4575_reg ( clk, reset, ex_wire62, n1471 );
not U_inv403 ( n19116, ex_wire62 );
dff g4540_reg ( clk, reset, g4540, n940 );
dff g4543_reg ( clk, reset, g4543, n945 );
dff g4567_reg ( clk, reset, g4567, n950 );
dff g4546_reg ( clk, reset, g4546, n955 );
dff g4549_reg ( clk, reset, ex_wire63, n960 );
not U_inv404 ( n19115, ex_wire63 );
dff g4552_reg ( clk, reset, n10940, n965 );
not U_inv405 ( n19114, n10940 );
dff g4570_reg ( clk, reset, g4570, n970 );
dff g4571_reg ( clk, reset, n979, g4570 );
dff g4555_reg ( clk, reset, ex_wire64, n979 );
not U_inv406 ( n19574, ex_wire64 );
dff g4558_reg ( clk, reset, ex_wire65, n984 );
not U_inv407 ( n19113, ex_wire65 );
dff g4561_reg ( clk, reset, ex_wire66, n989 );
not U_inv408 ( n19112, ex_wire66 );
dff g4564_reg ( clk, reset, g4564, n994 );
dff g4534_reg ( clk, reset, ex_wire67, n999 );
not U_inv409 ( n19513, ex_wire67 );
dff g4420_reg ( clk, reset, n10897, n1004 );
dff g2864_reg ( clk, reset, n10770, n7513 );
not U_inv410 ( n19478, n10770 );
dff g47_reg ( clk, reset, g47, new_g34975_ );
dff g8_reg ( clk, reset, ex_wire68, new_g34975_ );
not U_inv411 ( n19497, ex_wire68 );
dff g2994_reg ( clk, reset, n10517, n7448 );
not U_inv412 ( n20216, n10517 );
dff g2988_reg ( clk, reset, n10481, n7453 );
not U_inv413 ( n20217, n10481 );
dff g48_reg ( clk, reset, g48, new_g34976_ );
dff g9_reg ( clk, reset, ex_wire69, new_g34976_ );
not U_inv414 ( n19498, ex_wire69 );
dff g2894_reg ( clk, reset, n10542, n7488 );
dff g37_reg ( clk, reset, n10386, n7493 );
not U_inv415 ( g30327, n10386 );
dff g3863_reg ( clk, reset, n10463, n4250 );
not U_inv416 ( n19905, n10463 );
dff g3869_reg ( clk, reset, n10396, n4255 );
not U_inv417 ( n19906, n10396 );
dff g3873_reg ( clk, reset, n10272, n4260 );
not U_inv418 ( n19907, n10272 );
dff g3881_reg ( clk, reset, n10595, n4265 );
not U_inv419 ( n19908, n10595 );
dff g3794_reg ( clk, reset, g8344, n4137 );
not U_inv420 ( n19903, g8344 );
dff g3802_reg ( clk, reset, n10876, g8344 );
dff g3752_reg ( clk, reset, n10875, n4146 );
dff g3798_reg ( clk, reset, g8398, n4151 );
dff g3857_reg ( clk, reset, n10244, n4245 );
not U_inv421 ( n19904, n10244 );
dff g3512_reg ( clk, reset, n10464, n3891 );
not U_inv422 ( n19869, n10464 );
dff g3518_reg ( clk, reset, n10397, n3896 );
not U_inv423 ( n19870, n10397 );
dff g3522_reg ( clk, reset, n10273, n3901 );
not U_inv424 ( n19871, n10273 );
dff g3530_reg ( clk, reset, n10596, n3906 );
not U_inv425 ( n19872, n10596 );
dff g3443_reg ( clk, reset, g8279, n3778 );
not U_inv426 ( n19867, g8279 );
dff g3451_reg ( clk, reset, n10878, g8279 );
dff g3401_reg ( clk, reset, n10877, n3787 );
dff g3447_reg ( clk, reset, g8342, n3792 );
dff g3506_reg ( clk, reset, n10245, n3886 );
not U_inv427 ( n19868, n10245 );
dff g3155_reg ( clk, reset, n10276, n3527 );
not U_inv428 ( n19832, n10276 );
dff g3161_reg ( clk, reset, n10465, n3532 );
not U_inv429 ( n19833, n10465 );
dff g3167_reg ( clk, reset, n10336, n3537 );
not U_inv430 ( n19834, n10336 );
dff g3171_reg ( clk, reset, n10432, n3542 );
not U_inv431 ( n19835, n10432 );
dff g3179_reg ( clk, reset, n10266, n3547 );
not U_inv432 ( n19836, n10266 );
dff g3092_reg ( clk, reset, g8215, n3419 );
not U_inv433 ( n19831, g8215 );
dff g3100_reg ( clk, reset, n10880, g8215 );
dff g3050_reg ( clk, reset, n10879, n3428 );
dff g3096_reg ( clk, reset, g8277, n3433 );
dff g6555_reg ( clk, reset, n10466, n3173 );
not U_inv434 ( n19795, n10466 );
dff g6561_reg ( clk, reset, n10304, n3178 );
not U_inv435 ( n19796, n10304 );
dff g6565_reg ( clk, reset, n10434, n3183 );
not U_inv436 ( n19797, n10434 );
dff g6573_reg ( clk, reset, n10267, n3188 );
not U_inv437 ( n19798, n10267 );
dff g6486_reg ( clk, reset, g9743, n3060 );
not U_inv438 ( n19793, g9743 );
dff g6494_reg ( clk, reset, n10882, g9743 );
dff g6444_reg ( clk, reset, n10881, n3069 );
dff g6490_reg ( clk, reset, g9817, n3074 );
dff g6549_reg ( clk, reset, n10246, n3168 );
not U_inv439 ( n19794, n10246 );
dff g6209_reg ( clk, reset, n10467, n2814 );
not U_inv440 ( n19759, n10467 );
dff g6215_reg ( clk, reset, n10398, n2819 );
not U_inv441 ( n19760, n10398 );
dff g6219_reg ( clk, reset, n10274, n2824 );
not U_inv442 ( n19761, n10274 );
dff g6227_reg ( clk, reset, n10597, n2829 );
not U_inv443 ( n19762, n10597 );
dff g6140_reg ( clk, reset, g9682, n2701 );
not U_inv444 ( n19757, g9682 );
dff g6148_reg ( clk, reset, n10884, g9682 );
dff g6098_reg ( clk, reset, n10883, n2710 );
dff g6144_reg ( clk, reset, g9741, n2715 );
dff g6203_reg ( clk, reset, n10247, n2809 );
not U_inv445 ( n19758, n10247 );
dff g5863_reg ( clk, reset, n10468, n2455 );
not U_inv446 ( n19722, n10468 );
dff g5869_reg ( clk, reset, n10399, n2460 );
not U_inv447 ( n19723, n10399 );
dff g5873_reg ( clk, reset, n10275, n2465 );
not U_inv448 ( n19724, n10275 );
dff g5881_reg ( clk, reset, n10598, n2470 );
not U_inv449 ( n19725, n10598 );
dff g5794_reg ( clk, reset, g9617, n2342 );
not U_inv450 ( n19720, g9617 );
dff g5802_reg ( clk, reset, n10886, g9617 );
dff g5752_reg ( clk, reset, n10885, n2351 );
dff g5798_reg ( clk, reset, g9680, n2356 );
dff g5857_reg ( clk, reset, n10248, n2450 );
not U_inv451 ( n19721, n10248 );
dff g5517_reg ( clk, reset, n10469, n2096 );
not U_inv452 ( n19686, n10469 );
dff g5523_reg ( clk, reset, n10305, n2101 );
not U_inv453 ( n19687, n10305 );
dff g5527_reg ( clk, reset, n10435, n2106 );
not U_inv454 ( n19688, n10435 );
dff g5535_reg ( clk, reset, n10268, n2111 );
not U_inv455 ( n19689, n10268 );
dff g5448_reg ( clk, reset, g9555, n1983 );
not U_inv456 ( n19684, g9555 );
dff g5456_reg ( clk, reset, n10888, g9555 );
dff g5406_reg ( clk, reset, n10887, n1992 );
dff g5452_reg ( clk, reset, g9615, n1997 );
dff g5511_reg ( clk, reset, n10249, n2091 );
not U_inv457 ( n19685, n10249 );
dff g5170_reg ( clk, reset, n10470, n1737 );
not U_inv458 ( n19651, n10470 );
dff g5176_reg ( clk, reset, n10306, n1742 );
not U_inv459 ( n19652, n10306 );
dff g5180_reg ( clk, reset, n10436, n1747 );
not U_inv460 ( n19653, n10436 );
dff g5188_reg ( clk, reset, n10269, n1752 );
not U_inv461 ( n19654, n10269 );
dff g43_reg ( clk, reset, ex_wire70, new_g34663_ );
not U_inv462 ( n19425, ex_wire70 );
dff g5101_reg ( clk, reset, g9497, n1624 );
not U_inv463 ( n19633, g9497 );
dff g5109_reg ( clk, reset, n10890, g9497 );
dff g5062_reg ( clk, reset, n10236, n1633 );
not U_inv464 ( n19634, n10236 );
dff g5105_reg ( clk, reset, g9553, n1638 );
not U_inv465 ( n19635, g9553 );
dff g5112_reg ( clk, reset, n10889, g9553 );
dff g5022_reg ( clk, reset, n10603, n1647 );
not U_inv466 ( n19636, n10603 );
dff g5016_reg ( clk, reset, n10362, n1652 );
not U_inv467 ( n19637, n10362 );
dff g5033_reg ( clk, reset, n10594, n1662 );
not U_inv468 ( n19638, n10594 );
dff g5037_reg ( clk, reset, n10591, n1667 );
not U_inv469 ( n19639, n10591 );
dff g5041_reg ( clk, reset, n10583, n1672 );
not U_inv470 ( n19640, n10583 );
dff g5046_reg ( clk, reset, ex_wire71, n1677 );
not U_inv471 ( n19641, ex_wire71 );
dff g5052_reg ( clk, reset, n10447, n1682 );
not U_inv472 ( n19429, n10447 );
dff g5057_reg ( clk, reset, n10445, n1687 );
not U_inv473 ( n19642, n10445 );
dff g5069_reg ( clk, reset, n10579, n1692 );
not U_inv474 ( n19643, n10579 );
dff g5073_reg ( clk, reset, ex_wire72, n1697 );
not U_inv475 ( n19644, ex_wire72 );
dff g5077_reg ( clk, reset, ex_wire73, n1702 );
not U_inv476 ( n19645, ex_wire73 );
dff g5084_reg ( clk, reset, n10402, n1712 );
not U_inv477 ( n19647, n10402 );
dff g5092_reg ( clk, reset, ex_wire74, n1717 );
not U_inv478 ( n19427, ex_wire74 );
dff g5097_reg ( clk, reset, ex_wire75, n1722 );
not U_inv479 ( n19648, ex_wire75 );
dff g86_reg ( clk, reset, g20557, n1727 );
not U_inv480 ( n19649, g20557 );
dff g5080_reg ( clk, reset, n10923, n1707 );
not U_inv481 ( n19646, n10923 );
dff g5029_reg ( clk, reset, n10901, n1657 );
not U_inv482 ( n19428, n10901 );
dff g5164_reg ( clk, reset, n10250, n1732 );
not U_inv483 ( n19650, n10250 );
dff g4639_reg ( clk, reset, n10593, n40 );
not U_inv484 ( n19582, n10593 );
dff g4621_reg ( clk, reset, n10601, n1129 );
not U_inv485 ( n19583, n10601 );
dff g4628_reg ( clk, reset, n10666, n1134 );
not U_inv486 ( n19584, n10666 );
dff g4633_reg ( clk, reset, n10658, n1139 );
not U_inv487 ( n19585, n10658 );
dff g4643_reg ( clk, reset, ex_wire76, n1144 );
not U_inv488 ( n19586, ex_wire76 );
dff g4462_reg ( clk, reset, n10259, n832 );
not U_inv489 ( n19573, n10259 );
dff g4467_reg ( clk, reset, g4467, n842 );
not U_inv490 ( n19126, g4467 );
dff g4474_reg ( clk, reset, n852, g4467 );
not U_inv491 ( n19127, n852 );
dff g4477_reg ( clk, reset, ex_wire77, n852 );
not U_inv492 ( n19128, ex_wire77 );
dff g4459_reg ( clk, reset, ex_wire78, n817 );
not U_inv493 ( n19129, ex_wire78 );
dff g4507_reg ( clk, reset, ex_wire79, n812 );
not U_inv494 ( n19570, ex_wire79 );
dff g4473_reg ( clk, reset, n10254, n827 );
not U_inv495 ( n19572, n10254 );
dff g4369_reg ( clk, reset, ex_wire80, n822 );
not U_inv496 ( n19571, ex_wire80 );
dff g4581_reg ( clk, reset, n10636, n837 );
not U_inv497 ( n19125, n10636 );
dff g4340_reg ( clk, reset, n10302, n1149 );
not U_inv498 ( n19587, n10302 );
dff g4349_reg ( clk, reset, n10223, n1154 );
not U_inv499 ( n19588, n10223 );
dff g4358_reg ( clk, reset, n10292, n1159 );
not U_inv500 ( n19589, n10292 );
dff g4311_reg ( clk, reset, n10346, n1174 );
not U_inv501 ( n19590, n10346 );
dff g4322_reg ( clk, reset, n10227, n1179 );
not U_inv502 ( n19591, n10227 );
dff g4332_reg ( clk, reset, n10351, n1184 );
not U_inv503 ( n19592, n10351 );
dff g4864_reg ( clk, reset, n10812, n1229 );
not U_inv504 ( n19598, n10812 );
dff g4871_reg ( clk, reset, n10289, n1234 );
not U_inv505 ( n19599, n10289 );
dff g4878_reg ( clk, reset, n10460, n1239 );
not U_inv506 ( n19600, n10460 );
dff g4843_reg ( clk, reset, n10287, n1244 );
not U_inv507 ( n19601, n10287 );
dff g4849_reg ( clk, reset, n10610, n1249 );
not U_inv508 ( n19602, n10610 );
dff g4854_reg ( clk, reset, n10920, n1254 );
not U_inv509 ( n19603, n10920 );
dff g4859_reg ( clk, reset, n10767, n1259 );
not U_inv510 ( n19500, n10767 );
dff g4991_reg ( clk, reset, n10451, n1331 );
not U_inv511 ( n19605, n10451 );
dff g4966_reg ( clk, reset, n10308, n1336 );
not U_inv512 ( n19606, n10308 );
dff g4975_reg ( clk, reset, n10407, n1341 );
not U_inv513 ( n19607, n10407 );
dff g4899_reg ( clk, reset, n10443, n1346 );
not U_inv514 ( n19608, n10443 );
dff g4983_reg ( clk, reset, n10391, n1326 );
not U_inv515 ( n19457, n10391 );
dff g63_reg ( clk, reset, ex_wire81, new_g34783_ );
not U_inv516 ( n19499, ex_wire81 );
dff g4674_reg ( clk, reset, n10811, n1396 );
not U_inv517 ( n19613, n10811 );
dff g4681_reg ( clk, reset, n10290, n1401 );
not U_inv518 ( n19614, n10290 );
dff g4688_reg ( clk, reset, n10459, n1406 );
not U_inv519 ( n19615, n10459 );
dff g4653_reg ( clk, reset, n10288, n1411 );
not U_inv520 ( n19616, n10288 );
dff g4659_reg ( clk, reset, n10609, n1416 );
not U_inv521 ( n19617, n10609 );
dff g4664_reg ( clk, reset, n10919, n1421 );
not U_inv522 ( n19618, n10919 );
dff g4669_reg ( clk, reset, n10768, n1426 );
not U_inv523 ( n19447, n10768 );
dff g4801_reg ( clk, reset, n10450, n1498 );
not U_inv524 ( n19620, n10450 );
dff g4776_reg ( clk, reset, n10309, n1503 );
not U_inv525 ( n19621, n10309 );
dff g4785_reg ( clk, reset, n10406, n1508 );
not U_inv526 ( n19622, n10406 );
dff g4709_reg ( clk, reset, n10444, n1513 );
not U_inv527 ( n19623, n10444 );
dff g4793_reg ( clk, reset, n10392, n1493 );
not U_inv528 ( n19445, n10392 );
dff g4646_reg ( clk, reset, ex_wire82, n1391 );
not U_inv529 ( n19612, ex_wire82 );
dff g4836_reg ( clk, reset, ex_wire83, n1224 );
not U_inv530 ( n19597, ex_wire83 );
dff g4584_reg ( clk, reset, n10585, n1189 );
not U_inv531 ( n19593, n10585 );
dff g4593_reg ( clk, reset, n10584, n1194 );
not U_inv532 ( n19594, n10584 );
dff g4601_reg ( clk, reset, n10334, n1199 );
not U_inv533 ( n19504, n10334 );
dff g4608_reg ( clk, reset, n10430, n1204 );
not U_inv534 ( n19595, n10430 );
dff g4616_reg ( clk, reset, n10478, n1209 );
not U_inv535 ( n19596, n10478 );
dff g4366_reg ( clk, reset, n10895, n1214 );
dff g66_reg ( clk, reset, g29218, n1164 );
dff g65_reg ( clk, reset, g65, g29218 );
dff g4531_reg ( clk, reset, g4531, n1169 );
dff g4888_reg ( clk, reset, ex_wire84, n1356 );
not U_inv536 ( n19456, ex_wire84 );
dff g71_reg ( clk, reset, ex_wire85, new_g34649_ );
not U_inv537 ( n19450, ex_wire85 );
dff g4933_reg ( clk, reset, ex_wire86, n1366 );
not U_inv538 ( n19609, ex_wire86 );
dff g3352_reg ( clk, reset, n10243, n3409 );
not U_inv539 ( n19829, n10243 );
dff g3288_reg ( clk, reset, n10472, n3414 );
not U_inv540 ( n19830, n10472 );
dff g93_reg ( clk, reset, ex_wire87, new_g34809_ );
not U_inv541 ( n19430, ex_wire87 );
dff g4054_reg ( clk, reset, n10263, n4127 );
not U_inv542 ( n19902, n10263 );
dff g4961_reg ( clk, reset, n10554, n1381 );
dff g4955_reg ( clk, reset, ex_wire88, n1386 );
not U_inv543 ( n19611, ex_wire88 );
dff g3990_reg ( clk, reset, n10614, n4132 );
not U_inv544 ( n19448, n10614 );
dff g3703_reg ( clk, reset, n10264, n3768 );
not U_inv545 ( n19866, n10264 );
dff g4950_reg ( clk, reset, n10555, n1371 );
dff g4944_reg ( clk, reset, ex_wire89, n1376 );
not U_inv546 ( n19610, ex_wire89 );
dff g3639_reg ( clk, reset, n10615, n3773 );
not U_inv547 ( n19449, n10615 );
dff g6741_reg ( clk, reset, n10265, n3050 );
not U_inv548 ( n19792, n10265 );
dff g6682_reg ( clk, reset, n10616, n3055 );
not U_inv549 ( n19452, n10616 );
dff g4894_reg ( clk, reset, n10557, n1351 );
dff g5357_reg ( clk, reset, n10270, n1614 );
not U_inv550 ( n19632, n10270 );
dff g4704_reg ( clk, reset, n10553, n1518 );
dff g4698_reg ( clk, reset, ex_wire90, n1523 );
not U_inv551 ( n19444, ex_wire90 );
dff g5297_reg ( clk, reset, n10604, n1619 );
not U_inv552 ( n19441, n10604 );
dff g101_reg ( clk, reset, ex_wire91, new_g34657_ );
not U_inv553 ( n19439, ex_wire91 );
dff g4765_reg ( clk, reset, ex_wire92, n1553 );
not U_inv554 ( n19626, ex_wire92 );
dff g6395_reg ( clk, reset, n10261, n2691 );
not U_inv555 ( n19756, n10261 );
dff g6336_reg ( clk, reset, n10612, n2696 );
not U_inv556 ( n19436, n10612 );
dff g4771_reg ( clk, reset, n10550, n1548 );
dff g4754_reg ( clk, reset, ex_wire93, n1543 );
not U_inv557 ( n19625, ex_wire93 );
dff g6049_reg ( clk, reset, n10262, n2332 );
not U_inv558 ( n19719, n10262 );
dff g5990_reg ( clk, reset, n10613, n2337 );
not U_inv559 ( n19437, n10613 );
dff g4760_reg ( clk, reset, n10551, n1538 );
dff g4743_reg ( clk, reset, ex_wire94, n1533 );
not U_inv560 ( n19624, ex_wire94 );
dff g5703_reg ( clk, reset, n10242, n1973 );
not U_inv561 ( n19683, n10242 );
dff g5644_reg ( clk, reset, n10471, n1978 );
not U_inv562 ( n19438, n10471 );
dff g4749_reg ( clk, reset, n10552, n1528 );
dff g3106_reg ( clk, reset, n10486, n3667 );
not U_inv563 ( n19857, n10486 );
dff g3115_reg ( clk, reset, ex_wire95, n3672 );
not U_inv564 ( n19518, ex_wire95 );
dff g3119_reg ( clk, reset, n10566, n3677 );
not U_inv565 ( n19369, n10566 );
dff g3125_reg ( clk, reset, n10728, n3682 );
not U_inv566 ( n19368, n10728 );
dff g3129_reg ( clk, reset, n10778, n3687 );
not U_inv567 ( n19536, n10778 );
dff g3133_reg ( clk, reset, ex_wire96, n3692 );
not U_inv568 ( n19858, ex_wire96 );
dff g3139_reg ( clk, reset, n10727, n3697 );
not U_inv569 ( n19859, n10727 );
dff g3143_reg ( clk, reset, ex_wire97, n3702 );
not U_inv570 ( n19537, ex_wire97 );
dff g2898_reg ( clk, reset, n10771, n7518 );
not U_inv571 ( n19469, n10771 );
dff g2882_reg ( clk, reset, ex_wire98, n7523 );
not U_inv572 ( n20220, ex_wire98 );
dff g2878_reg ( clk, reset, ex_wire99, n7528 );
not U_inv573 ( n19338, ex_wire99 );
dff g50_reg ( clk, reset, ex_wire100, new_g34978_ );
not U_inv574 ( n19340, ex_wire100 );
dff g19_reg ( clk, reset, ex_wire101, new_g34978_ );
not U_inv575 ( n20235, ex_wire101 );
dff g1296_reg ( clk, reset, ex_wire102, n5837 );
not U_inv576 ( n20051, ex_wire102 );
dff g1283_reg ( clk, reset, n10785, n5842 );
not U_inv577 ( n19333, n10785 );
dff g51_reg ( clk, reset, ex_wire103, new_g34979_ );
not U_inv578 ( n19334, ex_wire103 );
dff g28_reg ( clk, reset, n10310, new_g34979_ );
not U_inv579 ( n20236, n10310 );
dff g136_reg ( clk, reset, g21292, n5428 );
not U_inv580 ( g30329, g21292 );
dff g199_reg ( clk, reset, ex_wire104, n5433 );
not U_inv581 ( n19319, ex_wire104 );
dff g52_reg ( clk, reset, ex_wire105, new_g34971_ );
not U_inv582 ( n19325, ex_wire105 );
dff g31_reg ( clk, reset, n10602, new_g34971_ );
not U_inv583 ( n20237, n10602 );
dff g2984_reg ( clk, reset, n10769, n7543 );
not U_inv584 ( n19322, n10769 );
dff g2907_reg ( clk, reset, n10508, n7548 );
not U_inv585 ( n20221, n10508 );
dff g2912_reg ( clk, reset, n10509, n7553 );
not U_inv586 ( n20222, n10509 );
dff g2922_reg ( clk, reset, n10674, n7558 );
not U_inv587 ( n20223, n10674 );
dff g2936_reg ( clk, reset, n10673, n7563 );
not U_inv588 ( n20224, n10673 );
dff g2950_reg ( clk, reset, n10562, n7568 );
not U_inv589 ( n20225, n10562 );
dff g2960_reg ( clk, reset, n10672, n7573 );
not U_inv590 ( n20226, n10672 );
dff g2970_reg ( clk, reset, n10671, n7578 );
not U_inv591 ( n20227, n10671 );
dff g2902_reg ( clk, reset, n10700, n7583 );
not U_inv592 ( n20228, n10700 );
dff g2917_reg ( clk, reset, n10665, n7588 );
not U_inv593 ( n20229, n10665 );
dff g46_reg ( clk, reset, g46, new_g34974_ );
dff g7_reg ( clk, reset, ex_wire106, new_g34974_ );
not U_inv594 ( n19496, ex_wire106 );
dff g34_reg ( clk, reset, n10939, n51 );
not U_inv595 ( n19493, n10939 );
dff g45_reg ( clk, reset, g45, new_g34970_ );
dff g6_reg ( clk, reset, ex_wire107, new_g34970_ );
not U_inv596 ( n19495, ex_wire107 );
dff g4172_reg ( clk, reset, n10832, n4555 );
not U_inv597 ( n19458, n10832 );
dff g4176_reg ( clk, reset, n10775, n4560 );
not U_inv598 ( n19339, n10775 );
dff g4146_reg ( clk, reset, n10385, n4565 );
not U_inv599 ( n19945, n10385 );
dff g4157_reg ( clk, reset, n10547, n4570 );
not U_inv600 ( n19946, n10547 );
dff g4145_reg ( clk, reset, n10905, n4500 );
not U_inv601 ( n19941, n10905 );
dff g4112_reg ( clk, reset, ex_wire108, n4505 );
not U_inv602 ( n19344, ex_wire108 );
dff g4116_reg ( clk, reset, ex_wire109, n4510 );
not U_inv603 ( n19942, ex_wire109 );
dff g4119_reg ( clk, reset, ex_wire110, n4515 );
not U_inv604 ( n19943, ex_wire110 );
dff g4122_reg ( clk, reset, n10872, n4520 );
dff g4153_reg ( clk, reset, n10291, n4525 );
not U_inv605 ( n19341, n10291 );
dff g4164_reg ( clk, reset, ex_wire111, n4530 );
not U_inv606 ( n19944, ex_wire111 );
dff g4185_reg ( clk, reset, g11770, n4694 );
not U_inv607 ( n19301, g11770 );
dff g4213_reg ( clk, reset, g8915, g11770 );
not U_inv608 ( n19302, g8915 );
dff g4216_reg ( clk, reset, g8916, g8915 );
not U_inv609 ( n19303, g8916 );
dff g4219_reg ( clk, reset, g8917, g8916 );
not U_inv610 ( n19299, g8917 );
dff g4222_reg ( clk, reset, g8870, g8917 );
not U_inv611 ( n19952, g8870 );
dff g4226_reg ( clk, reset, g8918, g8870 );
not U_inv612 ( n19300, g8918 );
dff g4229_reg ( clk, reset, g8919, g8918 );
dff g4232_reg ( clk, reset, g8920, g8919 );
not U_inv613 ( n19298, g8920 );
dff g4235_reg ( clk, reset, n10774, g8920 );
not U_inv614 ( n19953, n10774 );
dff g4242_reg ( clk, reset, ex_wire112, n4731 );
not U_inv615 ( n19315, ex_wire112 );
dff g4300_reg ( clk, reset, n10787, n4609 );
not U_inv616 ( n19460, n10787 );
dff g4253_reg ( clk, reset, n10366, n4614 );
not U_inv617 ( n19949, n10366 );
dff g4249_reg ( clk, reset, n10546, n4619 );
dff g4245_reg ( clk, reset, n10545, n4624 );
dff g4277_reg ( clk, reset, g8839, n4629 );
not U_inv618 ( n19313, g8839 );
dff g4281_reg ( clk, reset, ex_wire113, g8839 );
not U_inv619 ( n19314, ex_wire113 );
dff g4284_reg ( clk, reset, ex_wire114, n4638 );
not U_inv620 ( n19424, ex_wire114 );
dff g4287_reg ( clk, reset, g9019, n4643 );
not U_inv621 ( n19311, g9019 );
dff g4291_reg ( clk, reset, ex_wire115, g9019 );
not U_inv622 ( n19312, ex_wire115 );
dff g2946_reg ( clk, reset, ex_wire116, n4652 );
not U_inv623 ( n19310, ex_wire116 );
dff g4191_reg ( clk, reset, g11447, n4657 );
not U_inv624 ( n19307, g11447 );
dff g4188_reg ( clk, reset, g8783, g11447 );
not U_inv625 ( n19308, g8783 );
dff g4194_reg ( clk, reset, g8784, g8783 );
not U_inv626 ( n19309, g8784 );
dff g4197_reg ( clk, reset, g8785, g8784 );
not U_inv627 ( n19305, g8785 );
dff g4200_reg ( clk, reset, g8786, g8785 );
not U_inv628 ( n19950, g8786 );
dff g4204_reg ( clk, reset, g8787, g8786 );
not U_inv629 ( n19306, g8787 );
dff g4207_reg ( clk, reset, g8788, g8787 );
dff g4210_reg ( clk, reset, g8789, g8788 );
not U_inv630 ( n19304, g8789 );
dff g4180_reg ( clk, reset, n10457, g8789 );
not U_inv631 ( n19951, n10457 );
dff g3889_reg ( clk, reset, ex_wire117, n4270 );
not U_inv632 ( n19909, ex_wire117 );
dff g3538_reg ( clk, reset, ex_wire118, n3911 );
not U_inv633 ( n19873, ex_wire118 );
dff g3187_reg ( clk, reset, ex_wire119, n3552 );
not U_inv634 ( n19837, ex_wire119 );
dff g6581_reg ( clk, reset, ex_wire120, n3193 );
not U_inv635 ( n19799, ex_wire120 );
dff g6235_reg ( clk, reset, ex_wire121, n2834 );
not U_inv636 ( n19763, ex_wire121 );
dff g5889_reg ( clk, reset, ex_wire122, n2475 );
not U_inv637 ( n19726, ex_wire122 );
dff g5543_reg ( clk, reset, ex_wire123, n2116 );
not U_inv638 ( n19690, ex_wire123 );
dff g5196_reg ( clk, reset, ex_wire124, n1757 );
not U_inv639 ( n19655, ex_wire124 );
dff g3849_reg ( clk, reset, n10837, n4375 );
not U_inv640 ( n19350, n10837 );
dff g3813_reg ( clk, reset, n10373, n4380 );
dff g3917_reg ( clk, reset, ex_wire125, n4275 );
not U_inv641 ( n19910, ex_wire125 );
dff g3933_reg ( clk, reset, ex_wire126, n4280 );
not U_inv642 ( n19911, ex_wire126 );
dff g3949_reg ( clk, reset, ex_wire127, n4285 );
not U_inv643 ( n19912, ex_wire127 );
dff g3897_reg ( clk, reset, ex_wire128, n4290 );
not U_inv644 ( n19913, ex_wire128 );
dff g3893_reg ( clk, reset, n10796, n4295 );
not U_inv645 ( n19914, n10796 );
dff g3921_reg ( clk, reset, n10840, n4300 );
not U_inv646 ( n19915, n10840 );
dff g3937_reg ( clk, reset, ex_wire129, n4305 );
not U_inv647 ( n19916, ex_wire129 );
dff g3953_reg ( clk, reset, n10839, n4310 );
not U_inv648 ( n19917, n10839 );
dff g3905_reg ( clk, reset, ex_wire130, n4315 );
not U_inv649 ( n19918, ex_wire130 );
dff g3901_reg ( clk, reset, ex_wire131, n4320 );
not U_inv650 ( n19919, ex_wire131 );
dff g3925_reg ( clk, reset, ex_wire132, n4325 );
not U_inv651 ( n19920, ex_wire132 );
dff g3941_reg ( clk, reset, ex_wire133, n4330 );
not U_inv652 ( n19921, ex_wire133 );
dff g3957_reg ( clk, reset, ex_wire134, n4335 );
not U_inv653 ( n19922, ex_wire134 );
dff g3913_reg ( clk, reset, ex_wire135, n4340 );
not U_inv654 ( n19923, ex_wire135 );
dff g3909_reg ( clk, reset, n10795, n4345 );
not U_inv655 ( n19924, n10795 );
dff g3929_reg ( clk, reset, n10838, n4350 );
not U_inv656 ( n19925, n10838 );
dff g3945_reg ( clk, reset, ex_wire136, n4355 );
not U_inv657 ( n19926, ex_wire136 );
dff g3961_reg ( clk, reset, n10760, n4360 );
not U_inv658 ( n19927, n10760 );
dff g3965_reg ( clk, reset, ex_wire137, n4365 );
not U_inv659 ( n19928, ex_wire137 );
dff g3808_reg ( clk, reset, n10484, n4385 );
not U_inv660 ( n19929, n10484 );
dff g3817_reg ( clk, reset, n10698, n4390 );
not U_inv661 ( n19520, n10698 );
dff g3821_reg ( clk, reset, n10564, n4395 );
not U_inv662 ( n19349, n10564 );
dff g3827_reg ( clk, reset, n10724, n4400 );
not U_inv663 ( n19348, n10724 );
dff g3831_reg ( clk, reset, n10776, n4405 );
not U_inv664 ( n19524, n10776 );
dff g3835_reg ( clk, reset, ex_wire138, n4410 );
not U_inv665 ( n19930, ex_wire138 );
dff g3841_reg ( clk, reset, n10723, n4415 );
not U_inv666 ( n19931, n10723 );
dff g3845_reg ( clk, reset, ex_wire139, n4420 );
not U_inv667 ( n19525, ex_wire139 );
dff g4035_reg ( clk, reset, n10928, n4370 );
not U_inv668 ( n19455, n10928 );
dff g3498_reg ( clk, reset, n10841, n4016 );
not U_inv669 ( n19360, n10841 );
dff g3462_reg ( clk, reset, n10374, n4021 );
dff g3566_reg ( clk, reset, ex_wire140, n3916 );
not U_inv670 ( n19874, ex_wire140 );
dff g3582_reg ( clk, reset, ex_wire141, n3921 );
not U_inv671 ( n19875, ex_wire141 );
dff g3598_reg ( clk, reset, ex_wire142, n3926 );
not U_inv672 ( n19876, ex_wire142 );
dff g3546_reg ( clk, reset, ex_wire143, n3931 );
not U_inv673 ( n19877, ex_wire143 );
dff g3542_reg ( clk, reset, n10798, n3936 );
not U_inv674 ( n19878, n10798 );
dff g3570_reg ( clk, reset, n10844, n3941 );
not U_inv675 ( n19879, n10844 );
dff g3586_reg ( clk, reset, ex_wire144, n3946 );
not U_inv676 ( n19880, ex_wire144 );
dff g3602_reg ( clk, reset, n10843, n3951 );
not U_inv677 ( n19881, n10843 );
dff g3554_reg ( clk, reset, ex_wire145, n3956 );
not U_inv678 ( n19882, ex_wire145 );
dff g3550_reg ( clk, reset, ex_wire146, n3961 );
not U_inv679 ( n19883, ex_wire146 );
dff g3574_reg ( clk, reset, ex_wire147, n3966 );
not U_inv680 ( n19884, ex_wire147 );
dff g3590_reg ( clk, reset, ex_wire148, n3971 );
not U_inv681 ( n19885, ex_wire148 );
dff g3606_reg ( clk, reset, ex_wire149, n3976 );
not U_inv682 ( n19886, ex_wire149 );
dff g3562_reg ( clk, reset, ex_wire150, n3981 );
not U_inv683 ( n19887, ex_wire150 );
dff g3558_reg ( clk, reset, n10797, n3986 );
not U_inv684 ( n19888, n10797 );
dff g3578_reg ( clk, reset, n10842, n3991 );
not U_inv685 ( n19889, n10842 );
dff g3594_reg ( clk, reset, ex_wire151, n3996 );
not U_inv686 ( n19890, ex_wire151 );
dff g3610_reg ( clk, reset, n10761, n4001 );
not U_inv687 ( n19891, n10761 );
dff g3614_reg ( clk, reset, ex_wire152, n4006 );
not U_inv688 ( n19892, ex_wire152 );
dff g3457_reg ( clk, reset, n10485, n4026 );
not U_inv689 ( n19893, n10485 );
dff g3466_reg ( clk, reset, n10640, n4031 );
not U_inv690 ( n19519, n10640 );
dff g3470_reg ( clk, reset, n10565, n4036 );
not U_inv691 ( n19359, n10565 );
dff g3476_reg ( clk, reset, n10726, n4041 );
not U_inv692 ( n19358, n10726 );
dff g3480_reg ( clk, reset, n10777, n4046 );
not U_inv693 ( n19534, n10777 );
dff g3484_reg ( clk, reset, ex_wire153, n4051 );
not U_inv694 ( n19894, ex_wire153 );
dff g3490_reg ( clk, reset, n10725, n4056 );
not U_inv695 ( n19895, n10725 );
dff g3494_reg ( clk, reset, ex_wire154, n4061 );
not U_inv696 ( n19535, ex_wire154 );
dff g3684_reg ( clk, reset, n10938, n4011 );
not U_inv697 ( n19454, n10938 );
dff g3147_reg ( clk, reset, n10845, n3657 );
not U_inv698 ( n19370, n10845 );
dff g3111_reg ( clk, reset, n10375, n3662 );
dff g3215_reg ( clk, reset, ex_wire155, n3557 );
not U_inv699 ( n19838, ex_wire155 );
dff g3231_reg ( clk, reset, ex_wire156, n3562 );
not U_inv700 ( n19839, ex_wire156 );
dff g3247_reg ( clk, reset, ex_wire157, n3567 );
not U_inv701 ( n19840, ex_wire157 );
dff g3195_reg ( clk, reset, ex_wire158, n3572 );
not U_inv702 ( n19841, ex_wire158 );
dff g3191_reg ( clk, reset, n10800, n3577 );
not U_inv703 ( n19842, n10800 );
dff g3219_reg ( clk, reset, n10848, n3582 );
not U_inv704 ( n19843, n10848 );
dff g3235_reg ( clk, reset, ex_wire159, n3587 );
not U_inv705 ( n19844, ex_wire159 );
dff g3251_reg ( clk, reset, n10847, n3592 );
not U_inv706 ( n19845, n10847 );
dff g3203_reg ( clk, reset, ex_wire160, n3597 );
not U_inv707 ( n19846, ex_wire160 );
dff g3199_reg ( clk, reset, ex_wire161, n3602 );
not U_inv708 ( n19847, ex_wire161 );
dff g3223_reg ( clk, reset, ex_wire162, n3607 );
not U_inv709 ( n19848, ex_wire162 );
dff g3239_reg ( clk, reset, ex_wire163, n3612 );
not U_inv710 ( n19849, ex_wire163 );
dff g3255_reg ( clk, reset, ex_wire164, n3617 );
not U_inv711 ( n19850, ex_wire164 );
dff g3211_reg ( clk, reset, ex_wire165, n3622 );
not U_inv712 ( n19851, ex_wire165 );
dff g3207_reg ( clk, reset, n10799, n3627 );
not U_inv713 ( n19852, n10799 );
dff g3227_reg ( clk, reset, n10846, n3632 );
not U_inv714 ( n19853, n10846 );
dff g3243_reg ( clk, reset, ex_wire166, n3637 );
not U_inv715 ( n19854, ex_wire166 );
dff g3259_reg ( clk, reset, n10762, n3642 );
not U_inv716 ( n19855, n10762 );
dff g3263_reg ( clk, reset, ex_wire167, n3647 );
not U_inv717 ( n19856, ex_wire167 );
dff g3333_reg ( clk, reset, n10894, n3652 );
dff g6541_reg ( clk, reset, n10849, n3298 );
not U_inv718 ( n19380, n10849 );
dff g6505_reg ( clk, reset, n10376, n3303 );
dff g6609_reg ( clk, reset, ex_wire168, n3198 );
not U_inv719 ( n19800, ex_wire168 );
dff g6625_reg ( clk, reset, ex_wire169, n3203 );
not U_inv720 ( n19801, ex_wire169 );
dff g6641_reg ( clk, reset, ex_wire170, n3208 );
not U_inv721 ( n19802, ex_wire170 );
dff g6589_reg ( clk, reset, ex_wire171, n3213 );
not U_inv722 ( n19803, ex_wire171 );
dff g6585_reg ( clk, reset, n10802, n3218 );
not U_inv723 ( n19804, n10802 );
dff g6613_reg ( clk, reset, n10852, n3223 );
not U_inv724 ( n19805, n10852 );
dff g6629_reg ( clk, reset, ex_wire172, n3228 );
not U_inv725 ( n19806, ex_wire172 );
dff g6645_reg ( clk, reset, n10851, n3233 );
not U_inv726 ( n19807, n10851 );
dff g6597_reg ( clk, reset, ex_wire173, n3238 );
not U_inv727 ( n19808, ex_wire173 );
dff g6593_reg ( clk, reset, ex_wire174, n3243 );
not U_inv728 ( n19809, ex_wire174 );
dff g6617_reg ( clk, reset, ex_wire175, n3248 );
not U_inv729 ( n19810, ex_wire175 );
dff g6633_reg ( clk, reset, ex_wire176, n3253 );
not U_inv730 ( n19811, ex_wire176 );
dff g6649_reg ( clk, reset, ex_wire177, n3258 );
not U_inv731 ( n19812, ex_wire177 );
dff g6605_reg ( clk, reset, ex_wire178, n3263 );
not U_inv732 ( n19813, ex_wire178 );
dff g6601_reg ( clk, reset, n10801, n3268 );
not U_inv733 ( n19814, n10801 );
dff g6621_reg ( clk, reset, n10850, n3273 );
not U_inv734 ( n19815, n10850 );
dff g6637_reg ( clk, reset, ex_wire179, n3278 );
not U_inv735 ( n19816, ex_wire179 );
dff g6653_reg ( clk, reset, n10763, n3283 );
not U_inv736 ( n19817, n10763 );
dff g6657_reg ( clk, reset, ex_wire180, n3288 );
not U_inv737 ( n19818, ex_wire180 );
dff g6500_reg ( clk, reset, n10487, n3308 );
not U_inv738 ( n19820, n10487 );
dff g6509_reg ( clk, reset, ex_wire181, n3313 );
not U_inv739 ( n19521, ex_wire181 );
dff g6513_reg ( clk, reset, n10567, n3318 );
not U_inv740 ( n19379, n10567 );
dff g6519_reg ( clk, reset, n10730, n3323 );
not U_inv741 ( n19378, n10730 );
dff g6523_reg ( clk, reset, n10779, n3328 );
not U_inv742 ( n19532, n10779 );
dff g6527_reg ( clk, reset, ex_wire182, n3333 );
not U_inv743 ( n19821, ex_wire182 );
dff g6533_reg ( clk, reset, n10729, n3338 );
not U_inv744 ( n19822, n10729 );
dff g6537_reg ( clk, reset, ex_wire183, n3343 );
not U_inv745 ( n19533, ex_wire183 );
dff g5011_reg ( clk, reset, n10924, n3293 );
not U_inv746 ( n19819, n10924 );
dff g6195_reg ( clk, reset, n10853, n2939 );
not U_inv747 ( n19390, n10853 );
dff g6159_reg ( clk, reset, n10377, n2944 );
dff g6263_reg ( clk, reset, ex_wire184, n2839 );
not U_inv748 ( n19764, ex_wire184 );
dff g6279_reg ( clk, reset, ex_wire185, n2844 );
not U_inv749 ( n19765, ex_wire185 );
dff g6295_reg ( clk, reset, ex_wire186, n2849 );
not U_inv750 ( n19766, ex_wire186 );
dff g6243_reg ( clk, reset, ex_wire187, n2854 );
not U_inv751 ( n19767, ex_wire187 );
dff g6239_reg ( clk, reset, n10804, n2859 );
not U_inv752 ( n19768, n10804 );
dff g6267_reg ( clk, reset, n10856, n2864 );
not U_inv753 ( n19769, n10856 );
dff g6283_reg ( clk, reset, ex_wire188, n2869 );
not U_inv754 ( n19770, ex_wire188 );
dff g6299_reg ( clk, reset, n10855, n2874 );
not U_inv755 ( n19771, n10855 );
dff g6251_reg ( clk, reset, ex_wire189, n2879 );
not U_inv756 ( n19772, ex_wire189 );
dff g6247_reg ( clk, reset, ex_wire190, n2884 );
not U_inv757 ( n19773, ex_wire190 );
dff g6271_reg ( clk, reset, ex_wire191, n2889 );
not U_inv758 ( n19774, ex_wire191 );
dff g6287_reg ( clk, reset, ex_wire192, n2894 );
not U_inv759 ( n19775, ex_wire192 );
dff g6303_reg ( clk, reset, ex_wire193, n2899 );
not U_inv760 ( n19776, ex_wire193 );
dff g6259_reg ( clk, reset, ex_wire194, n2904 );
not U_inv761 ( n19777, ex_wire194 );
dff g6255_reg ( clk, reset, n10803, n2909 );
not U_inv762 ( n19778, n10803 );
dff g6275_reg ( clk, reset, n10854, n2914 );
not U_inv763 ( n19779, n10854 );
dff g6291_reg ( clk, reset, ex_wire195, n2919 );
not U_inv764 ( n19780, ex_wire195 );
dff g6307_reg ( clk, reset, n10764, n2924 );
not U_inv765 ( n19781, n10764 );
dff g6311_reg ( clk, reset, ex_wire196, n2929 );
not U_inv766 ( n19782, ex_wire196 );
dff g6154_reg ( clk, reset, n10488, n2949 );
not U_inv767 ( n19783, n10488 );
dff g6163_reg ( clk, reset, ex_wire197, n2954 );
not U_inv768 ( n19522, ex_wire197 );
dff g6167_reg ( clk, reset, n10568, n2959 );
not U_inv769 ( n19389, n10568 );
dff g6173_reg ( clk, reset, n10732, n2964 );
not U_inv770 ( n19388, n10732 );
dff g6177_reg ( clk, reset, n10279, n2969 );
dff g6181_reg ( clk, reset, ex_wire198, n2974 );
not U_inv771 ( n19784, ex_wire198 );
dff g6187_reg ( clk, reset, n10731, n2979 );
not U_inv772 ( n19785, n10731 );
dff g6191_reg ( clk, reset, n10896, n2984 );
dff g4826_reg ( clk, reset, n10929, n2934 );
not U_inv773 ( n19446, n10929 );
dff g5849_reg ( clk, reset, n10857, n2580 );
not U_inv774 ( n19400, n10857 );
dff g5813_reg ( clk, reset, n10378, n2585 );
dff g5917_reg ( clk, reset, ex_wire199, n2480 );
not U_inv775 ( n19727, ex_wire199 );
dff g5933_reg ( clk, reset, ex_wire200, n2485 );
not U_inv776 ( n19728, ex_wire200 );
dff g5949_reg ( clk, reset, ex_wire201, n2490 );
not U_inv777 ( n19729, ex_wire201 );
dff g5897_reg ( clk, reset, ex_wire202, n2495 );
not U_inv778 ( n19730, ex_wire202 );
dff g5893_reg ( clk, reset, n10806, n2500 );
not U_inv779 ( n19731, n10806 );
dff g5921_reg ( clk, reset, n10860, n2505 );
not U_inv780 ( n19732, n10860 );
dff g5937_reg ( clk, reset, ex_wire203, n2510 );
not U_inv781 ( n19733, ex_wire203 );
dff g5953_reg ( clk, reset, n10859, n2515 );
not U_inv782 ( n19734, n10859 );
dff g5905_reg ( clk, reset, ex_wire204, n2520 );
not U_inv783 ( n19735, ex_wire204 );
dff g5901_reg ( clk, reset, ex_wire205, n2525 );
not U_inv784 ( n19736, ex_wire205 );
dff g5925_reg ( clk, reset, ex_wire206, n2530 );
not U_inv785 ( n19737, ex_wire206 );
dff g5941_reg ( clk, reset, ex_wire207, n2535 );
not U_inv786 ( n19738, ex_wire207 );
dff g5957_reg ( clk, reset, ex_wire208, n2540 );
not U_inv787 ( n19739, ex_wire208 );
dff g5913_reg ( clk, reset, ex_wire209, n2545 );
not U_inv788 ( n19740, ex_wire209 );
dff g5909_reg ( clk, reset, n10805, n2550 );
not U_inv789 ( n19741, n10805 );
dff g5929_reg ( clk, reset, n10858, n2555 );
not U_inv790 ( n19742, n10858 );
dff g5945_reg ( clk, reset, ex_wire210, n2560 );
not U_inv791 ( n19743, ex_wire210 );
dff g5961_reg ( clk, reset, n10765, n2565 );
not U_inv792 ( n19744, n10765 );
dff g5965_reg ( clk, reset, ex_wire211, n2570 );
not U_inv793 ( n19745, ex_wire211 );
dff g5808_reg ( clk, reset, n10489, n2590 );
not U_inv794 ( n19747, n10489 );
dff g5817_reg ( clk, reset, ex_wire212, n2595 );
not U_inv795 ( n19516, ex_wire212 );
dff g5821_reg ( clk, reset, n10569, n2600 );
not U_inv796 ( n19399, n10569 );
dff g5827_reg ( clk, reset, n10734, n2605 );
not U_inv797 ( n19398, n10734 );
dff g5831_reg ( clk, reset, n10282, n2610 );
not U_inv798 ( n19530, n10282 );
dff g5835_reg ( clk, reset, ex_wire213, n2615 );
not U_inv799 ( n19748, ex_wire213 );
dff g5841_reg ( clk, reset, n10733, n2620 );
not U_inv800 ( n19749, n10733 );
dff g5845_reg ( clk, reset, n10759, n2625 );
not U_inv801 ( n19531, n10759 );
dff g4831_reg ( clk, reset, n10925, n2575 );
not U_inv802 ( n19746, n10925 );
dff g5503_reg ( clk, reset, n10861, n2221 );
not U_inv803 ( n19410, n10861 );
dff g5467_reg ( clk, reset, n10379, n2226 );
dff g5571_reg ( clk, reset, ex_wire214, n2121 );
not U_inv804 ( n19691, ex_wire214 );
dff g5587_reg ( clk, reset, ex_wire215, n2126 );
not U_inv805 ( n19692, ex_wire215 );
dff g5603_reg ( clk, reset, ex_wire216, n2131 );
not U_inv806 ( n19693, ex_wire216 );
dff g5551_reg ( clk, reset, ex_wire217, n2136 );
not U_inv807 ( n19694, ex_wire217 );
dff g5547_reg ( clk, reset, n10808, n2141 );
not U_inv808 ( n19695, n10808 );
dff g5575_reg ( clk, reset, n10864, n2146 );
not U_inv809 ( n19696, n10864 );
dff g5591_reg ( clk, reset, ex_wire218, n2151 );
not U_inv810 ( n19697, ex_wire218 );
dff g5607_reg ( clk, reset, n10863, n2156 );
not U_inv811 ( n19698, n10863 );
dff g5559_reg ( clk, reset, ex_wire219, n2161 );
not U_inv812 ( n19699, ex_wire219 );
dff g5555_reg ( clk, reset, ex_wire220, n2166 );
not U_inv813 ( n19700, ex_wire220 );
dff g5579_reg ( clk, reset, ex_wire221, n2171 );
not U_inv814 ( n19701, ex_wire221 );
dff g5595_reg ( clk, reset, ex_wire222, n2176 );
not U_inv815 ( n19702, ex_wire222 );
dff g5611_reg ( clk, reset, ex_wire223, n2181 );
not U_inv816 ( n19703, ex_wire223 );
dff g5567_reg ( clk, reset, ex_wire224, n2186 );
not U_inv817 ( n19704, ex_wire224 );
dff g5563_reg ( clk, reset, n10807, n2191 );
not U_inv818 ( n19705, n10807 );
dff g5583_reg ( clk, reset, n10862, n2196 );
not U_inv819 ( n19706, n10862 );
dff g5599_reg ( clk, reset, ex_wire225, n2201 );
not U_inv820 ( n19707, ex_wire225 );
dff g5615_reg ( clk, reset, n10766, n2206 );
not U_inv821 ( n19708, n10766 );
dff g5619_reg ( clk, reset, ex_wire226, n2211 );
not U_inv822 ( n19709, ex_wire226 );
dff g5462_reg ( clk, reset, n10490, n2231 );
not U_inv823 ( n19710, n10490 );
dff g5471_reg ( clk, reset, n10625, n2236 );
not U_inv824 ( n19514, n10625 );
dff g5475_reg ( clk, reset, n10623, n2241 );
not U_inv825 ( n19409, n10623 );
dff g5481_reg ( clk, reset, n10736, n2246 );
not U_inv826 ( n19408, n10736 );
dff g5485_reg ( clk, reset, n10780, n2251 );
not U_inv827 ( n19528, n10780 );
dff g5489_reg ( clk, reset, ex_wire227, n2256 );
not U_inv828 ( n19711, ex_wire227 );
dff g5495_reg ( clk, reset, n10735, n2261 );
not U_inv829 ( n19712, n10735 );
dff g5499_reg ( clk, reset, ex_wire228, n2266 );
not U_inv830 ( n19529, ex_wire228 );
dff g4821_reg ( clk, reset, n10892, n2216 );
dff g5156_reg ( clk, reset, n10865, n1862 );
not U_inv831 ( n19420, n10865 );
dff g5120_reg ( clk, reset, n10380, n1867 );
dff g5224_reg ( clk, reset, ex_wire229, n1762 );
not U_inv832 ( n19656, ex_wire229 );
dff g5240_reg ( clk, reset, ex_wire230, n1767 );
not U_inv833 ( n19657, ex_wire230 );
dff g5256_reg ( clk, reset, ex_wire231, n1772 );
not U_inv834 ( n19658, ex_wire231 );
dff g5204_reg ( clk, reset, ex_wire232, n1777 );
not U_inv835 ( n19659, ex_wire232 );
dff g5200_reg ( clk, reset, n10810, n1782 );
not U_inv836 ( n19660, n10810 );
dff g5228_reg ( clk, reset, n10868, n1787 );
not U_inv837 ( n19661, n10868 );
dff g5244_reg ( clk, reset, ex_wire233, n1792 );
not U_inv838 ( n19662, ex_wire233 );
dff g5260_reg ( clk, reset, n10867, n1797 );
not U_inv839 ( n19663, n10867 );
dff g5212_reg ( clk, reset, ex_wire234, n1802 );
not U_inv840 ( n19664, ex_wire234 );
dff g5208_reg ( clk, reset, ex_wire235, n1807 );
not U_inv841 ( n19665, ex_wire235 );
dff g5232_reg ( clk, reset, ex_wire236, n1812 );
not U_inv842 ( n19666, ex_wire236 );
dff g5248_reg ( clk, reset, ex_wire237, n1817 );
not U_inv843 ( n19667, ex_wire237 );
dff g5264_reg ( clk, reset, ex_wire238, n1822 );
not U_inv844 ( n19668, ex_wire238 );
dff g5220_reg ( clk, reset, ex_wire239, n1827 );
not U_inv845 ( n19669, ex_wire239 );
dff g5216_reg ( clk, reset, n10809, n1832 );
not U_inv846 ( n19670, n10809 );
dff g5236_reg ( clk, reset, n10866, n1837 );
not U_inv847 ( n19671, n10866 );
dff g5252_reg ( clk, reset, ex_wire240, n1842 );
not U_inv848 ( n19672, ex_wire240 );
dff g5268_reg ( clk, reset, n10563, n1847 );
dff g5272_reg ( clk, reset, ex_wire241, n1852 );
not U_inv849 ( n19673, ex_wire241 );
dff g5115_reg ( clk, reset, n10491, n1872 );
not U_inv850 ( n19674, n10491 );
dff g5124_reg ( clk, reset, ex_wire242, n1877 );
not U_inv851 ( n19515, ex_wire242 );
dff g5128_reg ( clk, reset, n10624, n1882 );
not U_inv852 ( n19419, n10624 );
dff g5134_reg ( clk, reset, n10738, n1887 );
not U_inv853 ( n19418, n10738 );
dff g5138_reg ( clk, reset, n10781, n1892 );
not U_inv854 ( n19526, n10781 );
dff g5142_reg ( clk, reset, ex_wire243, n1897 );
not U_inv855 ( n19675, ex_wire243 );
dff g5148_reg ( clk, reset, n10737, n1902 );
not U_inv856 ( n19676, n10737 );
dff g5152_reg ( clk, reset, ex_wire244, n1907 );
not U_inv857 ( n19527, ex_wire244 );
dff g128_reg ( clk, reset, g21245, n1857 );
not U_inv858 ( n19443, g21245 );
dff g94_reg ( clk, reset, g20652, n7498 );
not U_inv859 ( n20238, g20652 );
dff g2689_reg ( clk, reset, n10238, n7253 );
not U_inv860 ( n20196, n10238 );
dff g2697_reg ( clk, reset, n10296, n7258 );
dff g2704_reg ( clk, reset, n10383, n7263 );
not U_inv861 ( n20197, n10383 );
dff g2130_reg ( clk, reset, n10237, n6708 );
not U_inv862 ( n20141, n10237 );
dff g2138_reg ( clk, reset, n10295, n6713 );
dff g2145_reg ( clk, reset, n10382, n6718 );
not U_inv863 ( n20142, n10382 );
dff g2886_reg ( clk, reset, ex_wire245, n7533 );
not U_inv864 ( n19331, ex_wire245 );
dff g2980_reg ( clk, reset, n10772, n7538 );
not U_inv865 ( n19329, n10772 );
dff g947_reg ( clk, reset, n10586, n6158 );
not U_inv866 ( n20088, n10586 );
dff g952_reg ( clk, reset, ex_wire246, n6163 );
not U_inv867 ( n20089, ex_wire246 );
dff g939_reg ( clk, reset, n10784, n6168 );
not U_inv868 ( n19332, n10784 );
dff g2868_reg ( clk, reset, n10507, n7458 );
not U_inv869 ( n20218, n10507 );
dff g2873_reg ( clk, reset, n10364, n7463 );
dff g2890_reg ( clk, reset, ex_wire247, n7468 );
not U_inv870 ( n19321, ex_wire247 );
dff g1291_reg ( clk, reset, n10587, n5832 );
not U_inv871 ( n20050, n10587 );
dff g2153_reg ( clk, reset, n10320, n6733 );
not U_inv872 ( n19172, n10320 );
dff g2204_reg ( clk, reset, ex_wire248, n6738 );
not U_inv873 ( n20143, ex_wire248 );
dff g2197_reg ( clk, reset, n10298, n6743 );
not U_inv874 ( n20144, n10298 );
dff g2227_reg ( clk, reset, n10389, n6748 );
not U_inv875 ( n20145, n10389 );
dff g112_reg ( clk, reset, ex_wire249, new_g34843_ );
not U_inv876 ( n19565, ex_wire249 );
dff g2555_reg ( clk, reset, n10353, n7123 );
not U_inv877 ( n19149, n10353 );
dff g2606_reg ( clk, reset, ex_wire250, n7128 );
not U_inv878 ( n20183, ex_wire250 );
dff g2599_reg ( clk, reset, n10312, n7133 );
not U_inv879 ( n20184, n10312 );
dff g2629_reg ( clk, reset, n10438, n7138 );
not U_inv880 ( n20185, n10438 );
dff g2643_reg ( clk, reset, n10524, n7143 );
dff g2648_reg ( clk, reset, n10751, n7148 );
not U_inv881 ( n19148, n10751 );
dff g2567_reg ( clk, reset, ex_wire251, n7153 );
not U_inv882 ( n20186, ex_wire251 );
dff g2563_reg ( clk, reset, ex_wire252, n7158 );
not U_inv883 ( n20187, ex_wire252 );
dff g2571_reg ( clk, reset, ex_wire253, n7163 );
not U_inv884 ( n20188, ex_wire253 );
dff g2583_reg ( clk, reset, ex_wire254, n7168 );
not U_inv885 ( n20189, ex_wire254 );
dff g2579_reg ( clk, reset, ex_wire255, n7173 );
not U_inv886 ( n19147, ex_wire255 );
dff g2575_reg ( clk, reset, n10523, n7178 );
dff g2421_reg ( clk, reset, n10354, n6993 );
not U_inv887 ( n19157, n10354 );
dff g2472_reg ( clk, reset, ex_wire256, n6998 );
not U_inv888 ( n20170, ex_wire256 );
dff g2465_reg ( clk, reset, n10313, n7003 );
not U_inv889 ( n20171, n10313 );
dff g2495_reg ( clk, reset, n10439, n7008 );
not U_inv890 ( n20172, n10439 );
dff g2509_reg ( clk, reset, n10526, n7013 );
dff g2514_reg ( clk, reset, n10752, n7018 );
not U_inv891 ( n19156, n10752 );
dff g2433_reg ( clk, reset, ex_wire257, n7023 );
not U_inv892 ( n20173, ex_wire257 );
dff g2429_reg ( clk, reset, ex_wire258, n7028 );
not U_inv893 ( n20174, ex_wire258 );
dff g2437_reg ( clk, reset, ex_wire259, n7033 );
not U_inv894 ( n20175, ex_wire259 );
dff g2449_reg ( clk, reset, ex_wire260, n7038 );
not U_inv895 ( n20176, ex_wire260 );
dff g2445_reg ( clk, reset, ex_wire261, n7043 );
not U_inv896 ( n19155, ex_wire261 );
dff g2441_reg ( clk, reset, n10525, n7048 );
dff g2287_reg ( clk, reset, n10319, n6863 );
not U_inv897 ( n19165, n10319 );
dff g2338_reg ( clk, reset, ex_wire262, n6868 );
not U_inv898 ( n20157, ex_wire262 );
dff g2331_reg ( clk, reset, n10297, n6873 );
not U_inv899 ( n20158, n10297 );
dff g2361_reg ( clk, reset, n10388, n6878 );
not U_inv900 ( n20159, n10388 );
dff g2375_reg ( clk, reset, n10528, n6883 );
dff g2380_reg ( clk, reset, n10753, n6888 );
not U_inv901 ( n19164, n10753 );
dff g2299_reg ( clk, reset, ex_wire263, n6893 );
not U_inv902 ( n20160, ex_wire263 );
dff g2295_reg ( clk, reset, ex_wire264, n6898 );
not U_inv903 ( n20161, ex_wire264 );
dff g2303_reg ( clk, reset, ex_wire265, n6903 );
not U_inv904 ( n20162, ex_wire265 );
dff g2315_reg ( clk, reset, n10789, n6908 );
not U_inv905 ( n20163, n10789 );
dff g2311_reg ( clk, reset, ex_wire266, n6913 );
not U_inv906 ( n19163, ex_wire266 );
dff g2307_reg ( clk, reset, n10527, n6918 );
dff g1996_reg ( clk, reset, n10355, n6578 );
not U_inv907 ( n19180, n10355 );
dff g2047_reg ( clk, reset, ex_wire267, n6583 );
not U_inv908 ( n20128, ex_wire267 );
dff g2040_reg ( clk, reset, n10314, n6588 );
not U_inv909 ( n20129, n10314 );
dff g2070_reg ( clk, reset, n10440, n6593 );
not U_inv910 ( n20130, n10440 );
dff g2084_reg ( clk, reset, n10532, n6598 );
dff g2089_reg ( clk, reset, n10755, n6603 );
not U_inv911 ( n19179, n10755 );
dff g2008_reg ( clk, reset, ex_wire268, n6608 );
not U_inv912 ( n20131, ex_wire268 );
dff g2004_reg ( clk, reset, ex_wire269, n6613 );
not U_inv913 ( n20132, ex_wire269 );
dff g2012_reg ( clk, reset, ex_wire270, n6618 );
not U_inv914 ( n20133, ex_wire270 );
dff g2024_reg ( clk, reset, ex_wire271, n6623 );
not U_inv915 ( n20134, ex_wire271 );
dff g2020_reg ( clk, reset, ex_wire272, n6628 );
not U_inv916 ( n19178, ex_wire272 );
dff g2016_reg ( clk, reset, n10531, n6633 );
dff g1862_reg ( clk, reset, n10356, n6448 );
not U_inv917 ( n19188, n10356 );
dff g1913_reg ( clk, reset, ex_wire273, n6453 );
not U_inv918 ( n20115, ex_wire273 );
dff g1906_reg ( clk, reset, n10315, n6458 );
not U_inv919 ( n20116, n10315 );
dff g1936_reg ( clk, reset, n10441, n6463 );
not U_inv920 ( n20117, n10441 );
dff g1950_reg ( clk, reset, n10534, n6468 );
dff g1955_reg ( clk, reset, n10756, n6473 );
not U_inv921 ( n19187, n10756 );
dff g1874_reg ( clk, reset, ex_wire274, n6478 );
not U_inv922 ( n20118, ex_wire274 );
dff g1870_reg ( clk, reset, ex_wire275, n6483 );
not U_inv923 ( n20119, ex_wire275 );
dff g1878_reg ( clk, reset, ex_wire276, n6488 );
not U_inv924 ( n20120, ex_wire276 );
dff g1890_reg ( clk, reset, ex_wire277, n6493 );
not U_inv925 ( n20121, ex_wire277 );
dff g1886_reg ( clk, reset, ex_wire278, n6498 );
not U_inv926 ( n19186, ex_wire278 );
dff g1882_reg ( clk, reset, n10533, n6503 );
dff g1728_reg ( clk, reset, n10321, n6318 );
not U_inv927 ( n19196, n10321 );
dff g1779_reg ( clk, reset, ex_wire279, n6323 );
not U_inv928 ( n20102, ex_wire279 );
dff g1772_reg ( clk, reset, n10299, n6328 );
not U_inv929 ( n20103, n10299 );
dff g1802_reg ( clk, reset, n10390, n6333 );
not U_inv930 ( n20104, n10390 );
dff g1816_reg ( clk, reset, n10536, n6338 );
dff g1821_reg ( clk, reset, n10757, n6343 );
not U_inv931 ( n19195, n10757 );
dff g1740_reg ( clk, reset, ex_wire280, n6348 );
not U_inv932 ( n20105, ex_wire280 );
dff g1736_reg ( clk, reset, ex_wire281, n6353 );
not U_inv933 ( n20106, ex_wire281 );
dff g1744_reg ( clk, reset, ex_wire282, n6358 );
not U_inv934 ( n20107, ex_wire282 );
dff g1756_reg ( clk, reset, n10791, n6363 );
not U_inv935 ( n20108, n10791 );
dff g1752_reg ( clk, reset, ex_wire283, n6368 );
not U_inv936 ( n19194, ex_wire283 );
dff g1748_reg ( clk, reset, n10535, n6373 );
dff g1644_reg ( clk, reset, ex_wire284, n6193 );
not U_inv937 ( n20090, ex_wire284 );
dff g1636_reg ( clk, reset, n10316, n6198 );
not U_inv938 ( n20091, n10316 );
dff g1668_reg ( clk, reset, n10442, n6203 );
not U_inv939 ( n20092, n10442 );
dff g1592_reg ( clk, reset, n10357, n6188 );
not U_inv940 ( n19208, n10357 );
dff g1682_reg ( clk, reset, n10537, n6208 );
dff g1687_reg ( clk, reset, n10758, n6213 );
not U_inv941 ( n19207, n10758 );
dff g1604_reg ( clk, reset, ex_wire285, n6218 );
not U_inv942 ( n20093, ex_wire285 );
dff g1600_reg ( clk, reset, n10793, n6223 );
not U_inv943 ( n19206, n10793 );
dff g1608_reg ( clk, reset, ex_wire286, n6228 );
not U_inv944 ( n19205, ex_wire286 );
dff g1620_reg ( clk, reset, n10912, n6233 );
not U_inv945 ( n20094, n10912 );
dff g1616_reg ( clk, reset, ex_wire287, n6238 );
not U_inv946 ( n19204, ex_wire287 );
dff g1612_reg ( clk, reset, n10792, n6243 );
not U_inv947 ( n19203, n10792 );
dff g2241_reg ( clk, reset, n10530, n6753 );
dff g2246_reg ( clk, reset, n10754, n6758 );
not U_inv948 ( n19171, n10754 );
dff g2165_reg ( clk, reset, ex_wire288, n6763 );
not U_inv949 ( n20146, ex_wire288 );
dff g2161_reg ( clk, reset, ex_wire289, n6768 );
not U_inv950 ( n20147, ex_wire289 );
dff g2169_reg ( clk, reset, ex_wire290, n6773 );
not U_inv951 ( n20148, ex_wire290 );
dff g2181_reg ( clk, reset, n10790, n6778 );
not U_inv952 ( n20149, n10790 );
dff g2177_reg ( clk, reset, ex_wire291, n6783 );
not U_inv953 ( n19170, ex_wire291 );
dff g2173_reg ( clk, reset, n10529, n6788 );
dff g2193_reg ( clk, reset, n10826, n6793 );
not U_inv954 ( n19169, n10826 );
dff g2185_reg ( clk, reset, ex_wire292, n6798 );
not U_inv955 ( n20150, ex_wire292 );
dff g2208_reg ( clk, reset, n10234, n6803 );
not U_inv956 ( n20151, n10234 );
dff g2223_reg ( clk, reset, ex_wire293, n6808 );
not U_inv957 ( n20152, ex_wire293 );
dff g2217_reg ( clk, reset, n10411, n6813 );
not U_inv958 ( n20153, n10411 );
dff g110_reg ( clk, reset, ex_wire294, new_g34781_ );
not U_inv959 ( n19200, ex_wire294 );
dff g1894_reg ( clk, reset, ex_wire295, n6513 );
not U_inv960 ( n20122, ex_wire295 );
dff g1917_reg ( clk, reset, n10342, n6518 );
not U_inv961 ( n20123, n10342 );
dff g1932_reg ( clk, reset, ex_wire296, n6523 );
not U_inv962 ( n20124, ex_wire296 );
dff g1926_reg ( clk, reset, n10413, n6528 );
not U_inv963 ( n20125, n10413 );
dff g1902_reg ( clk, reset, n10828, n6508 );
not U_inv964 ( n19185, n10828 );
dff g2791_reg ( clk, reset, n10820, n7353 );
not U_inv965 ( n19137, n10820 );
dff g2795_reg ( clk, reset, n10819, n7358 );
not U_inv966 ( n19136, n10819 );
dff g2787_reg ( clk, reset, n10635, n7363 );
not U_inv967 ( n20207, n10635 );
dff g2066_reg ( clk, reset, ex_wire297, n6653 );
not U_inv968 ( n20137, ex_wire297 );
dff g2060_reg ( clk, reset, n10412, n6658 );
not U_inv969 ( n20138, n10412 );
dff g2036_reg ( clk, reset, n10827, n6638 );
not U_inv970 ( n19177, n10827 );
dff g2028_reg ( clk, reset, ex_wire298, n6643 );
not U_inv971 ( n20135, ex_wire298 );
dff g2051_reg ( clk, reset, n10341, n6648 );
not U_inv972 ( n20136, n10341 );
dff g2079_reg ( clk, reset, n10686, n6663 );
not U_inv973 ( n19176, n10686 );
dff g2093_reg ( clk, reset, n10426, n6668 );
not U_inv974 ( n19175, n10426 );
dff g2098_reg ( clk, reset, ex_wire299, n6673 );
not U_inv975 ( n19559, ex_wire299 );
dff g2102_reg ( clk, reset, n10574, n6678 );
not U_inv976 ( n20139, n10574 );
dff g2108_reg ( clk, reset, n10715, n6683 );
not U_inv977 ( n20140, n10715 );
dff g2112_reg ( clk, reset, ex_wire300, n6688 );
not U_inv978 ( n19549, ex_wire300 );
dff g2116_reg ( clk, reset, n10630, n6693 );
not U_inv979 ( n19174, n10630 );
dff g2122_reg ( clk, reset, n10714, n6698 );
not U_inv980 ( n19173, n10714 );
dff g2126_reg ( clk, reset, ex_wire301, n6703 );
not U_inv981 ( n19548, ex_wire301 );
dff g2783_reg ( clk, reset, ex_wire302, n7368 );
not U_inv982 ( n20208, ex_wire302 );
dff g2775_reg ( clk, reset, n10560, n7373 );
not U_inv983 ( n20209, n10560 );
dff g1768_reg ( clk, reset, n10829, n6378 );
not U_inv984 ( n19193, n10829 );
dff g1760_reg ( clk, reset, ex_wire303, n6383 );
not U_inv985 ( n20109, ex_wire303 );
dff g1783_reg ( clk, reset, n10235, n6388 );
not U_inv986 ( n20110, n10235 );
dff g1798_reg ( clk, reset, ex_wire304, n6393 );
not U_inv987 ( n20111, ex_wire304 );
dff g1792_reg ( clk, reset, n10414, n6398 );
not U_inv988 ( n20112, n10414 );
dff g1811_reg ( clk, reset, n10688, n6403 );
not U_inv989 ( n19192, n10688 );
dff g1825_reg ( clk, reset, n10428, n6408 );
not U_inv990 ( n19191, n10428 );
dff g1830_reg ( clk, reset, ex_wire305, n6413 );
not U_inv991 ( n19561, ex_wire305 );
dff g1834_reg ( clk, reset, n10576, n6418 );
not U_inv992 ( n20113, n10576 );
dff g1840_reg ( clk, reset, n10719, n6423 );
not U_inv993 ( n20114, n10719 );
dff g1844_reg ( clk, reset, ex_wire306, n6428 );
not U_inv994 ( n19553, ex_wire306 );
dff g1848_reg ( clk, reset, n10632, n6433 );
not U_inv995 ( n19190, n10632 );
dff g1854_reg ( clk, reset, n10718, n6438 );
not U_inv996 ( n19189, n10718 );
dff g1858_reg ( clk, reset, ex_wire307, n6443 );
not U_inv997 ( n19552, ex_wire307 );
dff g2771_reg ( clk, reset, n10369, n7378 );
not U_inv998 ( n20210, n10369 );
dff g85_reg ( clk, reset, ex_wire308, g33435 );
not U_inv999 ( n19135, ex_wire308 );
dff g1632_reg ( clk, reset, n10830, n6248 );
not U_inv1000 ( n19202, n10830 );
dff g2767_reg ( clk, reset, n10822, n7343 );
not U_inv1001 ( n19139, n10822 );
dff g2779_reg ( clk, reset, n10821, n7348 );
not U_inv1002 ( n19138, n10821 );
dff g1624_reg ( clk, reset, ex_wire309, n6253 );
not U_inv1003 ( n20095, ex_wire309 );
dff g1648_reg ( clk, reset, n10350, n6258 );
not U_inv1004 ( n20096, n10350 );
dff g1664_reg ( clk, reset, ex_wire310, n6263 );
not U_inv1005 ( n20097, ex_wire310 );
dff g1657_reg ( clk, reset, n10348, n6268 );
not U_inv1006 ( n20098, n10348 );
dff g1677_reg ( clk, reset, n10696, n6273 );
not U_inv1007 ( n20099, n10696 );
dff g1691_reg ( clk, reset, n10429, n6278 );
not U_inv1008 ( n19199, n10429 );
dff g1696_reg ( clk, reset, ex_wire311, n6283 );
not U_inv1009 ( n19560, ex_wire311 );
dff g1700_reg ( clk, reset, n10577, n6288 );
not U_inv1010 ( n20100, n10577 );
dff g1706_reg ( clk, reset, n10721, n6293 );
not U_inv1011 ( n20101, n10721 );
dff g1710_reg ( clk, reset, ex_wire312, n6298 );
not U_inv1012 ( n19551, ex_wire312 );
dff g1714_reg ( clk, reset, n10633, n6303 );
not U_inv1013 ( n19198, n10633 );
dff g1720_reg ( clk, reset, n10720, n6308 );
not U_inv1014 ( n19197, n10720 );
dff g1724_reg ( clk, reset, ex_wire313, n6313 );
not U_inv1015 ( n19550, ex_wire313 );
dff g1945_reg ( clk, reset, n10687, n6533 );
not U_inv1016 ( n19184, n10687 );
dff g2831_reg ( clk, reset, ex_wire314, n7383 );
not U_inv1017 ( g30331, ex_wire314 );
dff g121_reg ( clk, reset, g20654, n7388 );
dff g2799_reg ( clk, reset, n10818, n7393 );
not U_inv1018 ( n19134, n10818 );
dff g2811_reg ( clk, reset, n10817, n7398 );
not U_inv1019 ( n19133, n10817 );
dff g2823_reg ( clk, reset, n10816, n7403 );
not U_inv1020 ( n19132, n10816 );
dff g2827_reg ( clk, reset, n10815, n7408 );
not U_inv1021 ( n19131, n10815 );
dff g2819_reg ( clk, reset, n10634, n7413 );
not U_inv1022 ( n20211, n10634 );
dff g2625_reg ( clk, reset, ex_wire315, n7198 );
not U_inv1023 ( n20192, ex_wire315 );
dff g2619_reg ( clk, reset, n10408, n7203 );
not U_inv1024 ( n20193, n10408 );
dff g2595_reg ( clk, reset, n10823, n7183 );
not U_inv1025 ( n19146, n10823 );
dff g2587_reg ( clk, reset, ex_wire316, n7188 );
not U_inv1026 ( n20190, ex_wire316 );
dff g2610_reg ( clk, reset, n10339, n7193 );
not U_inv1027 ( n20191, n10339 );
dff g2638_reg ( clk, reset, n10683, n7208 );
not U_inv1028 ( n19145, n10683 );
dff g2652_reg ( clk, reset, n10422, n7213 );
not U_inv1029 ( n19144, n10422 );
dff g2657_reg ( clk, reset, ex_wire317, n7218 );
not U_inv1030 ( n19555, ex_wire317 );
dff g2661_reg ( clk, reset, n10570, n7223 );
not U_inv1031 ( n20194, n10570 );
dff g2667_reg ( clk, reset, n10707, n7228 );
not U_inv1032 ( n20195, n10707 );
dff g2671_reg ( clk, reset, ex_wire318, n7233 );
not U_inv1033 ( n19541, ex_wire318 );
dff g2675_reg ( clk, reset, n10626, n7238 );
not U_inv1034 ( n19143, n10626 );
dff g2681_reg ( clk, reset, n10706, n7243 );
not U_inv1035 ( n19142, n10706 );
dff g2685_reg ( clk, reset, ex_wire319, n7248 );
not U_inv1036 ( n19540, ex_wire319 );
dff g2815_reg ( clk, reset, ex_wire320, n7418 );
not U_inv1037 ( n20212, ex_wire320 );
dff g2491_reg ( clk, reset, ex_wire321, n7068 );
not U_inv1038 ( n20179, ex_wire321 );
dff g2485_reg ( clk, reset, n10409, n7073 );
not U_inv1039 ( n20180, n10409 );
dff g2461_reg ( clk, reset, n10824, n7053 );
not U_inv1040 ( n19154, n10824 );
dff g2453_reg ( clk, reset, ex_wire322, n7058 );
not U_inv1041 ( n20177, ex_wire322 );
dff g2476_reg ( clk, reset, n10340, n7063 );
not U_inv1042 ( n20178, n10340 );
dff g2504_reg ( clk, reset, n10684, n7078 );
not U_inv1043 ( n19153, n10684 );
dff g2518_reg ( clk, reset, n10423, n7083 );
not U_inv1044 ( n19152, n10423 );
dff g2523_reg ( clk, reset, ex_wire323, n7088 );
not U_inv1045 ( n19554, ex_wire323 );
dff g2527_reg ( clk, reset, n10571, n7093 );
not U_inv1046 ( n20181, n10571 );
dff g2533_reg ( clk, reset, n10709, n7098 );
not U_inv1047 ( n20182, n10709 );
dff g2537_reg ( clk, reset, ex_wire324, n7103 );
not U_inv1048 ( n19539, ex_wire324 );
dff g2541_reg ( clk, reset, n10627, n7108 );
not U_inv1049 ( n19151, n10627 );
dff g2547_reg ( clk, reset, n10708, n7113 );
not U_inv1050 ( n19150, n10708 );
dff g2551_reg ( clk, reset, ex_wire325, n7118 );
not U_inv1051 ( n19538, ex_wire325 );
dff g2807_reg ( clk, reset, n10559, n7423 );
not U_inv1052 ( n20213, n10559 );
dff g2357_reg ( clk, reset, ex_wire326, n6938 );
not U_inv1053 ( n20166, ex_wire326 );
dff g2351_reg ( clk, reset, n10410, n6943 );
not U_inv1054 ( n20167, n10410 );
dff g2327_reg ( clk, reset, n10825, n6923 );
not U_inv1055 ( n19162, n10825 );
dff g2319_reg ( clk, reset, ex_wire327, n6928 );
not U_inv1056 ( n20164, ex_wire327 );
dff g2342_reg ( clk, reset, n10233, n6933 );
not U_inv1057 ( n20165, n10233 );
dff g2370_reg ( clk, reset, n10685, n6948 );
not U_inv1058 ( n19161, n10685 );
dff g2384_reg ( clk, reset, n10424, n6953 );
not U_inv1059 ( n19160, n10424 );
dff g2389_reg ( clk, reset, ex_wire328, n6958 );
not U_inv1060 ( n19557, ex_wire328 );
dff g2393_reg ( clk, reset, n10572, n6963 );
not U_inv1061 ( n20168, n10572 );
dff g2399_reg ( clk, reset, n10711, n6968 );
not U_inv1062 ( n20169, n10711 );
dff g2403_reg ( clk, reset, ex_wire329, n6973 );
not U_inv1063 ( n19545, ex_wire329 );
dff g2407_reg ( clk, reset, n10628, n6978 );
not U_inv1064 ( n19159, n10628 );
dff g2413_reg ( clk, reset, n10710, n6983 );
not U_inv1065 ( n19158, n10710 );
dff g2417_reg ( clk, reset, ex_wire330, n6988 );
not U_inv1066 ( n19544, ex_wire330 );
dff g2803_reg ( clk, reset, n10358, n7428 );
not U_inv1067 ( n20214, n10358 );
dff g111_reg ( clk, reset, ex_wire331, g33079 );
not U_inv1068 ( n19130, ex_wire331 );
dff g1959_reg ( clk, reset, n10427, n6538 );
not U_inv1069 ( n19183, n10427 );
dff g1964_reg ( clk, reset, ex_wire332, n6543 );
not U_inv1070 ( n19558, ex_wire332 );
dff g1968_reg ( clk, reset, n10575, n6548 );
not U_inv1071 ( n20126, n10575 );
dff g1974_reg ( clk, reset, n10717, n6553 );
not U_inv1072 ( n20127, n10717 );
dff g1978_reg ( clk, reset, ex_wire333, n6558 );
not U_inv1073 ( n19547, ex_wire333 );
dff g1982_reg ( clk, reset, n10631, n6563 );
not U_inv1074 ( n19182, n10631 );
dff g1988_reg ( clk, reset, n10716, n6568 );
not U_inv1075 ( n19181, n10716 );
dff g1992_reg ( clk, reset, ex_wire334, n6573 );
not U_inv1076 ( n19546, ex_wire334 );
dff g2236_reg ( clk, reset, n10695, n6818 );
not U_inv1077 ( n20154, n10695 );
dff g2834_reg ( clk, reset, ex_wire335, n7433 );
not U_inv1078 ( g30330, ex_wire335 );
dff g117_reg ( clk, reset, g21270, n7438 );
dff g2250_reg ( clk, reset, n10425, n6823 );
not U_inv1079 ( n19168, n10425 );
dff g2255_reg ( clk, reset, ex_wire336, n6828 );
not U_inv1080 ( n19556, ex_wire336 );
dff g2259_reg ( clk, reset, n10573, n6833 );
not U_inv1081 ( n20155, n10573 );
dff g2265_reg ( clk, reset, n10713, n6838 );
not U_inv1082 ( n20156, n10713 );
dff g2269_reg ( clk, reset, ex_wire337, n6843 );
not U_inv1083 ( n19543, ex_wire337 );
dff g2273_reg ( clk, reset, n10629, n6848 );
not U_inv1084 ( n19167, n10629 );
dff g2279_reg ( clk, reset, n10712, n6853 );
not U_inv1085 ( n19166, n10712 );
dff g2283_reg ( clk, reset, ex_wire338, n6858 );
not U_inv1086 ( n19542, ex_wire338 );
dff g2848_reg ( clk, reset, n10782, n7503 );
not U_inv1087 ( n20219, n10782 );
dff g2844_reg ( clk, reset, n10539, n7473 );
dff g538_reg ( clk, reset, n10831, n5403 );
not U_inv1088 ( n19489, n10831 );
dff g546_reg ( clk, reset, ex_wire339, n5408 );
not U_inv1089 ( n19475, ex_wire339 );
dff g542_reg ( clk, reset, ex_wire340, n5413 );
not U_inv1090 ( n19466, ex_wire340 );
dff g534_reg ( clk, reset, ex_wire341, n5418 );
not U_inv1091 ( n19461, ex_wire341 );
dff g550_reg ( clk, reset, n10813, n5423 );
not U_inv1092 ( n19336, n10813 );
dff g3853_reg ( clk, reset, n10931, n4425 );
not U_inv1093 ( n19486, n10931 );
dff g6199_reg ( clk, reset, n10930, n2989 );
not U_inv1094 ( n19491, n10930 );
dff g4727_reg ( clk, reset, n10511, n1431 );
not U_inv1095 ( n19490, n10511 );
dff g4917_reg ( clk, reset, n10513, n1264 );
not U_inv1096 ( n19494, n10513 );
dff g55_reg ( clk, reset, g55, n51 );
dff g2856_reg ( clk, reset, n10783, n7508 );
not U_inv1097 ( n19484, n10783 );
dff g2852_reg ( clk, reset, n10540, n7478 );
dff g2860_reg ( clk, reset, n10541, n7483 );
dff g4732_reg ( clk, reset, n10367, n1436 );
dff g4717_reg ( clk, reset, n10515, n1441 );
not U_inv1098 ( n19479, n10515 );
dff g4922_reg ( clk, reset, n10368, n1269 );
dff g4907_reg ( clk, reset, n10516, n1274 );
not U_inv1099 ( n19480, n10516 );
dff g2999_reg ( clk, reset, n10833, n7443 );
not U_inv1100 ( n20215, n10833 );
dff g3502_reg ( clk, reset, n10933, n4066 );
not U_inv1101 ( n19483, n10933 );
dff g5853_reg ( clk, reset, n10932, n2630 );
not U_inv1102 ( n19485, n10932 );
dff g2927_reg ( clk, reset, n10677, n7593 );
not U_inv1103 ( n20230, n10677 );
dff g2941_reg ( clk, reset, n10705, n7598 );
not U_inv1104 ( n20231, n10705 );
dff g2955_reg ( clk, reset, n10281, n7603 );
not U_inv1105 ( n19465, n10281 );
dff g2965_reg ( clk, reset, ex_wire342, n7608 );
not U_inv1106 ( n20232, ex_wire342 );
dff g2975_reg ( clk, reset, ex_wire343, n7613 );
not U_inv1107 ( n20233, ex_wire343 );
dff g3003_reg ( clk, reset, ex_wire344, new_g18597_ );
not U_inv1108 ( n19110, ex_wire344 );
dff g943_reg ( clk, reset, n10926, n6173 );
not U_inv1109 ( n19323, n10926 );
dff g1287_reg ( clk, reset, n10927, n5847 );
not U_inv1110 ( n19324, n10927 );
dff g4939_reg ( clk, reset, n10556, n1361 );
dff g4722_reg ( clk, reset, n10510, n1446 );
not U_inv1111 ( n19470, n10510 );
dff g4912_reg ( clk, reset, n10512, n1279 );
not U_inv1112 ( n19471, n10512 );
dff g4572_reg ( clk, reset, ex_wire345, n177 );
not U_inv1113 ( n19453, ex_wire345 );
dff g4495_reg ( clk, reset, g4495, n862 );
dff g4498_reg ( clk, reset, g4498, n867 );
dff g4501_reg ( clk, reset, g4501, n872 );
dff g4504_reg ( clk, reset, ex_wire346, n877 );
not U_inv1114 ( n19123, ex_wire346 );
dff g4512_reg ( clk, reset, n10869, n882 );
dff g4521_reg ( clk, reset, n10284, n887 );
not U_inv1115 ( n19117, n10284 );
dff g4527_reg ( clk, reset, ex_wire347, n892 );
not U_inv1116 ( n19118, ex_wire347 );
dff g4515_reg ( clk, reset, n10835, n897 );
not U_inv1117 ( n19501, n10835 );
dff g4519_reg ( clk, reset, g4519, n902 );
dff g4520_reg ( clk, reset, n911, g4519 );
dff g4483_reg ( clk, reset, ex_wire348, n911 );
not U_inv1118 ( n19120, ex_wire348 );
dff g4486_reg ( clk, reset, ex_wire349, n916 );
not U_inv1119 ( n19119, ex_wire349 );
dff g4489_reg ( clk, reset, ex_wire350, n921 );
not U_inv1120 ( n19122, ex_wire350 );
dff g4492_reg ( clk, reset, ex_wire351, n926 );
not U_inv1121 ( n19121, ex_wire351 );
dff g4537_reg ( clk, reset, g10306, n931 );
dff g4423_reg ( clk, reset, ex_wire352, g10306 );
not U_inv1122 ( n19512, ex_wire352 );
dff g4438_reg ( clk, reset, n10907, n145 );
not U_inv1123 ( n19575, n10907 );
dff g4375_reg ( clk, reset, n10592, n1047 );
not U_inv1124 ( n19577, n10592 );
dff g4414_reg ( clk, reset, g7257, n1052 );
dff g4411_reg ( clk, reset, n10558, g7257 );
dff g4408_reg ( clk, reset, g7243, n1061 );
dff g4405_reg ( clk, reset, ex_wire353, g7243 );
not U_inv1125 ( n19578, ex_wire353 );
dff g4401_reg ( clk, reset, ex_wire354, n1070 );
not U_inv1126 ( n19508, ex_wire354 );
dff g4388_reg ( clk, reset, n10514, n1075 );
not U_inv1127 ( n19509, n10514 );
dff g4382_reg ( clk, reset, ex_wire355, n1080 );
not U_inv1128 ( n19579, ex_wire355 );
dff g4417_reg ( clk, reset, n10704, n1085 );
not U_inv1129 ( n19507, n10704 );
dff g4392_reg ( clk, reset, n10251, n1090 );
not U_inv1130 ( n19580, n10251 );
dff g4456_reg ( clk, reset, n1100, new_g24298_ );
dff g4455_reg ( clk, reset, g4455, n1100 );
dff g1_reg ( clk, reset, g12832, n1105 );
dff g4446_reg ( clk, reset, g7245, n1023 );
dff g4452_reg ( clk, reset, ex_wire356, g7245 );
not U_inv1131 ( n19576, ex_wire356 );
dff g4449_reg ( clk, reset, g7260, n1014 );
dff g4443_reg ( clk, reset, n10493, g7260 );
dff g4434_reg ( clk, reset, n10921, n1032 );
not U_inv1132 ( n19510, n10921 );
dff g4430_reg ( clk, reset, n10906, n1037 );
not U_inv1133 ( n19511, n10906 );
dff g4427_reg ( clk, reset, ex_wire357, n1042 );
not U_inv1134 ( n19517, ex_wire357 );
dff g4372_reg ( clk, reset, ex_wire358, n1219 );
not U_inv1135 ( n19124, ex_wire358 );
dff g4480_reg ( clk, reset, g4480, n857 );
dff g4578_reg ( clk, reset, g4578, n1304 );
dff g6545_reg ( clk, reset, n10937, n3348 );
not U_inv1136 ( n19468, n10937 );
dff g5160_reg ( clk, reset, n10936, n1912 );
not U_inv1137 ( n19472, n10936 );
dff g3151_reg ( clk, reset, n10935, n3707 );
not U_inv1138 ( n19477, n10935 );
dff g5507_reg ( clk, reset, n10934, n2271 );
not U_inv1139 ( n19481, n10934 );
dff g22_reg ( clk, reset, n10588, n137 );
not U_inv1140 ( n19111, n10588 );
dff g25_reg ( clk, reset, new_g10520_, new_g10520_ );
or U10125 ( n10301, n10965, n15649 );
not U10126 ( n15730, n10942 );
not U10127 ( n10942, n10301 );
not U10128 ( n10943, n10301 );
not U10129 ( n10944, n10301 );
nor U10130 ( n15240, n10954, n15328 );
buf U10131 ( n10945, n11051 );
buf U10132 ( n10946, n11051 );
buf U10133 ( n10947, n11050 );
buf U10134 ( n10948, n11050 );
buf U10135 ( n10949, n11050 );
buf U10136 ( n10950, n11049 );
buf U10137 ( n10951, n11049 );
buf U10138 ( n10952, n11049 );
buf U10139 ( n10953, n11048 );
buf U10140 ( n10954, n11048 );
buf U10141 ( n10955, n11048 );
buf U10142 ( n10956, n11047 );
buf U10143 ( n10957, n11047 );
buf U10144 ( n10958, n11047 );
buf U10145 ( n10959, n11046 );
buf U10146 ( n10960, n11046 );
buf U10147 ( n10961, n11046 );
buf U10148 ( n10962, n11045 );
buf U10149 ( n10963, n11045 );
buf U10150 ( n10964, n11045 );
buf U10151 ( n10965, n11044 );
buf U10152 ( n10966, n11044 );
buf U10153 ( n10967, n11044 );
buf U10154 ( n10968, n11043 );
buf U10155 ( n10969, n11043 );
buf U10156 ( n10970, n11043 );
buf U10157 ( n10971, n11042 );
buf U10158 ( n10972, n11042 );
buf U10159 ( n10973, n11042 );
buf U10160 ( n10974, n11041 );
buf U10161 ( n10975, n11041 );
buf U10162 ( n10976, n11041 );
buf U10163 ( n10977, n11040 );
buf U10164 ( n10978, n11040 );
buf U10165 ( n10979, n11040 );
buf U10166 ( n10980, n11039 );
buf U10167 ( n10981, n11039 );
buf U10168 ( n10982, n11039 );
buf U10169 ( n10983, n11038 );
buf U10170 ( n10984, n11038 );
buf U10171 ( n10985, n11038 );
buf U10172 ( n10986, n11037 );
buf U10173 ( n10987, n11037 );
buf U10174 ( n10988, n11037 );
buf U10175 ( n10989, n11036 );
buf U10176 ( n10990, n11036 );
buf U10177 ( n10991, n11036 );
buf U10178 ( n10992, n11035 );
buf U10179 ( n10993, n11035 );
buf U10180 ( n10994, n11035 );
buf U10181 ( n10995, n11034 );
buf U10182 ( n10996, n11034 );
buf U10183 ( n10997, n11034 );
buf U10184 ( n10998, n11033 );
buf U10185 ( n10999, n11033 );
buf U10186 ( n11000, n11033 );
buf U10187 ( n11001, n11032 );
buf U10188 ( n11002, n11032 );
buf U10189 ( n11003, n11032 );
buf U10190 ( n11004, n11031 );
buf U10191 ( n11005, n11031 );
buf U10192 ( n11006, n11031 );
buf U10193 ( n11007, n11030 );
buf U10194 ( n11008, n11030 );
buf U10195 ( n11009, n11030 );
buf U10196 ( n11010, n11029 );
buf U10197 ( n11011, n11029 );
buf U10198 ( n11012, n11029 );
buf U10199 ( n11013, n11028 );
buf U10200 ( n11014, n11028 );
buf U10201 ( n11015, n11028 );
buf U10202 ( n11016, n11027 );
buf U10203 ( n11017, n11027 );
buf U10204 ( n11018, n11027 );
buf U10205 ( n11019, n11026 );
buf U10206 ( n11020, n11026 );
buf U10207 ( n11021, n11026 );
buf U10208 ( n11022, n11025 );
buf U10209 ( n11023, n11025 );
buf U10210 ( n11024, n11025 );
buf U10211 ( n11025, n11226 );
buf U10212 ( n11026, n11226 );
buf U10213 ( n11027, n11226 );
buf U10214 ( n11028, n11226 );
buf U10215 ( n11029, n11226 );
buf U10216 ( n11030, n11226 );
buf U10217 ( n11031, n11226 );
buf U10218 ( n11032, n11226 );
buf U10219 ( n11033, n11226 );
buf U10220 ( n11034, n11226 );
buf U10221 ( n11035, n11226 );
buf U10222 ( n11036, n11226 );
buf U10223 ( n11037, n11226 );
buf U10224 ( n11038, n11226 );
buf U10225 ( n11039, n11226 );
buf U10226 ( n11040, n11226 );
buf U10227 ( n11041, n11226 );
buf U10228 ( n11042, n11226 );
buf U10229 ( n11043, n11226 );
buf U10230 ( n11044, n11226 );
buf U10231 ( n11045, n11226 );
buf U10232 ( n11046, n11226 );
buf U10233 ( n11047, n11226 );
buf U10234 ( n11048, n11226 );
buf U10235 ( n11049, n11226 );
buf U10236 ( n11050, n11226 );
buf U10237 ( n11051, n11226 );
nand U10238 ( g34972, n11052, n10588 );
or U10239 ( g34913, new_g34970_, n19111 );
or U10240 ( g34917, new_g34974_, n19111 );
or U10241 ( g34919, new_g34975_, n19111 );
or U10242 ( g34921, new_g34976_, n19111 );
or U10243 ( g34923, new_g34977_, n19111 );
or U10244 ( g34925, new_g34978_, n19111 );
or U10245 ( g34927, new_g34979_, n19111 );
or U10246 ( g34915, new_g34971_, n19111 );
nand U10247 ( g34383, n11053, n11054 );
nor U10248 ( n11053, new_g34843_, n11055 );
nor U10249 ( n11055, n11056, n11057 );
nand U10250 ( n11057, n11058, n11059 );
nor U10251 ( n11059, n11060, n11061 );
nor U10252 ( n11058, n11062, n11063 );
nand U10253 ( n11056, n11064, n11065 );
nor U10254 ( n11065, n11066, n11067 );
nor U10255 ( n11064, n11068, n11069 );
nand U10256 ( new_g34843_, n11070, n11071 );
nor U10257 ( n11071, n11072, n11073 );
nand U10258 ( n11073, n11074, n11075 );
nand U10259 ( n11075, n11076, n20103 );
nor U10260 ( n11076, n20104, n11077 );
nand U10261 ( n11074, n11069, n11078 );
nand U10262 ( n11072, n11079, n11080 );
nand U10263 ( n11080, n11081, n20158 );
nor U10264 ( n11081, n20159, n11082 );
nand U10265 ( n11079, n11083, n20144 );
nor U10266 ( n11083, n20145, n11084 );
nor U10267 ( n11070, n11085, n11086 );
nand U10268 ( n11086, n11087, n11088 );
nand U10269 ( n11088, n11063, n11089 );
nand U10270 ( n11087, g25259, n11066 );
nand U10271 ( n11085, n11090, n11091 );
nand U10272 ( n11091, n11060, n11092 );
nand U10273 ( n11090, n11062, n11093 );
nand U10274 ( g34425, n11094, n11095 );
not U10275 ( n11095, new_g34809_ );
nand U10276 ( new_g34809_, n11096, n11097 );
nand U10277 ( n11097, n11098, n10292 );
nand U10278 ( n11098, n11099, n11100 );
nor U10279 ( n11100, n11101, n11102 );
nor U10280 ( n11102, n11103, n11104 );
nor U10281 ( n11101, n11105, n11106 );
nor U10282 ( n11099, n11107, n11108 );
nor U10283 ( n11108, n11109, n11110 );
nor U10284 ( n11107, n11111, n11112 );
nand U10285 ( n11096, n19589, n11113 );
nand U10286 ( n11113, n11114, n11115 );
nor U10287 ( n11115, n11116, n11117 );
nor U10288 ( n11117, n11118, n11103 );
nor U10289 ( n11116, n11119, n11106 );
nand U10290 ( n11106, n11120, n10223 );
nor U10291 ( n11114, n11121, n11122 );
nor U10292 ( n11122, n11123, n11109 );
nor U10293 ( n11121, n11124, n11111 );
nand U10294 ( g34201, n11125, n11054 );
nor U10295 ( n11125, new_g34781_, n11126 );
nor U10296 ( n11126, n11127, n11128 );
nand U10297 ( n11128, n11129, n11130 );
nor U10298 ( n11130, n11131, n11132 );
nor U10299 ( n11129, n11133, n11134 );
nand U10300 ( n11127, n11135, n11136 );
nor U10301 ( n11136, n11137, n11138 );
nor U10302 ( n11135, n11139, n11140 );
nand U10303 ( new_g34781_, n11141, n11142 );
nor U10304 ( n11142, n11143, n11144 );
nand U10305 ( n11144, n11145, n11146 );
nand U10306 ( n11146, n11147, n20167 );
nor U10307 ( n11147, n20165, n11148 );
nand U10308 ( n11145, n11149, n20153 );
nor U10309 ( n11149, n20151, n11150 );
nand U10310 ( n11143, n11151, n11152 );
nand U10311 ( n11152, n11153, n20193 );
nor U10312 ( n11153, n20191, n11154 );
nand U10313 ( n11151, n11155, n20180 );
nor U10314 ( n11155, n20178, n11156 );
nor U10315 ( n11141, n11157, n11158 );
nand U10316 ( n11158, n11159, n11160 );
nand U10317 ( n11160, n11161, n20112 );
nor U10318 ( n11161, n20110, n11162 );
nand U10319 ( n11159, g25167, n11137 );
nand U10320 ( n11157, n11163, n11164 );
nand U10321 ( n11164, n11165, n20138 );
nor U10322 ( n11165, n20136, n11166 );
nand U10323 ( n11163, n11167, n20125 );
nor U10324 ( n11167, n20123, n11168 );
nand U10325 ( g34221, n11094, n11169 );
not U10326 ( n11169, new_g34783_ );
nand U10327 ( new_g34783_, n11170, n11171 );
nand U10328 ( n11171, n11172, n11173 );
nor U10329 ( n11172, n11174, n11175 );
nand U10330 ( n11170, n11176, n11177 );
nor U10331 ( n11176, n11178, n11179 );
and U10332 ( n11094, n11054, n11180 );
nand U10333 ( n11180, n11174, n11178 );
nand U10334 ( g33935, n11181, n11182 );
nor U10335 ( n11182, n19103, n19104 );
nor U10336 ( n11181, new_g34649_, n11183 );
nand U10337 ( g33636, n11184, n11185 );
nor U10338 ( n11185, n19105, n19106 );
nor U10339 ( n11184, new_g34657_, n11183 );
nand U10340 ( g33659, n11186, n11054 );
nor U10341 ( n11054, n19566, n11183 );
nor U10342 ( n11186, new_g34663_, n11187 );
nor U10343 ( new_g34663_, n11187, n11188 );
and U10344 ( n11188, n11189, n11190 );
nor U10345 ( n11190, n11191, n11192 );
nor U10346 ( n11192, n10293, n11193 );
nand U10347 ( n11193, n11194, n11195 );
nor U10348 ( n11191, n19939, n11196 );
nor U10349 ( n11196, n11197, n11198 );
nor U10350 ( n11198, n11199, n11200 );
nor U10351 ( n11197, n11201, n11202 );
nor U10352 ( n11189, n11203, n11204 );
nor U10353 ( n11204, n19938, n11205 );
nand U10354 ( n11205, n11206, n11207 );
nand U10355 ( n11207, n11208, n10232 );
nand U10356 ( n11208, n11209, n11210 );
nand U10357 ( n11210, n19939, n11211 );
nand U10358 ( n11209, n11212, n10293 );
nand U10359 ( n11206, n11213, n19937 );
nand U10360 ( n11213, n11214, n11215 );
nand U10361 ( n11215, n19939, n11216 );
nand U10362 ( n11214, n11217, n10293 );
nor U10363 ( n11203, n11218, n11219 );
nand U10364 ( g33874, n11220, n11221 );
nor U10365 ( n11220, g29218, n19570 );
nor U10366 ( g33894, n19976, n11222 );
nor U10367 ( n11222, n19263, n11223 );
nand U10368 ( new_g25690_, n11224, n11225 );
nand U10369 ( n11225, n11007, n10311 );
nand U10370 ( n11224, n11227, g35 );
nor U10371 ( n11227, n10701, n19107 );
nor U10372 ( new_g25688_, n19109, n10980 );
nand U10373 ( g31656, g113, n10364 );
nand U10374 ( g31665, g113, n10507 );
nor U10375 ( g31521, n11228, n11229 );
nand U10376 ( n11229, n19932, n19933 );
nand U10377 ( n11228, n19347, n11230 );
nand U10378 ( n11230, n11231, n11232 );
nand U10379 ( n11232, n11233, n11234 );
nor U10380 ( n11233, n19344, n19936 );
nor U10381 ( g33435, n11235, n11236 );
nand U10382 ( n11236, n11237, n11238 );
nand U10383 ( n11238, n11239, n10332 );
nor U10384 ( n11239, n20200, n20207 );
nand U10385 ( n11237, n11240, n20201 );
nand U10386 ( n11240, n11241, n11242 );
nand U10387 ( n11242, n10560, n10228 );
nand U10388 ( n11241, n20200, n10369 );
nor U10389 ( n11235, n20208, n11243 );
nor U10390 ( g33079, n11244, n11245 );
nand U10391 ( n11245, n11246, n11247 );
nand U10392 ( n11247, n11248, n10332 );
nor U10393 ( n11248, n20200, n20211 );
nand U10394 ( n11246, n11249, n20201 );
nand U10395 ( n11249, n11250, n11251 );
nand U10396 ( n11251, n10559, n10228 );
nand U10397 ( n11250, n20200, n10358 );
nor U10398 ( n11244, n20212, n11243 );
not U10399 ( n11243, n11252 );
nor U10400 ( new_g24298_, n19580, g35 );
nand U10401 ( new_g24266_, n11253, n11254 );
nand U10402 ( n11254, n10997, n10476 );
nand U10403 ( n11253, n11255, g35 );
nor U10404 ( n11255, n10922, n19108 );
nor U10405 ( g21727, n19110, g35 );
nor U10406 ( new_g18597_, n20233, g35 );
nor U10407 ( g23190, new_g10520_, n10588 );
nand U10408 ( n999, n11256, n11257 );
nand U10409 ( n11257, n11258, g35 );
nor U10410 ( n11258, n11259, n11260 );
nand U10411 ( n11256, n11261, g4564 );
nand U10412 ( n11261, g35, n11262 );
nand U10413 ( n11262, n11263, n11264 );
nor U10414 ( n11264, n19112, n19113 );
nor U10415 ( n11263, n19574, n11259 );
and U10416 ( n11259, n11265, n19114 );
nor U10417 ( n11265, n11266, n10636 );
nand U10418 ( n994, n11267, n11268 );
or U10419 ( n11267, g35, n19112 );
nand U10420 ( n989, n11269, n11270 );
or U10421 ( n11269, g35, n19113 );
nand U10422 ( n984, n11271, n11272 );
or U10423 ( n11271, g35, n19574 );
nand U10424 ( n970, n11273, n11274 );
nand U10425 ( n11274, n11275, n10940 );
or U10426 ( n11275, n11276, n11024 );
nand U10427 ( n11273, n11277, n11276 );
nand U10428 ( n11276, n11278, n19116 );
nand U10429 ( n965, n11279, n11280 );
nor U10430 ( n11279, n11281, n11282 );
nor U10431 ( n11282, n19115, n11277 );
nand U10432 ( n960, n11283, n11284 );
nand U10433 ( n11284, n11285, g4546 );
nor U10434 ( n11283, n11286, n11287 );
nand U10435 ( n955, n11288, n11289 );
nand U10436 ( n11289, n11285, g4567 );
nor U10437 ( n11288, n11286, n11290 );
nand U10438 ( n950, n11291, n11292 );
nand U10439 ( n11292, n11285, g4543 );
nor U10440 ( n11291, n11293, n11287 );
nand U10441 ( n945, n11294, n11295 );
nand U10442 ( n11295, n11285, g4540 );
nor U10443 ( n11294, n11293, n11290 );
not U10444 ( n11290, n11280 );
nand U10445 ( n11280, n11277, g4578 );
nand U10446 ( n940, n11296, n11297 );
nor U10447 ( n11296, n11287, n11298 );
nor U10448 ( n11298, n19512, g35 );
nor U10449 ( n11287, n11285, n19116 );
nand U10450 ( n931, n11299, n11300 );
nand U10451 ( n11300, n11301, n11302 );
nand U10452 ( n11302, n11260, n11303 );
nor U10453 ( n11260, n10481, n11304 );
nand U10454 ( n11301, n11305, n11306 );
nand U10455 ( n11306, n11266, g35 );
not U10456 ( n11305, n11307 );
or U10457 ( n11299, g35, n19121 );
nand U10458 ( n926, n11308, n11268 );
nand U10459 ( n11268, g6750, g35 );
or U10460 ( n11308, g35, n19122 );
nand U10461 ( n921, n11309, n11270 );
nand U10462 ( n11270, g6749, g35 );
or U10463 ( n11309, g35, n19119 );
nand U10464 ( n916, n11310, n11272 );
nand U10465 ( n11272, g6748, g35 );
or U10466 ( n11310, g35, n19120 );
nand U10467 ( n902, n11311, n11312 );
nand U10468 ( n11312, n11307, n11313 );
nand U10469 ( n11313, n11278, n19442 );
nor U10470 ( n11278, n19125, n11304 );
nand U10471 ( n11307, n11285, n11314 );
nand U10472 ( n11314, g35, n10869 );
nand U10473 ( n11311, n11002, n10835 );
nand U10474 ( n897, n11315, n11316 );
or U10475 ( n11316, g35, n19118 );
nand U10476 ( n11315, n11317, g35 );
nand U10477 ( n11317, n11318, n11319 );
nand U10478 ( n11319, n10835, n10284 );
or U10479 ( n11318, n10284, n11320 );
nand U10480 ( n892, n11321, n11322 );
nand U10481 ( n11322, n11323, n10284 );
nand U10482 ( n11323, g35, n11320 );
xnor U10483 ( n11320, n11303, n19118 );
nand U10484 ( n11303, n11324, n11325 );
nor U10485 ( n11325, n19119, n19120 );
nor U10486 ( n11324, n19121, n19122 );
nand U10487 ( n11321, n11326, n19117 );
nor U10488 ( n11326, n10972, n11327 );
nand U10489 ( n887, n11328, n11329 );
nand U10490 ( n11329, n10997, n10869 );
nand U10491 ( n11328, g35, n11330 );
nand U10492 ( n11330, g4531, n10636 );
nand U10493 ( n882, n11331, n11332 );
not U10494 ( n11332, n11333 );
nor U10495 ( n11331, n11281, n11334 );
nor U10496 ( n11334, n19123, n11277 );
nor U10497 ( n11281, n11266, n11285 );
nand U10498 ( n877, n11335, n11336 );
nand U10499 ( n11336, n11285, g4501 );
nor U10500 ( n11335, n11286, n11337 );
nand U10501 ( n872, n11338, n11339 );
nand U10502 ( n11339, n11285, g4498 );
nor U10503 ( n11338, n11286, n11333 );
and U10504 ( n11286, n11277, n11340 );
nand U10505 ( n11340, n19563, g72 );
nand U10506 ( n867, n11341, n11342 );
nand U10507 ( n11342, n11285, g4495 );
nor U10508 ( n11341, n11293, n11337 );
nand U10509 ( n862, n11343, n11344 );
nand U10510 ( n11344, n11285, g4480 );
nor U10511 ( n11343, n11293, n11333 );
nor U10512 ( n11333, n11285, n19453 );
and U10513 ( n11293, n11277, n11345 );
nand U10514 ( n11345, n19562, g73 );
nand U10515 ( n857, n11346, n11297 );
and U10516 ( n11297, n11347, n11348 );
nand U10517 ( n11348, n11349, n19125 );
nor U10518 ( n11349, n19124, n10980 );
nand U10519 ( n11347, n11277, n11350 );
nand U10520 ( n11350, g72, g73 );
nor U10521 ( n11346, n11337, n11351 );
nor U10522 ( n11351, n19128, g35 );
nor U10523 ( n11337, n11285, n19442 );
not U10524 ( n11285, n11277 );
nor U10525 ( n11277, n10972, n19125 );
nand U10526 ( n842, n11352, n11353 );
nor U10527 ( n11353, n11354, n11355 );
nor U10528 ( n11355, n19126, n19572 );
nor U10529 ( n11352, n10971, n10259 );
nand U10530 ( n837, n11356, n11357 );
nand U10531 ( n11357, n10998, n10259 );
nand U10532 ( n11356, n11358, g35 );
nor U10533 ( n11358, n10254, g4467 );
nand U10534 ( n832, n11359, n11360 );
nand U10535 ( n11360, n11361, n10254 );
nand U10536 ( n11361, n11362, n11363 );
nor U10537 ( n11363, n19573, n19586 );
nor U10538 ( n11362, n10971, g4467 );
nand U10539 ( n11359, n11354, g35 );
nand U10540 ( n827, n11364, n11365 );
or U10541 ( n11365, g35, n19571 );
nand U10542 ( n11364, g35, n11366 );
nand U10543 ( n11366, n11367, n19129 );
nor U10544 ( n11367, n11354, n11368 );
nor U10545 ( n11368, n19572, n10259 );
nand U10546 ( n822, n11369, n11370 );
nand U10547 ( n11370, g35, n10254 );
or U10548 ( n11369, g35, n19129 );
nor U10549 ( n817, n11371, n10980 );
nor U10550 ( n11371, n11354, n11372 );
nand U10551 ( n11372, n10259, g4467 );
and U10552 ( n11354, n11373, n19128 );
nor U10553 ( n11373, n19127, n11374 );
nor U10554 ( n11374, n11375, n11304 );
and U10555 ( n11375, n11221, n19570 );
nand U10556 ( n812, n11376, g35 );
nor U10557 ( n11376, n11377, n11378 );
nor U10558 ( n11378, n19570, n11379 );
not U10559 ( n11379, n11380 );
nor U10560 ( n11377, n19566, n11380 );
nand U10561 ( n11380, n19129, n10254 );
nand U10562 ( n7613, n11381, n11382 );
or U10563 ( n11382, g35, n20232 );
nand U10564 ( n11381, g35, n11383 );
nand U10565 ( n11383, n11384, n20233 );
nor U10566 ( n11384, n19523, n20070 );
nand U10567 ( n7608, n11385, n11386 );
nand U10568 ( n11386, n10998, n10281 );
nand U10569 ( n11385, g35, n11387 );
nand U10570 ( n11387, n11388, n20232 );
and U10571 ( n11388, g91, n11389 );
nand U10572 ( n7603, n11390, n11391 );
nand U10573 ( n11391, n10998, n10705 );
nand U10574 ( n11390, g35, n11392 );
nand U10575 ( n11392, n11393, n11394 );
nor U10576 ( n11394, n11395, n11396 );
nand U10577 ( n11396, n11397, n11398 );
not U10578 ( n11397, n11399 );
nand U10579 ( n11395, n11400, n11401 );
nor U10580 ( n11393, n11402, n11403 );
nand U10581 ( n11403, n19310, n19465 );
or U10582 ( n11402, n11404, n11405 );
nand U10583 ( n7598, n11406, n11407 );
nand U10584 ( n11407, n10998, n10677 );
nand U10585 ( n11406, g35, n11408 );
nand U10586 ( n11408, n11409, n19341 );
and U10587 ( n11409, n20231, n19345 );
nand U10588 ( n7593, n11410, n11411 );
nand U10589 ( n11411, n10998, n10665 );
nand U10590 ( n11410, g35, n11412 );
nand U10591 ( n11412, n11413, n19581 );
nor U10592 ( n11413, n19568, n10677 );
nand U10593 ( n7588, n11414, n11415 );
nand U10594 ( n11415, n10998, n10700 );
nand U10595 ( n11414, g35, n11416 );
nand U10596 ( n11416, n11417, n20229 );
and U10597 ( n11417, n11418, n11419 );
nand U10598 ( n7583, n11420, n11421 );
nand U10599 ( n11421, n10998, n10671 );
nand U10600 ( n11420, g35, n11422 );
nand U10601 ( n11422, n11423, n19262 );
and U10602 ( n11423, n11424, n20228 );
nand U10603 ( n7578, n11425, n11426 );
nand U10604 ( n11426, g35, n10671 );
nand U10605 ( n11425, n10998, n10672 );
nand U10606 ( n7573, n11427, n11428 );
nand U10607 ( n11428, g35, n10672 );
nand U10608 ( n11427, n10998, n10562 );
nand U10609 ( n7568, n11429, n11430 );
nand U10610 ( n11430, g35, n10562 );
nand U10611 ( n11429, n10998, n10673 );
nand U10612 ( n7563, n11431, n11432 );
nand U10613 ( n11432, g35, n10673 );
nand U10614 ( n11431, n10999, n10674 );
nand U10615 ( n7558, n11433, n11434 );
nand U10616 ( n11434, g35, n10674 );
nand U10617 ( n11433, n10999, n10509 );
nand U10618 ( n7553, n11435, n11436 );
nand U10619 ( n11436, g35, n10509 );
nand U10620 ( n11435, n10999, n10508 );
nand U10621 ( n7548, n11437, n11438 );
nand U10622 ( n11438, g35, n10508 );
nand U10623 ( n11437, n10999, n10769 );
nand U10624 ( n7543, n11439, n11440 );
nand U10625 ( n11440, n10999, n10772 );
nand U10626 ( n11439, g35, n11441 );
nand U10627 ( n11441, n19322, n11442 );
nand U10628 ( n11442, n11443, n11444 );
and U10629 ( n11444, n19569, n19492 );
nor U10630 ( n11443, g54, n11052 );
nand U10631 ( n7538, n11445, n11446 );
or U10632 ( n11446, g35, n19331 );
nand U10633 ( n11445, g35, n11447 );
nand U10634 ( n11447, n19329, n19493 );
nand U10635 ( n7533, n11448, n11449 );
or U10636 ( n11449, g35, n19338 );
nand U10637 ( n11448, g35, n11450 );
nand U10638 ( n11450, n19331, n19310 );
nand U10639 ( n7528, n11451, n11452 );
or U10640 ( n11452, g35, n20220 );
nand U10641 ( n11451, g35, n11453 );
nand U10642 ( n11453, n19338, g91 );
nand U10643 ( n7523, n11454, n11455 );
nand U10644 ( n11455, n10999, n10771 );
nand U10645 ( n11454, g35, n11456 );
nand U10646 ( n11456, n20220, n11389 );
nor U10647 ( n11389, n11457, n11458 );
nand U10648 ( n7518, n11459, n11460 );
nand U10649 ( n11460, n10999, n10770 );
nand U10650 ( n11459, g35, n11461 );
nand U10651 ( n11461, n19469, n11398 );
and U10652 ( n11398, n11462, n11463 );
nor U10653 ( n11463, n11464, n11465 );
nand U10654 ( n11465, n11466, n11467 );
nor U10655 ( n11462, n11468, n11469 );
nand U10656 ( n7513, n11470, n11471 );
nand U10657 ( n11471, n10999, n10783 );
nand U10658 ( n11470, g35, n11472 );
nand U10659 ( n11472, n19478, n11400 );
and U10660 ( n11400, n11473, n11474 );
nor U10661 ( n11473, n11475, n11476 );
nand U10662 ( n7508, n11477, n11478 );
nand U10663 ( n11478, n10999, n10782 );
nand U10664 ( n11477, g35, n11479 );
nand U10665 ( n11479, n11480, n19484 );
nor U10666 ( n11480, n11399, n11405 );
nand U10667 ( n7503, n11481, n11482 );
nand U10668 ( n11482, n10999, g20652 );
nand U10669 ( n11481, g35, n11483 );
nand U10670 ( n11483, n11484, n20219 );
nor U10671 ( n11484, n11485, n11404 );
nand U10672 ( n7498, n11486, n11487 );
nand U10673 ( n11487, g35, g20652 );
nand U10674 ( n11486, n10999, n10386 );
nand U10675 ( n7493, n11488, n11489 );
nand U10676 ( n11489, g35, n10386 );
nand U10677 ( n11488, n10999, n10542 );
nand U10678 ( n7488, n11490, n11491 );
nand U10679 ( n11491, g35, n10542 );
nand U10680 ( n11490, n11000, n10541 );
nand U10681 ( n7483, n11492, n11493 );
nand U10682 ( n11493, g35, n10541 );
nand U10683 ( n11492, n11000, n10540 );
nand U10684 ( n7478, n11494, n11495 );
nand U10685 ( n11495, g35, n10540 );
nand U10686 ( n11494, n11000, n10539 );
nand U10687 ( n7473, n11496, n11497 );
nand U10688 ( n11497, g35, n10539 );
or U10689 ( n11496, g35, n19321 );
nand U10690 ( n7468, n11498, n11499 );
nand U10691 ( n11499, n11000, n10364 );
nand U10692 ( n11498, g35, n11500 );
nand U10693 ( n11500, n19321, g44 );
nand U10694 ( n7463, n11501, n11502 );
nand U10695 ( n11502, g35, n10364 );
nand U10696 ( n11501, n11000, n10507 );
nand U10697 ( n7458, n11503, n11504 );
nand U10698 ( n11504, g35, n10507 );
nand U10699 ( n11503, n11000, n10481 );
nand U10700 ( n7453, n11505, n11506 );
nand U10701 ( n11506, g35, n10481 );
nand U10702 ( n11505, n11000, n10517 );
nand U10703 ( n7448, n11507, n11508 );
nand U10704 ( n11508, g35, n10517 );
nand U10705 ( n11507, n11000, n10833 );
nor U10706 ( n7443, n11509, n10981 );
and U10707 ( n11509, n19581, n20215 );
nand U10708 ( n7438, n11510, n11511 );
or U10709 ( n11511, g35, g30330 );
nand U10710 ( n7433, n11510, n11512 );
nand U10711 ( n11512, n11000, n10358 );
nand U10712 ( n11510, n11513, g35 );
nand U10713 ( n11513, n11514, n11515 );
nand U10714 ( n11515, n11516, n11517 );
nor U10715 ( n11516, n11518, n11519 );
nand U10716 ( n11519, n11520, n11521 );
nand U10717 ( n11521, n19153, n11522 );
nand U10718 ( n11520, n19161, n11523 );
nand U10719 ( n11518, n11524, n11525 );
nand U10720 ( n11525, n11526, n20154 );
nand U10721 ( n11524, n19145, n11527 );
nand U10722 ( n11514, n11528, n11529 );
nor U10723 ( n11528, n11530, n11531 );
nand U10724 ( n11531, n11532, n11533 );
nand U10725 ( n11533, n11534, n20199 );
nor U10726 ( n11534, n11535, n11536 );
nor U10727 ( n11536, n10358, n10225 );
nor U10728 ( n11535, n20198, n10559 );
nand U10729 ( n11532, n11527, n10634 );
nor U10730 ( n11530, n20212, n11537 );
nand U10731 ( n7428, n11538, n11539 );
nand U10732 ( n11539, n11000, n10559 );
nor U10733 ( n11538, n11540, n11541 );
nor U10734 ( n11541, n20214, n11542 );
nor U10735 ( n11540, n11543, n11544 );
nor U10736 ( n11543, n11545, n11546 );
nor U10737 ( n11545, n11547, n10818 );
nand U10738 ( n7423, n11548, n11549 );
or U10739 ( n11549, g35, n20212 );
nor U10740 ( n11548, n11550, n11551 );
nor U10741 ( n11551, n20213, n11552 );
nor U10742 ( n11550, n11553, n11554 );
nor U10743 ( n11553, n11555, n11546 );
nor U10744 ( n11555, n11547, n10817 );
nand U10745 ( n7418, n11556, n11557 );
nand U10746 ( n11557, n11000, n10634 );
nor U10747 ( n11556, n11558, n11559 );
nor U10748 ( n11559, n20212, n11560 );
nor U10749 ( n11558, n11561, n11562 );
nor U10750 ( n11561, n11563, n11546 );
nor U10751 ( n11563, n11547, n10816 );
nand U10752 ( n7413, n11564, n11565 );
nand U10753 ( n11565, n11000, n10815 );
nor U10754 ( n11564, n11566, n11567 );
nor U10755 ( n11567, n20211, n11568 );
nor U10756 ( n11566, n11569, n11570 );
nor U10757 ( n11569, n11571, n11546 );
and U10758 ( n11546, n19130, n11572 );
nor U10759 ( n11571, n11547, n10815 );
nand U10760 ( n7408, n11573, n11574 );
nand U10761 ( n11574, n11001, n10816 );
nor U10762 ( n11573, n11575, n11576 );
nor U10763 ( n11576, n19131, n11577 );
nor U10764 ( n11575, n11578, n10823 );
nand U10765 ( n7403, n11579, n11580 );
nand U10766 ( n11580, n11001, n10817 );
nor U10767 ( n11579, n11581, n11582 );
nor U10768 ( n11582, n19132, n11577 );
nor U10769 ( n11581, n11578, n10824 );
nand U10770 ( n7398, n11583, n11584 );
nand U10771 ( n11584, n11001, n10818 );
nor U10772 ( n11583, n11585, n11586 );
nor U10773 ( n11586, n19133, n11577 );
nor U10774 ( n11585, n11578, n10825 );
nand U10775 ( n7393, n11587, n11588 );
nand U10776 ( n11588, n11001, g20654 );
nor U10777 ( n11587, n11589, n11590 );
nor U10778 ( n11590, n19134, n11577 );
nor U10779 ( n11589, n11578, n10826 );
nand U10780 ( n7388, n11591, n11592 );
or U10781 ( n11592, g35, g30331 );
nand U10782 ( n7383, n11591, n11593 );
nand U10783 ( n11593, n11001, n10369 );
nand U10784 ( n11591, n11594, g35 );
nand U10785 ( n11594, n11595, n11596 );
nand U10786 ( n11596, n11597, n11517 );
nor U10787 ( n11597, n11598, n11599 );
nand U10788 ( n11599, n11600, n11601 );
nand U10789 ( n11601, n19184, n11522 );
nand U10790 ( n11600, n19192, n11523 );
nand U10791 ( n11598, n11602, n11603 );
nand U10792 ( n11603, n11526, n20099 );
nor U10793 ( n11526, n10225, n10420 );
nand U10794 ( n11602, n19176, n11527 );
nand U10795 ( n11595, n11604, n11529 );
not U10796 ( n11529, n11517 );
nand U10797 ( n11517, n11605, n20202 );
nor U10798 ( n11605, n11606, n11607 );
nor U10799 ( n11604, n11608, n11609 );
nand U10800 ( n11609, n11610, n11611 );
nand U10801 ( n11611, n11612, n20199 );
nor U10802 ( n11612, n11613, n11614 );
nor U10803 ( n11614, n10225, n10369 );
nor U10804 ( n11613, n20198, n10560 );
nand U10805 ( n11610, n11527, n10635 );
nor U10806 ( n11608, n20208, n11537 );
nand U10807 ( n7378, n11615, n11616 );
nand U10808 ( n11616, n11001, n10560 );
nor U10809 ( n11615, n11617, n11618 );
nor U10810 ( n11618, n20210, n11542 );
nand U10811 ( n11542, g35, n11544 );
nor U10812 ( n11617, n11619, n11544 );
nand U10813 ( n11544, n11620, n11621 );
nor U10814 ( n11619, n11622, n11623 );
nor U10815 ( n11622, n11547, n10822 );
nand U10816 ( n7373, n11624, n11625 );
or U10817 ( n11625, g35, n20208 );
nor U10818 ( n11624, n11626, n11627 );
nor U10819 ( n11627, n20209, n11552 );
nand U10820 ( n11552, g35, n11554 );
nor U10821 ( n11626, n11628, n11554 );
nand U10822 ( n11554, n11629, n20201 );
nor U10823 ( n11628, n11630, n11623 );
nor U10824 ( n11630, n11547, n10821 );
nand U10825 ( n7368, n11631, n11632 );
nand U10826 ( n11632, n11001, n10635 );
nor U10827 ( n11631, n11633, n11634 );
nor U10828 ( n11634, n20208, n11560 );
nand U10829 ( n11560, g35, n11562 );
nor U10830 ( n11633, n11635, n11562 );
nand U10831 ( n11562, n11620, n11252 );
nor U10832 ( n11252, n10228, n20201 );
nor U10833 ( n11635, n11636, n11623 );
nor U10834 ( n11636, n11547, n10820 );
nand U10835 ( n7363, n11637, n11638 );
nand U10836 ( n11638, n11001, n10819 );
nor U10837 ( n11637, n11639, n11640 );
nor U10838 ( n11640, n20207, n11568 );
nand U10839 ( n11568, g35, n11570 );
nor U10840 ( n11639, n11641, n11570 );
nand U10841 ( n11570, n11629, n10332 );
and U10842 ( n11629, n11620, n10228 );
nor U10843 ( n11641, n11642, n11623 );
and U10844 ( n11623, n19135, n11572 );
nor U10845 ( n11642, n11547, n10819 );
nand U10846 ( n7358, n11643, n11644 );
nand U10847 ( n11644, n11001, n10820 );
nor U10848 ( n11643, n11645, n11646 );
nor U10849 ( n11646, n19136, n11577 );
nor U10850 ( n11645, n11578, n10827 );
nand U10851 ( n7353, n11647, n11648 );
nand U10852 ( n11648, n11001, n10821 );
nor U10853 ( n11647, n11649, n11650 );
nor U10854 ( n11650, n19137, n11577 );
nor U10855 ( n11649, n11578, n10828 );
nand U10856 ( n7348, n11651, n11652 );
nand U10857 ( n11652, n11001, n10822 );
nor U10858 ( n11651, n11653, n11654 );
nor U10859 ( n11654, n19138, n11577 );
nor U10860 ( n11653, n11578, n10829 );
nand U10861 ( n7343, n11655, n11656 );
nand U10862 ( n11656, n11006, n10474 );
nor U10863 ( n11655, n11657, n11658 );
nor U10864 ( n11658, n19139, n11577 );
nor U10865 ( n11657, n11578, n10830 );
nand U10866 ( n11578, n11659, n11660 );
not U10867 ( n11660, n11577 );
nand U10868 ( n11577, g35, n11661 );
nand U10869 ( n11661, n11662, n20204 );
nor U10870 ( n11659, n11620, n11663 );
nor U10871 ( n11663, n10222, n10405 );
and U10872 ( n11620, n11664, n11665 );
nor U10873 ( n11665, n20202, n20203 );
nor U10874 ( n11664, n20204, n20205 );
nand U10875 ( n7338, n11666, n11667 );
nor U10876 ( n11667, n11668, n11669 );
nor U10877 ( n11669, n20206, g35 );
nor U10878 ( n11668, n10971, n11670 );
nand U10879 ( n11670, n11671, n10474 );
nor U10880 ( n11666, n11672, n11673 );
nor U10881 ( n11673, n10474, n11671 );
nand U10882 ( n11671, n11674, n10461 );
nand U10883 ( n7333, n11675, n11676 );
nor U10884 ( n11676, n11677, n11678 );
nor U10885 ( n11678, n20205, g35 );
nor U10886 ( n11677, n10971, n11679 );
nand U10887 ( n11679, n11680, n10461 );
nor U10888 ( n11675, n11672, n11681 );
nor U10889 ( n11681, n10461, n11680 );
not U10890 ( n11680, n11674 );
nor U10891 ( n11674, n11682, n20205 );
nand U10892 ( n7328, n11683, n11684 );
nor U10893 ( n11683, n11685, n11686 );
nor U10894 ( n11686, n10971, n11687 );
xnor U10895 ( n11687, n20205, n11682 );
nand U10896 ( n11682, n11688, n10222 );
nor U10897 ( n11685, n20204, g35 );
nand U10898 ( n7323, n11689, n11690 );
nand U10899 ( n11690, n11002, n10231 );
nor U10900 ( n11689, n11691, n11692 );
nor U10901 ( n11692, n10222, n11693 );
nand U10902 ( n11693, n11688, n10476 );
not U10903 ( n11688, n11694 );
nor U10904 ( n11691, n20204, n11695 );
nand U10905 ( n11695, n11696, n11694 );
nand U10906 ( n11694, n11697, n10231 );
nand U10907 ( n7318, n11698, n11699 );
nand U10908 ( n11699, n11700, n11696 );
xnor U10909 ( n11700, n11697, n20203 );
nor U10910 ( n11697, n11701, n20202 );
nand U10911 ( n11698, n11002, n10437 );
nand U10912 ( n7313, n11702, n11703 );
nor U10913 ( n11703, n11704, n11705 );
nor U10914 ( n11705, n20201, g35 );
nor U10915 ( n11704, n10971, n11706 );
nand U10916 ( n11706, n11701, n10437 );
nor U10917 ( n11702, n11672, n11707 );
nor U10918 ( n11707, n10437, n11701 );
or U10919 ( n11701, n11708, n20201 );
nand U10920 ( n7308, n11709, n11684 );
nor U10921 ( n11709, n11710, n11711 );
nor U10922 ( n11711, n10971, n11712 );
xnor U10923 ( n11712, n20201, n11708 );
nand U10924 ( n11708, n11527, n10228 );
nor U10925 ( n11710, n20200, g35 );
nand U10926 ( n7303, n11713, n11714 );
nand U10927 ( n11714, n11715, n11696 );
nor U10928 ( n11696, n10971, n19141 );
xnor U10929 ( n11715, n20200, n11527 );
nand U10930 ( n11713, n11002, n10420 );
nand U10931 ( n7298, n11716, n11717 );
nor U10932 ( n11717, n11718, n11719 );
nor U10933 ( n11719, n10971, n11537 );
not U10934 ( n11537, n11522 );
nor U10935 ( n11718, n20198, g35 );
nor U10936 ( n11716, n11523, n11672 );
nand U10937 ( n7293, n11720, n11684 );
not U10938 ( n11684, n11672 );
nor U10939 ( n11672, n10476, n10981 );
nor U10940 ( n11720, n11721, n11722 );
nor U10941 ( n11722, n19140, g35 );
nor U10942 ( n11721, n10970, n10225 );
nand U10943 ( n7263, n11723, n11724 );
nand U10944 ( n11724, g35, n10383 );
nand U10945 ( n11723, n11002, n10296 );
nand U10946 ( n7258, n11725, n11726 );
nand U10947 ( n11726, g35, n10296 );
nand U10948 ( n11725, n11003, n10238 );
nor U10949 ( n7253, n20196, n10982 );
nand U10950 ( n7248, n11727, n11728 );
or U10951 ( n11728, n11729, n19540 );
nor U10952 ( n11727, n11730, n11731 );
nor U10953 ( n11731, n10706, n11732 );
nand U10954 ( n11732, n11733, n19143 );
nor U10955 ( n11733, n10970, n11734 );
nor U10956 ( n11730, n19142, n11735 );
nor U10957 ( n11735, n11736, n10982 );
nor U10958 ( n11736, n19143, n11734 );
nand U10959 ( n7243, n11737, n11738 );
nand U10960 ( n11738, n11739, n10706 );
nand U10961 ( n11737, n11729, n10626 );
nand U10962 ( n7238, n11740, n11741 );
nand U10963 ( n11741, n11742, n10626 );
nor U10964 ( n11740, n11743, n11744 );
nor U10965 ( n11744, n19541, g35 );
nor U10966 ( n11743, n10970, n11745 );
nand U10967 ( n11745, n11746, n19143 );
nand U10968 ( n7233, n11747, n11748 );
or U10969 ( n11748, n11749, n19541 );
nor U10970 ( n11747, n11750, n11751 );
nor U10971 ( n11751, n10707, n11752 );
nand U10972 ( n11752, n11753, n20194 );
nor U10973 ( n11753, n10970, n11754 );
nor U10974 ( n11750, n20195, n11755 );
nor U10975 ( n11755, n11756, n10982 );
nor U10976 ( n11756, n20194, n11754 );
nand U10977 ( n7228, n11757, n11758 );
nand U10978 ( n11758, n11742, n10707 );
nand U10979 ( n11757, n11749, n10570 );
nand U10980 ( n7223, n11759, n11760 );
nand U10981 ( n11760, n11739, n10570 );
not U10982 ( n11739, n11729 );
nand U10983 ( n11729, g35, n11734 );
nor U10984 ( n11759, n11761, n11762 );
nor U10985 ( n11762, n19555, g35 );
nor U10986 ( n11761, n10970, n11763 );
or U10987 ( n11763, n10570, n11734 );
nand U10988 ( n7218, n11764, n11765 );
nand U10989 ( n11765, n11003, n10422 );
nand U10990 ( n11764, n11766, g35 );
nand U10991 ( n11766, n11767, n11768 );
or U10992 ( n11768, n11769, n19555 );
nand U10993 ( n11767, n11770, n11769 );
nor U10994 ( n11769, n11771, n11772 );
xnor U10995 ( n11770, n10422, n19148 );
nand U10996 ( n7213, n11773, n11774 );
nand U10997 ( n11774, n11775, g35 );
nor U10998 ( n11775, n19144, n11776 );
nor U10999 ( n11776, n11777, n11772 );
nor U11000 ( n11777, n11778, n10683 );
nand U11001 ( n11773, n11779, n10683 );
nand U11002 ( n11779, g35, n11780 );
nand U11003 ( n11780, n11781, n11782 );
nand U11004 ( n11782, n10422, n11771 );
nand U11005 ( n7208, n11783, n11784 );
nand U11006 ( n11784, n11003, n10408 );
nand U11007 ( n11783, g35, n11785 );
nand U11008 ( n11785, n11786, n11787 );
or U11009 ( n11787, n11734, n20186 );
nand U11010 ( n11734, n11788, n11781 );
nor U11011 ( n11788, n20190, n20193 );
nor U11012 ( n11786, n11789, n11790 );
nor U11013 ( n11790, n11791, n11772 );
nor U11014 ( n11791, n11792, n11793 );
nand U11015 ( n11793, n11794, n11795 );
nand U11016 ( n11795, n20193, n11796 );
nand U11017 ( n11796, n11797, n11798 );
or U11018 ( n11798, n20191, n20189 );
nand U11019 ( n11797, n20190, n10523 );
nand U11020 ( n11794, n20191, n11799 );
nand U11021 ( n11799, n11800, n11801 );
or U11022 ( n11801, n20193, n20188 );
or U11023 ( n11800, n20190, n19147 );
nor U11024 ( n11792, n20187, n11771 );
nor U11025 ( n11789, n19145, n11781 );
nand U11026 ( n7203, n11802, n11803 );
nor U11027 ( n11803, n11804, n11805 );
nor U11028 ( n11805, n10970, n11806 );
nand U11029 ( n11806, n11781, n10339 );
nor U11030 ( n11804, n20192, g35 );
nor U11031 ( n11802, n11807, n11808 );
nor U11032 ( n11808, n20193, n11809 );
nand U11033 ( n7198, n11810, n11811 );
nand U11034 ( n11811, n11003, n10339 );
nor U11035 ( n11810, n11812, n11813 );
nor U11036 ( n11813, n20192, n11814 );
nor U11037 ( n11814, n11815, n11816 );
nand U11038 ( n11816, n11809, n11547 );
nor U11039 ( n11815, n11134, n10982 );
nor U11040 ( n11812, n11817, n11818 );
nand U11041 ( n11817, n11819, n11820 );
nand U11042 ( n11820, n11821, n11822 );
nand U11043 ( n11819, n11823, n11824 );
not U11044 ( n11823, n11821 );
nor U11045 ( n11821, n10339, n20193 );
nand U11046 ( n7193, n11825, n11826 );
not U11047 ( n11826, n11807 );
nor U11048 ( n11825, n11827, n11828 );
nor U11049 ( n11828, n20190, n11829 );
nor U11050 ( n11827, n20191, n11809 );
nand U11051 ( n7188, n11830, n11831 );
nor U11052 ( n11831, n11832, n11833 );
nor U11053 ( n11833, n10970, n11834 );
nand U11054 ( n11834, n11835, n11781 );
nor U11055 ( n11835, n11778, n10408 );
not U11056 ( n11778, n11771 );
nand U11057 ( n11771, n20190, n10339 );
nor U11058 ( n11832, n19146, g35 );
nor U11059 ( n11830, n11807, n11836 );
nor U11060 ( n11836, n20190, n11809 );
not U11061 ( n11809, n11829 );
nor U11062 ( n11829, n10970, n11781 );
nor U11063 ( n11807, n11818, n11837 );
nand U11064 ( n11818, n11781, n11134 );
not U11065 ( n11134, n11154 );
nand U11066 ( n11154, n11838, n11839 );
nor U11067 ( n11838, n20203, n20204 );
nand U11068 ( n7183, n11840, n11841 );
nand U11069 ( n11841, n11004, n10523 );
nand U11070 ( n11840, n11842, g35 );
nand U11071 ( n11842, n11843, n11844 );
nand U11072 ( n11844, n11845, n10823 );
nand U11073 ( n11843, n11846, n11847 );
nand U11074 ( n11847, n19149, n10312 );
not U11075 ( n11846, n11845 );
nand U11076 ( n11845, n11848, n11781 );
not U11077 ( n11781, n11772 );
nand U11078 ( n11772, n11849, n11527 );
nor U11079 ( n11849, n11850, n11851 );
nor U11080 ( n11851, n20211, n11607 );
nor U11081 ( n11848, n20191, n10408 );
nand U11082 ( n7178, n11852, n11853 );
or U11083 ( n11853, n11854, n11855 );
nor U11084 ( n11852, n11856, n11857 );
nor U11085 ( n11857, n19147, g35 );
nor U11086 ( n11856, n10970, n11858 );
nand U11087 ( n11858, n11855, n10523 );
nand U11088 ( n11855, n11859, n10438 );
nand U11089 ( n7173, n11860, n11861 );
nand U11090 ( n11861, n11862, n11863 );
nor U11091 ( n11860, n11864, n11865 );
nor U11092 ( n11865, n20189, g35 );
nor U11093 ( n11864, n10970, n11866 );
or U11094 ( n11866, n11862, n19147 );
nor U11095 ( n11862, n11867, n10353 );
nand U11096 ( n7168, n11868, n11869 );
nand U11097 ( n11869, n11870, n11863 );
nor U11098 ( n11868, n11871, n11872 );
nor U11099 ( n11872, n20188, g35 );
nor U11100 ( n11871, n10970, n11873 );
or U11101 ( n11873, n11870, n20189 );
nor U11102 ( n11870, n11874, n11875 );
not U11103 ( n11874, n11089 );
nand U11104 ( n7163, n11876, n11877 );
nand U11105 ( n11877, n11878, n11863 );
nor U11106 ( n11876, n11879, n11880 );
nor U11107 ( n11880, n20187, g35 );
nor U11108 ( n11879, n10970, n11881 );
or U11109 ( n11881, n11878, n20188 );
nor U11110 ( n11878, n11867, n10438 );
nand U11111 ( n7158, n11882, n11883 );
nand U11112 ( n11883, n11884, n11863 );
not U11113 ( n11863, n11854 );
nor U11114 ( n11882, n11885, n11886 );
nor U11115 ( n11886, n20186, g35 );
nor U11116 ( n11885, n10969, n11887 );
or U11117 ( n11887, n11884, n20187 );
and U11118 ( n11884, n11859, n20184 );
nand U11119 ( n7153, n11888, n11889 );
nand U11120 ( n11889, n11004, n10751 );
nor U11121 ( n11888, n11890, n11891 );
nor U11122 ( n11891, n20186, n11749 );
nor U11123 ( n11890, n11754, n11854 );
nand U11124 ( n11854, n11892, g35 );
nor U11125 ( n11892, n11893, n11894 );
nor U11126 ( n11894, n11895, n11896 );
nor U11127 ( n11893, n20025, n11897 );
not U11128 ( n11754, n11746 );
nand U11129 ( n7148, n11898, n11899 );
nand U11130 ( n11899, n11742, n10751 );
nand U11131 ( n11898, n11749, n10524 );
not U11132 ( n11749, n11742 );
nor U11133 ( n11742, n10969, n11746 );
nor U11134 ( n11746, n11900, n11875 );
nand U11135 ( n7143, n11901, n11902 );
nand U11136 ( n11902, n11903, n10524 );
nor U11137 ( n11901, n11904, n11905 );
nor U11138 ( n11905, n10969, n11906 );
nand U11139 ( n11906, n11907, n11908 );
nand U11140 ( n11908, n11909, n11910 );
nor U11141 ( n11909, n11911, n11912 );
nor U11142 ( n11912, n11895, n11913 );
nor U11143 ( n11911, n11897, n10337 );
nor U11144 ( n11907, n11875, n11914 );
nor U11145 ( n11914, n11915, n11910 );
nand U11146 ( n11910, n11900, n10524 );
nand U11147 ( n11900, n19149, n20185 );
nand U11148 ( n11915, n11916, n11917 );
nand U11149 ( n11917, n11895, n10337 );
not U11150 ( n11895, n11897 );
nand U11151 ( n11916, n11913, n11897 );
not U11152 ( n11913, n11896 );
nand U11153 ( n11896, n11918, n11919 );
nor U11154 ( n11904, n20185, g35 );
nand U11155 ( n7138, n11920, n11921 );
nand U11156 ( n11921, n11004, n10312 );
nor U11157 ( n11920, n11922, n11923 );
nor U11158 ( n11923, n11924, n11867 );
or U11159 ( n11867, n20184, n11875 );
nor U11160 ( n11922, n20185, n11925 );
nand U11161 ( n7133, n11926, n11927 );
nand U11162 ( n11927, n11903, n10312 );
nor U11163 ( n11926, n11928, n11929 );
nor U11164 ( n11929, n10969, n11930 );
nand U11165 ( n11930, n11859, n11931 );
nor U11166 ( n11859, n19149, n11875 );
nor U11167 ( n11928, n20183, g35 );
nand U11168 ( n7128, n11932, n11933 );
nand U11169 ( n11933, n11004, n10353 );
nor U11170 ( n11932, n11934, n11935 );
nor U11171 ( n11935, n20183, n11936 );
nor U11172 ( n11936, n11937, n11938 );
nor U11173 ( n11937, n11939, n10983 );
nor U11174 ( n11939, n11940, n11941 );
nor U11175 ( n11934, n11942, n11943 );
nand U11176 ( n11943, n11944, n11945 );
xnor U11177 ( n11944, n11089, n19565 );
nor U11178 ( n11089, n10312, n20185 );
nand U11179 ( n11942, n11572, n11063 );
nand U11180 ( n7123, n11946, n11947 );
nand U11181 ( n11947, n11903, n10353 );
not U11182 ( n11903, n11925 );
nand U11183 ( n11925, n11875, g35 );
nand U11184 ( n11946, n11948, n11949 );
nor U11185 ( n11949, n11924, n11950 );
nor U11186 ( n11950, n11951, n10353 );
nor U11187 ( n11951, n11875, n10312 );
nor U11188 ( n11875, n11897, n11945 );
not U11189 ( n11945, n11941 );
nand U11190 ( n11941, n10590, n11952 );
nand U11191 ( n11952, n11953, n20031 );
nor U11192 ( n11953, n11954, n10303 );
nand U11193 ( n11897, n11955, n11919 );
nand U11194 ( n11919, n20050, n10622 );
nor U11195 ( n11955, n11956, n11957 );
nor U11196 ( n11957, n20197, n11958 );
not U11197 ( n11924, n11931 );
nand U11198 ( n11931, n11959, n11063 );
not U11199 ( n11063, n11940 );
nand U11200 ( n11940, n11960, n19996 );
nor U11201 ( n11960, n19997, n11961 );
nor U11202 ( n11948, n10969, n10438 );
nand U11203 ( n7118, n11962, n11963 );
or U11204 ( n11963, n11964, n19538 );
nor U11205 ( n11962, n11965, n11966 );
nor U11206 ( n11966, n10708, n11967 );
nand U11207 ( n11967, n11968, n19151 );
nor U11208 ( n11968, n10969, n11969 );
nor U11209 ( n11965, n19150, n11970 );
nor U11210 ( n11970, n11971, n10983 );
nor U11211 ( n11971, n19151, n11969 );
nand U11212 ( n7113, n11972, n11973 );
nand U11213 ( n11973, n11974, n10708 );
nand U11214 ( n11972, n11964, n10627 );
nand U11215 ( n7108, n11975, n11976 );
nand U11216 ( n11976, n11977, n10627 );
nor U11217 ( n11975, n11978, n11979 );
nor U11218 ( n11979, n19539, g35 );
nor U11219 ( n11978, n10969, n11980 );
nand U11220 ( n11980, n11981, n19151 );
nand U11221 ( n7103, n11982, n11983 );
or U11222 ( n11983, n11984, n19539 );
nor U11223 ( n11982, n11985, n11986 );
nor U11224 ( n11986, n10709, n11987 );
nand U11225 ( n11987, n11988, n20181 );
nor U11226 ( n11988, n10968, n11989 );
nor U11227 ( n11985, n20182, n11990 );
nor U11228 ( n11990, n11991, n10983 );
nor U11229 ( n11991, n20181, n11989 );
nand U11230 ( n7098, n11992, n11993 );
nand U11231 ( n11993, n11977, n10709 );
nand U11232 ( n11992, n11984, n10571 );
nand U11233 ( n7093, n11994, n11995 );
nand U11234 ( n11995, n11974, n10571 );
not U11235 ( n11974, n11964 );
nand U11236 ( n11964, g35, n11969 );
nor U11237 ( n11994, n11996, n11997 );
nor U11238 ( n11997, n19554, g35 );
nor U11239 ( n11996, n10968, n11998 );
or U11240 ( n11998, n10571, n11969 );
nand U11241 ( n7088, n11999, n12000 );
nand U11242 ( n12000, n11005, n10423 );
nand U11243 ( n11999, n12001, g35 );
nand U11244 ( n12001, n12002, n12003 );
or U11245 ( n12003, n12004, n19554 );
nand U11246 ( n12002, n12005, n12004 );
nor U11247 ( n12004, n12006, n12007 );
xnor U11248 ( n12005, n10423, n19156 );
nand U11249 ( n7083, n12008, n12009 );
nand U11250 ( n12009, n12010, g35 );
nor U11251 ( n12010, n19152, n12011 );
nor U11252 ( n12011, n12012, n12007 );
nor U11253 ( n12012, n12013, n10684 );
nand U11254 ( n12008, n12014, n10684 );
nand U11255 ( n12014, g35, n12015 );
nand U11256 ( n12015, n12016, n12017 );
nand U11257 ( n12017, n10423, n12006 );
nand U11258 ( n7078, n12018, n12019 );
nand U11259 ( n12019, n11005, n10409 );
nand U11260 ( n12018, g35, n12020 );
nand U11261 ( n12020, n12021, n12022 );
or U11262 ( n12022, n11969, n20173 );
nand U11263 ( n11969, n12023, n12016 );
nor U11264 ( n12023, n20177, n20180 );
nor U11265 ( n12021, n12024, n12025 );
nor U11266 ( n12025, n12026, n12007 );
nor U11267 ( n12026, n12027, n12028 );
nand U11268 ( n12028, n12029, n12030 );
nand U11269 ( n12030, n20180, n12031 );
nand U11270 ( n12031, n12032, n12033 );
or U11271 ( n12033, n20178, n20176 );
nand U11272 ( n12032, n20177, n10525 );
nand U11273 ( n12029, n20178, n12034 );
nand U11274 ( n12034, n12035, n12036 );
or U11275 ( n12036, n20180, n20175 );
or U11276 ( n12035, n20177, n19155 );
nor U11277 ( n12027, n20174, n12006 );
nor U11278 ( n12024, n19153, n12016 );
nand U11279 ( n7073, n12037, n12038 );
nor U11280 ( n12038, n12039, n12040 );
nor U11281 ( n12040, n10968, n12041 );
nand U11282 ( n12041, n12016, n10340 );
nor U11283 ( n12039, n20179, g35 );
nor U11284 ( n12037, n12042, n12043 );
nor U11285 ( n12043, n20180, n12044 );
nand U11286 ( n7068, n12045, n12046 );
nand U11287 ( n12046, n11005, n10340 );
nor U11288 ( n12045, n12047, n12048 );
nor U11289 ( n12048, n20179, n12049 );
nor U11290 ( n12049, n12050, n12051 );
nand U11291 ( n12051, n12044, n11547 );
nor U11292 ( n12050, n11133, n10984 );
nor U11293 ( n12047, n12052, n12053 );
nand U11294 ( n12053, n12016, n11133 );
not U11295 ( n11133, n11156 );
nand U11296 ( n12052, n12054, n12055 );
nand U11297 ( n12055, n12056, n11822 );
nand U11298 ( n12054, n12057, n11824 );
not U11299 ( n12057, n12056 );
nor U11300 ( n12056, n10340, n20180 );
nand U11301 ( n7063, n12058, n12059 );
nor U11302 ( n12058, n12060, n12061 );
nor U11303 ( n12061, n20177, n12062 );
nor U11304 ( n12060, n20178, n12044 );
nand U11305 ( n7058, n12063, n12064 );
nor U11306 ( n12064, n12065, n12066 );
nor U11307 ( n12066, n10968, n12067 );
nand U11308 ( n12067, n12068, n12016 );
nor U11309 ( n12068, n12013, n10409 );
not U11310 ( n12013, n12006 );
nand U11311 ( n12006, n20177, n10340 );
nor U11312 ( n12065, n19154, g35 );
nor U11313 ( n12063, n12042, n12069 );
nor U11314 ( n12069, n20177, n12044 );
not U11315 ( n12044, n12062 );
nor U11316 ( n12062, n10968, n12016 );
not U11317 ( n12042, n12059 );
nand U11318 ( n12059, n12070, n12016 );
nor U11319 ( n12070, n11156, n11837 );
nand U11320 ( n11156, n12071, n20203 );
nor U11321 ( n12071, n20204, n12072 );
nand U11322 ( n7053, n12073, n12074 );
nand U11323 ( n12074, n11005, n10525 );
nand U11324 ( n12073, n12075, g35 );
nand U11325 ( n12075, n12076, n12077 );
nand U11326 ( n12077, n12078, n10824 );
nand U11327 ( n12076, n12079, n12080 );
nand U11328 ( n12080, n19157, n10313 );
not U11329 ( n12079, n12078 );
nand U11330 ( n12078, n12081, n12016 );
not U11331 ( n12016, n12007 );
nand U11332 ( n12007, n12082, n11522 );
nor U11333 ( n12082, n11850, n12083 );
nor U11334 ( n12083, n20212, n11607 );
nor U11335 ( n12081, n20178, n10409 );
nand U11336 ( n7048, n12084, n12085 );
or U11337 ( n12085, n12086, n12087 );
nor U11338 ( n12084, n12088, n12089 );
nor U11339 ( n12089, n19155, g35 );
nor U11340 ( n12088, n10968, n12090 );
nand U11341 ( n12090, n12087, n10525 );
nand U11342 ( n12087, n12091, n10439 );
nand U11343 ( n7043, n12092, n12093 );
nand U11344 ( n12093, n12094, n12095 );
nor U11345 ( n12092, n12096, n12097 );
nor U11346 ( n12097, n20176, g35 );
nor U11347 ( n12096, n10968, n12098 );
or U11348 ( n12098, n12094, n19155 );
nor U11349 ( n12094, n12099, n10354 );
nand U11350 ( n7038, n12100, n12101 );
nand U11351 ( n12101, n12102, n12095 );
nor U11352 ( n12100, n12103, n12104 );
nor U11353 ( n12104, n20175, g35 );
nor U11354 ( n12103, n10968, n12105 );
or U11355 ( n12105, n12102, n20176 );
nor U11356 ( n12102, n12106, n12107 );
not U11357 ( n12106, n11093 );
nand U11358 ( n7033, n12108, n12109 );
nand U11359 ( n12109, n12110, n12095 );
nor U11360 ( n12108, n12111, n12112 );
nor U11361 ( n12112, n20174, g35 );
nor U11362 ( n12111, n10967, n12113 );
or U11363 ( n12113, n12110, n20175 );
nor U11364 ( n12110, n12099, n10439 );
nand U11365 ( n7028, n12114, n12115 );
nand U11366 ( n12115, n12116, n12095 );
not U11367 ( n12095, n12086 );
nor U11368 ( n12114, n12117, n12118 );
nor U11369 ( n12118, n20173, g35 );
nor U11370 ( n12117, n10967, n12119 );
or U11371 ( n12119, n12116, n20174 );
and U11372 ( n12116, n12091, n20171 );
nand U11373 ( n7023, n12120, n12121 );
nand U11374 ( n12121, n11005, n10752 );
nor U11375 ( n12120, n12122, n12123 );
nor U11376 ( n12123, n20173, n11984 );
nor U11377 ( n12122, n11989, n12086 );
nand U11378 ( n12086, n12124, g35 );
nor U11379 ( n12124, n12125, n12126 );
nor U11380 ( n12126, n12127, n10473 );
nor U11381 ( n12125, n12128, n12129 );
not U11382 ( n11989, n11981 );
nand U11383 ( n7018, n12130, n12131 );
nand U11384 ( n12131, n11977, n10752 );
nand U11385 ( n12130, n11984, n10526 );
not U11386 ( n11984, n11977 );
nor U11387 ( n11977, n10967, n11981 );
nor U11388 ( n11981, n12132, n12107 );
nand U11389 ( n7013, n12133, n12134 );
nand U11390 ( n12134, n12135, n10526 );
nor U11391 ( n12133, n12136, n12137 );
nor U11392 ( n12137, n10967, n12138 );
nand U11393 ( n12138, n12139, n12140 );
nand U11394 ( n12140, n12141, n12142 );
nor U11395 ( n12141, n12143, n12144 );
nor U11396 ( n12144, n12128, n12145 );
nor U11397 ( n12143, n20026, n12127 );
nor U11398 ( n12139, n12107, n12146 );
nor U11399 ( n12146, n12147, n12142 );
nand U11400 ( n12142, n12132, n10526 );
nand U11401 ( n12132, n19157, n20172 );
nand U11402 ( n12147, n12148, n12149 );
nand U11403 ( n12149, n12145, n12127 );
not U11404 ( n12145, n12129 );
nand U11405 ( n12129, n11918, n12150 );
nand U11406 ( n12148, n12128, n20026 );
not U11407 ( n12128, n12127 );
nor U11408 ( n12136, n20172, g35 );
nand U11409 ( n7008, n12151, n12152 );
nand U11410 ( n12152, n11006, n10313 );
nor U11411 ( n12151, n12153, n12154 );
nor U11412 ( n12154, n12155, n12099 );
or U11413 ( n12099, n20171, n12107 );
nor U11414 ( n12153, n20172, n12156 );
nand U11415 ( n7003, n12157, n12158 );
nand U11416 ( n12158, n12135, n10313 );
nor U11417 ( n12157, n12159, n12160 );
nor U11418 ( n12160, n10967, n12161 );
nand U11419 ( n12161, n12091, n12162 );
nor U11420 ( n12091, n19157, n12107 );
nor U11421 ( n12159, n20170, g35 );
nand U11422 ( n6998, n12163, n12164 );
nand U11423 ( n12164, n11006, n10354 );
nor U11424 ( n12163, n12165, n12166 );
nor U11425 ( n12166, n20170, n12167 );
nor U11426 ( n12167, n12168, n11938 );
nor U11427 ( n12168, n12169, n10984 );
nor U11428 ( n12169, n12170, n12171 );
nor U11429 ( n12165, n12172, n12173 );
nand U11430 ( n12173, n12174, n12175 );
xnor U11431 ( n12174, n11093, n19565 );
nor U11432 ( n11093, n10313, n20172 );
nand U11433 ( n12172, n11572, n11062 );
nand U11434 ( n6993, n12176, n12177 );
nand U11435 ( n12177, n12135, n10354 );
not U11436 ( n12135, n12156 );
nand U11437 ( n12156, n12107, g35 );
nand U11438 ( n12176, n12178, n12179 );
nor U11439 ( n12179, n12155, n12180 );
nor U11440 ( n12180, n12181, n10354 );
nor U11441 ( n12181, n12107, n10313 );
nor U11442 ( n12107, n12127, n12175 );
not U11443 ( n12175, n12171 );
nand U11444 ( n12171, g17423, n12182 );
nand U11445 ( n12182, n12183, n12184 );
not U11446 ( n12184, n11954 );
nor U11447 ( n12183, n20031, n20032 );
nand U11448 ( n12127, n12185, n12150 );
nand U11449 ( n12150, n20050, n10453 );
nor U11450 ( n12185, n11956, n12186 );
nor U11451 ( n12186, n10383, n11958 );
nand U11452 ( n11958, n10296, n10238 );
not U11453 ( n12155, n12162 );
nand U11454 ( n12162, n11959, n11062 );
not U11455 ( n11062, n12170 );
nand U11456 ( n12170, n12187, n12188 );
nor U11457 ( n12178, n10967, n10439 );
nand U11458 ( n6988, n12189, n12190 );
or U11459 ( n12190, n12191, n19544 );
nor U11460 ( n12189, n12192, n12193 );
nor U11461 ( n12193, n10710, n12194 );
nand U11462 ( n12194, n12195, n19159 );
nor U11463 ( n12195, n10967, n12196 );
nor U11464 ( n12192, n19158, n12197 );
nor U11465 ( n12197, n12198, n10984 );
nor U11466 ( n12198, n19159, n12196 );
nand U11467 ( n6983, n12199, n12200 );
nand U11468 ( n12200, n12201, n10710 );
nand U11469 ( n12199, n12191, n10628 );
nand U11470 ( n6978, n12202, n12203 );
nand U11471 ( n12203, n12204, n10628 );
nor U11472 ( n12202, n12205, n12206 );
nor U11473 ( n12206, n19545, g35 );
nor U11474 ( n12205, n10966, n12207 );
nand U11475 ( n12207, n12208, n19159 );
nand U11476 ( n6973, n12209, n12210 );
or U11477 ( n12210, n12211, n19545 );
nor U11478 ( n12209, n12212, n12213 );
nor U11479 ( n12213, n10711, n12214 );
nand U11480 ( n12214, n12215, n20168 );
nor U11481 ( n12215, n10966, n12216 );
nor U11482 ( n12212, n20169, n12217 );
nor U11483 ( n12217, n12218, n10984 );
nor U11484 ( n12218, n20168, n12216 );
nand U11485 ( n6968, n12219, n12220 );
nand U11486 ( n12220, n12204, n10711 );
nand U11487 ( n12219, n12211, n10572 );
nand U11488 ( n6963, n12221, n12222 );
nand U11489 ( n12222, n12201, n10572 );
not U11490 ( n12201, n12191 );
nand U11491 ( n12191, g35, n12196 );
nor U11492 ( n12221, n12223, n12224 );
nor U11493 ( n12224, n19557, g35 );
nor U11494 ( n12223, n10966, n12225 );
or U11495 ( n12225, n10572, n12196 );
nand U11496 ( n6958, n12226, n12227 );
nand U11497 ( n12227, n11006, n10424 );
nand U11498 ( n12226, n12228, g35 );
nand U11499 ( n12228, n12229, n12230 );
or U11500 ( n12230, n12231, n19557 );
nand U11501 ( n12229, n12232, n12231 );
nor U11502 ( n12231, n12233, n12234 );
xnor U11503 ( n12232, n10424, n19164 );
nand U11504 ( n6953, n12235, n12236 );
nand U11505 ( n12236, n12237, g35 );
nor U11506 ( n12237, n19160, n12238 );
nor U11507 ( n12238, n12239, n12234 );
nor U11508 ( n12239, n12240, n10685 );
nand U11509 ( n12235, n12241, n10685 );
nand U11510 ( n12241, g35, n12242 );
nand U11511 ( n12242, n12243, n12244 );
nand U11512 ( n12244, n10424, n12233 );
nand U11513 ( n6948, n12245, n12246 );
nand U11514 ( n12246, n11006, n10410 );
nand U11515 ( n12245, g35, n12247 );
nand U11516 ( n12247, n12248, n12249 );
or U11517 ( n12249, n12196, n20160 );
nand U11518 ( n12196, n12250, n12243 );
nor U11519 ( n12250, n20164, n20167 );
nor U11520 ( n12248, n12251, n12252 );
nor U11521 ( n12252, n12253, n12234 );
nor U11522 ( n12253, n12254, n12255 );
nand U11523 ( n12255, n12256, n12257 );
nand U11524 ( n12257, n20167, n12258 );
nand U11525 ( n12258, n12259, n12260 );
nand U11526 ( n12260, n10233, n10789 );
nand U11527 ( n12259, n20164, n10527 );
nand U11528 ( n12256, n20165, n12261 );
nand U11529 ( n12261, n12262, n12263 );
or U11530 ( n12263, n20167, n20162 );
or U11531 ( n12262, n20164, n19163 );
nor U11532 ( n12254, n20161, n12233 );
nor U11533 ( n12251, n19161, n12243 );
nand U11534 ( n6943, n12264, n12265 );
nor U11535 ( n12265, n12266, n12267 );
nor U11536 ( n12267, n10965, n12268 );
nand U11537 ( n12268, n12243, n10233 );
nor U11538 ( n12266, n20166, g35 );
nor U11539 ( n12264, n12269, n12270 );
nor U11540 ( n12270, n20167, n12271 );
nand U11541 ( n6938, n12272, n12273 );
nand U11542 ( n12273, n11006, n10233 );
nor U11543 ( n12272, n12274, n12275 );
nor U11544 ( n12275, n20166, n12276 );
nor U11545 ( n12276, n12277, n12278 );
nand U11546 ( n12278, n12271, n11547 );
nor U11547 ( n12277, n11132, n10984 );
nor U11548 ( n12274, n12279, n12280 );
nand U11549 ( n12280, n12243, n11132 );
not U11550 ( n11132, n11148 );
nand U11551 ( n12279, n12281, n12282 );
nand U11552 ( n12282, n12283, n11822 );
nand U11553 ( n12281, n12284, n11824 );
not U11554 ( n12284, n12283 );
nor U11555 ( n12283, n10233, n20167 );
nand U11556 ( n6933, n12285, n12286 );
nor U11557 ( n12285, n12287, n12288 );
nor U11558 ( n12288, n20164, n12289 );
nor U11559 ( n12287, n20165, n12271 );
nand U11560 ( n6928, n12290, n12291 );
nor U11561 ( n12291, n12292, n12293 );
nor U11562 ( n12293, n10965, n12294 );
nand U11563 ( n12294, n12295, n12243 );
nor U11564 ( n12295, n12240, n10410 );
not U11565 ( n12240, n12233 );
nand U11566 ( n12233, n20164, n10233 );
nor U11567 ( n12292, n19162, g35 );
nor U11568 ( n12290, n12269, n12296 );
nor U11569 ( n12296, n20164, n12271 );
not U11570 ( n12271, n12289 );
nor U11571 ( n12289, n10965, n12243 );
not U11572 ( n12269, n12286 );
nand U11573 ( n12286, n12297, n12243 );
nor U11574 ( n12297, n11148, n11837 );
nand U11575 ( n11148, n12298, n20204 );
nor U11576 ( n12298, n20203, n12072 );
nand U11577 ( n6923, n12299, n12300 );
nand U11578 ( n12300, n10997, n10527 );
nand U11579 ( n12299, n12301, g35 );
nand U11580 ( n12301, n12302, n12303 );
nand U11581 ( n12303, n12304, n10825 );
nand U11582 ( n12302, n12305, n12306 );
nand U11583 ( n12306, n19165, n10297 );
not U11584 ( n12305, n12304 );
nand U11585 ( n12304, n12307, n12243 );
not U11586 ( n12243, n12234 );
nand U11587 ( n12234, n12308, n11523 );
nor U11588 ( n12308, n11850, n12309 );
nor U11589 ( n12309, n20213, n11607 );
nor U11590 ( n12307, n20165, n10410 );
nand U11591 ( n6918, n12310, n12311 );
or U11592 ( n12311, n12312, n12313 );
nor U11593 ( n12310, n12314, n12315 );
nor U11594 ( n12315, n19163, g35 );
nor U11595 ( n12314, n10965, n12316 );
nand U11596 ( n12316, n12313, n10527 );
nand U11597 ( n12313, n12317, n12318 );
nor U11598 ( n12317, n19165, n20159 );
nand U11599 ( n6913, n12319, n12320 );
nand U11600 ( n12320, n12321, n12322 );
nor U11601 ( n12319, n12323, n12324 );
nor U11602 ( n12324, n20163, g35 );
nor U11603 ( n12323, n10965, n12325 );
or U11604 ( n12325, n12321, n19163 );
nor U11605 ( n12321, n12326, n10319 );
nand U11606 ( n6908, n12327, n12328 );
or U11607 ( n12328, n12329, n12312 );
nor U11608 ( n12327, n12330, n12331 );
nor U11609 ( n12331, n20162, g35 );
nor U11610 ( n12330, n10977, n12332 );
nand U11611 ( n12332, n12329, n10789 );
nand U11612 ( n12329, n12333, n10388 );
nand U11613 ( n6903, n12334, n12335 );
nand U11614 ( n12335, n12336, n12322 );
nor U11615 ( n12334, n12337, n12338 );
nor U11616 ( n12338, n20161, g35 );
nor U11617 ( n12337, n10979, n12339 );
or U11618 ( n12339, n12336, n20162 );
nor U11619 ( n12336, n12326, n10388 );
nand U11620 ( n6898, n12340, n12341 );
nand U11621 ( n12341, n12342, n12322 );
not U11622 ( n12322, n12312 );
nor U11623 ( n12340, n12343, n12344 );
nor U11624 ( n12344, n20160, g35 );
nor U11625 ( n12343, n10979, n12345 );
or U11626 ( n12345, n12342, n20161 );
and U11627 ( n12342, n12333, n10319 );
nand U11628 ( n6893, n12346, n12347 );
nand U11629 ( n12347, n10996, n10753 );
nor U11630 ( n12346, n12348, n12349 );
nor U11631 ( n12349, n20160, n12211 );
nor U11632 ( n12348, n12216, n12312 );
nand U11633 ( n12312, n12350, g35 );
nor U11634 ( n12350, n12351, n12352 );
nor U11635 ( n12352, n12353, n12354 );
nor U11636 ( n12351, n20025, n12355 );
not U11637 ( n12216, n12208 );
nand U11638 ( n6888, n12356, n12357 );
nand U11639 ( n12357, n12204, n10753 );
nand U11640 ( n12356, n12211, n10528 );
not U11641 ( n12211, n12204 );
nor U11642 ( n12204, n10979, n12208 );
nor U11643 ( n12208, n12358, n12359 );
nand U11644 ( n6883, n12360, n12361 );
nand U11645 ( n12361, n12362, n10528 );
nor U11646 ( n12360, n12363, n12364 );
nor U11647 ( n12364, n10979, n12365 );
nand U11648 ( n12365, n12366, n12367 );
nand U11649 ( n12367, n12368, n12369 );
nor U11650 ( n12368, n12370, n12371 );
nor U11651 ( n12371, n12353, n12372 );
nor U11652 ( n12370, n10337, n12355 );
nor U11653 ( n12366, n12359, n12373 );
nor U11654 ( n12373, n12374, n12369 );
nand U11655 ( n12369, n12358, n10528 );
nand U11656 ( n12358, n19165, n20159 );
nand U11657 ( n12374, n12375, n12376 );
nand U11658 ( n12376, n12353, n10337 );
nand U11659 ( n12375, n12372, n12355 );
not U11660 ( n12372, n12354 );
nand U11661 ( n12354, n11918, n12377 );
nor U11662 ( n12363, n20159, g35 );
nand U11663 ( n6878, n12378, n12379 );
nand U11664 ( n12379, n10996, n10297 );
nor U11665 ( n12378, n12380, n12381 );
nor U11666 ( n12381, n12382, n12326 );
nand U11667 ( n12326, n10297, n12318 );
and U11668 ( n12380, n10388, n12362 );
nand U11669 ( n6873, n12383, n12384 );
nand U11670 ( n12384, n12362, n10297 );
nor U11671 ( n12383, n12385, n12386 );
nor U11672 ( n12386, n10979, n12387 );
nand U11673 ( n12387, n12388, n12389 );
nor U11674 ( n12388, n19165, n12359 );
nor U11675 ( n12385, n20157, g35 );
nand U11676 ( n6868, n12390, n12391 );
nand U11677 ( n12391, n10996, n10319 );
nor U11678 ( n12390, n12392, n12393 );
nor U11679 ( n12393, n12394, n12395 );
nand U11680 ( n12395, n12396, n11572 );
xor U11681 ( n12394, n19565, n12397 );
nor U11682 ( n12397, n20159, n10297 );
nor U11683 ( n12392, n20157, n12398 );
nor U11684 ( n12398, n12399, n11938 );
nor U11685 ( n12399, n12396, n10985 );
and U11686 ( n12396, n12400, n11061 );
nor U11687 ( n12400, n19247, n12401 );
nand U11688 ( n6863, n12402, n12403 );
nand U11689 ( n12403, n12362, n10319 );
nor U11690 ( n12362, n12318, n10985 );
nand U11691 ( n12402, n12404, n12405 );
nor U11692 ( n12405, n12382, n12406 );
nor U11693 ( n12406, n12333, n10319 );
nor U11694 ( n12333, n10297, n12359 );
not U11695 ( n12359, n12318 );
nand U11696 ( n12318, n12353, n12407 );
or U11697 ( n12407, n12401, n19247 );
nor U11698 ( n12401, n12408, n11954 );
not U11699 ( n12353, n12355 );
nand U11700 ( n12355, n12409, n12377 );
nand U11701 ( n12377, n20050, n10323 );
nor U11702 ( n12409, n11956, n12410 );
nor U11703 ( n12410, n10296, n12411 );
nand U11704 ( n12411, n10383, n10238 );
not U11705 ( n12382, n12389 );
nand U11706 ( n12389, n11959, n11061 );
not U11707 ( n11061, n11082 );
nand U11708 ( n11082, n12412, n19997 );
nor U11709 ( n12412, n19996, n11961 );
nor U11710 ( n12404, n10978, n10388 );
nand U11711 ( n6858, n12413, n12414 );
or U11712 ( n12414, n12415, n19542 );
nor U11713 ( n12413, n12416, n12417 );
nor U11714 ( n12417, n10712, n12418 );
nand U11715 ( n12418, n12419, n19167 );
nor U11716 ( n12419, n10979, n12420 );
nor U11717 ( n12416, n19166, n12421 );
nor U11718 ( n12421, n12422, n10985 );
nor U11719 ( n12422, n19167, n12420 );
nand U11720 ( n6853, n12423, n12424 );
nand U11721 ( n12424, n12425, n10712 );
nand U11722 ( n12423, n12415, n10629 );
nand U11723 ( n6848, n12426, n12427 );
nand U11724 ( n12427, n12428, n10629 );
nor U11725 ( n12426, n12429, n12430 );
nor U11726 ( n12430, n19543, g35 );
nor U11727 ( n12429, n10978, n12431 );
nand U11728 ( n12431, n12432, n19167 );
nand U11729 ( n6843, n12433, n12434 );
or U11730 ( n12434, n12435, n19543 );
nor U11731 ( n12433, n12436, n12437 );
nor U11732 ( n12437, n10713, n12438 );
nand U11733 ( n12438, n12439, n20155 );
nor U11734 ( n12439, n10978, n12440 );
nor U11735 ( n12436, n20156, n12441 );
nor U11736 ( n12441, n12442, n10985 );
nor U11737 ( n12442, n20155, n12440 );
nand U11738 ( n6838, n12443, n12444 );
nand U11739 ( n12444, n12428, n10713 );
nand U11740 ( n12443, n12435, n10573 );
nand U11741 ( n6833, n12445, n12446 );
nand U11742 ( n12446, n12425, n10573 );
not U11743 ( n12425, n12415 );
nand U11744 ( n12415, g35, n12420 );
nor U11745 ( n12445, n12447, n12448 );
nor U11746 ( n12448, n19556, g35 );
nor U11747 ( n12447, n10978, n12449 );
or U11748 ( n12449, n10573, n12420 );
nand U11749 ( n6828, n12450, n12451 );
nand U11750 ( n12451, n10995, n10425 );
nand U11751 ( n12450, n12452, g35 );
nand U11752 ( n12452, n12453, n12454 );
or U11753 ( n12454, n12455, n19556 );
nand U11754 ( n12453, n12456, n12455 );
nor U11755 ( n12455, n12457, n12458 );
xnor U11756 ( n12456, n10425, n19171 );
nand U11757 ( n6823, n12459, n12460 );
nand U11758 ( n12460, n12461, g35 );
nor U11759 ( n12461, n19168, n12462 );
nor U11760 ( n12462, n12463, n12458 );
nor U11761 ( n12463, n12464, n10695 );
nand U11762 ( n12459, n12465, n10695 );
nand U11763 ( n12465, g35, n12466 );
nand U11764 ( n12466, n12467, n12468 );
nand U11765 ( n12468, n10425, n12457 );
nand U11766 ( n6818, n12469, n12470 );
nand U11767 ( n12470, n10994, n10411 );
nand U11768 ( n12469, g35, n12471 );
nand U11769 ( n12471, n12472, n12473 );
or U11770 ( n12473, n12420, n20146 );
nand U11771 ( n12420, n12474, n12467 );
nor U11772 ( n12474, n20150, n20153 );
nor U11773 ( n12472, n12475, n12476 );
nor U11774 ( n12476, n12477, n12458 );
nor U11775 ( n12477, n12478, n12479 );
nand U11776 ( n12479, n12480, n12481 );
nand U11777 ( n12481, n20153, n12482 );
nand U11778 ( n12482, n12483, n12484 );
nand U11779 ( n12484, n10234, n10790 );
nand U11780 ( n12483, n20150, n10529 );
nand U11781 ( n12480, n20151, n12485 );
nand U11782 ( n12485, n12486, n12487 );
or U11783 ( n12487, n20153, n20148 );
or U11784 ( n12486, n20150, n19170 );
nor U11785 ( n12478, n20147, n12457 );
nor U11786 ( n12475, n20154, n12467 );
nand U11787 ( n6813, n12488, n12489 );
nor U11788 ( n12489, n12490, n12491 );
nor U11789 ( n12491, n10978, n12492 );
nand U11790 ( n12492, n12467, n10234 );
nor U11791 ( n12490, n20152, g35 );
nor U11792 ( n12488, n12493, n12494 );
nor U11793 ( n12494, n20153, n12495 );
nand U11794 ( n6808, n12496, n12497 );
nand U11795 ( n12497, n10995, n10234 );
nor U11796 ( n12496, n12498, n12499 );
nor U11797 ( n12499, n20152, n12500 );
nor U11798 ( n12500, n12501, n12502 );
nand U11799 ( n12502, n12495, n11547 );
nor U11800 ( n12501, n11131, n10985 );
nor U11801 ( n12498, n12503, n12504 );
nand U11802 ( n12504, n12467, n11131 );
not U11803 ( n11131, n11150 );
nand U11804 ( n12503, n12505, n12506 );
nand U11805 ( n12506, n12507, n11822 );
nand U11806 ( n12505, n12508, n11824 );
not U11807 ( n12508, n12507 );
nor U11808 ( n12507, n10234, n20153 );
nand U11809 ( n6803, n12509, n12510 );
nor U11810 ( n12509, n12511, n12512 );
nor U11811 ( n12512, n20150, n12513 );
nor U11812 ( n12511, n20151, n12495 );
nand U11813 ( n6798, n12514, n12515 );
nor U11814 ( n12515, n12516, n12517 );
nor U11815 ( n12517, n10978, n12518 );
nand U11816 ( n12518, n12519, n12467 );
nor U11817 ( n12519, n12464, n10411 );
not U11818 ( n12464, n12457 );
nand U11819 ( n12457, n20150, n10234 );
nor U11820 ( n12516, n19169, g35 );
nor U11821 ( n12514, n12493, n12520 );
nor U11822 ( n12520, n20150, n12495 );
not U11823 ( n12495, n12513 );
nor U11824 ( n12513, n10976, n12467 );
not U11825 ( n12493, n12510 );
nand U11826 ( n12510, n12521, n12467 );
nor U11827 ( n12521, n11150, n11837 );
nand U11828 ( n11150, n12522, n20204 );
nor U11829 ( n12522, n12072, n10231 );
not U11830 ( n12072, n11839 );
nor U11831 ( n11839, n12523, n20205 );
nand U11832 ( n6793, n12524, n12525 );
nand U11833 ( n12525, n10993, n10529 );
nand U11834 ( n12524, n12526, g35 );
nand U11835 ( n12526, n12527, n12528 );
nand U11836 ( n12528, n12529, n10826 );
nand U11837 ( n12527, n12530, n12531 );
nand U11838 ( n12531, n19172, n10298 );
not U11839 ( n12530, n12529 );
nand U11840 ( n12529, n12532, n12467 );
not U11841 ( n12467, n12458 );
nand U11842 ( n12458, n12533, n12534 );
nand U11843 ( n12534, n11621, n10358 );
nor U11844 ( n12532, n20151, n10411 );
nand U11845 ( n6788, n12535, n12536 );
or U11846 ( n12536, n12537, n12538 );
nor U11847 ( n12535, n12539, n12540 );
nor U11848 ( n12540, n19170, g35 );
nor U11849 ( n12539, n10975, n12541 );
nand U11850 ( n12541, n12538, n10529 );
nand U11851 ( n12538, n12542, n12543 );
nor U11852 ( n12542, n19172, n20145 );
nand U11853 ( n6783, n12544, n12545 );
nand U11854 ( n12545, n12546, n12547 );
nor U11855 ( n12544, n12548, n12549 );
nor U11856 ( n12549, n20149, g35 );
nor U11857 ( n12548, n10975, n12550 );
or U11858 ( n12550, n12546, n19170 );
nor U11859 ( n12546, n12551, n10320 );
nand U11860 ( n6778, n12552, n12553 );
or U11861 ( n12553, n12554, n12537 );
nor U11862 ( n12552, n12555, n12556 );
nor U11863 ( n12556, n20148, g35 );
nor U11864 ( n12555, n10975, n12557 );
nand U11865 ( n12557, n12554, n10790 );
nand U11866 ( n12554, n12558, n10389 );
nand U11867 ( n6773, n12559, n12560 );
nand U11868 ( n12560, n12561, n12547 );
nor U11869 ( n12559, n12562, n12563 );
nor U11870 ( n12563, n20147, g35 );
nor U11871 ( n12562, n10975, n12564 );
or U11872 ( n12564, n12561, n20148 );
nor U11873 ( n12561, n12551, n10389 );
nand U11874 ( n6768, n12565, n12566 );
nand U11875 ( n12566, n12567, n12547 );
not U11876 ( n12547, n12537 );
nor U11877 ( n12565, n12568, n12569 );
nor U11878 ( n12569, n20146, g35 );
nor U11879 ( n12568, n10975, n12570 );
or U11880 ( n12570, n12567, n20147 );
and U11881 ( n12567, n12558, n10320 );
nand U11882 ( n6763, n12571, n12572 );
nand U11883 ( n12572, n10994, n10754 );
nor U11884 ( n12571, n12573, n12574 );
nor U11885 ( n12574, n20146, n12435 );
nor U11886 ( n12573, n12440, n12537 );
nand U11887 ( n12537, n12575, g35 );
nor U11888 ( n12575, n12576, n12577 );
nor U11889 ( n12577, n10473, n12578 );
nor U11890 ( n12576, n12579, n12580 );
not U11891 ( n12440, n12432 );
nand U11892 ( n6758, n12581, n12582 );
nand U11893 ( n12582, n12428, n10754 );
nand U11894 ( n12581, n12435, n10530 );
not U11895 ( n12435, n12428 );
nor U11896 ( n12428, n10975, n12432 );
nor U11897 ( n12432, n12583, n12584 );
nand U11898 ( n6753, n12585, n12586 );
nand U11899 ( n12586, n12587, n10530 );
nor U11900 ( n12585, n12588, n12589 );
nor U11901 ( n12589, n10975, n12590 );
nand U11902 ( n12590, n12591, n12592 );
nand U11903 ( n12592, n12593, n12594 );
nor U11904 ( n12593, n12595, n12596 );
nor U11905 ( n12596, n12579, n12597 );
nor U11906 ( n12595, n20026, n12578 );
nor U11907 ( n12591, n12584, n12598 );
nor U11908 ( n12598, n12599, n12594 );
nand U11909 ( n12594, n12583, n10530 );
nand U11910 ( n12583, n19172, n20145 );
nand U11911 ( n12599, n12600, n12601 );
nand U11912 ( n12601, n12597, n12578 );
not U11913 ( n12597, n12580 );
nand U11914 ( n12580, n11918, n12602 );
nor U11915 ( n11918, n19951, n11956 );
nand U11916 ( n12600, n12579, n20026 );
not U11917 ( n12579, n12578 );
nor U11918 ( n12588, n20145, g35 );
nand U11919 ( n6748, n12603, n12604 );
nand U11920 ( n12604, n10993, n10298 );
nor U11921 ( n12603, n12605, n12606 );
nor U11922 ( n12606, n12607, n12551 );
nand U11923 ( n12551, n10298, n12543 );
and U11924 ( n12605, n10389, n12587 );
nand U11925 ( n6743, n12608, n12609 );
nand U11926 ( n12609, n12587, n10298 );
nor U11927 ( n12608, n12610, n12611 );
nor U11928 ( n12611, n10975, n12612 );
nand U11929 ( n12612, n12613, n12614 );
nor U11930 ( n12613, n19172, n12584 );
nor U11931 ( n12610, n20143, g35 );
nand U11932 ( n6738, n12615, n12616 );
nand U11933 ( n12616, n10993, n10320 );
nor U11934 ( n12615, n12617, n12618 );
nor U11935 ( n12618, n20143, n12619 );
nor U11936 ( n12619, n12620, n11938 );
nor U11937 ( n12620, n12621, n10984 );
nor U11938 ( n12617, n12622, n12623 );
nand U11939 ( n12623, n12621, n11572 );
and U11940 ( n12621, n12624, n11067 );
xor U11941 ( n12622, n19565, n12625 );
nor U11942 ( n12625, n20145, n10298 );
nand U11943 ( n6733, n12626, n12627 );
nand U11944 ( n12627, n12587, n10320 );
nor U11945 ( n12587, n12543, n10983 );
not U11946 ( n12543, n12584 );
nand U11947 ( n12626, n12628, n12629 );
nor U11948 ( n12629, n12607, n12630 );
nor U11949 ( n12630, n12558, n10320 );
nor U11950 ( n12558, n10298, n12584 );
nor U11951 ( n12584, n12578, n12624 );
nor U11952 ( n12624, n20023, n12631 );
and U11953 ( n12631, n12632, n20032 );
nor U11954 ( n12632, n20031, n11954 );
nand U11955 ( n11954, n12633, n12634 );
nor U11956 ( n12634, n10660, n12635 );
nand U11957 ( n12635, n10642, n10286 );
nor U11958 ( n12633, n10480, n12636 );
nand U11959 ( n12636, n19243, n19244 );
nand U11960 ( n12578, n12637, n12602 );
nand U11961 ( n12602, n20050, n10455 );
nor U11962 ( n12637, n11956, n12638 );
nor U11963 ( n12638, n10296, n12639 );
nand U11964 ( n12639, n20197, n10238 );
and U11965 ( n11956, n19567, n12640 );
nand U11966 ( n12640, n11424, n11418 );
not U11967 ( n12607, n12614 );
nand U11968 ( n12614, n11959, n11067 );
not U11969 ( n11067, n11084 );
nand U11970 ( n11084, n12641, n19996 );
nor U11971 ( n12641, n11961, n10224 );
not U11972 ( n11961, n12188 );
nor U11973 ( n12188, n12642, n12643 );
or U11974 ( n12642, n19998, n12644 );
nor U11975 ( n12628, n10974, n10389 );
nand U11976 ( n6718, n12645, n12646 );
nand U11977 ( n12646, g35, n10382 );
nand U11978 ( n12645, n10994, n10295 );
nand U11979 ( n6713, n12647, n12648 );
nand U11980 ( n12648, g35, n10295 );
nand U11981 ( n12647, n10994, n10237 );
nor U11982 ( n6708, n20141, n10983 );
nand U11983 ( n6703, n12649, n12650 );
or U11984 ( n12650, n12651, n19548 );
nor U11985 ( n12649, n12652, n12653 );
nor U11986 ( n12653, n10714, n12654 );
nand U11987 ( n12654, n12655, n19174 );
nor U11988 ( n12655, n10974, n12656 );
nor U11989 ( n12652, n19173, n12657 );
nor U11990 ( n12657, n12658, n10983 );
nor U11991 ( n12658, n19174, n12656 );
nand U11992 ( n6698, n12659, n12660 );
nand U11993 ( n12660, n12661, n10714 );
nand U11994 ( n12659, n12651, n10630 );
nand U11995 ( n6693, n12662, n12663 );
nand U11996 ( n12663, n12664, n10630 );
nor U11997 ( n12662, n12665, n12666 );
nor U11998 ( n12666, n19549, g35 );
nor U11999 ( n12665, n10974, n12667 );
nand U12000 ( n12667, n12668, n19174 );
nand U12001 ( n6688, n12669, n12670 );
or U12002 ( n12670, n12671, n19549 );
nor U12003 ( n12669, n12672, n12673 );
nor U12004 ( n12673, n10715, n12674 );
nand U12005 ( n12674, n12675, n20139 );
nor U12006 ( n12675, n10974, n12676 );
nor U12007 ( n12672, n20140, n12677 );
nor U12008 ( n12677, n12678, n10981 );
nor U12009 ( n12678, n20139, n12676 );
nand U12010 ( n6683, n12679, n12680 );
nand U12011 ( n12680, n12664, n10715 );
nand U12012 ( n12679, n12671, n10574 );
nand U12013 ( n6678, n12681, n12682 );
nand U12014 ( n12682, n12661, n10574 );
not U12015 ( n12661, n12651 );
nand U12016 ( n12651, g35, n12656 );
nor U12017 ( n12681, n12683, n12684 );
nor U12018 ( n12684, n19559, g35 );
nor U12019 ( n12683, n10974, n12685 );
or U12020 ( n12685, n10574, n12656 );
nand U12021 ( n6673, n12686, n12687 );
nand U12022 ( n12687, n10995, n10426 );
nand U12023 ( n12686, n12688, g35 );
nand U12024 ( n12688, n12689, n12690 );
or U12025 ( n12690, n12691, n19559 );
nand U12026 ( n12689, n12692, n12691 );
nor U12027 ( n12691, n12693, n12694 );
xnor U12028 ( n12692, n10426, n19179 );
nand U12029 ( n6668, n12695, n12696 );
nand U12030 ( n12696, n12697, g35 );
nor U12031 ( n12697, n19175, n12698 );
nor U12032 ( n12698, n12699, n12694 );
nor U12033 ( n12699, n12700, n10686 );
nand U12034 ( n12695, n12701, n10686 );
nand U12035 ( n12701, g35, n12702 );
nand U12036 ( n12702, n12703, n12704 );
nand U12037 ( n12704, n10426, n12693 );
nand U12038 ( n6663, n12705, n12706 );
nand U12039 ( n12706, n10994, n10412 );
nand U12040 ( n12705, g35, n12707 );
nand U12041 ( n12707, n12708, n12709 );
or U12042 ( n12709, n12656, n20131 );
nand U12043 ( n12656, n12710, n12703 );
nor U12044 ( n12710, n20135, n20138 );
nor U12045 ( n12708, n12711, n12712 );
nor U12046 ( n12712, n12713, n12694 );
nor U12047 ( n12713, n12714, n12715 );
nand U12048 ( n12715, n12716, n12717 );
nand U12049 ( n12717, n20138, n12718 );
nand U12050 ( n12718, n12719, n12720 );
or U12051 ( n12720, n20136, n20134 );
nand U12052 ( n12719, n20135, n10531 );
nand U12053 ( n12716, n20136, n12721 );
nand U12054 ( n12721, n12722, n12723 );
or U12055 ( n12723, n20138, n20133 );
or U12056 ( n12722, n20135, n19178 );
nor U12057 ( n12714, n20132, n12693 );
nor U12058 ( n12711, n19176, n12703 );
nand U12059 ( n6658, n12724, n12725 );
nor U12060 ( n12725, n12726, n12727 );
nor U12061 ( n12727, n10974, n12728 );
nand U12062 ( n12728, n12703, n10341 );
nor U12063 ( n12726, n20137, g35 );
nor U12064 ( n12724, n12729, n12730 );
nor U12065 ( n12730, n20138, n12731 );
nand U12066 ( n6653, n12732, n12733 );
nand U12067 ( n12733, n10995, n10341 );
nor U12068 ( n12732, n12734, n12735 );
nor U12069 ( n12735, n20137, n12736 );
nor U12070 ( n12736, n12737, n12738 );
nand U12071 ( n12738, n12731, n11547 );
nor U12072 ( n12737, n11140, n10981 );
nor U12073 ( n12734, n12739, n12740 );
nand U12074 ( n12740, n12703, n11140 );
not U12075 ( n11140, n11166 );
nand U12076 ( n12739, n12741, n12742 );
nand U12077 ( n12742, n12743, n11822 );
nand U12078 ( n12741, n12744, n11824 );
not U12079 ( n12744, n12743 );
nor U12080 ( n12743, n10341, n20138 );
nand U12081 ( n6648, n12745, n12746 );
nor U12082 ( n12745, n12747, n12748 );
nor U12083 ( n12748, n20135, n12749 );
nor U12084 ( n12747, n20136, n12731 );
nand U12085 ( n6643, n12750, n12751 );
nor U12086 ( n12751, n12752, n12753 );
nor U12087 ( n12753, n10976, n12754 );
nand U12088 ( n12754, n12755, n12703 );
nor U12089 ( n12755, n12700, n10412 );
not U12090 ( n12700, n12693 );
nand U12091 ( n12693, n20135, n10341 );
nor U12092 ( n12752, n19177, g35 );
nor U12093 ( n12750, n12729, n12756 );
nor U12094 ( n12756, n20135, n12731 );
not U12095 ( n12731, n12749 );
nor U12096 ( n12749, n10976, n12703 );
not U12097 ( n12729, n12746 );
nand U12098 ( n12746, n12757, n12703 );
nor U12099 ( n12757, n11166, n11837 );
nand U12100 ( n11166, n12758, n11662 );
nand U12101 ( n6638, n12759, n12760 );
nand U12102 ( n12760, n10995, n10531 );
nand U12103 ( n12759, n12761, g35 );
nand U12104 ( n12761, n12762, n12763 );
nand U12105 ( n12763, n12764, n10827 );
nand U12106 ( n12762, n12765, n12766 );
nand U12107 ( n12766, n19180, n10314 );
not U12108 ( n12765, n12764 );
nand U12109 ( n12764, n12767, n12703 );
not U12110 ( n12703, n12694 );
nand U12111 ( n12694, n12768, n11527 );
nor U12112 ( n11527, n20199, n20198 );
nor U12113 ( n12768, n11850, n12769 );
nor U12114 ( n12769, n20207, n11607 );
nor U12115 ( n12767, n20136, n10412 );
nand U12116 ( n6633, n12770, n12771 );
or U12117 ( n12771, n12772, n12773 );
nor U12118 ( n12770, n12774, n12775 );
nor U12119 ( n12775, n19178, g35 );
nor U12120 ( n12774, n10977, n12776 );
nand U12121 ( n12776, n12773, n10531 );
nand U12122 ( n12773, n12777, n10440 );
nand U12123 ( n6628, n12778, n12779 );
nand U12124 ( n12779, n12780, n12781 );
nor U12125 ( n12778, n12782, n12783 );
nor U12126 ( n12783, n20134, g35 );
nor U12127 ( n12782, n10979, n12784 );
or U12128 ( n12784, n12780, n19178 );
nor U12129 ( n12780, n12785, n10355 );
nand U12130 ( n6623, n12786, n12787 );
nand U12131 ( n12787, n12788, n12781 );
nor U12132 ( n12786, n12789, n12790 );
nor U12133 ( n12790, n20133, g35 );
nor U12134 ( n12789, n10978, n12791 );
or U12135 ( n12791, n12788, n20134 );
nor U12136 ( n12788, n12792, n12793 );
not U12137 ( n12792, n11092 );
nand U12138 ( n6618, n12794, n12795 );
nand U12139 ( n12795, n12796, n12781 );
nor U12140 ( n12794, n12797, n12798 );
nor U12141 ( n12798, n20132, g35 );
nor U12142 ( n12797, n10954, n12799 );
or U12143 ( n12799, n12796, n20133 );
nor U12144 ( n12796, n12785, n10440 );
nand U12145 ( n6613, n12800, n12801 );
nand U12146 ( n12801, n12802, n12781 );
not U12147 ( n12781, n12772 );
nor U12148 ( n12800, n12803, n12804 );
nor U12149 ( n12804, n20131, g35 );
nor U12150 ( n12803, n10954, n12805 );
or U12151 ( n12805, n12802, n20132 );
and U12152 ( n12802, n12777, n20129 );
nand U12153 ( n6608, n12806, n12807 );
nand U12154 ( n12807, n10996, n10755 );
nor U12155 ( n12806, n12808, n12809 );
nor U12156 ( n12809, n20131, n12671 );
nor U12157 ( n12808, n12676, n12772 );
nand U12158 ( n12772, n12810, g35 );
nor U12159 ( n12810, n12811, n12812 );
nor U12160 ( n12812, n12813, n12814 );
nor U12161 ( n12811, n20061, n12815 );
not U12162 ( n12676, n12668 );
nand U12163 ( n6603, n12816, n12817 );
nand U12164 ( n12817, n12664, n10755 );
nand U12165 ( n12816, n12671, n10532 );
not U12166 ( n12671, n12664 );
nor U12167 ( n12664, n10954, n12668 );
nor U12168 ( n12668, n12818, n12793 );
nand U12169 ( n6598, n12819, n12820 );
nand U12170 ( n12820, n12821, n10532 );
nor U12171 ( n12819, n12822, n12823 );
nor U12172 ( n12823, n10954, n12824 );
nand U12173 ( n12824, n12825, n12826 );
nand U12174 ( n12826, n12827, n12828 );
nor U12175 ( n12827, n12829, n12830 );
nor U12176 ( n12830, n12813, n12831 );
nor U12177 ( n12829, n12815, n10338 );
nor U12178 ( n12825, n12793, n12832 );
nor U12179 ( n12832, n12833, n12828 );
nand U12180 ( n12828, n12818, n10532 );
nand U12181 ( n12818, n19180, n20130 );
nand U12182 ( n12833, n12834, n12835 );
nand U12183 ( n12835, n12813, n10338 );
not U12184 ( n12813, n12815 );
nand U12185 ( n12834, n12831, n12815 );
not U12186 ( n12831, n12814 );
nand U12187 ( n12814, n12836, n12837 );
nor U12188 ( n12822, n20130, g35 );
nand U12189 ( n6593, n12838, n12839 );
nand U12190 ( n12839, n10996, n10314 );
nor U12191 ( n12838, n12840, n12841 );
nor U12192 ( n12841, n12842, n12785 );
or U12193 ( n12785, n20129, n12793 );
nor U12194 ( n12840, n20130, n12843 );
nand U12195 ( n6588, n12844, n12845 );
nand U12196 ( n12845, n12821, n10314 );
nor U12197 ( n12844, n12846, n12847 );
nor U12198 ( n12847, n10953, n12848 );
nand U12199 ( n12848, n12777, n12849 );
nor U12200 ( n12777, n19180, n12793 );
nor U12201 ( n12846, n20128, g35 );
nand U12202 ( n6583, n12850, n12851 );
nand U12203 ( n12851, n10996, n10355 );
nor U12204 ( n12850, n12852, n12853 );
nor U12205 ( n12853, n20128, n12854 );
nor U12206 ( n12854, n12855, n11938 );
nor U12207 ( n12855, n12856, n10980 );
nor U12208 ( n12856, n12857, n12858 );
nor U12209 ( n12852, n12859, n12860 );
nand U12210 ( n12860, n12861, n12862 );
xnor U12211 ( n12861, n11092, n19565 );
nor U12212 ( n11092, n10314, n20130 );
nand U12213 ( n12859, n11572, n11060 );
nand U12214 ( n6578, n12863, n12864 );
nand U12215 ( n12864, n12821, n10355 );
not U12216 ( n12821, n12843 );
nand U12217 ( n12843, n12793, g35 );
nand U12218 ( n12863, n12865, n12866 );
nor U12219 ( n12866, n12842, n12867 );
nor U12220 ( n12867, n12868, n10355 );
nor U12221 ( n12868, n12793, n10314 );
nor U12222 ( n12793, n12815, n12862 );
not U12223 ( n12862, n12858 );
nand U12224 ( n12858, n10589, n12869 );
nand U12225 ( n12869, n12870, n20067 );
nor U12226 ( n12870, n10294, n12871 );
nand U12227 ( n12815, n12872, n12837 );
nand U12228 ( n12837, n20088, n10621 );
nor U12229 ( n12872, n12873, n12874 );
nor U12230 ( n12874, n20142, n12875 );
not U12231 ( n12842, n12849 );
nand U12232 ( n12849, n11959, n11060 );
not U12233 ( n11060, n12857 );
nand U12234 ( n12857, n12876, n12877 );
nor U12235 ( n12876, n19997, n10404 );
nor U12236 ( n12865, n10953, n10440 );
nand U12237 ( n6573, n12878, n12879 );
or U12238 ( n12879, n12880, n19546 );
nor U12239 ( n12878, n12881, n12882 );
nor U12240 ( n12882, n10716, n12883 );
nand U12241 ( n12883, n12884, n19182 );
nor U12242 ( n12884, n10952, n12885 );
nor U12243 ( n12881, n19181, n12886 );
nor U12244 ( n12886, n12887, n10983 );
nor U12245 ( n12887, n19182, n12885 );
nand U12246 ( n6568, n12888, n12889 );
nand U12247 ( n12889, n12890, n10716 );
nand U12248 ( n12888, n12880, n10631 );
nand U12249 ( n6563, n12891, n12892 );
nand U12250 ( n12892, n12893, n10631 );
nor U12251 ( n12891, n12894, n12895 );
nor U12252 ( n12895, n19547, g35 );
nor U12253 ( n12894, n10951, n12896 );
nand U12254 ( n12896, n12897, n19182 );
nand U12255 ( n6558, n12898, n12899 );
or U12256 ( n12899, n12900, n19547 );
nor U12257 ( n12898, n12901, n12902 );
nor U12258 ( n12902, n10717, n12903 );
nand U12259 ( n12903, n12904, n20126 );
nor U12260 ( n12904, n10951, n12905 );
nor U12261 ( n12901, n20127, n12906 );
nor U12262 ( n12906, n12907, n10983 );
nor U12263 ( n12907, n20126, n12905 );
nand U12264 ( n6553, n12908, n12909 );
nand U12265 ( n12909, n12893, n10717 );
nand U12266 ( n12908, n12900, n10575 );
nand U12267 ( n6548, n12910, n12911 );
nand U12268 ( n12911, n12890, n10575 );
not U12269 ( n12890, n12880 );
nand U12270 ( n12880, g35, n12885 );
nor U12271 ( n12910, n12912, n12913 );
nor U12272 ( n12913, n19558, g35 );
nor U12273 ( n12912, n10951, n12914 );
or U12274 ( n12914, n10575, n12885 );
nand U12275 ( n6543, n12915, n12916 );
nand U12276 ( n12916, n11015, n10427 );
nand U12277 ( n12915, n12917, g35 );
nand U12278 ( n12917, n12918, n12919 );
or U12279 ( n12919, n12920, n19558 );
nand U12280 ( n12918, n12921, n12920 );
nor U12281 ( n12920, n12922, n12923 );
xnor U12282 ( n12921, n10427, n19187 );
nand U12283 ( n6538, n12924, n12925 );
nand U12284 ( n12925, n12926, g35 );
nor U12285 ( n12926, n19183, n12927 );
nor U12286 ( n12927, n12928, n12923 );
nor U12287 ( n12928, n12929, n10687 );
nand U12288 ( n12924, n12930, n10687 );
nand U12289 ( n12930, g35, n12931 );
nand U12290 ( n12931, n12932, n12933 );
nand U12291 ( n12933, n10427, n12922 );
nand U12292 ( n6533, n12934, n12935 );
nand U12293 ( n12935, n11015, n10413 );
nand U12294 ( n12934, g35, n12936 );
nand U12295 ( n12936, n12937, n12938 );
or U12296 ( n12938, n12885, n20118 );
nand U12297 ( n12885, n12939, n12932 );
nor U12298 ( n12939, n20122, n20125 );
nor U12299 ( n12937, n12940, n12941 );
nor U12300 ( n12941, n12942, n12923 );
nor U12301 ( n12942, n12943, n12944 );
nand U12302 ( n12944, n12945, n12946 );
nand U12303 ( n12946, n20125, n12947 );
nand U12304 ( n12947, n12948, n12949 );
or U12305 ( n12949, n20123, n20121 );
nand U12306 ( n12948, n20122, n10533 );
nand U12307 ( n12945, n20123, n12950 );
nand U12308 ( n12950, n12951, n12952 );
or U12309 ( n12952, n20125, n20120 );
or U12310 ( n12951, n20122, n19186 );
nor U12311 ( n12943, n20119, n12922 );
nor U12312 ( n12940, n19184, n12932 );
nand U12313 ( n6528, n12953, n12954 );
nor U12314 ( n12954, n12955, n12956 );
nor U12315 ( n12956, n10951, n12957 );
nand U12316 ( n12957, n12932, n10342 );
nor U12317 ( n12955, n20124, g35 );
nor U12318 ( n12953, n12958, n12959 );
nor U12319 ( n12959, n20125, n12960 );
nand U12320 ( n6523, n12961, n12962 );
nand U12321 ( n12962, n11015, n10342 );
nor U12322 ( n12961, n12963, n12964 );
nor U12323 ( n12964, n20124, n12965 );
nor U12324 ( n12965, n12966, n12967 );
nand U12325 ( n12967, n12960, n11547 );
nor U12326 ( n12966, n11139, n10983 );
nor U12327 ( n12963, n12968, n12969 );
nand U12328 ( n12969, n12932, n11139 );
not U12329 ( n11139, n11168 );
nand U12330 ( n12968, n12970, n12971 );
nand U12331 ( n12971, n12972, n11822 );
nand U12332 ( n12970, n12973, n11824 );
not U12333 ( n12973, n12972 );
nor U12334 ( n12972, n10342, n20125 );
nand U12335 ( n6518, n12974, n12975 );
nor U12336 ( n12974, n12976, n12977 );
nor U12337 ( n12977, n20122, n12978 );
nor U12338 ( n12976, n20123, n12960 );
nand U12339 ( n6513, n12979, n12980 );
nor U12340 ( n12980, n12981, n12982 );
nor U12341 ( n12982, n10951, n12983 );
nand U12342 ( n12983, n12984, n12932 );
nor U12343 ( n12984, n12929, n10413 );
not U12344 ( n12929, n12922 );
nand U12345 ( n12922, n20122, n10342 );
nor U12346 ( n12981, n19185, g35 );
nor U12347 ( n12979, n12958, n12985 );
nor U12348 ( n12985, n20122, n12960 );
not U12349 ( n12960, n12978 );
nor U12350 ( n12978, n10951, n12932 );
not U12351 ( n12958, n12975 );
nand U12352 ( n12975, n12986, n12932 );
nor U12353 ( n12986, n11168, n11837 );
nand U12354 ( n11168, n12987, n12758 );
nor U12355 ( n12758, n20204, n12523 );
nor U12356 ( n12987, n10231, n10405 );
nand U12357 ( n6508, n12988, n12989 );
nand U12358 ( n12989, n11016, n10533 );
nand U12359 ( n12988, n12990, g35 );
nand U12360 ( n12990, n12991, n12992 );
nand U12361 ( n12992, n12993, n10828 );
nand U12362 ( n12991, n12994, n12995 );
nand U12363 ( n12995, n19188, n10315 );
not U12364 ( n12994, n12993 );
nand U12365 ( n12993, n12996, n12932 );
not U12366 ( n12932, n12923 );
nand U12367 ( n12923, n12997, n11522 );
nor U12368 ( n11522, n10225, n20199 );
nor U12369 ( n12997, n11850, n12998 );
nor U12370 ( n12998, n20208, n11607 );
nor U12371 ( n12996, n20123, n10413 );
nand U12372 ( n6503, n12999, n13000 );
or U12373 ( n13000, n13001, n13002 );
nor U12374 ( n12999, n13003, n13004 );
nor U12375 ( n13004, n19186, g35 );
nor U12376 ( n13003, n10951, n13005 );
nand U12377 ( n13005, n13002, n10533 );
nand U12378 ( n13002, n13006, n10441 );
nand U12379 ( n6498, n13007, n13008 );
nand U12380 ( n13008, n13009, n13010 );
nor U12381 ( n13007, n13011, n13012 );
nor U12382 ( n13012, n20121, g35 );
nor U12383 ( n13011, n10951, n13013 );
or U12384 ( n13013, n13009, n19186 );
nor U12385 ( n13009, n13014, n10356 );
nand U12386 ( n6493, n13015, n13016 );
nand U12387 ( n13016, n13017, n13010 );
nor U12388 ( n13015, n13018, n13019 );
nor U12389 ( n13019, n20120, g35 );
nor U12390 ( n13018, n10950, n13020 );
or U12391 ( n13020, n13017, n20121 );
nor U12392 ( n13017, n13021, n13022 );
not U12393 ( n13021, n11078 );
nand U12394 ( n6488, n13023, n13024 );
nand U12395 ( n13024, n13025, n13010 );
nor U12396 ( n13023, n13026, n13027 );
nor U12397 ( n13027, n20119, g35 );
nor U12398 ( n13026, n10950, n13028 );
or U12399 ( n13028, n13025, n20120 );
nor U12400 ( n13025, n13014, n10441 );
nand U12401 ( n6483, n13029, n13030 );
nand U12402 ( n13030, n13031, n13010 );
not U12403 ( n13010, n13001 );
nor U12404 ( n13029, n13032, n13033 );
nor U12405 ( n13033, n20118, g35 );
nor U12406 ( n13032, n10950, n13034 );
or U12407 ( n13034, n13031, n20119 );
and U12408 ( n13031, n13006, n20116 );
nand U12409 ( n6478, n13035, n13036 );
nand U12410 ( n13036, n11016, n10756 );
nor U12411 ( n13035, n13037, n13038 );
nor U12412 ( n13038, n20118, n12900 );
nor U12413 ( n13037, n12905, n13001 );
nand U12414 ( n13001, n13039, g35 );
nor U12415 ( n13039, n13040, n13041 );
nor U12416 ( n13041, n13042, g23683 );
nor U12417 ( n13040, n13043, n13044 );
not U12418 ( n12905, n12897 );
nand U12419 ( n6473, n13045, n13046 );
nand U12420 ( n13046, n12893, n10756 );
nand U12421 ( n13045, n12900, n10534 );
not U12422 ( n12900, n12893 );
nor U12423 ( n12893, n10950, n12897 );
nor U12424 ( n12897, n13047, n13022 );
nand U12425 ( n6468, n13048, n13049 );
nand U12426 ( n13049, n13050, n10534 );
nor U12427 ( n13048, n13051, n13052 );
nor U12428 ( n13052, n10950, n13053 );
nand U12429 ( n13053, n13054, n13055 );
nand U12430 ( n13055, n13056, n13057 );
nor U12431 ( n13056, n13058, n13059 );
nor U12432 ( n13059, n13043, n13060 );
nor U12433 ( n13058, n20062, n13042 );
nor U12434 ( n13054, n13022, n13061 );
nor U12435 ( n13061, n13062, n13057 );
nand U12436 ( n13057, n13047, n10534 );
nand U12437 ( n13047, n19188, n20117 );
nand U12438 ( n13062, n13063, n13064 );
nand U12439 ( n13064, n13060, n13042 );
not U12440 ( n13060, n13044 );
nand U12441 ( n13044, n12836, n13065 );
nand U12442 ( n13063, n13043, n20062 );
not U12443 ( n13043, n13042 );
nor U12444 ( n13051, n20117, g35 );
nand U12445 ( n6463, n13066, n13067 );
nand U12446 ( n13067, n11016, n10315 );
nor U12447 ( n13066, n13068, n13069 );
nor U12448 ( n13069, n13070, n13014 );
or U12449 ( n13014, n20116, n13022 );
nor U12450 ( n13068, n20117, n13071 );
nand U12451 ( n6458, n13072, n13073 );
nand U12452 ( n13073, n13050, n10315 );
nor U12453 ( n13072, n13074, n13075 );
nor U12454 ( n13075, n10948, n13076 );
nand U12455 ( n13076, n13006, n13077 );
nor U12456 ( n13006, n19188, n13022 );
nor U12457 ( n13074, n20115, g35 );
nand U12458 ( n6453, n13078, n13079 );
nand U12459 ( n13079, n11016, n10356 );
nor U12460 ( n13078, n13080, n13081 );
nor U12461 ( n13081, n20115, n13082 );
nor U12462 ( n13082, n13083, n11938 );
nor U12463 ( n13083, n13084, n10984 );
nor U12464 ( n13084, n13085, n13086 );
nor U12465 ( n13080, n13087, n13088 );
nand U12466 ( n13088, n13089, n13090 );
xnor U12467 ( n13089, n11078, n19565 );
nor U12468 ( n11078, n10315, n20117 );
nand U12469 ( n13087, n11572, n11069 );
nand U12470 ( n6448, n13091, n13092 );
nand U12471 ( n13092, n13050, n10356 );
not U12472 ( n13050, n13071 );
nand U12473 ( n13071, n13022, g35 );
nand U12474 ( n13091, n13093, n13094 );
nor U12475 ( n13094, n13070, n13095 );
nor U12476 ( n13095, n13096, n10356 );
nor U12477 ( n13096, n13022, n10315 );
nor U12478 ( n13022, n13042, n13090 );
not U12479 ( n13090, n13086 );
nand U12480 ( n13086, g17400, n13097 );
nand U12481 ( n13097, n13098, n13099 );
nor U12482 ( n13098, n20067, n20068 );
nand U12483 ( n13042, n13100, n13065 );
nand U12484 ( n13065, n20088, n10452 );
nor U12485 ( n13100, n12873, n13101 );
nor U12486 ( n13101, n10382, n12875 );
nand U12487 ( n12875, n10295, n10237 );
not U12488 ( n13070, n13077 );
nand U12489 ( n13077, n11959, n11069 );
not U12490 ( n11069, n13085 );
nand U12491 ( n13085, n12187, n12877 );
nor U12492 ( n12187, n19996, n19997 );
nor U12493 ( n13093, n10948, n10441 );
nand U12494 ( n6443, n13102, n13103 );
or U12495 ( n13103, n13104, n19552 );
nor U12496 ( n13102, n13105, n13106 );
nor U12497 ( n13106, n10718, n13107 );
nand U12498 ( n13107, n13108, n19190 );
nor U12499 ( n13108, n10948, n13109 );
nor U12500 ( n13105, n19189, n13110 );
nor U12501 ( n13110, n13111, n10984 );
nor U12502 ( n13111, n19190, n13109 );
nand U12503 ( n6438, n13112, n13113 );
nand U12504 ( n13113, n13114, n10718 );
nand U12505 ( n13112, n13104, n10632 );
nand U12506 ( n6433, n13115, n13116 );
nand U12507 ( n13116, n13117, n10632 );
nor U12508 ( n13115, n13118, n13119 );
nor U12509 ( n13119, n19553, g35 );
nor U12510 ( n13118, n10948, n13120 );
nand U12511 ( n13120, n13121, n19190 );
nand U12512 ( n6428, n13122, n13123 );
or U12513 ( n13123, n13124, n19553 );
nor U12514 ( n13122, n13125, n13126 );
nor U12515 ( n13126, n10719, n13127 );
nand U12516 ( n13127, n13128, n20113 );
nor U12517 ( n13128, n10948, n13129 );
nor U12518 ( n13125, n20114, n13130 );
nor U12519 ( n13130, n13131, n10984 );
nor U12520 ( n13131, n20113, n13129 );
nand U12521 ( n6423, n13132, n13133 );
nand U12522 ( n13133, n13117, n10719 );
nand U12523 ( n13132, n13124, n10576 );
nand U12524 ( n6418, n13134, n13135 );
nand U12525 ( n13135, n13114, n10576 );
not U12526 ( n13114, n13104 );
nand U12527 ( n13104, g35, n13109 );
nor U12528 ( n13134, n13136, n13137 );
nor U12529 ( n13137, n19561, g35 );
nor U12530 ( n13136, n10948, n13138 );
or U12531 ( n13138, n10576, n13109 );
nand U12532 ( n6413, n13139, n13140 );
nand U12533 ( n13140, n11017, n10428 );
nand U12534 ( n13139, n13141, g35 );
nand U12535 ( n13141, n13142, n13143 );
or U12536 ( n13143, n13144, n19561 );
nand U12537 ( n13142, n13145, n13144 );
nor U12538 ( n13144, n13146, n13147 );
xnor U12539 ( n13145, n10428, n19195 );
nand U12540 ( n6408, n13148, n13149 );
nand U12541 ( n13149, n13150, g35 );
nor U12542 ( n13150, n19191, n13151 );
nor U12543 ( n13151, n13152, n13147 );
nor U12544 ( n13152, n13153, n10688 );
nand U12545 ( n13148, n13154, n10688 );
nand U12546 ( n13154, g35, n13155 );
nand U12547 ( n13155, n13156, n13157 );
nand U12548 ( n13157, n10428, n13146 );
nand U12549 ( n6403, n13158, n13159 );
nand U12550 ( n13159, n11017, n10414 );
nand U12551 ( n13158, g35, n13160 );
nand U12552 ( n13160, n13161, n13162 );
or U12553 ( n13162, n13109, n20105 );
nand U12554 ( n13109, n13163, n13156 );
nor U12555 ( n13163, n20109, n20112 );
nor U12556 ( n13161, n13164, n13165 );
nor U12557 ( n13165, n13166, n13147 );
nor U12558 ( n13166, n13167, n13168 );
nand U12559 ( n13168, n13169, n13170 );
nand U12560 ( n13170, n20112, n13171 );
nand U12561 ( n13171, n13172, n13173 );
nand U12562 ( n13173, n10235, n10791 );
nand U12563 ( n13172, n20109, n10535 );
nand U12564 ( n13169, n20110, n13174 );
nand U12565 ( n13174, n13175, n13176 );
or U12566 ( n13176, n20112, n20107 );
or U12567 ( n13175, n20109, n19194 );
nor U12568 ( n13167, n20106, n13146 );
nor U12569 ( n13164, n19192, n13156 );
nand U12570 ( n6398, n13177, n13178 );
nor U12571 ( n13178, n13179, n13180 );
nor U12572 ( n13180, n10948, n13181 );
nand U12573 ( n13181, n13156, n10235 );
nor U12574 ( n13179, n20111, g35 );
nor U12575 ( n13177, n13182, n13183 );
nor U12576 ( n13183, n20112, n13184 );
nand U12577 ( n6393, n13185, n13186 );
nand U12578 ( n13186, n11017, n10235 );
nor U12579 ( n13185, n13187, n13188 );
nor U12580 ( n13188, n20111, n13189 );
nor U12581 ( n13189, n13190, n13191 );
nand U12582 ( n13191, n13184, n11547 );
nor U12583 ( n13190, n11138, n10985 );
nor U12584 ( n13187, n13192, n13193 );
nand U12585 ( n13193, n13156, n11138 );
not U12586 ( n11138, n11162 );
nand U12587 ( n13192, n13194, n13195 );
nand U12588 ( n13195, n13196, n11822 );
nand U12589 ( n13194, n13197, n11824 );
not U12590 ( n13197, n13196 );
nor U12591 ( n13196, n10235, n20112 );
nand U12592 ( n6388, n13198, n13199 );
nor U12593 ( n13198, n13200, n13201 );
nor U12594 ( n13201, n20109, n13202 );
nor U12595 ( n13200, n20110, n13184 );
nand U12596 ( n6383, n13203, n13204 );
nor U12597 ( n13204, n13205, n13206 );
nor U12598 ( n13206, n10947, n13207 );
nand U12599 ( n13207, n13208, n13156 );
nor U12600 ( n13208, n13153, n10414 );
not U12601 ( n13153, n13146 );
nand U12602 ( n13146, n20109, n10235 );
nor U12603 ( n13205, n19193, g35 );
nor U12604 ( n13203, n13182, n13209 );
nor U12605 ( n13209, n20109, n13184 );
not U12606 ( n13184, n13202 );
nor U12607 ( n13202, n10947, n13156 );
not U12608 ( n13182, n13199 );
nand U12609 ( n13199, n13210, n13156 );
nor U12610 ( n13210, n11162, n11837 );
nand U12611 ( n11162, n13211, n11662 );
nor U12612 ( n11662, n10405, n20203 );
nor U12613 ( n13211, n12523, n10222 );
nand U12614 ( n6378, n13212, n13213 );
nand U12615 ( n13213, n11017, n10535 );
nand U12616 ( n13212, n13214, g35 );
nand U12617 ( n13214, n13215, n13216 );
nand U12618 ( n13216, n13217, n10829 );
nand U12619 ( n13215, n13218, n13219 );
nand U12620 ( n13219, n19196, n10299 );
not U12621 ( n13218, n13217 );
nand U12622 ( n13217, n13220, n13156 );
not U12623 ( n13156, n13147 );
nand U12624 ( n13147, n13221, n11523 );
nor U12625 ( n11523, n10420, n20198 );
nor U12626 ( n13221, n11850, n13222 );
nor U12627 ( n13222, n20209, n11607 );
not U12628 ( n11607, n11621 );
nor U12629 ( n13220, n20110, n10414 );
nand U12630 ( n6373, n13223, n13224 );
or U12631 ( n13224, n13225, n13226 );
nor U12632 ( n13223, n13227, n13228 );
nor U12633 ( n13228, n19194, g35 );
nor U12634 ( n13227, n10947, n13229 );
nand U12635 ( n13229, n13226, n10535 );
nand U12636 ( n13226, n13230, n13231 );
nor U12637 ( n13230, n19196, n20104 );
nand U12638 ( n6368, n13232, n13233 );
nand U12639 ( n13233, n13234, n13235 );
nor U12640 ( n13232, n13236, n13237 );
nor U12641 ( n13237, n20108, g35 );
nor U12642 ( n13236, n10947, n13238 );
or U12643 ( n13238, n13234, n19194 );
nor U12644 ( n13234, n13239, n10321 );
nand U12645 ( n6363, n13240, n13241 );
or U12646 ( n13241, n13242, n13225 );
nor U12647 ( n13240, n13243, n13244 );
nor U12648 ( n13244, n20107, g35 );
nor U12649 ( n13243, n10947, n13245 );
nand U12650 ( n13245, n13242, n10791 );
nand U12651 ( n13242, n13246, n10390 );
nand U12652 ( n6358, n13247, n13248 );
nand U12653 ( n13248, n13249, n13235 );
nor U12654 ( n13247, n13250, n13251 );
nor U12655 ( n13251, n20106, g35 );
nor U12656 ( n13250, n10947, n13252 );
or U12657 ( n13252, n13249, n20107 );
nor U12658 ( n13249, n13239, n10390 );
nand U12659 ( n6353, n13253, n13254 );
nand U12660 ( n13254, n13255, n13235 );
not U12661 ( n13235, n13225 );
nor U12662 ( n13253, n13256, n13257 );
nor U12663 ( n13257, n20105, g35 );
nor U12664 ( n13256, n10945, n13258 );
or U12665 ( n13258, n13255, n20106 );
and U12666 ( n13255, n13246, n10321 );
nand U12667 ( n6348, n13259, n13260 );
nand U12668 ( n13260, n11018, n10757 );
nor U12669 ( n13259, n13261, n13262 );
nor U12670 ( n13262, n20105, n13124 );
nor U12671 ( n13261, n13129, n13225 );
nand U12672 ( n13225, n13263, g35 );
nor U12673 ( n13263, n13264, n13265 );
nor U12674 ( n13265, n13266, n13267 );
nor U12675 ( n13264, n20061, n13268 );
not U12676 ( n13129, n13121 );
nand U12677 ( n6343, n13269, n13270 );
nand U12678 ( n13270, n13117, n10757 );
nand U12679 ( n13269, n13124, n10536 );
not U12680 ( n13124, n13117 );
nor U12681 ( n13117, n10945, n13121 );
nor U12682 ( n13121, n13271, n13272 );
nand U12683 ( n6338, n13273, n13274 );
nand U12684 ( n13274, n13275, n10536 );
nor U12685 ( n13273, n13276, n13277 );
nor U12686 ( n13277, n10945, n13278 );
nand U12687 ( n13278, n13279, n13280 );
nand U12688 ( n13280, n13281, n13282 );
nor U12689 ( n13281, n13283, n13284 );
nor U12690 ( n13284, n13266, n13285 );
nor U12691 ( n13283, n10338, n13268 );
nor U12692 ( n13279, n13272, n13286 );
nor U12693 ( n13286, n13287, n13282 );
nand U12694 ( n13282, n13271, n10536 );
nand U12695 ( n13271, n19196, n20104 );
nand U12696 ( n13287, n13288, n13289 );
nand U12697 ( n13289, n13266, n10338 );
nand U12698 ( n13288, n13285, n13268 );
not U12699 ( n13285, n13267 );
nand U12700 ( n13267, n12836, n13290 );
nor U12701 ( n13276, n20104, g35 );
nand U12702 ( n6333, n13291, n13292 );
nand U12703 ( n13292, n11018, n10299 );
nor U12704 ( n13291, n13293, n13294 );
nor U12705 ( n13294, n13295, n13239 );
nand U12706 ( n13239, n10299, n13231 );
and U12707 ( n13293, n10390, n13275 );
nand U12708 ( n6328, n13296, n13297 );
nand U12709 ( n13297, n13275, n10299 );
nor U12710 ( n13296, n13298, n13299 );
nor U12711 ( n13299, n10945, n13300 );
nand U12712 ( n13300, n13301, n13302 );
nor U12713 ( n13301, n19196, n13272 );
nor U12714 ( n13298, n20102, g35 );
nand U12715 ( n6323, n13303, n13304 );
nand U12716 ( n13304, n11018, n10321 );
nor U12717 ( n13303, n13305, n13306 );
nor U12718 ( n13306, n13307, n13308 );
nand U12719 ( n13308, n13309, n11572 );
xor U12720 ( n13307, n19565, n13310 );
nor U12721 ( n13310, n20104, n10299 );
nor U12722 ( n13305, n20102, n13311 );
nor U12723 ( n13311, n13312, n11938 );
nor U12724 ( n13312, n13309, n10981 );
and U12725 ( n13309, n13313, n11068 );
nor U12726 ( n13313, n19226, n13314 );
nand U12727 ( n6318, n13315, n13316 );
nand U12728 ( n13316, n13275, n10321 );
nor U12729 ( n13275, n13231, n10985 );
nand U12730 ( n13315, n13317, n13318 );
nor U12731 ( n13318, n13295, n13319 );
nor U12732 ( n13319, n13246, n10321 );
nor U12733 ( n13246, n10299, n13272 );
not U12734 ( n13272, n13231 );
nand U12735 ( n13231, n13266, n13320 );
or U12736 ( n13320, n13314, n19226 );
nor U12737 ( n13314, n13321, n12871 );
not U12738 ( n13266, n13268 );
nand U12739 ( n13268, n13322, n13290 );
nand U12740 ( n13290, n20088, n10322 );
nor U12741 ( n13322, n12873, n13323 );
nor U12742 ( n13323, n10295, n13324 );
nand U12743 ( n13324, n10382, n10237 );
not U12744 ( n13295, n13302 );
nand U12745 ( n13302, n11959, n11068 );
not U12746 ( n11068, n11077 );
nand U12747 ( n11077, n13325, n12877 );
nor U12748 ( n13325, n19996, n10224 );
nor U12749 ( n13317, n10945, n10390 );
nand U12750 ( n6313, n13326, n13327 );
or U12751 ( n13327, n13328, n19550 );
nor U12752 ( n13326, n13329, n13330 );
nor U12753 ( n13330, n10720, n13331 );
nand U12754 ( n13331, n13332, n19198 );
nor U12755 ( n13332, n10945, n13333 );
nor U12756 ( n13329, n19197, n13334 );
nor U12757 ( n13334, n13335, n10985 );
nor U12758 ( n13335, n19198, n13333 );
nand U12759 ( n6308, n13336, n13337 );
nand U12760 ( n13337, n13338, n10720 );
nand U12761 ( n13336, n13328, n10633 );
nand U12762 ( n6303, n13339, n13340 );
nand U12763 ( n13340, n13341, n10633 );
nor U12764 ( n13339, n13342, n13343 );
nor U12765 ( n13343, n19551, g35 );
nor U12766 ( n13342, n10945, n13344 );
nand U12767 ( n13344, n13345, n19198 );
nand U12768 ( n6298, n13346, n13347 );
or U12769 ( n13347, n13348, n19551 );
nor U12770 ( n13346, n13349, n13350 );
nor U12771 ( n13350, n10721, n13351 );
nand U12772 ( n13351, n13352, n20100 );
nor U12773 ( n13352, n10963, n13353 );
nor U12774 ( n13349, n20101, n13354 );
nor U12775 ( n13354, n13355, n10985 );
nor U12776 ( n13355, n20100, n13353 );
nand U12777 ( n6293, n13356, n13357 );
nand U12778 ( n13357, n13341, n10721 );
nand U12779 ( n13356, n13348, n10577 );
nand U12780 ( n6288, n13358, n13359 );
nand U12781 ( n13359, n13338, n10577 );
not U12782 ( n13338, n13328 );
nand U12783 ( n13328, g35, n13333 );
nor U12784 ( n13358, n13360, n13361 );
nor U12785 ( n13361, n19560, g35 );
nor U12786 ( n13360, n10963, n13362 );
or U12787 ( n13362, n10577, n13333 );
nand U12788 ( n6283, n13363, n13364 );
nand U12789 ( n13364, n11018, n10429 );
nand U12790 ( n13363, n13365, g35 );
nand U12791 ( n13365, n13366, n13367 );
or U12792 ( n13367, n13368, n19560 );
nand U12793 ( n13366, n13369, n13368 );
nor U12794 ( n13368, n13370, n13371 );
xnor U12795 ( n13369, n10429, n19207 );
nand U12796 ( n6278, n13372, n13373 );
nand U12797 ( n13373, n13374, g35 );
nor U12798 ( n13374, n19199, n13375 );
nor U12799 ( n13375, n13376, n13371 );
nor U12800 ( n13376, n13377, n10696 );
nand U12801 ( n13372, n13378, n10696 );
nand U12802 ( n13378, g35, n13379 );
nand U12803 ( n13379, n13380, n13381 );
nand U12804 ( n13381, n10429, n13370 );
nand U12805 ( n6273, n13382, n13383 );
nand U12806 ( n13383, n11018, n10348 );
nand U12807 ( n13382, g35, n13384 );
nand U12808 ( n13384, n13385, n13386 );
or U12809 ( n13386, n13333, n20093 );
nand U12810 ( n13333, n13387, n13380 );
nor U12811 ( n13387, n20095, n20098 );
nor U12812 ( n13385, n13388, n13389 );
nor U12813 ( n13389, n13390, n13371 );
nor U12814 ( n13390, n13391, n13392 );
nand U12815 ( n13392, n13393, n13394 );
nand U12816 ( n13394, n13377, n10793 );
nand U12817 ( n13393, g25167, n10912 );
nand U12818 ( n13391, n13395, n13396 );
nand U12819 ( n13396, n13397, n20095 );
nor U12820 ( n13397, n19203, n10348 );
nand U12821 ( n13395, n20096, n13398 );
nand U12822 ( n13398, n13399, n13400 );
or U12823 ( n13400, n20098, n19205 );
or U12824 ( n13399, n20095, n19204 );
nor U12825 ( n13388, n20099, n13380 );
nand U12826 ( n6268, n13401, n13402 );
nor U12827 ( n13402, n13403, n13404 );
nor U12828 ( n13404, n10963, n13405 );
nand U12829 ( n13405, n13380, n10350 );
nor U12830 ( n13403, n20097, g35 );
nor U12831 ( n13401, n13406, n13407 );
nor U12832 ( n13407, n20098, n13408 );
nand U12833 ( n6263, n13409, n13410 );
nand U12834 ( n13410, n11019, n10350 );
nor U12835 ( n13409, n13411, n13412 );
nor U12836 ( n13412, n20097, n13413 );
nor U12837 ( n13413, n13414, n13415 );
nand U12838 ( n13415, n13408, n11547 );
not U12839 ( n11547, n11938 );
nor U12840 ( n13414, n11137, n10985 );
nor U12841 ( n13411, n13416, n13417 );
nand U12842 ( n13417, n13380, n11137 );
nand U12843 ( n13416, n13418, n13419 );
nand U12844 ( n13419, n13420, n11822 );
nand U12845 ( n11822, n19200, n11572 );
nand U12846 ( n13418, n13421, n11824 );
or U12847 ( n11824, n13422, n19200 );
not U12848 ( n13421, n13420 );
nor U12849 ( n13420, n10350, n20098 );
nand U12850 ( n6258, n13423, n13424 );
nor U12851 ( n13423, n13425, n13426 );
nor U12852 ( n13426, n20095, n13427 );
nor U12853 ( n13425, n20096, n13408 );
nand U12854 ( n6253, n13428, n13429 );
nor U12855 ( n13429, n13430, n13431 );
nor U12856 ( n13431, n10963, n13432 );
nand U12857 ( n13432, n13433, n13380 );
nor U12858 ( n13433, n13377, n10348 );
not U12859 ( n13377, n13370 );
nand U12860 ( n13370, n20095, n10350 );
nor U12861 ( n13430, n19202, g35 );
nor U12862 ( n13428, n13406, n13434 );
nor U12863 ( n13434, n20095, n13408 );
not U12864 ( n13408, n13427 );
nor U12865 ( n13427, n10963, n13380 );
not U12866 ( n13406, n13424 );
nand U12867 ( n13424, n13435, n13380 );
nor U12868 ( n13435, n13436, n11837 );
nand U12869 ( n11837, n13437, n13438 );
nor U12870 ( n13437, n19200, n10984 );
not U12871 ( n13436, n11137 );
nor U12872 ( n11137, n11606, n12523 );
nand U12873 ( n12523, n13439, n13440 );
xnor U12874 ( n13440, n20206, n19562 );
xnor U12875 ( n13439, n19201, n19563 );
nand U12876 ( n6248, n13441, n13442 );
nand U12877 ( n13442, n11019, n10792 );
nand U12878 ( n13441, n13443, g35 );
nand U12879 ( n13443, n13444, n13445 );
nand U12880 ( n13445, n13446, n10830 );
nand U12881 ( n13444, n13447, n13448 );
nand U12882 ( n13448, n19208, n10316 );
not U12883 ( n13447, n13446 );
nand U12884 ( n13446, n13380, g25167 );
nor U12885 ( g25167, n10348, n20096 );
not U12886 ( n13380, n13371 );
nand U12887 ( n13371, n12533, n13449 );
nand U12888 ( n13449, n11621, n10369 );
and U12889 ( n12533, n13450, n20199 );
nor U12890 ( n13450, n11850, n10225 );
and U12891 ( n11850, n11621, n13451 );
or U12892 ( n13451, n11606, n20202 );
nand U12893 ( n11606, n13452, n20205 );
nor U12894 ( n13452, n10231, n10222 );
nor U12895 ( n11621, n10332, n10228 );
nand U12896 ( n6243, n13453, n13454 );
or U12897 ( n13454, n13455, n13456 );
nor U12898 ( n13453, n13457, n13458 );
nor U12899 ( n13458, n19204, g35 );
nor U12900 ( n13457, n10961, n13459 );
nand U12901 ( n13459, n13456, n10792 );
nand U12902 ( n13456, n13460, n10442 );
nand U12903 ( n6238, n13461, n13462 );
nand U12904 ( n13462, n13463, n13464 );
nor U12905 ( n13461, n13465, n13466 );
nor U12906 ( n13466, n20094, g35 );
nor U12907 ( n13465, n10961, n13467 );
or U12908 ( n13467, n13463, n19204 );
nor U12909 ( n13463, n13468, n10357 );
nand U12910 ( n6233, n13469, n13470 );
nand U12911 ( n13470, n13471, n13464 );
nor U12912 ( n13469, n13472, n13473 );
nor U12913 ( n13473, n19205, g35 );
nor U12914 ( n13472, n10961, n13474 );
or U12915 ( n13474, n13471, n20094 );
nor U12916 ( n13471, n13475, n13476 );
not U12917 ( n13475, g25259 );
nand U12918 ( n6228, n13477, n13478 );
nand U12919 ( n13478, n13479, n13464 );
not U12920 ( n13464, n13455 );
nor U12921 ( n13477, n13480, n13481 );
nor U12922 ( n13481, n19206, g35 );
nor U12923 ( n13480, n10961, n13482 );
or U12924 ( n13482, n13479, n19205 );
nor U12925 ( n13479, n13468, n10442 );
nand U12926 ( n6223, n13483, n13484 );
or U12927 ( n13484, n13485, n13455 );
nor U12928 ( n13483, n13486, n13487 );
nor U12929 ( n13487, n20093, g35 );
nor U12930 ( n13486, n10960, n13488 );
nand U12931 ( n13488, n13485, n10793 );
nand U12932 ( n13485, n13460, n20091 );
nand U12933 ( n6218, n13489, n13490 );
nand U12934 ( n13490, n11019, n10758 );
nor U12935 ( n13489, n13491, n13492 );
nor U12936 ( n13492, n20093, n13348 );
nor U12937 ( n13491, n13353, n13455 );
nand U12938 ( n13455, n13493, g35 );
nor U12939 ( n13493, n13494, n13495 );
nor U12940 ( n13495, g23683, n13496 );
nor U12941 ( n13494, n13497, n13498 );
not U12942 ( n13353, n13345 );
nand U12943 ( n6213, n13499, n13500 );
nand U12944 ( n13500, n13341, n10758 );
nand U12945 ( n13499, n13348, n10537 );
not U12946 ( n13348, n13341 );
nor U12947 ( n13341, n10960, n13345 );
nor U12948 ( n13345, n13501, n13476 );
nand U12949 ( n6208, n13502, n13503 );
nand U12950 ( n13503, n13504, n10537 );
nor U12951 ( n13502, n13505, n13506 );
nor U12952 ( n13506, n10960, n13507 );
nand U12953 ( n13507, n13508, n13509 );
nand U12954 ( n13509, n13510, n13511 );
nor U12955 ( n13510, n13512, n13513 );
nor U12956 ( n13513, n13497, n13514 );
nor U12957 ( n13512, n20062, n13496 );
nor U12958 ( n13508, n13476, n13515 );
nor U12959 ( n13515, n13516, n13511 );
nand U12960 ( n13511, n13501, n10537 );
nand U12961 ( n13501, n19208, n20092 );
nand U12962 ( n13516, n13517, n13518 );
nand U12963 ( n13518, n13514, n13496 );
not U12964 ( n13514, n13498 );
nand U12965 ( n13498, n12836, n13519 );
nor U12966 ( n12836, n19951, n12873 );
nand U12967 ( n13517, n13497, n20062 );
not U12968 ( n13497, n13496 );
nor U12969 ( n13505, n20092, g35 );
nand U12970 ( n6203, n13520, n13521 );
nand U12971 ( n13521, n11019, n10316 );
nor U12972 ( n13520, n13522, n13523 );
nor U12973 ( n13523, n13524, n13468 );
or U12974 ( n13468, n20091, n13476 );
nor U12975 ( n13522, n20092, n13525 );
nand U12976 ( n6198, n13526, n13527 );
nand U12977 ( n13527, n13504, n10316 );
nor U12978 ( n13526, n13528, n13529 );
nor U12979 ( n13529, n10960, n13530 );
nand U12980 ( n13530, n13460, n13531 );
nor U12981 ( n13460, n19208, n13476 );
nor U12982 ( n13528, n20090, g35 );
nand U12983 ( n6193, n13532, n13533 );
nand U12984 ( n13533, n11019, n10357 );
nor U12985 ( n13532, n13534, n13535 );
nor U12986 ( n13535, n20090, n13536 );
nor U12987 ( n13536, n13537, n11938 );
nor U12988 ( n11938, n10960, n13438 );
nor U12989 ( n13537, n13538, n10984 );
and U12990 ( n13538, n11066, g27831 );
nor U12991 ( n13534, n13539, n13540 );
nand U12992 ( n13540, n13541, g27831 );
xnor U12993 ( n13541, g25259, n19565 );
nor U12994 ( g25259, n10316, n20092 );
nand U12995 ( n13539, n11572, n11066 );
nand U12996 ( n6188, n13542, n13543 );
nand U12997 ( n13543, n13504, n10357 );
not U12998 ( n13504, n13525 );
nand U12999 ( n13525, n13476, g35 );
nand U13000 ( n13542, n13544, n13545 );
nor U13001 ( n13545, n13524, n13546 );
nor U13002 ( n13546, n13547, n10357 );
nor U13003 ( n13547, n13476, n10316 );
nor U13004 ( n13476, n13496, g27831 );
nor U13005 ( g27831, n13548, n20059 );
and U13006 ( n13548, n13099, n13549 );
not U13007 ( n13099, n12871 );
nand U13008 ( n12871, n13550, n13551 );
nor U13009 ( n13551, n10659, n13552 );
nand U13010 ( n13552, n10641, n10285 );
nor U13011 ( n13550, n10479, n13553 );
nand U13012 ( n13553, n19222, n19223 );
nand U13013 ( n13496, n13554, n13519 );
nand U13014 ( n13519, n20088, n10454 );
nor U13015 ( n13554, n12873, n13555 );
nor U13016 ( n13555, n10295, n13556 );
nand U13017 ( n13556, n20142, n10237 );
and U13018 ( n12873, n19567, n13557 );
nand U13019 ( n13557, n11424, n11419 );
nor U13020 ( n11424, n10252, n19991 );
not U13021 ( n13524, n13531 );
nand U13022 ( n13531, n11959, n11066 );
and U13023 ( n11066, n13558, n12877 );
not U13024 ( n12877, n11223 );
nand U13025 ( n11223, n13559, n19998 );
nor U13026 ( n13559, n12644, n12643 );
xnor U13027 ( n12643, n19270, g73 );
xnor U13028 ( n12644, n19999, g72 );
nor U13029 ( n13558, n10224, n10404 );
nor U13030 ( n11959, n13560, n19565 );
nor U13031 ( n13544, n10960, n10442 );
nand U13032 ( n6173, n13561, n13562 );
nand U13033 ( n13562, n11020, n10784 );
nand U13034 ( n13561, g35, n13563 );
nand U13035 ( n13563, n19323, n11419 );
nand U13036 ( n6168, n13564, n13565 );
or U13037 ( n13565, g35, n20089 );
nand U13038 ( n13564, g35, n13566 );
nand U13039 ( n13566, n19209, n19332 );
nand U13040 ( n6163, n13567, n13568 );
nand U13041 ( n13568, n11020, n10586 );
nand U13042 ( n13567, g35, n13569 );
nand U13043 ( n13569, n20089, n10381 );
nor U13044 ( n6158, n20088, n10984 );
nand U13045 ( n6153, n13570, n13571 );
nand U13046 ( n13571, n20087, n13572 );
nor U13047 ( n13570, n13573, n13574 );
nor U13048 ( n13574, n19210, g35 );
nor U13049 ( n13573, n10960, n13575 );
or U13050 ( n13575, n13572, n20087 );
nor U13051 ( n13572, n13576, n13577 );
or U13052 ( n13576, n19210, n13578 );
nand U13053 ( n6148, n13579, n13580 );
nand U13054 ( n13580, n11020, n10452 );
nand U13055 ( n13579, n13581, g35 );
nor U13056 ( n13581, n13582, n13583 );
nor U13057 ( n13583, n13584, n10913 );
nor U13058 ( n13584, n13577, n13585 );
nor U13059 ( n13582, n13586, n13577 );
xnor U13060 ( n13586, n20087, n13587 );
nand U13061 ( n6143, n13588, n13589 );
nand U13062 ( n13589, n20086, n13590 );
nor U13063 ( n13588, n13591, n13592 );
nor U13064 ( n13592, n19211, g35 );
nor U13065 ( n13591, n10960, n13593 );
or U13066 ( n13593, n13590, n20086 );
nor U13067 ( n13590, n13594, n13595 );
or U13068 ( n13594, n19211, n13578 );
nand U13069 ( n6138, n13596, n13597 );
nand U13070 ( n13597, n11020, n10322 );
nand U13071 ( n13596, n13598, g35 );
nor U13072 ( n13598, n13599, n13600 );
nor U13073 ( n13600, n13601, n10914 );
nor U13074 ( n13601, n13585, n13595 );
nor U13075 ( n13599, n13602, n13595 );
nand U13076 ( n13595, n13603, n10294 );
nor U13077 ( n13603, n19218, n20067 );
xnor U13078 ( n13602, n20086, n13587 );
nand U13079 ( n6133, n13604, n13605 );
or U13080 ( n13605, n10322, n13606 );
nor U13081 ( n13604, n13607, n13608 );
nor U13082 ( n13608, n19212, g35 );
nor U13083 ( n13607, n10959, n13609 );
nand U13084 ( n13609, n13606, n10322 );
nand U13085 ( n13606, n13610, n13611 );
nor U13086 ( n13610, n19212, n13578 );
nand U13087 ( n6128, n13612, n13613 );
nand U13088 ( n13613, n11021, n10454 );
nand U13089 ( n13612, n13614, g35 );
nor U13090 ( n13614, n13615, n13616 );
nor U13091 ( n13616, n13617, n10908 );
nor U13092 ( n13617, n13585, n13618 );
nor U13093 ( n13615, n13619, n13618 );
not U13094 ( n13618, n13611 );
nor U13095 ( n13611, n13321, n19218 );
xnor U13096 ( n13619, n20085, n13587 );
nand U13097 ( n6123, n13620, n13621 );
nand U13098 ( n13621, n20084, n13622 );
nor U13099 ( n13620, n13623, n13624 );
nor U13100 ( n13624, n19213, g35 );
nor U13101 ( n13623, n10958, n13625 );
or U13102 ( n13625, n13622, n20084 );
nor U13103 ( n13622, n13626, n13627 );
or U13104 ( n13626, n19213, n13578 );
nand U13105 ( n13578, n20083, n10370 );
nand U13106 ( n6118, n13628, n13629 );
nand U13107 ( n13629, n11021, n10370 );
nand U13108 ( n13628, n13630, g35 );
nor U13109 ( n13630, n13631, n13632 );
nor U13110 ( n13632, n13633, n10915 );
nor U13111 ( n13633, n13585, n13627 );
nand U13112 ( n13585, n19215, n20082 );
nor U13113 ( n13631, n13634, n13627 );
nand U13114 ( n13627, n13549, g13259 );
nor U13115 ( n13549, n10294, n20067 );
xnor U13116 ( n13634, n20084, n13587 );
and U13117 ( n13587, n19214, n11419 );
nand U13118 ( n6113, n13635, n13636 );
nand U13119 ( n13636, n13637, n10370 );
nand U13120 ( n13635, n13638, n10667 );
nand U13121 ( n6108, n13639, n13640 );
nand U13122 ( n13640, n13637, n10667 );
or U13123 ( n13639, n13637, n20082 );
not U13124 ( n13637, n13638 );
nand U13125 ( n13638, g35, n13577 );
nor U13126 ( n6103, n13641, n10983 );
nor U13127 ( n13641, n13642, n13643 );
nor U13128 ( n13643, n13577, n10370 );
nor U13129 ( n13642, n20082, n13644 );
nor U13130 ( n13644, n20083, n13577 );
nand U13131 ( n13577, n13645, n20067 );
nor U13132 ( n13645, n19218, n10294 );
nand U13133 ( n6098, n13646, n13647 );
nand U13134 ( n13647, n13648, g35 );
nor U13135 ( n13648, n20081, n13649 );
nor U13136 ( n13649, n13650, n13651 );
nor U13137 ( n13650, n20075, n10518 );
nand U13138 ( n13646, n13652, n10518 );
nand U13139 ( n13652, g35, n13653 );
nand U13140 ( n13653, n13654, n20081 );
nand U13141 ( n6093, n13655, n13656 );
nand U13142 ( n13656, n11020, n10637 );
nand U13143 ( n13655, n13657, g35 );
nand U13144 ( n13657, n13658, n13659 );
nand U13145 ( n13659, n13651, n10518 );
nand U13146 ( n13658, n13654, n20080 );
nor U13147 ( n13654, n20075, n13651 );
nand U13148 ( n6088, n13660, n13661 );
nand U13149 ( n13661, n13662, g35 );
nor U13150 ( n13662, n19217, n13663 );
nor U13151 ( n13663, n13664, n13665 );
nor U13152 ( n13664, n13666, n10317 );
nand U13153 ( n13660, n13667, n10317 );
nand U13154 ( n13667, g35, n13668 );
nand U13155 ( n13668, n13669, n19217 );
nor U13156 ( n13669, n13666, n13665 );
nand U13157 ( n6083, n13670, n13671 );
nand U13158 ( n13671, n13672, n13673 );
nor U13159 ( n13672, n10317, n13665 );
nor U13160 ( n13670, n13674, n13675 );
nor U13161 ( n13675, n20078, g35 );
nor U13162 ( n13674, n10957, n13676 );
nand U13163 ( n13676, n13665, n10317 );
nand U13164 ( n13665, n13677, n13678 );
nand U13165 ( n13678, n20078, n13679 );
not U13166 ( n13677, n13680 );
nand U13167 ( n6078, n13681, n13682 );
nand U13168 ( n13682, n13683, n13673 );
nor U13169 ( n13683, n10393, n13680 );
nor U13170 ( n13681, n13684, n13685 );
nor U13171 ( n13685, n20077, g35 );
nor U13172 ( n13684, n10957, n13686 );
nand U13173 ( n13686, n13680, n10393 );
nand U13174 ( n13680, n13687, n13688 );
nand U13175 ( n13688, n20077, n13679 );
nand U13176 ( n6073, n13689, n13690 );
nand U13177 ( n13690, n13691, g35 );
nor U13178 ( n13691, n20077, n13687 );
and U13179 ( n13687, n13692, n13693 );
nand U13180 ( n13693, n20076, n13679 );
not U13181 ( n13679, n13666 );
nand U13182 ( n13689, n13694, n10257 );
nand U13183 ( n13694, g35, n13695 );
nand U13184 ( n13695, n13696, n20077 );
nor U13185 ( n13696, n13697, n13666 );
nand U13186 ( n6068, n13698, n13699 );
nand U13187 ( n13699, n13700, n13673 );
nor U13188 ( n13673, n13666, n10983 );
nand U13189 ( n13666, n13701, n20074 );
nor U13190 ( n13701, n13702, n13703 );
nor U13191 ( n13703, n13704, n13705 );
nor U13192 ( n13702, n13706, n13707 );
nor U13193 ( n13706, n20075, n10617 );
nor U13194 ( n13700, n13697, n10257 );
nor U13195 ( n13698, n13708, n13709 );
nor U13196 ( n13709, n20075, g35 );
nor U13197 ( n13708, n10957, n13710 );
nand U13198 ( n13710, n13697, n10257 );
nand U13199 ( n6063, n13711, n13712 );
nand U13200 ( n13712, n13713, n10606 );
nand U13201 ( n13713, g35, n13651 );
nand U13202 ( n13711, n13714, n13715 );
nor U13203 ( n13715, n20075, n13716 );
nor U13204 ( n13716, n13697, n13717 );
or U13205 ( n13717, n20079, n20077 );
nor U13206 ( n13714, n13718, n10983 );
nor U13207 ( n13718, n20081, n13651 );
nor U13208 ( n6058, n10957, n13719 );
nand U13209 ( n13719, n13720, n13721 );
nand U13210 ( n13721, n13722, n13692 );
nor U13211 ( n13722, n13723, n13724 );
nor U13212 ( n13724, n13725, n13705 );
nor U13213 ( n13725, n10606, n13726 );
nand U13214 ( n13726, n13727, n13704 );
nand U13215 ( n13727, n13728, n13729 );
nor U13216 ( n13729, n19217, n20076 );
and U13217 ( n13728, n10393, n20075 );
nor U13218 ( n13723, n10617, n13704 );
nand U13219 ( n13704, n13730, n10317 );
nor U13220 ( n13730, n20075, n20077 );
nand U13221 ( n13720, n13697, n20074 );
nand U13222 ( n6053, n13731, n13732 );
nand U13223 ( n13732, g35, n13733 );
nand U13224 ( n13733, g19334, n13734 );
nand U13225 ( n13734, n20073, n13735 );
nand U13226 ( n13735, n20072, g12919 );
nand U13227 ( n13731, n13736, n10641 );
nand U13228 ( n13736, n20060, g35 );
nand U13229 ( n6048, n13737, n13738 );
nand U13230 ( n13738, n13739, n20066 );
nor U13231 ( n13739, n13740, n13741 );
nor U13232 ( n13741, n13742, n13743 );
nor U13233 ( n13743, n20073, n10982 );
not U13234 ( n13742, n13744 );
nor U13235 ( n13740, n20073, n13744 );
nand U13236 ( n13744, n13745, n10416 );
nand U13237 ( n13737, n11021, n10416 );
nor U13238 ( n6043, n13746, n13747 );
nand U13239 ( n13747, n20066, g35 );
xnor U13240 ( n13746, n10416, n13745 );
and U13241 ( n13745, g12919, n13748 );
nand U13242 ( n13748, n13749, n19219 );
nor U13243 ( n13749, n10400, g7916 );
nand U13244 ( n6038, n13750, n13751 );
nand U13245 ( n13751, n13752, n13753 );
nor U13246 ( n13752, n13754, n13755 );
nor U13247 ( n13755, n13756, n13757 );
nor U13248 ( n13757, n19216, n10982 );
not U13249 ( n13756, n13758 );
nor U13250 ( n13754, n19216, n13758 );
nand U13251 ( n13750, n11021, n10418 );
nand U13252 ( n6033, n13759, n13760 );
nand U13253 ( n13760, n11021, n10675 );
nand U13254 ( n13759, n13761, g35 );
nor U13255 ( n13761, n13762, n13763 );
xnor U13256 ( n13763, n10418, n13764 );
nand U13257 ( n6028, n13765, n13766 );
nand U13258 ( n13766, n11021, n10360 );
nand U13259 ( n13765, g35, n13767 );
nand U13260 ( n13767, n13768, n13769 );
nand U13261 ( n13769, n13770, n10675 );
or U13262 ( n13770, n13758, n19216 );
nand U13263 ( n13758, n13764, n10418 );
and U13264 ( n13764, n13771, n13772 );
nor U13265 ( n13771, n20064, n13773 );
nor U13266 ( n13773, n10360, n13774 );
nand U13267 ( n13774, n10387, n10239 );
nand U13268 ( n6023, n13775, n13776 );
nand U13269 ( n13776, n11021, n10381 );
nand U13270 ( n13775, n13777, g35 );
nand U13271 ( n13777, n13778, n13779 );
nand U13272 ( n13779, n10387, g7916 );
nand U13273 ( n13778, n20064, n10360 );
nand U13274 ( n6018, n13780, n13781 );
nand U13275 ( n13781, n11022, n10387 );
nand U13276 ( n13780, n13782, g35 );
nand U13277 ( n13782, n13783, n13784 );
or U13278 ( n13784, n13785, n20063 );
nand U13279 ( n13783, n13785, n10381 );
nand U13280 ( n13785, n13786, n10294 );
nor U13281 ( n13786, n20064, n20067 );
nand U13282 ( n6013, n13787, n13788 );
nand U13283 ( n13788, n11022, n10294 );
nand U13284 ( n13787, n13789, g35 );
nand U13285 ( n13789, n13790, n13791 );
nand U13286 ( n13790, n20064, n10387 );
nand U13287 ( n6008, n13792, n13793 );
nand U13288 ( n13793, g35, n13794 );
nand U13289 ( n13794, n13321, n13753 );
not U13290 ( n13753, n13762 );
not U13291 ( n13321, n13772 );
nand U13292 ( n13792, n13795, n10580 );
nand U13293 ( n13795, n13796, g35 );
xnor U13294 ( n13796, n20068, n20064 );
nor U13295 ( n6003, n13797, n10982 );
nor U13296 ( n13797, n13762, n13798 );
xnor U13297 ( n13798, g7916, n20067 );
nor U13298 ( n13762, n13768, n13799 );
nor U13299 ( n13799, n20071, n13772 );
nor U13300 ( n13772, n10580, n20068 );
nand U13301 ( n13768, n13800, n13801 );
nor U13302 ( n13801, n20069, n13791 );
nand U13303 ( n13791, g7916, n10239 );
nor U13304 ( n13800, n13802, n10360 );
nor U13305 ( n13802, n13803, n13804 );
nor U13306 ( n13803, n13805, n13806 );
nand U13307 ( n13806, n13707, n10393 );
not U13308 ( n13707, n13705 );
nand U13309 ( n13805, n10257, n10637 );
xnor U13310 ( n5990, n13807, n10400 );
or U13311 ( n13807, n13808, n11024 );
nand U13312 ( n5977, n13809, n13810 );
nand U13313 ( n13810, n11022, n10239 );
nand U13314 ( n13809, n13811, g35 );
xor U13315 ( n13811, n13808, n13812 );
nand U13316 ( n13812, n13813, n13814 );
nor U13317 ( n13814, g19334, n13815 );
nand U13318 ( n13815, n20064, n20065 );
nor U13319 ( n13813, g13259, g8416 );
nand U13320 ( n13808, n13816, n13817 );
nor U13321 ( n13816, n13818, n13651 );
xnor U13322 ( n13818, n19220, n20066 );
nand U13323 ( n5972, n13819, n13820 );
or U13324 ( n13820, g35, n19220 );
nand U13325 ( n5963, n13821, n13822 );
nand U13326 ( n13822, n13823, g17400 );
nor U13327 ( n13821, n13824, n13825 );
nor U13328 ( n13825, n20062, g35 );
nor U13329 ( n13824, n10957, n13826 );
nand U13330 ( n13826, n19227, g10500 );
nand U13331 ( n5958, n13819, n13827 );
nand U13332 ( n13827, n11022, g23683 );
nand U13333 ( n5949, n13828, n13829 );
nand U13334 ( n13829, g35, g20901 );
nand U13335 ( n13828, n11022, n10448 );
nand U13336 ( n5944, n13830, n13831 );
nand U13337 ( n13831, n13832, g35 );
nor U13338 ( n13832, n19222, n13833 );
nand U13339 ( n13830, n13834, n10479 );
nand U13340 ( n13834, g35, n13835 );
nand U13341 ( n13835, n13833, n19222 );
nand U13342 ( n5939, n13836, n13837 );
nand U13343 ( n13837, n11022, n10619 );
nand U13344 ( n13836, n13838, g35 );
nand U13345 ( n13838, n13839, n13840 );
nand U13346 ( n13840, n13841, n10479 );
nand U13347 ( n13839, n13842, n19221 );
nor U13348 ( n13842, n10448, n13841 );
nand U13349 ( n5934, n13843, n13844 );
nand U13350 ( n13844, n13845, n19223 );
nor U13351 ( n13843, n13846, n13847 );
nor U13352 ( n13847, n19224, g35 );
nor U13353 ( n13846, n10957, n13848 );
nand U13354 ( n13848, n13849, n10619 );
xnor U13355 ( n5929, n13850, n10589 );
nand U13356 ( n13850, g35, n10659 );
nor U13357 ( n5912, n13851, n13852 );
nand U13358 ( n13852, n19226, n20059 );
nand U13359 ( n13851, n13853, n19227 );
nor U13360 ( n13853, n13854, n10982 );
nor U13361 ( n13854, n13841, n13855 );
nand U13362 ( n13855, n13856, n10448 );
or U13363 ( n13856, n13804, n13651 );
nand U13364 ( n13651, n13705, n13692 );
not U13365 ( n13692, n13697 );
nor U13366 ( n13697, n10400, n10285 );
xnor U13367 ( n13705, n20066, n10239 );
not U13368 ( n13841, n13833 );
nor U13369 ( n13833, n13849, n19223 );
not U13370 ( n13849, n13845 );
nor U13371 ( n13845, n19224, n19225 );
nor U13372 ( n5907, n20058, n13857 );
nor U13373 ( n13857, n13858, n10982 );
nor U13374 ( n13858, n11419, n13859 );
nand U13375 ( n5902, n13860, n13861 );
nand U13376 ( n13861, n11023, n10520 );
nor U13377 ( n13860, n13862, n13863 );
nor U13378 ( n13863, n13859, n10909 );
nor U13379 ( n13862, n20058, n13864 );
nand U13380 ( n13864, n13823, n13859 );
nand U13381 ( n13859, n13865, n10520 );
nand U13382 ( n5897, n13866, n13867 );
nand U13383 ( n13867, n11022, n10678 );
nor U13384 ( n13866, n13868, n13869 );
nor U13385 ( n13869, n13870, n10520 );
nor U13386 ( n13868, n20057, n13871 );
nand U13387 ( n13871, n13823, n13870 );
not U13388 ( n13870, n13865 );
nor U13389 ( n13865, n13872, n20056 );
nand U13390 ( n5892, n13873, n13874 );
nand U13391 ( n13874, n11023, n10741 );
nor U13392 ( n13873, n13875, n13876 );
nor U13393 ( n13876, n13872, n10678 );
nor U13394 ( n13875, n20056, n13877 );
nand U13395 ( n13877, n13823, n13872 );
or U13396 ( n13872, n13878, n20055 );
nand U13397 ( n5887, n13879, n13880 );
nand U13398 ( n13880, n11023, n10742 );
nor U13399 ( n13879, n13881, n13882 );
nor U13400 ( n13882, n13878, n10741 );
nor U13401 ( n13881, n20055, n13883 );
nand U13402 ( n13883, n13823, n13878 );
or U13403 ( n13878, n13884, n20054 );
nand U13404 ( n5882, n13885, n13886 );
nand U13405 ( n13886, n11023, n10743 );
nor U13406 ( n13885, n13887, n13888 );
nor U13407 ( n13888, n13884, n10742 );
nor U13408 ( n13887, n20054, n13889 );
nand U13409 ( n13889, n13823, n13884 );
or U13410 ( n13884, n13890, n20053 );
nand U13411 ( n5877, n13891, n13892 );
nand U13412 ( n13892, n11023, n10654 );
nor U13413 ( n13891, n13893, n13894 );
nor U13414 ( n13894, n13890, n10743 );
nor U13415 ( n13893, n20053, n13895 );
nand U13416 ( n13895, n13823, n13890 );
nand U13417 ( n13890, n13896, n13897 );
nor U13418 ( n13896, n19229, n20052 );
nand U13419 ( n5872, n13898, n13899 );
nand U13420 ( n13899, n11022, n10668 );
nor U13421 ( n13898, n13900, n13901 );
nor U13422 ( n13901, n10654, n13902 );
nand U13423 ( n13902, n13897, n10482 );
nor U13424 ( n13900, n20052, n13903 );
nor U13425 ( n13903, n13904, n5862 );
nor U13426 ( n13904, n13897, n13819 );
nor U13427 ( n13897, n19228, n20060 );
nand U13428 ( n5867, n13905, n13906 );
nand U13429 ( n13906, n13907, n10482 );
nand U13430 ( n13907, g35, n13908 );
nand U13431 ( n13908, n19228, g12919 );
nand U13432 ( n13905, n5862, n10668 );
nor U13433 ( n5862, n10482, n13819 );
not U13434 ( n13819, n13823 );
nor U13435 ( n13823, n10956, n20060 );
nand U13436 ( n5847, n13909, n13910 );
nand U13437 ( n13910, n11023, n10785 );
nand U13438 ( n13909, g35, n13911 );
nand U13439 ( n13911, n19324, n11418 );
nand U13440 ( n5842, n13912, n13913 );
or U13441 ( n13913, g35, n20051 );
nand U13442 ( n13912, g35, n13914 );
nand U13443 ( n13914, n19230, n19333 );
nand U13444 ( n5837, n13915, n13916 );
nand U13445 ( n13916, n11023, n10587 );
nand U13446 ( n13915, g35, n13917 );
nand U13447 ( n13917, n20051, n10492 );
nor U13448 ( n5832, n20050, n10982 );
nand U13449 ( n5827, n13918, n13919 );
nand U13450 ( n13919, n20049, n13920 );
nor U13451 ( n13918, n13921, n13922 );
nor U13452 ( n13922, n19231, g35 );
nor U13453 ( n13921, n10956, n13923 );
or U13454 ( n13923, n13920, n20049 );
nor U13455 ( n13920, n13924, n13925 );
or U13456 ( n13924, n19231, n13926 );
nand U13457 ( n5822, n13927, n13928 );
nand U13458 ( n13928, n11023, n10453 );
nand U13459 ( n13927, n13929, g35 );
nor U13460 ( n13929, n13930, n13931 );
nor U13461 ( n13931, n13932, n10916 );
nor U13462 ( n13932, n13925, n13933 );
nor U13463 ( n13930, n13934, n13925 );
xnor U13464 ( n13934, n20049, n13935 );
nand U13465 ( n5817, n13936, n13937 );
nand U13466 ( n13937, n20048, n13938 );
nor U13467 ( n13936, n13939, n13940 );
nor U13468 ( n13940, n19232, g35 );
nor U13469 ( n13939, n10956, n13941 );
or U13470 ( n13941, n13938, n20048 );
nor U13471 ( n13938, n13942, n13943 );
or U13472 ( n13942, n19232, n13926 );
nand U13473 ( n5812, n13944, n13945 );
nand U13474 ( n13945, n11023, n10323 );
nand U13475 ( n13944, n13946, g35 );
nor U13476 ( n13946, n13947, n13948 );
nor U13477 ( n13948, n13949, n10917 );
nor U13478 ( n13949, n13933, n13943 );
nor U13479 ( n13947, n13950, n13943 );
nand U13480 ( n13943, n13951, n10303 );
xnor U13481 ( n13950, n20048, n13935 );
nand U13482 ( n5807, n13952, n13953 );
or U13483 ( n13953, n10323, n13954 );
nor U13484 ( n13952, n13955, n13956 );
nor U13485 ( n13956, n19233, g35 );
nor U13486 ( n13955, n10956, n13957 );
nand U13487 ( n13957, n13954, n10323 );
nand U13488 ( n13954, n13958, n13959 );
nor U13489 ( n13958, n19233, n13926 );
nand U13490 ( n5802, n13960, n13961 );
nand U13491 ( n13961, n11023, n10455 );
nand U13492 ( n13960, n13962, g35 );
nor U13493 ( n13962, n13963, n13964 );
nor U13494 ( n13964, n13965, n10910 );
nor U13495 ( n13965, n13933, n13966 );
nor U13496 ( n13963, n13967, n13966 );
not U13497 ( n13966, n13959 );
nor U13498 ( n13959, n12408, n19239 );
xnor U13499 ( n13967, n20047, n13935 );
nand U13500 ( n5797, n13968, n13969 );
nand U13501 ( n13969, n20046, n13970 );
nor U13502 ( n13968, n13971, n13972 );
nor U13503 ( n13972, n19234, g35 );
nor U13504 ( n13971, n10956, n13973 );
or U13505 ( n13973, n13970, n20046 );
nor U13506 ( n13970, n13974, n13975 );
or U13507 ( n13974, n19234, n13926 );
nand U13508 ( n13926, n20045, n10371 );
nand U13509 ( n5792, n13976, n13977 );
nand U13510 ( n13977, n11011, n10371 );
nand U13511 ( n13976, n13978, g35 );
nor U13512 ( n13978, n13979, n13980 );
nor U13513 ( n13980, n13981, n10918 );
nor U13514 ( n13981, n13933, n13975 );
nand U13515 ( n13933, n19236, n20044 );
nor U13516 ( n13979, n13982, n13975 );
nand U13517 ( n13975, n13951, n20032 );
nor U13518 ( n13951, n19239, n20031 );
xnor U13519 ( n13982, n20046, n13935 );
and U13520 ( n13935, n19235, n11418 );
nand U13521 ( n5787, n13983, n13984 );
nand U13522 ( n13984, n13985, n10371 );
nand U13523 ( n13983, n13986, n10669 );
nand U13524 ( n5782, n13987, n13988 );
nand U13525 ( n13988, n13985, n10669 );
or U13526 ( n13987, n13985, n20044 );
not U13527 ( n13985, n13986 );
nand U13528 ( n13986, g35, n13925 );
nor U13529 ( n5777, n13989, n10981 );
nor U13530 ( n13989, n13990, n13991 );
nor U13531 ( n13991, n13925, n10371 );
nor U13532 ( n13990, n20044, n13992 );
nor U13533 ( n13992, n20045, n13925 );
nand U13534 ( n13925, n13993, n20031 );
nor U13535 ( n13993, n19239, n10303 );
nand U13536 ( n5772, n13994, n13995 );
nand U13537 ( n13995, n13996, g35 );
nor U13538 ( n13996, n20043, n13997 );
nor U13539 ( n13997, n13998, n13999 );
nor U13540 ( n13998, n20037, n10519 );
nand U13541 ( n13994, n14000, n10519 );
nand U13542 ( n14000, g35, n14001 );
nand U13543 ( n14001, n14002, n20043 );
nand U13544 ( n5767, n14003, n14004 );
nand U13545 ( n14004, n11007, n10638 );
nand U13546 ( n14003, n14005, g35 );
nand U13547 ( n14005, n14006, n14007 );
nand U13548 ( n14007, n13999, n10519 );
nand U13549 ( n14006, n14002, n20042 );
nor U13550 ( n14002, n20037, n13999 );
nand U13551 ( n5762, n14008, n14009 );
nand U13552 ( n14009, n14010, g35 );
nor U13553 ( n14010, n19238, n14011 );
nor U13554 ( n14011, n14012, n14013 );
nor U13555 ( n14012, n14014, n10318 );
nand U13556 ( n14008, n14015, n10318 );
nand U13557 ( n14015, g35, n14016 );
nand U13558 ( n14016, n14017, n19238 );
nor U13559 ( n14017, n14014, n14013 );
nand U13560 ( n5757, n14018, n14019 );
nand U13561 ( n14019, n14020, n14021 );
nor U13562 ( n14020, n10318, n14013 );
nor U13563 ( n14018, n14022, n14023 );
nor U13564 ( n14023, n20040, g35 );
nor U13565 ( n14022, n10955, n14024 );
nand U13566 ( n14024, n14013, n10318 );
nand U13567 ( n14013, n14025, n14026 );
nand U13568 ( n14026, n20040, n14027 );
not U13569 ( n14025, n14028 );
nand U13570 ( n5752, n14029, n14030 );
nand U13571 ( n14030, n14031, n14021 );
nor U13572 ( n14031, n10394, n14028 );
nor U13573 ( n14029, n14032, n14033 );
nor U13574 ( n14033, n20039, g35 );
nor U13575 ( n14032, n10955, n14034 );
nand U13576 ( n14034, n14028, n10394 );
nand U13577 ( n14028, n14035, n14036 );
nand U13578 ( n14036, n20039, n14027 );
nand U13579 ( n5747, n14037, n14038 );
nand U13580 ( n14038, n14039, g35 );
nor U13581 ( n14039, n20039, n14035 );
and U13582 ( n14035, n14040, n14041 );
nand U13583 ( n14041, n20038, n14027 );
not U13584 ( n14027, n14014 );
nand U13585 ( n14037, n14042, n10258 );
nand U13586 ( n14042, g35, n14043 );
nand U13587 ( n14043, n14044, n20039 );
nor U13588 ( n14044, n14045, n14014 );
nand U13589 ( n5742, n14046, n14047 );
nand U13590 ( n14047, n14048, n14021 );
nor U13591 ( n14021, n14014, n10985 );
nand U13592 ( n14014, n14049, n20036 );
nor U13593 ( n14049, n14050, n14051 );
nor U13594 ( n14051, n14052, n14053 );
nor U13595 ( n14050, n14054, n14055 );
nor U13596 ( n14054, n20037, n10618 );
nor U13597 ( n14048, n14045, n10258 );
nor U13598 ( n14046, n14056, n14057 );
nor U13599 ( n14057, n20037, g35 );
nor U13600 ( n14056, n10955, n14058 );
nand U13601 ( n14058, n14045, n10258 );
nand U13602 ( n5737, n14059, n14060 );
nand U13603 ( n14060, n14061, n10607 );
nand U13604 ( n14061, g35, n13999 );
nand U13605 ( n14059, n14062, n14063 );
nor U13606 ( n14063, n20037, n14064 );
nor U13607 ( n14064, n14045, n14065 );
or U13608 ( n14065, n20041, n20039 );
nor U13609 ( n14062, n14066, n10981 );
nor U13610 ( n14066, n20043, n13999 );
nor U13611 ( n5732, n10955, n14067 );
nand U13612 ( n14067, n14068, n14069 );
nand U13613 ( n14069, n14070, n14040 );
nor U13614 ( n14070, n14071, n14072 );
nor U13615 ( n14072, n14073, n14053 );
nor U13616 ( n14073, n10607, n14074 );
nand U13617 ( n14074, n14075, n14052 );
nand U13618 ( n14075, n14076, n14077 );
nor U13619 ( n14077, n19238, n20038 );
and U13620 ( n14076, n10394, n20037 );
nor U13621 ( n14071, n10618, n14052 );
nand U13622 ( n14052, n14078, n10318 );
nor U13623 ( n14078, n20037, n20039 );
nand U13624 ( n14068, n14045, n20036 );
nand U13625 ( n5727, n14079, n14080 );
nand U13626 ( n14080, g35, n14081 );
nand U13627 ( n14081, g19357, n14082 );
nand U13628 ( n14082, n20035, n14083 );
nand U13629 ( n14083, n20034, g12923 );
nand U13630 ( n14079, n14084, n10642 );
nand U13631 ( n14084, n20024, g35 );
nand U13632 ( n5722, n14085, n14086 );
nand U13633 ( n14086, n14087, n20030 );
nor U13634 ( n14087, n14088, n14089 );
nor U13635 ( n14089, n14090, n14091 );
nor U13636 ( n14091, n20035, n10981 );
not U13637 ( n14090, n14092 );
nor U13638 ( n14088, n20035, n14092 );
nand U13639 ( n14092, n14093, n10417 );
nand U13640 ( n14085, n11007, n10417 );
nor U13641 ( n5717, n14094, n14095 );
nand U13642 ( n14095, n20030, g35 );
xnor U13643 ( n14094, n10417, n14093 );
and U13644 ( n14093, g12923, n14096 );
nand U13645 ( n14096, n14097, n19240 );
nor U13646 ( n14097, n10401, g7946 );
nand U13647 ( n5712, n14098, n14099 );
nand U13648 ( n14099, n14100, n14101 );
nor U13649 ( n14100, n14102, n14103 );
nor U13650 ( n14103, n14104, n14105 );
nor U13651 ( n14105, n19237, n10981 );
not U13652 ( n14104, n14106 );
nor U13653 ( n14102, n19237, n14106 );
nand U13654 ( n14098, n11007, n10419 );
nand U13655 ( n5707, n14107, n14108 );
nand U13656 ( n14108, n11007, n10676 );
nand U13657 ( n14107, n14109, g35 );
nor U13658 ( n14109, n14110, n14111 );
xnor U13659 ( n14111, n10419, n14112 );
nand U13660 ( n5702, n14113, n14114 );
nand U13661 ( n14114, n11008, n10361 );
nand U13662 ( n14113, g35, n14115 );
nand U13663 ( n14115, n14116, n14117 );
nand U13664 ( n14117, n14118, n10676 );
or U13665 ( n14118, n14106, n19237 );
nand U13666 ( n14106, n14112, n10419 );
and U13667 ( n14112, n14119, n14120 );
nor U13668 ( n14119, n20028, n14121 );
nor U13669 ( n14121, n10361, n14122 );
nand U13670 ( n5697, n14123, n14124 );
nand U13671 ( n14124, n11008, n10492 );
nand U13672 ( n14123, n14125, g35 );
nand U13673 ( n14125, n14126, n14127 );
nand U13674 ( n14127, n20028, n10361 );
nand U13675 ( n14126, g7946, n10363 );
nand U13676 ( n5692, n14128, n14129 );
nand U13677 ( n14129, n11008, n10363 );
nand U13678 ( n14128, n14130, g35 );
nand U13679 ( n14130, n14131, n14132 );
or U13680 ( n14132, n14133, n20027 );
nand U13681 ( n14131, n14133, n10492 );
nand U13682 ( n14133, n14134, n10303 );
nor U13683 ( n14134, n20028, n20031 );
nand U13684 ( n5687, n14135, n14136 );
nand U13685 ( n14136, n11008, n10303 );
nand U13686 ( n14135, n14137, g35 );
nand U13687 ( n14137, n14138, n14139 );
nand U13688 ( n14139, n20028, n10363 );
nand U13689 ( n14138, g7946, n10240 );
nand U13690 ( n5682, n14140, n14141 );
nand U13691 ( n14141, g35, n14142 );
nand U13692 ( n14142, n12408, n14101 );
not U13693 ( n14101, n14110 );
not U13694 ( n12408, n14120 );
nand U13695 ( n14140, n14143, n10582 );
nand U13696 ( n14143, n14144, g35 );
xnor U13697 ( n14144, n20032, n20028 );
nor U13698 ( n5677, n14145, n10982 );
nor U13699 ( n14145, n14110, n14146 );
xnor U13700 ( n14146, g7946, n20031 );
nor U13701 ( n14110, n14116, n14147 );
nor U13702 ( n14147, n20033, n14120 );
nor U13703 ( n14120, n10582, n20032 );
nand U13704 ( n14116, n14148, n14149 );
nor U13705 ( n14149, n20028, n14122 );
nand U13706 ( n14122, n10240, n10363 );
nor U13707 ( n14148, n14150, n10361 );
nor U13708 ( n14150, n14151, n14152 );
nor U13709 ( n14151, n14153, n14154 );
nand U13710 ( n14154, n14055, n10394 );
not U13711 ( n14055, n14053 );
nand U13712 ( n14153, n10258, n10638 );
xnor U13713 ( n5664, n14155, n10401 );
or U13714 ( n14155, n14156, n11024 );
nand U13715 ( n5651, n14157, n14158 );
nand U13716 ( n14158, n11008, n10240 );
nand U13717 ( n14157, n14159, g35 );
xor U13718 ( n14159, n14156, n14160 );
nand U13719 ( n14160, n14161, n14162 );
nor U13720 ( n14162, g19357, n14163 );
nand U13721 ( n14163, n20028, n20029 );
nor U13722 ( n14161, g13272, g8475 );
nand U13723 ( n14156, n14164, n14165 );
nor U13724 ( n14164, n14166, n13999 );
xnor U13725 ( n14166, n19241, n20030 );
nand U13726 ( n5646, n14167, n14168 );
or U13727 ( n14168, g35, n19241 );
nand U13728 ( n5637, n14169, n14170 );
nand U13729 ( n14170, n14171, g17423 );
nor U13730 ( n14169, n14172, n14173 );
nor U13731 ( n14173, n20026, g35 );
nor U13732 ( n14172, n10955, n14174 );
nand U13733 ( n14174, n19248, g10527 );
nand U13734 ( n5632, n14167, n14175 );
nand U13735 ( n14175, n11008, n10473 );
nand U13736 ( n5623, n14176, n14177 );
nand U13737 ( n14177, g35, g496 );
nand U13738 ( n14176, n11008, n10449 );
nand U13739 ( n5618, n14178, n14179 );
nand U13740 ( n14179, n14180, g35 );
nor U13741 ( n14180, n19243, n14181 );
nand U13742 ( n14178, n14182, n10480 );
nand U13743 ( n14182, g35, n14183 );
nand U13744 ( n14183, n14181, n19243 );
nand U13745 ( n5613, n14184, n14185 );
nand U13746 ( n14185, n11008, n10620 );
nand U13747 ( n14184, n14186, g35 );
nand U13748 ( n14186, n14187, n14188 );
nand U13749 ( n14188, n14189, n10480 );
nand U13750 ( n14187, n14190, n19242 );
nor U13751 ( n14190, n10449, n14189 );
nand U13752 ( n5608, n14191, n14192 );
nand U13753 ( n14192, n14193, n19244 );
nor U13754 ( n14191, n14194, n14195 );
nor U13755 ( n14195, n19245, g35 );
nor U13756 ( n14194, n10955, n14196 );
nand U13757 ( n14196, n14197, n10620 );
xnor U13758 ( n5603, n14198, n10590 );
nand U13759 ( n14198, g35, n10660 );
nor U13760 ( n5586, n14199, n14200 );
nand U13761 ( n14200, n19247, n20023 );
nand U13762 ( n14199, n14201, n19248 );
nor U13763 ( n14201, n14202, n10980 );
nor U13764 ( n14202, n14189, n14203 );
nand U13765 ( n14203, n14204, n10449 );
or U13766 ( n14204, n14152, n13999 );
nand U13767 ( n13999, n14053, n14040 );
not U13768 ( n14040, n14045 );
nor U13769 ( n14045, n10401, n10286 );
xnor U13770 ( n14053, n20030, n10240 );
not U13771 ( n14189, n14181 );
nor U13772 ( n14181, n14197, n19244 );
not U13773 ( n14197, n14193 );
nor U13774 ( n14193, n19245, n19246 );
nor U13775 ( n5581, n20022, n14205 );
nor U13776 ( n14205, n14206, n10981 );
nor U13777 ( n14206, n11418, n14207 );
nand U13778 ( n5576, n14208, n14209 );
nand U13779 ( n14209, n11009, n10521 );
nor U13780 ( n14208, n14210, n14211 );
nor U13781 ( n14211, n14207, n10911 );
nor U13782 ( n14210, n20022, n14212 );
nand U13783 ( n14212, n14171, n14207 );
nand U13784 ( n14207, n14213, n10521 );
nand U13785 ( n5571, n14214, n14215 );
nand U13786 ( n14215, n11009, n10679 );
nor U13787 ( n14214, n14216, n14217 );
nor U13788 ( n14217, n14218, n10521 );
nor U13789 ( n14216, n20021, n14219 );
nand U13790 ( n14219, n14171, n14218 );
not U13791 ( n14218, n14213 );
nor U13792 ( n14213, n14220, n20020 );
nand U13793 ( n5566, n14221, n14222 );
nand U13794 ( n14222, n11009, n10744 );
nor U13795 ( n14221, n14223, n14224 );
nor U13796 ( n14224, n14220, n10679 );
nor U13797 ( n14223, n20020, n14225 );
nand U13798 ( n14225, n14171, n14220 );
or U13799 ( n14220, n14226, n20019 );
nand U13800 ( n5561, n14227, n14228 );
nand U13801 ( n14228, n11009, n10745 );
nor U13802 ( n14227, n14229, n14230 );
nor U13803 ( n14230, n14226, n10744 );
nor U13804 ( n14229, n20019, n14231 );
nand U13805 ( n14231, n14171, n14226 );
or U13806 ( n14226, n14232, n20018 );
nand U13807 ( n5556, n14233, n14234 );
nand U13808 ( n14234, n11009, n10746 );
nor U13809 ( n14233, n14235, n14236 );
nor U13810 ( n14236, n14232, n10745 );
nor U13811 ( n14235, n20018, n14237 );
nand U13812 ( n14237, n14171, n14232 );
or U13813 ( n14232, n14238, n20017 );
nand U13814 ( n5551, n14239, n14240 );
nand U13815 ( n14240, n11009, n10655 );
nor U13816 ( n14239, n14241, n14242 );
nor U13817 ( n14242, n14238, n10746 );
nor U13818 ( n14241, n20017, n14243 );
nand U13819 ( n14243, n14171, n14238 );
nand U13820 ( n14238, n14244, n14245 );
nor U13821 ( n14244, n19250, n20016 );
nand U13822 ( n5546, n14246, n14247 );
nand U13823 ( n14247, n11009, n10670 );
nor U13824 ( n14246, n14248, n14249 );
nor U13825 ( n14249, n10655, n14250 );
nand U13826 ( n14250, n14245, n10483 );
nor U13827 ( n14248, n20016, n14251 );
nor U13828 ( n14251, n14252, n5536 );
nor U13829 ( n14252, n14245, n14167 );
nor U13830 ( n14245, n19249, n20024 );
nand U13831 ( n5541, n14253, n14254 );
nand U13832 ( n14254, n14255, n10483 );
nand U13833 ( n14255, g35, n14256 );
nand U13834 ( n14256, n19249, g12923 );
nand U13835 ( n14253, n5536, n10670 );
nor U13836 ( n5536, n10483, n14167 );
not U13837 ( n14167, n14171 );
nor U13838 ( n14171, n10955, n20024 );
nand U13839 ( n5527, n14257, n14258 );
nand U13840 ( n14258, n19253, g35 );
nand U13841 ( n14257, n11009, n10252 );
nand U13842 ( n5522, n14259, n14260 );
or U13843 ( n14260, g35, n19252 );
nand U13844 ( n14259, n14261, g35 );
nand U13845 ( n14261, n14262, n14263 );
nand U13846 ( n14263, n14264, n10252 );
nand U13847 ( n14262, n14265, n14266 );
nand U13848 ( n5513, n14267, n14268 );
or U13849 ( n14268, g35, n19261 );
nand U13850 ( n14267, n14269, g35 );
xnor U13851 ( n14269, n19251, n14270 );
nor U13852 ( n14270, n14264, n14265 );
xor U13853 ( n14265, n19252, n19251 );
not U13854 ( n14264, n14266 );
nor U13855 ( n14266, n19253, n10941 );
nand U13856 ( n5508, n14271, n14272 );
or U13857 ( n14272, g35, n19262 );
nand U13858 ( n14271, n14273, g35 );
nor U13859 ( n14273, n19257, n14274 );
nor U13860 ( n5503, n20015, n14275 );
nor U13861 ( n14275, n14276, n10980 );
nand U13862 ( n5498, n14277, n14278 );
nand U13863 ( n14278, n11009, n10680 );
nor U13864 ( n14277, n14279, n14280 );
and U13865 ( n14280, n20015, n14276 );
nor U13866 ( n14279, n20015, n14281 );
nand U13867 ( n14281, n14282, n14283 );
not U13868 ( n14283, n14276 );
nor U13869 ( n14276, n14284, n19254 );
nand U13870 ( n5493, n14285, n14286 );
nand U13871 ( n14286, n11009, n10747 );
nor U13872 ( n14285, n14287, n14288 );
nor U13873 ( n14288, n14284, n10680 );
nor U13874 ( n14287, n19254, n14289 );
nand U13875 ( n14289, n14282, n14284 );
or U13876 ( n14284, n14290, n20014 );
nand U13877 ( n5488, n14291, n14292 );
nand U13878 ( n14292, n11009, n10748 );
nor U13879 ( n14291, n14293, n14294 );
nor U13880 ( n14294, n14290, n10747 );
nor U13881 ( n14293, n20014, n14295 );
nand U13882 ( n14295, n14282, n14290 );
or U13883 ( n14290, n14296, n19255 );
nand U13884 ( n5483, n14297, n14298 );
nand U13885 ( n14298, n11009, n10749 );
nor U13886 ( n14297, n14299, n14300 );
nor U13887 ( n14300, n14296, n10748 );
nor U13888 ( n14299, n19255, n14301 );
nand U13889 ( n14301, n14282, n14296 );
or U13890 ( n14296, n14302, n20013 );
nand U13891 ( n5478, n14303, n14304 );
or U13892 ( n14304, g35, n19256 );
nor U13893 ( n14303, n14305, n14306 );
nor U13894 ( n14306, n14302, n10749 );
nor U13895 ( n14305, n20013, n14307 );
nand U13896 ( n14307, n14282, n14302 );
nand U13897 ( n14302, n14308, n14309 );
nor U13898 ( n14308, n19256, n14310 );
nand U13899 ( n5473, n14311, n14312 );
nand U13900 ( n14312, n14313, n14282 );
and U13901 ( n14282, n14309, g35 );
and U13902 ( n14309, n14314, n14315 );
nand U13903 ( n14315, n14316, n14317 );
or U13904 ( n14317, n10578, n14318 );
xnor U13905 ( n14313, n14316, n19256 );
not U13906 ( n14316, n14310 );
nand U13907 ( n14311, n11010, n10699 );
nand U13908 ( n5468, n14319, n14320 );
nand U13909 ( n14320, n11010, n10522 );
nor U13910 ( n14319, n14321, n14322 );
nor U13911 ( n14322, n14274, n10699 );
nor U13912 ( n14321, n19257, n14323 );
nand U13913 ( n14323, n14324, n14274 );
nand U13914 ( n14274, n14325, n10522 );
nand U13915 ( n5463, n14326, n14327 );
nand U13916 ( n14327, n11010, n10681 );
nor U13917 ( n14326, n14328, n14329 );
nor U13918 ( n14329, n14330, n10522 );
nor U13919 ( n14328, n19258, n14331 );
nand U13920 ( n14331, n14324, n14330 );
not U13921 ( n14330, n14325 );
nor U13922 ( n14325, n14332, n19259 );
nand U13923 ( n5458, n14333, n14334 );
nand U13924 ( n14334, n11010, n10750 );
nor U13925 ( n14333, n14335, n14336 );
nor U13926 ( n14336, n14332, n10681 );
nor U13927 ( n14335, n19259, n14337 );
nand U13928 ( n14337, n14324, n14332 );
or U13929 ( n14332, n14338, n20012 );
nand U13930 ( n5453, n14339, n14340 );
or U13931 ( n14340, g35, n19260 );
nor U13932 ( n14339, n14341, n14342 );
nor U13933 ( n14342, n14338, n10750 );
nor U13934 ( n14341, n20012, n14343 );
nand U13935 ( n14343, n14324, n14338 );
nand U13936 ( n14338, n14344, n14345 );
nor U13937 ( n14344, n19260, n20011 );
nand U13938 ( n5448, n14346, n14347 );
nand U13939 ( n14347, n14348, n10902 );
nand U13940 ( n14348, g35, n14349 );
nand U13941 ( n14349, n19260, n14345 );
nand U13942 ( n14346, n14350, n20011 );
nor U13943 ( n14350, n19260, n14351 );
nand U13944 ( n5443, n14352, n14353 );
nand U13945 ( n14353, n20011, n14324 );
not U13946 ( n14324, n14351 );
nand U13947 ( n14351, n14345, g35 );
and U13948 ( n14345, n14354, n14314 );
nor U13949 ( n14314, n19991, n14355 );
nor U13950 ( n14354, n14356, n14357 );
and U13951 ( n14357, n10900, n14358 );
not U13952 ( n14356, n14359 );
nand U13953 ( n14352, n11010, n10900 );
nor U13954 ( n5438, n10955, n14360 );
nand U13955 ( n14360, n14359, n14358 );
nand U13956 ( n14358, n14361, n14362 );
nor U13957 ( n14362, n14363, n14364 );
nand U13958 ( n14364, n10349, n10241 );
nand U13959 ( n14363, n10335, n10230 );
nor U13960 ( n14361, n10253, n14365 );
nand U13961 ( n14365, n19971, n19973 );
nand U13962 ( n14359, n20010, n14366 );
nand U13963 ( n14366, n14367, n14368 );
nor U13964 ( n14368, n14369, n14370 );
nand U13965 ( n14370, n19974, n10431 );
nand U13966 ( n14369, n10458, n10253 );
nor U13967 ( n14367, n10230, n14371 );
nand U13968 ( n14371, n19970, n19972 );
nand U13969 ( n5433, n14372, n14373 );
nand U13970 ( n14373, n11010, g21292 );
nand U13971 ( n14372, g35, n14374 );
nand U13972 ( n14374, n19261, n19319 );
nand U13973 ( n5428, n14375, n14376 );
nand U13974 ( n14376, g35, g21292 );
nand U13975 ( n14375, n11010, n10813 );
nand U13976 ( n5423, n14377, n14378 );
or U13977 ( n14378, g35, n19461 );
nand U13978 ( n14377, g35, n14379 );
nand U13979 ( n14379, n19336, g20899 );
nand U13980 ( n5418, n14380, n14381 );
or U13981 ( n14381, g35, n19466 );
nand U13982 ( n14380, g35, n14382 );
nand U13983 ( n14382, n19461, n19262 );
nand U13984 ( n5413, n14383, n14384 );
nand U13985 ( n14384, n14385, n14386 );
nand U13986 ( n14386, n19466, n10307 );
or U13987 ( n14383, g35, n19475 );
nand U13988 ( n5408, n14387, n14388 );
nand U13989 ( n14388, n11010, n10831 );
nand U13990 ( n14387, g35, n14389 );
nand U13991 ( n14389, n19475, n10307 );
nor U13992 ( n5403, n14390, n10980 );
nor U13993 ( n14390, n10252, n10831 );
nand U13994 ( n5398, n14391, n14392 );
nand U13995 ( n14392, n14393, n10608 );
nand U13996 ( n14393, g35, n14394 );
nand U13997 ( n14391, n14385, n10794 );
nand U13998 ( n5393, n14395, n14396 );
nand U13999 ( n14396, n11010, n10495 );
nor U14000 ( n14395, n14397, n14398 );
nor U14001 ( n14398, n10608, n14394 );
nor U14002 ( n14397, n20008, n14399 );
nand U14003 ( n14399, n14385, n14394 );
nand U14004 ( n14394, n14400, n10495 );
nand U14005 ( n5388, n14401, n14402 );
nand U14006 ( n14402, n11010, n10494 );
nor U14007 ( n14401, n14403, n14404 );
nor U14008 ( n14404, n14405, n10495 );
nor U14009 ( n14403, n19462, n14406 );
nand U14010 ( n14406, n14385, n14405 );
not U14011 ( n14405, n14400 );
nor U14012 ( n14400, n14407, n19337 );
nand U14013 ( n5383, n14408, n14409 );
nand U14014 ( n14409, n11011, n10643 );
nor U14015 ( n14408, n14410, n14411 );
nor U14016 ( n14411, n14407, n10494 );
nor U14017 ( n14410, n19337, n14412 );
nand U14018 ( n14412, n14385, n14407 );
or U14019 ( n14407, n14413, n19326 );
nand U14020 ( n5378, n14414, n14415 );
nand U14021 ( n14415, n11011, n10497 );
nor U14022 ( n14414, n14416, n14417 );
nor U14023 ( n14417, n14413, n10643 );
nor U14024 ( n14416, n19326, n14418 );
nand U14025 ( n14418, n14385, n14413 );
or U14026 ( n14413, n14419, n19320 );
nand U14027 ( n5373, n14420, n14421 );
nand U14028 ( n14421, n11011, n10496 );
nor U14029 ( n14420, n14422, n14423 );
nor U14030 ( n14423, n14419, n10497 );
nor U14031 ( n14422, n19320, n14424 );
nand U14032 ( n14424, n14385, n14419 );
or U14033 ( n14419, n14425, n19488 );
nand U14034 ( n5368, n14426, n14427 );
nand U14035 ( n14427, n11011, n10498 );
nor U14036 ( n14426, n14428, n14429 );
nor U14037 ( n14429, n14425, n10496 );
nor U14038 ( n14428, n19488, n14430 );
nand U14039 ( n14430, n14385, n14425 );
or U14040 ( n14425, n14431, n19482 );
nand U14041 ( n5363, n14432, n14433 );
nand U14042 ( n14433, n11015, n10499 );
nor U14043 ( n14432, n14434, n14435 );
nor U14044 ( n14435, n14431, n10498 );
nor U14045 ( n14434, n19482, n14436 );
nand U14046 ( n14436, n14385, n14431 );
or U14047 ( n14431, n14437, n19476 );
nand U14048 ( n5358, n14438, n14439 );
nand U14049 ( n14439, n11011, n10644 );
nor U14050 ( n14438, n14440, n14441 );
nor U14051 ( n14441, n14437, n10499 );
nor U14052 ( n14440, n19476, n14442 );
nand U14053 ( n14442, n14385, n14437 );
or U14054 ( n14437, n14443, n19467 );
nand U14055 ( n5353, n14444, n14445 );
nand U14056 ( n14445, n11011, n10645 );
nor U14057 ( n14444, n14446, n14447 );
nor U14058 ( n14447, n14443, n10644 );
nor U14059 ( n14446, n19467, n14448 );
nand U14060 ( n14448, n14385, n14443 );
or U14061 ( n14443, n14449, n20007 );
nand U14062 ( n5348, n14450, n14451 );
nand U14063 ( n14451, n11011, n10500 );
nor U14064 ( n14450, n14452, n14453 );
nor U14065 ( n14453, n14449, n10645 );
nor U14066 ( n14452, n20007, n14454 );
nand U14067 ( n14454, n14385, n14449 );
or U14068 ( n14449, n14455, n19335 );
nand U14069 ( n5343, n14456, n14457 );
nand U14070 ( n14457, n11011, n10501 );
nor U14071 ( n14456, n14458, n14459 );
nor U14072 ( n14459, n14455, n10500 );
nor U14073 ( n14458, n19335, n14460 );
nand U14074 ( n14460, n14385, n14455 );
or U14075 ( n14455, n14461, n20006 );
nand U14076 ( n5338, n14462, n14463 );
or U14077 ( n14463, g35, n20005 );
nor U14078 ( n14462, n14464, n14465 );
nor U14079 ( n14465, n14461, n10501 );
nor U14080 ( n14464, n20006, n14466 );
nand U14081 ( n14466, n14385, n14461 );
nand U14082 ( n14461, n14467, n14468 );
nor U14083 ( n14467, n20005, n14469 );
nor U14084 ( n14469, n20004, n10581 );
nand U14085 ( n5333, n14470, n14471 );
nand U14086 ( n14471, n14472, n14385 );
and U14087 ( n14385, g35, n14473 );
or U14088 ( n14473, n10581, n20004 );
xnor U14089 ( n14472, n20005, n14468 );
and U14090 ( n14468, n14355, n14474 );
nand U14091 ( n14474, n20004, g12184 );
and U14092 ( n14355, n14475, n14476 );
nor U14093 ( n14476, n14477, n14478 );
nor U14094 ( n14478, n10333, n14479 );
nand U14095 ( n14479, n19274, n20003 );
nor U14096 ( n14477, n19273, n14480 );
nand U14097 ( n14480, n10814, n10277 );
nor U14098 ( n14475, n14481, n14482 );
nor U14099 ( n14481, n20009, n20008 );
nand U14100 ( n14470, n11011, n10581 );
nand U14101 ( n5320, n14483, n14484 );
nand U14102 ( n14484, n11011, n10814 );
nand U14103 ( n5315, n14485, n14486 );
or U14104 ( n14486, n14487, n20003 );
nand U14105 ( n14485, n14487, n10898 );
nand U14106 ( n14487, g35, n14482 );
nor U14107 ( n5310, n10955, n14488 );
xor U14108 ( n14488, n14489, n14490 );
xor U14109 ( n14490, n14491, n14492 );
xnor U14110 ( n14492, n19974, n14493 );
nand U14111 ( n14493, n10898, n14482 );
nand U14112 ( n14482, n14494, n14495 );
nor U14113 ( n14495, n10345, n14496 );
nand U14114 ( n14496, n19999, n19270 );
and U14115 ( n14494, n14497, n14498 );
xnor U14116 ( n14491, n10241, n19973 );
xor U14117 ( n14489, n14499, n14500 );
xnor U14118 ( n14500, n10335, n19971 );
xnor U14119 ( n14499, n10230, n19969 );
nand U14120 ( n5305, n14501, n14502 );
nand U14121 ( n14502, n11011, g20901 );
nand U14122 ( n14501, g35, n14503 );
nand U14123 ( n14503, n14504, n14505 );
nand U14124 ( n14505, n11266, n10431 );
nor U14125 ( n14504, n14506, n14507 );
and U14126 ( n14507, n14508, n19563 );
nor U14127 ( n14506, g72, n14509 );
nand U14128 ( n14509, n14508, n10253 );
nand U14129 ( n14508, n19563, n14510 );
nand U14130 ( n14510, n10458, g72 );
nand U14131 ( n5300, n14511, n14512 );
or U14132 ( n14512, g35, n19263 );
nand U14133 ( n14511, n14513, g35 );
nand U14134 ( n14513, n14514, n14515 );
nand U14135 ( n14515, n14516, g73 );
nand U14136 ( n14516, n14517, n14518 );
nand U14137 ( n14518, n10230, g72 );
nand U14138 ( n14517, n19562, n10335 );
nand U14139 ( n14514, n14519, n19563 );
nand U14140 ( n14519, n14520, n14521 );
nand U14141 ( n14521, n10241, g72 );
nand U14142 ( n14520, n19562, n10349 );
nor U14143 ( n5295, n14310, n14522 );
nand U14144 ( n14522, g35, n14523 );
nand U14145 ( n14523, n14524, n14525 );
nand U14146 ( n14525, n14318, n10578 );
nand U14147 ( n14310, n14526, n19268 );
nor U14148 ( n14526, n19264, n19997 );
nand U14149 ( n5270, n14527, n14528 );
or U14150 ( n14528, n14529, n19283 );
nand U14151 ( n14527, n14529, n10870 );
nand U14152 ( n5265, n14530, n14531 );
nand U14153 ( n14531, n14532, n10870 );
nor U14154 ( n14530, n14533, n14534 );
nor U14155 ( n14534, n10955, n14535 );
nand U14156 ( n14535, n14498, n10349 );
nor U14157 ( n14533, n19265, g35 );
nand U14158 ( n5260, n14536, n14537 );
nand U14159 ( n14537, n14532, n10578 );
nand U14160 ( n14536, n14529, n10561 );
nand U14161 ( n5255, n14538, n14539 );
nand U14162 ( n14539, n14532, n10561 );
nand U14163 ( n14538, n14529, n10278 );
not U14164 ( n14529, n14532 );
nand U14165 ( n5250, n14540, n14541 );
nand U14166 ( n14541, n14532, n10278 );
nor U14167 ( n14532, n10954, n14498 );
nor U14168 ( n14540, n14542, n14543 );
nor U14169 ( n14543, n10954, n14544 );
nand U14170 ( n14544, n14498, n10365 );
nor U14171 ( n14542, n19284, g35 );
nand U14172 ( n5245, n14545, n14546 );
nand U14173 ( n14546, n14547, n10415 );
nand U14174 ( n14545, n14548, n10271 );
nand U14175 ( n5240, n14549, n14550 );
nand U14176 ( n14550, n11012, n10544 );
nor U14177 ( n14549, n14551, n14552 );
nor U14178 ( n14552, n20002, n14548 );
nor U14179 ( n14551, n10300, n14553 );
nand U14180 ( n14553, n14554, n10773 );
nand U14181 ( n5235, n14555, n14556 );
nand U14182 ( n14556, n14547, n10544 );
nand U14183 ( n14555, n14548, n10871 );
nand U14184 ( n5230, n14557, n14558 );
nand U14185 ( n14558, n14547, n10871 );
or U14186 ( n14557, n14547, n19266 );
nand U14187 ( n5225, n14559, n14560 );
nand U14188 ( n14560, n11012, n10543 );
nor U14189 ( n14559, n14561, n14562 );
nor U14190 ( n14562, n19266, n14548 );
nor U14191 ( n14561, n19973, n14563 );
nand U14192 ( n5220, n14564, n14565 );
nand U14193 ( n14565, n14547, n10543 );
nand U14194 ( n14564, n14548, n10548 );
nand U14195 ( n5215, n14566, n14567 );
nand U14196 ( n14567, n14547, n10548 );
or U14197 ( n14566, n14547, n19267 );
nand U14198 ( n5210, n14568, n14569 );
nand U14199 ( n14569, n11012, n10506 );
nor U14200 ( n14568, n14570, n14571 );
nor U14201 ( n14571, n19267, n14548 );
nor U14202 ( n14570, n19974, n14563 );
nand U14203 ( n5205, n14572, n14573 );
nand U14204 ( n14573, n14547, n10506 );
nand U14205 ( n14572, n14548, n10352 );
nand U14206 ( n5200, n14574, n14575 );
nand U14207 ( n14575, n14547, n10352 );
nor U14208 ( n14574, n14576, n14577 );
nor U14209 ( n14577, n10229, n14578 );
nand U14210 ( n14578, n14554, n14579 );
nor U14211 ( n14576, n20000, n14580 );
nor U14212 ( n14580, n14581, n10980 );
nor U14213 ( n14581, n14579, n14582 );
nand U14214 ( n5195, n14583, n14584 );
nand U14215 ( n14584, n14554, n10365 );
nand U14216 ( n14583, n14547, n10229 );
nand U14217 ( n5190, n14585, n14586 );
nand U14218 ( n14586, n14587, n19270 );
nor U14219 ( n14585, n14588, n14589 );
nor U14220 ( n14589, n14590, n10980 );
nor U14221 ( n14590, n14591, n14592 );
nor U14222 ( n14591, n19270, n14587 );
nor U14223 ( n14587, n14593, n19999 );
nor U14224 ( n14588, n19999, g35 );
nand U14225 ( n5185, n14594, n14595 );
nand U14226 ( n14595, n11012, n10345 );
nand U14227 ( n14594, g35, n14596 );
nand U14228 ( n14596, n14597, n14598 );
xnor U14229 ( n14597, n19999, n14593 );
nand U14230 ( n14593, n14599, n14600 );
nand U14231 ( n14600, n19998, n14601 );
nand U14232 ( n5180, n14602, n14603 );
nand U14233 ( n14603, n11012, n10224 );
nand U14234 ( n14602, n14604, g35 );
nor U14235 ( n14604, n14592, n14605 );
nand U14236 ( n14605, n14606, n14607 );
nand U14237 ( n14607, n14599, n10345 );
nand U14238 ( n14606, n19998, n14608 );
nand U14239 ( n14608, n14599, n14601 );
and U14240 ( n14599, n14609, n14610 );
nor U14241 ( n14609, n19997, n10384 );
not U14242 ( n14592, n14598 );
nand U14243 ( n5175, n14611, n14612 );
nand U14244 ( n14612, n14613, n10384 );
nand U14245 ( n14611, n14614, n10224 );
nand U14246 ( n5170, n14615, n14616 );
nand U14247 ( n14616, n14613, n10404 );
nand U14248 ( n14613, g35, n14617 );
nand U14249 ( n14617, n14610, n14598 );
nand U14250 ( n14615, n14614, n10384 );
nand U14251 ( n5165, n14618, n14619 );
not U14252 ( n14619, n14620 );
nor U14253 ( n14618, n14621, n14622 );
nor U14254 ( n14622, n19995, n14614 );
nor U14255 ( n14621, n19996, n14623 );
nand U14256 ( n5160, n14624, n14625 );
nand U14257 ( n14625, n14626, n19997 );
nor U14258 ( n14624, n14620, n14627 );
nor U14259 ( n14627, n19995, n14628 );
nor U14260 ( n14628, n14629, n14614 );
nor U14261 ( n14629, n10954, n10384 );
nor U14262 ( n14620, n14630, n14598 );
nand U14263 ( n14598, n19992, n10538 );
nand U14264 ( n5155, n14631, n14632 );
nand U14265 ( n14632, n11012, n10656 );
nor U14266 ( n14631, n14633, n14634 );
nor U14267 ( n14634, n10663, n14635 );
nand U14268 ( n14635, n14636, n14637 );
nor U14269 ( n14633, n19994, n14638 );
nand U14270 ( n14638, n14639, n14640 );
not U14271 ( n14640, n14637 );
nor U14272 ( n14637, n14641, n19993 );
nand U14273 ( n5150, n14642, n14643 );
or U14274 ( n14643, g35, n19269 );
nor U14275 ( n14642, n14644, n14645 );
nor U14276 ( n14645, n10656, n14646 );
nand U14277 ( n14646, n14636, n14647 );
nor U14278 ( n14644, n19993, n14648 );
nand U14279 ( n14648, n14639, n14641 );
not U14280 ( n14641, n14647 );
nor U14281 ( n14647, n14649, n19269 );
nand U14282 ( n5145, n14650, n14651 );
nand U14283 ( n14651, n14652, n14639 );
and U14284 ( n14639, n14636, g35 );
and U14285 ( n14636, n14653, n10300 );
or U14286 ( n14653, n14649, n14654 );
xnor U14287 ( n14652, n14655, n19269 );
nand U14288 ( n14650, n11013, n10538 );
nand U14289 ( n5140, n14656, n14657 );
nand U14290 ( n14657, n14614, n10538 );
or U14291 ( n14656, n14614, n19992 );
nand U14292 ( n5135, n14658, n14659 );
nand U14293 ( n14659, n11013, n10307 );
nor U14294 ( n14658, n14660, n14661 );
nor U14295 ( n14661, n19992, n14623 );
not U14296 ( n14623, n14614 );
and U14297 ( n14660, n14662, n14626 );
nand U14298 ( n5130, n14663, n14664 );
nand U14299 ( n14664, n11013, g20899 );
nor U14300 ( n14663, n14665, n14666 );
nor U14301 ( n14666, n14630, n14662 );
nand U14302 ( n14662, n14667, n19991 );
nor U14303 ( n14667, n19982, n14654 );
nand U14304 ( n14654, n14668, n14669 );
nor U14305 ( n14669, n10722, n14670 );
nand U14306 ( n14670, n10836, n10260 );
nor U14307 ( n14668, n14671, n14672 );
nand U14308 ( n14672, n14673, n19988 );
xnor U14309 ( n14673, n19271, n19272 );
xnor U14310 ( n14671, n10333, n19274 );
not U14311 ( n14630, n14626 );
nor U14312 ( n14626, n14674, n10980 );
nor U14313 ( n14665, n19991, n14675 );
nor U14314 ( n14675, n14676, n14614 );
nor U14315 ( n14614, n10954, n14610 );
not U14316 ( n14610, n14674 );
nand U14317 ( n14674, n14677, n19978 );
nor U14318 ( n14677, n19278, n19979 );
nor U14319 ( n14676, n10663, n14678 );
nand U14320 ( n14678, g35, n10300 );
nand U14321 ( n5125, n14679, n14680 );
nand U14322 ( n14680, n14681, n14655 );
nor U14323 ( n14681, n19272, n10980 );
nor U14324 ( n14679, n14682, n14683 );
nor U14325 ( n14683, n19271, n14684 );
and U14326 ( n14682, g20899, n14684 );
nor U14327 ( n14684, n10954, n14655 );
not U14328 ( n14655, n14649 );
nand U14329 ( n14649, n14685, n14686 );
nor U14330 ( n14686, n10345, n14687 );
nand U14331 ( n14687, n19996, n10661 );
nor U14332 ( n14685, n14582, n14601 );
or U14333 ( n14601, n19270, n19999 );
nand U14334 ( n5120, n14688, n14689 );
or U14335 ( n14689, n14690, n19271 );
nand U14336 ( n14688, n14690, n10662 );
nand U14337 ( n5115, n14691, n14692 );
nand U14338 ( n14692, n14693, n10662 );
nand U14339 ( n14691, n14690, n10333 );
nand U14340 ( n5110, n14694, n14695 );
nand U14341 ( n14695, n14693, n10333 );
nand U14342 ( n14694, n14690, n10277 );
nand U14343 ( n5105, n14696, n14697 );
nand U14344 ( n14697, n14693, n10277 );
nand U14345 ( n14696, n14690, n10722 );
nand U14346 ( n5100, n14698, n14699 );
nand U14347 ( n14699, n11013, n10836 );
nor U14348 ( n14698, n14700, n14701 );
nor U14349 ( n14701, n19990, n14690 );
and U14350 ( n14700, n10260, n14702 );
not U14351 ( n51, n11052 );
xnor U14352 ( n11052, n14703, n14704 );
xor U14353 ( n14704, n14705, n14706 );
xor U14354 ( n14706, n14707, n14708 );
xor U14355 ( n14708, new_g34971_, new_g34970_ );
nand U14356 ( new_g34970_, n14709, n14710 );
nor U14357 ( n14710, n14711, n14712 );
nand U14358 ( n14712, n14713, n14714 );
nand U14359 ( n14714, n137, n14715 );
nand U14360 ( n14715, n14716, n14717 );
nor U14361 ( n14717, n14718, n14719 );
nand U14362 ( n14719, n14720, n14721 );
nand U14363 ( n14721, n14722, n10657 );
nand U14364 ( n14720, n14723, n10496 );
nand U14365 ( n14718, n14724, n14725 );
nand U14366 ( n14725, n14726, n10503 );
nor U14367 ( n14724, n14727, n14728 );
nor U14368 ( n14727, n19489, n14729 );
nor U14369 ( n14716, n14730, n14731 );
nand U14370 ( n14731, n14732, n14733 );
nand U14371 ( n14733, n14734, n10782 );
nand U14372 ( n14732, n14735, n10539 );
nand U14373 ( n14730, n14736, n14737 );
nand U14374 ( n14737, n14738, n10700 );
nand U14375 ( n14736, n14739, n10508 );
nand U14376 ( n14713, n14740, n10511 );
nand U14377 ( n14711, n14741, n14742 );
nand U14378 ( n14742, n14743, n10621 );
nand U14379 ( n14741, n14744, n10622 );
nor U14380 ( n14709, n14745, n14746 );
nand U14381 ( n14746, n14747, n14748 );
nand U14382 ( n14748, n14749, n10930 );
nand U14383 ( n14747, n14750, g45 );
nand U14384 ( n14745, n14751, n14752 );
nand U14385 ( n14752, n14753, n10513 );
nand U14386 ( n14751, n14754, n10931 );
nand U14387 ( new_g34971_, n14755, n14756 );
nor U14388 ( n14756, n14757, n14758 );
nand U14389 ( n14758, n14759, n14760 );
nand U14390 ( n14760, n14749, n10382 );
nand U14391 ( n14759, n14761, n10545 );
nand U14392 ( n14757, n14762, n14763 );
nand U14393 ( n14763, n137, n14764 );
nand U14394 ( n14764, n14765, n14766 );
nor U14395 ( n14766, n14767, n14768 );
nand U14396 ( n14768, n14769, n14770 );
nand U14397 ( n14770, n14726, n10403 );
nand U14398 ( n14769, n14722, n10502 );
nand U14399 ( n14767, n14771, n14772 );
nand U14400 ( n14772, n14773, n10497 );
nor U14401 ( n14771, n14774, n14775 );
nor U14402 ( n14775, n19319, n14729 );
nor U14403 ( n14774, n14776, n14777 );
nand U14404 ( n14777, n20237, n10769 );
nor U14405 ( n14765, n14778, n14779 );
nand U14406 ( n14779, n14780, n14781 );
nand U14407 ( n14781, n14735, n10547 );
nand U14408 ( n14778, n14782, n14783 );
nand U14409 ( n14783, n14784, g100 );
nor U14410 ( n14782, n14785, n14786 );
nor U14411 ( n14786, n19321, n14787 );
nor U14412 ( n14785, n20005, n14788 );
nand U14413 ( n14762, n14754, n10383 );
nor U14414 ( n14755, n14789, n14790 );
nand U14415 ( n14790, n14791, n14792 );
nand U14416 ( n14792, n14793, n10926 );
nand U14417 ( n14791, n14794, n10927 );
nor U14418 ( n14789, n19325, n14795 );
xor U14419 ( n14707, new_g34975_, new_g34974_ );
nand U14420 ( new_g34974_, n14796, n14797 );
nor U14421 ( n14797, n14798, n14799 );
nand U14422 ( n14799, n14800, n14801 );
nand U14423 ( n14801, n137, n14802 );
nand U14424 ( n14802, n14803, n14804 );
nor U14425 ( n14804, n14805, n14806 );
nand U14426 ( n14806, n14807, n14808 );
nand U14427 ( n14808, n14723, n10498 );
nand U14428 ( n14807, n14738, n10665 );
nand U14429 ( n14805, n14809, n14810 );
nand U14430 ( n14810, n14722, n10372 );
not U14431 ( n14722, n14811 );
nor U14432 ( n14809, n14728, n14812 );
nor U14433 ( n14812, n19962, n14813 );
nor U14434 ( n14728, g35, n14814 );
nor U14435 ( n14803, n14815, n14816 );
nand U14436 ( n14816, n14817, n14818 );
nand U14437 ( n14818, n14734, n10783 );
nand U14438 ( n14817, n14735, n10540 );
nand U14439 ( n14815, n14819, n14820 );
nand U14440 ( n14820, n14739, n10509 );
nand U14441 ( n14819, n14821, n10833 );
nand U14442 ( n14800, n14740, n10367 );
nand U14443 ( n14798, n14822, n14823 );
nand U14444 ( n14823, n14743, n10452 );
nand U14445 ( n14822, n14744, n10453 );
nor U14446 ( n14796, n14824, n14825 );
nand U14447 ( n14825, n14826, n14827 );
nand U14448 ( n14827, n14749, n10932 );
nand U14449 ( n14826, n14750, g46 );
nand U14450 ( n14824, n14828, n14829 );
nand U14451 ( n14829, n14753, n10368 );
nand U14452 ( n14828, n14754, n10933 );
nand U14453 ( new_g34975_, n14830, n14831 );
nor U14454 ( n14831, n14832, n14833 );
nand U14455 ( n14833, n14834, n14835 );
nand U14456 ( n14835, n137, n14836 );
nand U14457 ( n14836, n14837, n14838 );
nor U14458 ( n14838, n14839, n14840 );
nand U14459 ( n14840, n14841, n14842 );
nand U14460 ( n14842, n14723, n10499 );
nor U14461 ( n14841, n14843, n14844 );
nor U14462 ( n14844, n19474, n14811 );
nor U14463 ( n14843, n19473, n14813 );
nand U14464 ( n14839, n14845, n14846 );
nand U14465 ( n14846, n14773, n10794 );
nor U14466 ( n14845, n14847, n14848 );
nor U14467 ( n14848, n19475, n14729 );
nor U14468 ( n14837, n14849, n14850 );
nand U14469 ( n14850, n14851, n14852 );
nand U14470 ( n14852, n14734, n10770 );
nand U14471 ( n14851, n14735, n10541 );
nand U14472 ( n14849, n14853, n14854 );
nand U14473 ( n14854, n20216, n14821 );
nor U14474 ( n14853, n14855, n14856 );
nor U14475 ( n14856, n20223, n14857 );
nor U14476 ( n14855, n20230, n14858 );
nand U14477 ( n14834, n14740, n10515 );
nand U14478 ( n14832, n14859, n14860 );
nand U14479 ( n14860, n14743, n10322 );
nand U14480 ( n14859, n14744, n10323 );
nor U14481 ( n14830, n14861, n14862 );
nand U14482 ( n14862, n14863, n14864 );
nand U14483 ( n14864, n14749, n10934 );
nand U14484 ( n14863, n14750, g47 );
nand U14485 ( n14861, n14865, n14866 );
nand U14486 ( n14866, n14753, n10516 );
nand U14487 ( n14865, n14754, n10935 );
xor U14488 ( n14705, n14867, n14868 );
xor U14489 ( n14868, new_g34977_, new_g34976_ );
nand U14490 ( new_g34976_, n14869, n14870 );
nor U14491 ( n14870, n14871, n14872 );
nand U14492 ( n14872, n14873, n14874 );
nand U14493 ( n14874, n137, n14875 );
nand U14494 ( n14875, n14876, n14877 );
nor U14495 ( n14877, n14878, n14879 );
nand U14496 ( n14879, n14880, n14881 );
nand U14497 ( n14881, n14738, n10705 );
nor U14498 ( n14880, n14882, n14883 );
nor U14499 ( n14883, n19467, n14788 );
nor U14500 ( n14882, n19965, n14811 );
nand U14501 ( n14878, n14884, n14885 );
nand U14502 ( n14885, n14726, n10504 );
nor U14503 ( n14884, n14886, n14887 );
nor U14504 ( n14887, n20008, n14888 );
nor U14505 ( n14886, n19466, n14729 );
nor U14506 ( n14876, n14889, n14890 );
nand U14507 ( n14890, n14780, n14891 );
nand U14508 ( n14891, n14735, n10542 );
nand U14509 ( n14889, n14892, n14893 );
nand U14510 ( n14893, n14734, n10771 );
nor U14511 ( n14892, n14894, n14895 );
nor U14512 ( n14895, n20217, n14787 );
nor U14513 ( n14894, n20224, n14857 );
nand U14514 ( n14873, n14740, n10510 );
nand U14515 ( n14871, n14896, n14897 );
nand U14516 ( n14897, n14743, n10454 );
and U14517 ( n14743, n20088, n14793 );
nand U14518 ( n14896, n14744, n10455 );
and U14519 ( n14744, n20050, n14794 );
nor U14520 ( n14869, n14898, n14899 );
nand U14521 ( n14899, n14900, n14901 );
nand U14522 ( n14901, n14749, n10936 );
nand U14523 ( n14900, n14750, g48 );
nand U14524 ( n14898, n14902, n14903 );
nand U14525 ( n14903, n14753, n10512 );
nand U14526 ( n14902, n14754, n10937 );
nand U14527 ( new_g34977_, n14904, n14905 );
nor U14528 ( n14905, n14906, n14907 );
nand U14529 ( n14907, n14908, n14909 );
nand U14530 ( n14909, n19604, n14753 );
nor U14531 ( n14753, n14910, n14911 );
nand U14532 ( n14908, n14761, n10787 );
nand U14533 ( n14906, n14912, n14913 );
nand U14534 ( n14913, n137, n14914 );
nand U14535 ( n14914, n14915, n14916 );
nor U14536 ( n14916, n14917, n14918 );
nand U14537 ( n14918, n14919, n14920 );
nand U14538 ( n14920, n14738, n10281 );
not U14539 ( n14738, n14858 );
nor U14540 ( n14919, n14921, n14922 );
nor U14541 ( n14922, n20007, n14788 );
nor U14542 ( n14921, n19463, n14811 );
nand U14543 ( n14917, n14923, n14924 );
nand U14544 ( n14924, n14726, n10505 );
nor U14545 ( n14923, n14925, n14926 );
nor U14546 ( n14926, n19462, n14888 );
nor U14547 ( n14925, n19461, n14729 );
nor U14548 ( n14915, n14927, n14928 );
nand U14549 ( n14928, n14929, n14780 );
and U14550 ( n14780, n14930, n14931 );
nand U14551 ( n14931, n14932, n14933 );
nor U14552 ( n14933, n20235, n20236 );
nor U14553 ( n14932, n14934, n14935 );
nor U14554 ( n14929, n14936, n14937 );
nor U14555 ( n14937, n19458, n14938 );
nor U14556 ( n14936, n20220, n14939 );
nand U14557 ( n14927, n14940, n14941 );
nand U14558 ( n14941, n14784, n10386 );
not U14559 ( n14784, n14942 );
nor U14560 ( n14940, n14943, n14944 );
nor U14561 ( n14944, n20218, n14787 );
not U14562 ( n14787, n14821 );
nor U14563 ( n14943, n20225, n14857 );
nand U14564 ( n14912, n19619, n14740 );
and U14565 ( n14740, n14945, n14946 );
nor U14566 ( n14945, n10310, n14911 );
nor U14567 ( n14904, n14947, n14948 );
nand U14568 ( n14948, n14949, n14950 );
nand U14569 ( n14950, n14793, n10586 );
nand U14570 ( n14949, n14794, n10587 );
nor U14571 ( n14947, n19459, n14795 );
xor U14572 ( n14867, new_g34979_, new_g34978_ );
nand U14573 ( new_g34978_, n14951, n14952 );
nor U14574 ( n14952, n14953, n14954 );
nand U14575 ( n14954, n14955, n14956 );
nand U14576 ( n14956, n14749, n10237 );
nand U14577 ( n14955, n14761, n10366 );
nand U14578 ( n14953, n14957, n14958 );
nand U14579 ( n14958, n137, n14959 );
nand U14580 ( n14959, n14960, n14961 );
nor U14581 ( n14961, n14962, n14963 );
nand U14582 ( n14963, n14964, n14965 );
nand U14583 ( n14965, n14723, n10500 );
nor U14584 ( n14964, n14966, n14967 );
nor U14585 ( n14967, n19964, n14811 );
nor U14586 ( n14966, n19960, n14813 );
nand U14587 ( n14962, n14968, n14969 );
nand U14588 ( n14969, n14773, n10494 );
nor U14589 ( n14968, n14847, n14970 );
nor U14590 ( n14970, n14729, n10813 );
nor U14591 ( n14960, n14971, n14972 );
nand U14592 ( n14972, n14973, n14974 );
nand U14593 ( n14974, n14735, n10775 );
nor U14594 ( n14973, n14975, n14976 );
nor U14595 ( n14976, n19338, n14939 );
nor U14596 ( n14975, n20238, n14942 );
nand U14597 ( n14971, n14977, n14978 );
nand U14598 ( n14978, n14821, n10364 );
nor U14599 ( n14977, n14979, n14980 );
nor U14600 ( n14980, n20226, n14857 );
nor U14601 ( n14979, n20232, n14858 );
nand U14602 ( n14957, n14754, n10238 );
nor U14603 ( n14951, n14981, n14982 );
nand U14604 ( n14982, n14983, n14984 );
nand U14605 ( n14984, n20089, n14793 );
nand U14606 ( n14983, n20051, n14794 );
nor U14607 ( n14981, n19340, n14795 );
nand U14608 ( new_g34979_, n14985, n14986 );
nor U14609 ( n14986, n14987, n14988 );
nand U14610 ( n14988, n14989, n14990 );
nand U14611 ( n14990, n14749, n10295 );
nor U14612 ( n14749, n14991, n14935 );
nand U14613 ( n14989, n14761, n10546 );
nor U14614 ( n14761, n14992, n14910 );
or U14615 ( n14992, n14993, n14935 );
nand U14616 ( n14987, n14994, n14995 );
nand U14617 ( n14995, n137, n14996 );
nand U14618 ( n14996, n14997, n14998 );
nor U14619 ( n14998, n14999, n15000 );
nand U14620 ( n15000, n15001, n15002 );
nand U14621 ( n15002, n14723, n10501 );
nor U14622 ( n15001, n15003, n15004 );
nor U14623 ( n15004, n19327, n14811 );
nor U14624 ( n15003, n19328, n14813 );
nand U14625 ( n14999, n15005, n15006 );
nor U14626 ( n15006, n14847, n15007 );
nor U14627 ( n15007, n14776, n15008 );
nand U14628 ( n15008, n20237, n10772 );
nand U14629 ( n14776, n15009, n15010 );
nor U14630 ( n15010, n19498, n20234 );
not U14631 ( n14847, n14930 );
nand U14632 ( n14930, n11013, n15011 );
nand U14633 ( n15011, n14814, n14888 );
and U14634 ( n14814, n15012, n14811 );
nand U14635 ( n14811, n15013, n20236 );
nor U14636 ( n15013, n20235, n15014 );
nor U14637 ( n15012, n14723, n14726 );
not U14638 ( n14726, n14813 );
nand U14639 ( n14813, n15015, n15016 );
nor U14640 ( n15016, n20235, n10343 );
nor U14641 ( n15015, n15017, n10310 );
not U14642 ( n14723, n14788 );
nand U14643 ( n14788, n15018, n15019 );
nor U14644 ( n15018, n10343, n15020 );
nor U14645 ( n15005, n15021, n15022 );
nor U14646 ( n15022, n19326, n14888 );
not U14647 ( n14888, n14773 );
nor U14648 ( n14773, n15020, n15014 );
nor U14649 ( n15021, g30329, n14729 );
or U14650 ( n14729, n15023, n15014 );
nor U14651 ( n14997, n15024, n15025 );
nand U14652 ( n15025, n15026, n15027 );
nand U14653 ( n15027, n14735, n10385 );
not U14654 ( n14735, n14938 );
nand U14655 ( n14938, n15028, n15029 );
nor U14656 ( n15028, n14993, n15023 );
nor U14657 ( n15026, n15030, n15031 );
nor U14658 ( n15031, n19331, n14939 );
not U14659 ( n14939, n14734 );
nor U14660 ( n14734, n15032, n14993 );
nor U14661 ( n15030, n19330, n14942 );
nand U14662 ( n14942, n15033, n15019 );
not U14663 ( n15019, n15017 );
nand U14664 ( n15017, n15034, n19498 );
nor U14665 ( n15034, n20237, n14993 );
nor U14666 ( n15033, n20234, n15020 );
nand U14667 ( n15024, n15035, n15036 );
nand U14668 ( n15036, n14821, g127 );
nor U14669 ( n14821, n14911, n15020 );
nor U14670 ( n15035, n15037, n15038 );
nor U14671 ( n15038, n20227, n14857 );
not U14672 ( n14857, n14739 );
nor U14673 ( n14739, n15032, n14934 );
or U14674 ( n15032, n14935, n15020 );
nand U14675 ( n15020, n20235, n10310 );
nor U14676 ( n15037, n20233, n14858 );
nand U14677 ( n14858, n15009, n15029 );
not U14678 ( n15029, n14935 );
nand U14679 ( n14935, n15039, n20234 );
nor U14680 ( n15039, n19498, n10602 );
nor U14681 ( n15009, n14934, n15023 );
or U14682 ( n14934, n15040, n19497 );
or U14683 ( n15040, n19495, n19496 );
nand U14684 ( n14994, n14754, n10296 );
and U14685 ( n14754, n15041, n15042 );
nor U14686 ( n15042, n19498, n20237 );
nor U14687 ( n15041, n10343, n14991 );
nand U14688 ( n14991, n15043, n14946 );
nor U14689 ( n15043, n14993, n10310 );
nor U14690 ( n14985, n15044, n15045 );
nand U14691 ( n15045, n15046, n15047 );
nand U14692 ( n15047, n14793, n10784 );
nor U14693 ( n14793, n14910, n15014 );
nand U14694 ( n15014, n20234, n15048 );
nand U14695 ( n14910, n14946, n10310 );
nor U14696 ( n14946, n15049, n20235 );
nand U14697 ( n15046, n14794, n10785 );
and U14698 ( n14794, n15050, n137 );
nor U14699 ( n15050, n15023, n14911 );
nand U14700 ( n14911, n15048, n10343 );
and U14701 ( n15048, n15051, n19498 );
nor U14702 ( n15051, n14993, n10602 );
nand U14703 ( n14993, n15052, n19495 );
and U14704 ( n15052, n19497, n19496 );
nand U14705 ( n15023, n20236, n20235 );
nor U14706 ( n15044, n19334, n14795 );
not U14707 ( n14795, n14750 );
nor U14708 ( n14750, g53, n137 );
nand U14709 ( n14703, g55, n15053 );
nand U14710 ( n5095, n15054, n15055 );
nand U14711 ( n15055, n11013, n10260 );
nor U14712 ( n15054, n14702, n15056 );
nor U14713 ( n15056, n19989, n14548 );
nand U14714 ( n5090, n15057, n15058 );
nand U14715 ( n15058, n14693, n10260 );
nand U14716 ( n15057, n14690, n10786 );
nand U14717 ( n5085, n15059, n15060 );
nand U14718 ( n15060, n14702, n10365 );
nor U14719 ( n14702, n15061, n10980 );
nand U14720 ( n15059, n14693, n10786 );
not U14721 ( n14693, n14690 );
nand U14722 ( n14690, g35, n15061 );
nand U14723 ( n15061, n15062, n14498 );
and U14724 ( n14498, n15063, n19280 );
nor U14725 ( n15063, n19979, n15064 );
nor U14726 ( n15062, n15065, n15066 );
nor U14727 ( n15066, n15067, n10307 );
nor U14728 ( n15067, n10352, n15068 );
nand U14729 ( n15068, n20001, n10229 );
nor U14730 ( n15065, n19991, n14497 );
nor U14731 ( n14497, n10661, n10224 );
nand U14732 ( n5080, n15069, n15070 );
nand U14733 ( n15070, n11013, n10605 );
nor U14734 ( n15069, n15071, n15072 );
nor U14735 ( n15072, n10904, n15073 );
nand U14736 ( n15073, n15074, n15075 );
nor U14737 ( n15071, n19987, n15076 );
nand U14738 ( n15076, n15077, n15078 );
not U14739 ( n15078, n15074 );
nor U14740 ( n15074, n15079, n19986 );
nand U14741 ( n5075, n15080, n15081 );
nand U14742 ( n15081, n11014, n10664 );
nor U14743 ( n15080, n15082, n15083 );
nor U14744 ( n15083, n10605, n15084 );
or U14745 ( n15084, n15079, n15085 );
nor U14746 ( n15082, n19986, n15086 );
nand U14747 ( n15086, n15077, n15079 );
nand U14748 ( n15079, n15087, n10664 );
nand U14749 ( n5070, n15088, n15089 );
nand U14750 ( n15089, n15090, n15077 );
nor U14751 ( n15077, n10954, n15085 );
xnor U14752 ( n15090, n19277, n15087 );
and U14753 ( n15087, n15091, n15092 );
nor U14754 ( n15091, n19276, n19985 );
or U14755 ( n15088, g35, n19276 );
nand U14756 ( n5065, n15093, n15094 );
nand U14757 ( n15094, n15095, n15096 );
nand U14758 ( n15096, n14548, n15097 );
nand U14759 ( n15097, n19985, g35 );
nor U14760 ( n15095, n19276, n15085 );
nand U14761 ( n15093, n15098, n10599 );
nand U14762 ( n15098, g35, n15099 );
nand U14763 ( n15099, n15100, n19276 );
nor U14764 ( n15100, n15085, n14582 );
not U14765 ( n15085, n15075 );
nand U14766 ( n5060, n15101, n15102 );
nand U14767 ( n15102, n15103, n15075 );
nand U14768 ( n15075, n15104, n10433 );
nand U14769 ( n15104, n19984, n10256 );
nor U14770 ( n15103, n15105, n15106 );
nor U14771 ( n15106, n19985, n14547 );
nor U14772 ( n15105, n14554, n10599 );
nand U14773 ( n15101, n11014, n10456 );
nand U14774 ( n5055, n15107, n15108 );
nand U14775 ( n15108, n15109, n10256 );
nor U14776 ( n15109, n15110, n15111 );
nor U14777 ( n15111, n19984, n15112 );
nand U14778 ( n15112, n15113, n15114 );
nand U14779 ( n15114, n19275, g35 );
nor U14780 ( n15110, n15115, n10456 );
and U14781 ( n15115, n10899, n15116 );
nand U14782 ( n15107, n11014, n10899 );
nor U14783 ( n5050, n19983, n15117 );
nor U14784 ( n15117, n15118, n10981 );
xnor U14785 ( n15118, n19275, n15116 );
nand U14786 ( n5045, n15119, n15120 );
nand U14787 ( n15120, n15121, n10256 );
nand U14788 ( n15121, n14548, n15122 );
nand U14789 ( n15122, n15123, g35 );
nor U14790 ( n15123, n15124, n15125 );
nor U14791 ( n15125, n19981, n19984 );
nor U14792 ( n15124, n19276, n19986 );
nand U14793 ( n15119, n15126, n10300 );
nand U14794 ( n15126, g35, n15127 );
nand U14795 ( n15127, n19983, n15116 );
nor U14796 ( n15116, n14582, n19981 );
nand U14797 ( n5040, n15128, n15129 );
nand U14798 ( n15129, n15130, n10300 );
nand U14799 ( n15130, n15113, n15131 );
nand U14800 ( n15131, g35, n15132 );
nand U14801 ( n15132, n10256, n10456 );
and U14802 ( n15113, n14548, n15133 );
nand U14803 ( n15133, n19981, g35 );
nor U14804 ( n15128, n15134, n15135 );
nor U14805 ( n15135, n10433, n15136 );
nand U14806 ( n15136, n15137, n15138 );
nor U14807 ( n15138, n19277, n19985 );
nor U14808 ( n15137, n19987, n14563 );
not U14809 ( n14563, n14554 );
nor U14810 ( n14554, n14582, n10981 );
nor U14811 ( n15134, n19981, g35 );
nand U14812 ( n5035, n15139, n15140 );
nand U14813 ( n15140, n14547, n10433 );
nand U14814 ( n15139, n14548, n10773 );
not U14815 ( n14548, n14547 );
nor U14816 ( n14547, n10959, n15092 );
not U14817 ( n15092, n14582 );
nand U14818 ( n14582, n15141, n15142 );
nor U14819 ( n15141, n19280, n19979 );
nor U14820 ( n5030, n10945, n15143 );
nand U14821 ( n15143, n15144, n15145 );
nand U14822 ( n15145, n19980, n15146 );
nand U14823 ( n15144, n15147, n15148 );
nand U14824 ( n5025, n15149, n15150 );
nand U14825 ( n15150, n11014, n10347 );
nand U14826 ( n5020, n15151, n15152 );
nand U14827 ( n15152, n19979, n15142 );
nor U14828 ( n15151, n15153, n15154 );
nor U14829 ( n15154, n19978, g35 );
nor U14830 ( n15153, n10952, n15155 );
nand U14831 ( n15155, n15064, n10347 );
not U14832 ( n15064, n15142 );
nor U14833 ( n15142, n19278, n19978 );
nand U14834 ( n5015, n15156, n15157 );
or U14835 ( n15157, g35, n19280 );
nand U14836 ( n15156, n15158, g35 );
xor U14837 ( n15158, n19278, n19978 );
nand U14838 ( n5010, n15159, n15160 );
or U14839 ( n15160, g35, n19278 );
nand U14840 ( n15159, n15161, g35 );
xor U14841 ( n15161, n15149, n19280 );
nor U14842 ( n5001, g8719, n15162 );
nand U14843 ( n15162, n19278, g35 );
xnor U14844 ( n4986, n15163, n10331 );
nand U14845 ( n15163, n19976, g35 );
nand U14846 ( n4981, n15164, n15165 );
nand U14847 ( n15165, n11014, n10600 );
nand U14848 ( n15164, n15166, g35 );
nand U14849 ( n15166, n15167, n15168 );
nand U14850 ( n15168, n19977, n10331 );
nand U14851 ( n15167, n19976, n10283 );
nand U14852 ( n4976, n15169, n15170 );
nand U14853 ( n15170, n11014, n10365 );
nand U14854 ( n15169, g35, n15171 );
nand U14855 ( n15171, n15172, n15173 );
nand U14856 ( n15173, n15174, n10331 );
nand U14857 ( n15174, n10283, n15175 );
nand U14858 ( n15175, n15176, n15149 );
nand U14859 ( n15149, n15177, n10347 );
nor U14860 ( n15177, n19279, n19978 );
nand U14861 ( n15176, n15178, n15148 );
not U14862 ( n15148, n15146 );
nand U14863 ( n15146, n15179, n15180 );
nor U14864 ( n15180, n19279, n19280 );
nor U14865 ( n15179, n19978, n10347 );
nor U14866 ( n15178, n15147, n10300 );
nor U14867 ( n15147, n14579, n15181 );
and U14868 ( n15181, n15182, n15183 );
nor U14869 ( n15183, n15184, n15185 );
nor U14870 ( n15185, n20002, n15186 );
nor U14871 ( n15186, n15187, n10548 );
xnor U14872 ( n15187, n19283, n19281 );
nor U14873 ( n15184, n15188, n10271 );
nor U14874 ( n15188, n10352, n15189 );
nand U14875 ( n15189, n14524, n14318 );
nand U14876 ( n14318, n19281, n19282 );
nand U14877 ( n14524, n10561, n10278 );
nor U14878 ( n15182, n10229, n10307 );
xnor U14879 ( n14579, n15190, n10229 );
nand U14880 ( n15190, n15191, n15192 );
nand U14881 ( n15192, n15193, n10543 );
xnor U14882 ( n15193, n10415, n20002 );
nor U14883 ( n15191, n15194, n15195 );
nor U14884 ( n15195, n10415, n15196 );
nand U14885 ( n15196, n20002, n10506 );
nor U14886 ( n15194, n19284, n15197 );
nand U14887 ( n15197, n10271, n10544 );
nand U14888 ( n15172, n10283, n10600 );
nand U14889 ( n4971, n15198, n15199 );
nand U14890 ( n15199, n11014, n10349 );
nor U14891 ( n15198, n15200, n15201 );
nor U14892 ( n15201, n19975, n15202 );
nor U14893 ( n15200, n19291, n15203 );
nand U14894 ( n4966, n15204, n15205 );
nand U14895 ( n15205, n11015, n10431 );
nor U14896 ( n15204, n15206, n15207 );
nor U14897 ( n15207, n19974, n15202 );
nor U14898 ( n15206, n19285, n15203 );
nand U14899 ( n4961, n15208, n15209 );
nand U14900 ( n15209, n11015, n10241 );
nor U14901 ( n15208, n15210, n15211 );
nor U14902 ( n15211, n19973, n15202 );
nor U14903 ( n15210, n19286, n15203 );
nand U14904 ( n4956, n15212, n15213 );
nand U14905 ( n15213, n11015, n10458 );
nor U14906 ( n15212, n15214, n15215 );
nor U14907 ( n15215, n19972, n15202 );
nor U14908 ( n15214, n19287, n15203 );
nand U14909 ( n4951, n15216, n15217 );
nand U14910 ( n15217, n11015, n10335 );
nor U14911 ( n15216, n15218, n15219 );
nor U14912 ( n15219, n19971, n15202 );
nor U14913 ( n15218, n19288, n15203 );
nand U14914 ( n4946, n15220, n15221 );
nand U14915 ( n15221, n11015, n10253 );
nor U14916 ( n15220, n15222, n15223 );
nor U14917 ( n15223, n19970, n15202 );
nor U14918 ( n15222, n19289, n15203 );
nand U14919 ( n4941, n15224, n15225 );
nand U14920 ( n15225, n11015, n10230 );
nor U14921 ( n15224, n15226, n15227 );
nor U14922 ( n15227, n19969, n15202 );
nor U14923 ( n15226, n19290, n15203 );
nand U14924 ( n4936, n15228, n15229 );
or U14925 ( n15229, g35, n19291 );
nor U14926 ( n15228, n15230, n15231 );
nor U14927 ( n15231, n19968, n15202 );
nand U14928 ( n15202, g35, n15232 );
nor U14929 ( n15230, n19292, n15203 );
or U14930 ( n15203, n15232, n11024 );
nand U14931 ( n15232, n15233, n19977 );
nor U14932 ( n15233, n19976, n10331 );
nor U14933 ( n4903, n19293, n10991 );
nand U14934 ( n4898, n15234, n15235 );
nand U14935 ( n15235, n11014, n10372 );
nor U14936 ( n15234, n15236, n15237 );
nor U14937 ( n15237, n10657, n15238 );
nor U14938 ( n15236, n19967, n15239 );
nand U14939 ( n15239, n15240, n15238 );
nand U14940 ( n15238, n15241, n10372 );
nand U14941 ( n4893, n15242, n15243 );
nand U14942 ( n15243, n11014, n10639 );
nor U14943 ( n15242, n15244, n15245 );
nor U14944 ( n15245, n15246, n10372 );
nor U14945 ( n15244, n19966, n15247 );
nand U14946 ( n15247, n15240, n15246 );
not U14947 ( n15246, n15241 );
nor U14948 ( n15241, n15248, n19474 );
nand U14949 ( n4888, n15249, n15250 );
nand U14950 ( n15250, n11014, n10646 );
nor U14951 ( n15249, n15251, n15252 );
nor U14952 ( n15252, n15248, n10639 );
nor U14953 ( n15251, n19474, n15253 );
nand U14954 ( n15253, n15240, n15248 );
or U14955 ( n15248, n15254, n19965 );
nand U14956 ( n4883, n15255, n15256 );
nand U14957 ( n15256, n11014, n10647 );
nor U14958 ( n15255, n15257, n15258 );
nor U14959 ( n15258, n15254, n10646 );
nor U14960 ( n15257, n19965, n15259 );
nand U14961 ( n15259, n15240, n15254 );
or U14962 ( n15254, n15260, n19463 );
nand U14963 ( n4878, n15261, n15262 );
nand U14964 ( n15262, n11014, n10648 );
nor U14965 ( n15261, n15263, n15264 );
nor U14966 ( n15264, n15260, n10647 );
nor U14967 ( n15263, n19463, n15265 );
nand U14968 ( n15265, n15240, n15260 );
or U14969 ( n15260, n15266, n19964 );
nand U14970 ( n4873, n15267, n15268 );
nand U14971 ( n15268, n11013, n10649 );
nor U14972 ( n15267, n15269, n15270 );
nor U14973 ( n15270, n15266, n10648 );
nor U14974 ( n15269, n19964, n15271 );
nand U14975 ( n15271, n15240, n15266 );
or U14976 ( n15266, n15272, n19327 );
nand U14977 ( n4868, n15273, n15274 );
nand U14978 ( n15274, n11013, n10502 );
nor U14979 ( n15273, n15275, n15276 );
nor U14980 ( n15276, n15272, n10649 );
nor U14981 ( n15275, n19327, n15277 );
nand U14982 ( n15277, n15240, n15272 );
or U14983 ( n15272, n15278, n19963 );
nand U14984 ( n4863, n15279, n15280 );
nand U14985 ( n15280, n11013, n10503 );
nor U14986 ( n15279, n15281, n15282 );
nor U14987 ( n15282, n15278, n10502 );
nor U14988 ( n15281, n19963, n15283 );
nand U14989 ( n15283, n15240, n15278 );
or U14990 ( n15278, n15284, n19487 );
nand U14991 ( n4858, n15285, n15286 );
nand U14992 ( n15286, n11013, n10650 );
nor U14993 ( n15285, n15287, n15288 );
nor U14994 ( n15288, n15284, n10503 );
nor U14995 ( n15287, n19487, n15289 );
nand U14996 ( n15289, n15240, n15284 );
or U14997 ( n15284, n15290, n19962 );
nand U14998 ( n4853, n15291, n15292 );
nand U14999 ( n15292, n11013, n10651 );
nor U15000 ( n15291, n15293, n15294 );
nor U15001 ( n15294, n15290, n10650 );
nor U15002 ( n15293, n19962, n15295 );
nand U15003 ( n15295, n15240, n15290 );
or U15004 ( n15290, n15296, n19473 );
nand U15005 ( n4848, n15297, n15298 );
nand U15006 ( n15298, n11012, n10504 );
nor U15007 ( n15297, n15299, n15300 );
nor U15008 ( n15300, n15296, n10651 );
nor U15009 ( n15299, n19473, n15301 );
nand U15010 ( n15301, n15240, n15296 );
or U15011 ( n15296, n15302, n19961 );
nand U15012 ( n4843, n15303, n15304 );
nand U15013 ( n15304, n11012, n10505 );
nor U15014 ( n15303, n15305, n15306 );
nor U15015 ( n15306, n15302, n10504 );
nor U15016 ( n15305, n19961, n15307 );
nand U15017 ( n15307, n15240, n15302 );
or U15018 ( n15302, n15308, n19464 );
nand U15019 ( n4838, n15309, n15310 );
nand U15020 ( n15310, n11012, n10652 );
nor U15021 ( n15309, n15311, n15312 );
nor U15022 ( n15312, n15308, n10505 );
nor U15023 ( n15311, n19464, n15313 );
nand U15024 ( n15313, n15240, n15308 );
or U15025 ( n15308, n15314, n19960 );
nand U15026 ( n4833, n15315, n15316 );
nand U15027 ( n15316, n11012, n10653 );
nor U15028 ( n15315, n15317, n15318 );
nor U15029 ( n15318, n15314, n10652 );
nor U15030 ( n15317, n19960, n15319 );
nand U15031 ( n15319, n15240, n15314 );
or U15032 ( n15314, n15320, n19328 );
nand U15033 ( n4828, n15321, n15322 );
nand U15034 ( n15322, n11012, n10403 );
nor U15035 ( n15321, n15323, n15324 );
nor U15036 ( n15324, n15320, n10653 );
nor U15037 ( n15323, n19328, n15325 );
nand U15038 ( n15325, n15240, n15320 );
or U15039 ( n15320, n15326, n15327 );
or U15040 ( n15326, n19959, n15328 );
nand U15041 ( n4823, n15329, n15330 );
nand U15042 ( n15330, n11012, n10834 );
nand U15043 ( n15329, n15331, n15332 );
xnor U15044 ( n15332, n15327, n10403 );
nand U15045 ( n15327, g20763, n15333 );
nand U15046 ( n15333, n19958, g12368 );
nor U15047 ( n15331, n15334, n15335 );
not U15048 ( n15335, n15240 );
nor U15049 ( n15328, n10834, n19958 );
nor U15050 ( n15334, n19966, n19967 );
nand U15051 ( n4805, n15336, n15337 );
or U15052 ( n15337, n11024, n19297 );
or U15053 ( n15336, g35, n19293 );
nand U15054 ( n4800, n15338, n15339 );
nand U15055 ( n15339, n11010, g20763 );
nand U15056 ( n15338, n15340, g35 );
nor U15057 ( n15340, g341, n15341 );
nand U15058 ( n15341, n15342, n10549 );
nand U15059 ( n4795, n15343, n15344 );
nand U15060 ( n15344, n15345, g35 );
nor U15061 ( n15345, n15346, n15347 );
nor U15062 ( n15347, n19294, n10280 );
nand U15063 ( n15343, n15348, n10873 );
nand U15064 ( n15348, n15346, g35 );
nor U15065 ( n15346, g20763, n10697 );
nand U15066 ( n4790, n15349, n15350 );
nand U15067 ( n15350, n11010, n10697 );
nand U15068 ( n15349, n15351, n19294 );
nor U15069 ( n15351, n15352, n10989 );
nor U15070 ( n15352, n10280, n10873 );
nand U15071 ( n4785, n15353, n15354 );
or U15072 ( n15354, g35, n19296 );
nand U15073 ( n15353, n15355, n19296 );
nor U15074 ( n15355, n19295, n10989 );
nand U15075 ( n4776, n15356, n15357 );
nand U15076 ( n15357, n19296, g35 );
nand U15077 ( n15356, n11008, n10280 );
nand U15078 ( n4771, n15358, n15359 );
nand U15079 ( n15359, n11008, n10549 );
nand U15080 ( n15358, g35, n15360 );
nand U15081 ( n15360, n15361, n15362 );
nand U15082 ( n15362, n15363, n15364 );
and U15083 ( n15364, n19957, n19955 );
nor U15084 ( n15363, n10255, n10549 );
nand U15085 ( n15361, n15365, n15366 );
nand U15086 ( n15366, n15367, n19957 );
nor U15087 ( n15367, n15368, n15369 );
nor U15088 ( n15369, n19954, n19956 );
nor U15089 ( n15368, n19955, n10682 );
nand U15090 ( n4761, n15370, n15371 );
nor U15091 ( n15370, n15372, n15373 );
nor U15092 ( n15373, n19297, g35 );
nor U15093 ( n15372, n19955, n10988 );
nand U15094 ( n4756, n15374, n15375 );
nand U15095 ( n15375, n11008, n10395 );
nand U15096 ( n15374, n15365, g35 );
nand U15097 ( n4751, n15376, n15371 );
nor U15098 ( n15376, n15377, n15378 );
nor U15099 ( n15378, n10955, n15379 );
nand U15100 ( n15379, n19955, n10395 );
nor U15101 ( n15377, n19956, g35 );
nand U15102 ( n4746, n15380, n15381 );
or U15103 ( n15381, n15371, n15342 );
nand U15104 ( n15371, g35, n10255 );
nor U15105 ( n15380, n15382, n15383 );
nor U15106 ( n15383, n19955, g35 );
nor U15107 ( n15382, n10955, n15384 );
nand U15108 ( n15384, n15342, n10682 );
not U15109 ( n15342, n15365 );
nand U15110 ( n15365, n15385, n15386 );
nand U15111 ( n15386, n10255, n10395 );
or U15112 ( n15385, n10395, n19955 );
nand U15113 ( n4741, n15387, n15388 );
nand U15114 ( n15388, g6744, g35 );
nand U15115 ( n15387, n11008, n10255 );
and U15116 ( n4736, g6745, g35 );
nand U15117 ( n4731, n15389, n15390 );
nand U15118 ( n15390, n11007, n10774 );
nand U15119 ( n15389, n15391, g35 );
xor U15120 ( n15391, n15392, n15393 );
nand U15121 ( n15393, n15394, n15395 );
nand U15122 ( n15395, n19952, n10774 );
nand U15123 ( n15394, n19953, n15396 );
nand U15124 ( n15396, n19952, n15397 );
nand U15125 ( n15397, n15398, n15399 );
nor U15126 ( n15399, n15400, n15401 );
nand U15127 ( n15401, n19300, n19301 );
nand U15128 ( n15400, n19302, n19303 );
nor U15129 ( n15398, g8919, n15402 );
nand U15130 ( n15402, n19298, n19299 );
nand U15131 ( n4694, n15403, n15404 );
nand U15132 ( n15404, n11007, n10457 );
nand U15133 ( n15403, n15392, g35 );
nand U15134 ( n15392, n15405, n15406 );
nand U15135 ( n15406, n19944, n10366 );
nand U15136 ( n15405, n19941, n19949 );
nand U15137 ( n4657, n15407, n15408 );
or U15138 ( n15408, g35, n19310 );
nand U15139 ( n15407, n15409, g35 );
nand U15140 ( n15409, n15410, n15411 );
nand U15141 ( n15411, n19950, n10457 );
nand U15142 ( n15410, n19951, n15412 );
nand U15143 ( n15412, n19950, n15413 );
nand U15144 ( n15413, n15414, n15415 );
nor U15145 ( n15415, n15416, n15417 );
nand U15146 ( n15417, n19306, n19307 );
nand U15147 ( n15416, n19308, n19309 );
nor U15148 ( n15414, g8788, n15418 );
nand U15149 ( n15418, n19304, n19305 );
nand U15150 ( n4652, n15419, n15420 );
or U15151 ( n15420, g35, n19312 );
nand U15152 ( n15419, n15421, g35 );
nand U15153 ( n4643, n15422, n15423 );
or U15154 ( n15423, g35, n19424 );
nand U15155 ( n15422, n15424, g35 );
xor U15156 ( n15424, n19311, n15421 );
xor U15157 ( n15421, n19312, n19311 );
nand U15158 ( n4638, n15425, n15426 );
or U15159 ( n15426, g35, n19314 );
nand U15160 ( n15425, n15427, g35 );
nand U15161 ( n4629, n15428, n15429 );
nand U15162 ( n15429, n11007, n10545 );
nand U15163 ( n15428, n15430, g35 );
xor U15164 ( n15430, n19313, n15427 );
xor U15165 ( n15427, n19314, n19313 );
nand U15166 ( n4624, n15431, n15432 );
nand U15167 ( n15432, g35, n10545 );
nand U15168 ( n15431, n11007, n10546 );
nand U15169 ( n4619, n15433, n15434 );
nand U15170 ( n15434, g35, n10546 );
nand U15171 ( n15433, n11007, n10366 );
nand U15172 ( n4614, n15435, n15436 );
nand U15173 ( n15436, g35, n10366 );
nand U15174 ( n15435, n11007, n10787 );
nand U15175 ( n4609, n15437, n15438 );
nand U15176 ( n15438, n11007, n10874 );
nand U15177 ( n15437, g35, n15439 );
nand U15178 ( n15439, n19315, n19460 );
nand U15179 ( n4600, n15440, n15441 );
or U15180 ( n15441, g35, n19316 );
nand U15181 ( n15440, n15442, g35 );
nor U15182 ( n15442, g10122, n10874 );
nand U15183 ( n4595, n15443, n15444 );
nand U15184 ( n15444, n19316, g35 );
nand U15185 ( n15443, n11006, n10788 );
nand U15186 ( n4590, n15445, n15446 );
nand U15187 ( n15446, n15447, n10903 );
nand U15188 ( n15447, g35, n15448 );
nand U15189 ( n15448, n15449, n19317 );
nor U15190 ( n15449, n19318, n19947 );
nand U15191 ( n15445, n15450, n10788 );
nand U15192 ( n15450, n15451, n15452 );
nand U15193 ( n15452, n19948, g35 );
nand U15194 ( n4585, n15453, n15454 );
nand U15195 ( n15454, n15455, n10359 );
nand U15196 ( n15455, g35, n15456 );
nand U15197 ( n15456, n19948, n10477 );
or U15198 ( n15453, n15451, n19948 );
nor U15199 ( n15451, n4575, n15457 );
nor U15200 ( n15457, n10359, n10987 );
nand U15201 ( n4580, n15458, n15459 );
nand U15202 ( n15459, n15460, n10477 );
nand U15203 ( n15460, g35, n10359 );
nand U15204 ( n15458, n4575, n10359 );
nor U15205 ( n4575, n10477, n10987 );
nand U15206 ( n4570, n15461, n15462 );
nand U15207 ( n15462, g35, n10547 );
nand U15208 ( n15461, n11023, n10385 );
nand U15209 ( n4565, n15463, n15464 );
nand U15210 ( n15464, g35, n10385 );
nand U15211 ( n15463, n11022, n10775 );
nand U15212 ( n4560, n15465, n15466 );
nand U15213 ( n15466, n11023, n10832 );
nand U15214 ( n15465, g35, n15467 );
nand U15215 ( n15467, n19339, n19345 );
nor U15216 ( n4555, n15468, n10986 );
nor U15217 ( n15468, n10291, n10832 );
nand U15218 ( n4530, n15469, n15470 );
nand U15219 ( n15470, n11022, n10291 );
nand U15220 ( n15469, n15471, g35 );
nand U15221 ( n4525, n15472, n15473 );
nand U15222 ( n15473, n11022, n10872 );
nand U15223 ( n15472, g35, n15474 );
nand U15224 ( n15474, n15475, n15476 );
nand U15225 ( n15476, n19946, n15477 );
xor U15226 ( n15477, n15471, n19342 );
nand U15227 ( n15471, n15478, n15479 );
nand U15228 ( n15479, n19946, g114 );
nand U15229 ( n15478, n10547, g116 );
nand U15230 ( n15475, n19945, n15480 );
xor U15231 ( n15480, n15481, n19343 );
nand U15232 ( n4520, n15482, n15483 );
nand U15233 ( n15483, n15484, n15485 );
not U15234 ( n15485, n15486 );
nor U15235 ( n15482, n15487, n15488 );
nor U15236 ( n15488, n19943, g35 );
nor U15237 ( n15487, n10956, n15489 );
nand U15238 ( n15489, n15486, n10872 );
nand U15239 ( n15486, n15490, n10446 );
nand U15240 ( n4515, n15491, n15492 );
nand U15241 ( n15492, n15493, n15484 );
nor U15242 ( n15491, n15494, n15495 );
nor U15243 ( n15495, n19942, g35 );
nor U15244 ( n15494, n10956, n15496 );
or U15245 ( n15496, n15493, n19943 );
and U15246 ( n15493, n15497, n10446 );
nand U15247 ( n4510, n15498, n15499 );
nand U15248 ( n15499, n15500, n15484 );
nor U15249 ( n15484, n10956, n19941 );
nor U15250 ( n15498, n15501, n15502 );
nor U15251 ( n15502, n19344, g35 );
nor U15252 ( n15501, n10956, n15503 );
or U15253 ( n15503, n15500, n19942 );
and U15254 ( n15500, n15490, n19933 );
and U15255 ( n15490, n15504, n15505 );
nor U15256 ( n15505, n19932, n11218 );
nor U15257 ( n15504, n15506, n10226 );
nand U15258 ( n4505, n15507, n15508 );
or U15259 ( n15508, n15509, n19344 );
nand U15260 ( n15507, n15509, n10905 );
nand U15261 ( n15509, g35, n15510 );
nand U15262 ( n15510, n15497, n19933 );
and U15263 ( n15497, n15511, n15512 );
nor U15264 ( n15512, n11218, n15506 );
not U15265 ( n11218, n11234 );
nor U15266 ( n11234, n10293, n11199 );
not U15267 ( n11199, n15513 );
nor U15268 ( n15511, n10344, n10226 );
nand U15269 ( n4500, n15514, n15515 );
nand U15270 ( n15515, n11021, n10475 );
nand U15271 ( n15514, n15481, g35 );
nand U15272 ( n15481, n15516, n15517 );
nand U15273 ( n15517, n19945, g120 );
nand U15274 ( n15516, n10385, g124 );
nand U15275 ( n4495, n15518, n15519 );
nor U15276 ( n15519, n15520, n15521 );
nor U15277 ( n15521, n19940, g35 );
nor U15278 ( n15520, n10956, n15522 );
nand U15279 ( n15522, n15523, n10475 );
nor U15280 ( n15518, n15524, n15525 );
nor U15281 ( n15525, n10475, n15523 );
nand U15282 ( n15523, n15526, n10462 );
nand U15283 ( n4490, n15527, n15528 );
nor U15284 ( n15528, n15529, n15530 );
nor U15285 ( n15530, n19939, g35 );
nor U15286 ( n15529, n10956, n15531 );
nand U15287 ( n15531, n15532, n10462 );
nor U15288 ( n15527, n15524, n15533 );
nor U15289 ( n15533, n10462, n15532 );
not U15290 ( n15532, n15526 );
nor U15291 ( n15526, n15534, n19939 );
nand U15292 ( n4485, n15535, n15536 );
nor U15293 ( n15535, n15537, n15538 );
nor U15294 ( n15538, n10956, n15539 );
xnor U15295 ( n15539, n19939, n15534 );
or U15296 ( n15534, n15540, n19938 );
nor U15297 ( n15537, n19938, g35 );
nand U15298 ( n4480, n15541, n15542 );
nand U15299 ( n15542, n11021, n10232 );
nor U15300 ( n15541, n15543, n15544 );
nor U15301 ( n15544, n15545, n15546 );
nand U15302 ( n15546, n11194, n10311 );
not U15303 ( n15545, n15547 );
nor U15304 ( n15543, n15548, n15549 );
nand U15305 ( n15549, n15540, n10421 );
nand U15306 ( n15540, n15547, n10232 );
nand U15307 ( n4475, n15550, n15551 );
nand U15308 ( n15551, n15552, n15553 );
xnor U15309 ( n15552, n15547, n19937 );
nor U15310 ( n15547, n15554, n19936 );
nand U15311 ( n15550, n11022, n10226 );
nand U15312 ( n4470, n15555, n15556 );
nor U15313 ( n15556, n15557, n15558 );
nor U15314 ( n15558, n19935, g35 );
nor U15315 ( n15557, n10957, n15559 );
nand U15316 ( n15559, n15554, n10226 );
nor U15317 ( n15555, n15524, n15560 );
nor U15318 ( n15560, n10226, n15554 );
or U15319 ( n15554, n15561, n19935 );
nand U15320 ( n4465, n15562, n15536 );
nor U15321 ( n15562, n15563, n15564 );
nor U15322 ( n15564, n10957, n15565 );
xnor U15323 ( n15565, n19935, n15561 );
nand U15324 ( n15561, n15566, n10611 );
nor U15325 ( n15563, n19934, g35 );
nand U15326 ( n4460, n15567, n15568 );
nand U15327 ( n15568, n11021, n10446 );
nor U15328 ( n15567, n15569, n15570 );
nor U15329 ( n15570, n10611, n15571 );
nand U15330 ( n15571, n15566, n10311 );
nor U15331 ( n15569, n19934, n15572 );
or U15332 ( n15572, n15548, n15566 );
nor U15333 ( n15566, n19932, n19933 );
nand U15334 ( n4455, n15573, n15574 );
nand U15335 ( n15574, n15575, n10344 );
nand U15336 ( n15575, g35, n15576 );
nand U15337 ( n15576, n19933, n10311 );
nand U15338 ( n15573, n15577, n19932 );
nor U15339 ( n15577, n19933, n15548 );
not U15340 ( n15548, n15553 );
nor U15341 ( n15553, n10957, n19346 );
nand U15342 ( n4450, n15578, n15536 );
not U15343 ( n15536, n15524 );
nor U15344 ( n15578, n15579, n15580 );
nor U15345 ( n15580, n19345, g35 );
nor U15346 ( n15579, n10957, n10344 );
nand U15347 ( n4445, n15581, n15582 );
nand U15348 ( n15582, n15524, n15583 );
nand U15349 ( n15583, n15584, n15585 );
nor U15350 ( n15585, n11201, n15586 );
nand U15351 ( n15586, n10293, n10226 );
not U15352 ( n11201, n11194 );
nor U15353 ( n15584, n10344, n15587 );
nand U15354 ( n15587, n19933, n11231 );
not U15355 ( n11231, n15506 );
nand U15356 ( n15506, n19934, n19935 );
nor U15357 ( n15524, n10311, n10986 );
nand U15358 ( n15581, n11021, n10701 );
nor U15359 ( n4425, n19486, n10986 );
nand U15360 ( n4420, n15588, n15589 );
or U15361 ( n15589, n15590, n19525 );
nor U15362 ( n15588, n15591, n15592 );
nor U15363 ( n15592, n10723, n15593 );
nand U15364 ( n15593, n15594, n19930 );
nor U15365 ( n15594, n10957, n11212 );
nor U15366 ( n15591, n19931, n15595 );
nor U15367 ( n15595, n15596, n10986 );
nor U15368 ( n15596, n19930, n11212 );
nand U15369 ( n4415, n15597, n15598 );
nand U15370 ( n15598, n15599, n10723 );
or U15371 ( n15597, n15599, n19930 );
nand U15372 ( n4410, n15600, n15601 );
nand U15373 ( n15601, n11021, n10776 );
nor U15374 ( n15600, n15602, n15603 );
and U15375 ( n15603, n19930, n15604 );
nor U15376 ( n15602, n19930, n15605 );
nand U15377 ( n4405, n15606, n15607 );
nand U15378 ( n15607, n15608, n10776 );
nor U15379 ( n15606, n15609, n15610 );
nor U15380 ( n15610, n10724, n15611 );
nand U15381 ( n15611, n19349, n15604 );
nor U15382 ( n15609, n19348, n15612 );
nor U15383 ( n15612, n15613, n10987 );
nor U15384 ( n15613, n19349, n15614 );
nand U15385 ( n4400, n15615, n15616 );
nand U15386 ( n15616, n15608, n10724 );
nand U15387 ( n15615, n15605, n10564 );
nand U15388 ( n4395, n15617, n15618 );
nand U15389 ( n15618, n15599, n10564 );
nor U15390 ( n15617, n15619, n15620 );
nor U15391 ( n15620, n19520, g35 );
nor U15392 ( n15619, n10957, n15621 );
or U15393 ( n15621, n10564, n11212 );
nand U15394 ( n4390, n15622, n15623 );
nand U15395 ( n15623, n15608, n10698 );
not U15396 ( n15608, n15605 );
nand U15397 ( n15605, g35, n15614 );
nor U15398 ( n15622, n15624, n15625 );
nor U15399 ( n15625, n10484, n15626 );
nand U15400 ( n15626, n15604, n10373 );
nor U15401 ( n15604, n15614, n10987 );
nor U15402 ( n15624, n19929, n15627 );
nor U15403 ( n15627, n15628, n10987 );
nor U15404 ( n15628, n15614, n10373 );
nand U15405 ( n4385, n15629, n15630 );
nand U15406 ( n15630, n11020, n10373 );
nand U15407 ( n15629, n15631, g35 );
nor U15408 ( n15631, n15632, n15633 );
nand U15409 ( n15633, n15634, n15635 );
nand U15410 ( n15635, n15636, n15614 );
nor U15411 ( n15636, n15637, n15638 );
nand U15412 ( n15638, n15639, n10484 );
or U15413 ( n15634, n15639, n15614 );
nand U15414 ( n15614, n15640, n15641 );
nor U15415 ( n15641, n19356, n19899 );
nor U15416 ( n15640, n11105, n15637 );
nor U15417 ( n15632, n15642, n10484 );
and U15418 ( n15642, n15639, n15643 );
nand U15419 ( n4380, n15644, n15645 );
nand U15420 ( n15645, n15599, n10373 );
not U15421 ( n15599, n15590 );
nand U15422 ( n15644, n15590, n10837 );
nand U15423 ( n4375, n15646, n15647 );
nand U15424 ( n15647, n15648, n15649 );
nor U15425 ( n15648, n19350, n15590 );
nand U15426 ( n15646, n10944, n15650 );
nand U15427 ( n15650, n10837, n11212 );
nand U15428 ( n4370, n15651, n15652 );
nand U15429 ( n15652, n15653, n10928 );
nor U15430 ( n15651, n15654, n15655 );
nor U15431 ( n15655, n10958, n15656 );
nand U15432 ( n15656, n15643, n15639 );
nand U15433 ( n15639, n15657, n15658 );
nand U15434 ( n15658, n19899, n15659 );
nand U15435 ( n15659, n15660, n15661 );
nor U15436 ( n15661, n15662, n15663 );
nand U15437 ( n15663, n15664, n15665 );
nand U15438 ( n15665, n15666, n15667 );
nor U15439 ( n15666, n19353, n19921 );
nand U15440 ( n15664, n15668, n15669 );
nor U15441 ( n15668, n19351, n19920 );
nor U15442 ( n15662, n15670, n15671 );
nor U15443 ( n15670, n15672, n15673 );
nor U15444 ( n15673, n19356, n19918 );
nor U15445 ( n15672, n19352, n19922 );
nor U15446 ( n15660, n15674, n15675 );
nand U15447 ( n15675, n15676, n15677 );
nand U15448 ( n15677, n19355, n15678 );
nand U15449 ( n15676, n15679, g11418 );
nand U15450 ( n15679, n15680, n15681 );
nand U15451 ( n15681, n15669, n10795 );
not U15452 ( n15680, n15682 );
nor U15453 ( n15674, n15683, n15684 );
nor U15454 ( n15683, n15685, n15686 );
nor U15455 ( n15686, n19357, n19919 );
nor U15456 ( n15685, n19354, n19923 );
nand U15457 ( n15657, n15687, n10324 );
nand U15458 ( n15687, n15688, n15689 );
nor U15459 ( n15689, n15690, n15691 );
nand U15460 ( n15691, n15692, n15693 );
nand U15461 ( n15693, n15694, n15695 );
nor U15462 ( n15694, n19351, n19910 );
nand U15463 ( n15692, n15696, n15697 );
nor U15464 ( n15696, n19353, n19911 );
nor U15465 ( n15690, n15698, n15699 );
nor U15466 ( n15698, n15700, n15701 );
nor U15467 ( n15701, n19357, n19909 );
nor U15468 ( n15700, n19354, n19913 );
nor U15469 ( n15688, n15702, n15703 );
nand U15470 ( n15703, n15704, n15705 );
nand U15471 ( n15705, n19355, n15682 );
nand U15472 ( n15682, n15706, n15707 );
nand U15473 ( n15707, n15708, n15697 );
nor U15474 ( n15708, n19898, n19927 );
nor U15475 ( n15706, n15709, n15710 );
nor U15476 ( n15710, n15699, n15711 );
nand U15477 ( n15711, n10838, g13966 );
nor U15478 ( n15709, n15671, n15712 );
or U15479 ( n15712, n19926, n19897 );
not U15480 ( n15671, n15695 );
nand U15481 ( n15704, n15713, g11418 );
nand U15482 ( n15713, n15714, n15715 );
nand U15483 ( n15715, n15695, n10796 );
not U15484 ( n15714, n15678 );
nand U15485 ( n15678, n15716, n15717 );
nand U15486 ( n15717, n15718, n15669 );
nor U15487 ( n15718, n19897, n19916 );
nor U15488 ( n15716, n15719, n15720 );
nor U15489 ( n15720, n15684, n15721 );
nand U15490 ( n15721, n10840, g13966 );
nor U15491 ( n15719, n15699, n15722 );
nand U15492 ( n15722, n10839, g16659 );
not U15493 ( n15699, n15667 );
nor U15494 ( n15702, n15723, n11105 );
not U15495 ( n11105, n15669 );
nor U15496 ( n15723, n15724, n15725 );
nor U15497 ( n15725, n19352, n19912 );
nor U15498 ( n15724, n19356, n19928 );
nor U15499 ( n15654, n19928, g35 );
nand U15500 ( n4365, n15726, n15727 );
nand U15501 ( n15727, n11020, n10760 );
nor U15502 ( n15726, n15728, n15729 );
nor U15503 ( n15729, n11212, n15730 );
nor U15504 ( n15728, n19928, n15590 );
nand U15505 ( n15590, g35, n11212 );
nand U15506 ( n11212, n15731, n10396 );
nand U15507 ( n4360, n15732, n15733 );
or U15508 ( n15733, n15734, n15730 );
nor U15509 ( n15732, n15735, n15736 );
nor U15510 ( n15736, n19926, g35 );
nor U15511 ( n15735, n10958, n15737 );
nand U15512 ( n15737, n15734, n10760 );
nand U15513 ( n15734, n15738, n15731 );
nand U15514 ( n4355, n15739, n15740 );
nand U15515 ( n15740, n15741, n10942 );
nor U15516 ( n15739, n15742, n15743 );
nor U15517 ( n15743, n19925, g35 );
nor U15518 ( n15742, n10958, n15744 );
or U15519 ( n15744, n15741, n19926 );
and U15520 ( n15741, n15745, n15731 );
nand U15521 ( n4350, n15746, n15747 );
or U15522 ( n15747, n15748, n15730 );
nor U15523 ( n15746, n15749, n15750 );
nor U15524 ( n15750, n19924, g35 );
nor U15525 ( n15749, n10958, n15751 );
nand U15526 ( n15751, n15748, n10838 );
nand U15527 ( n15748, n15752, n15731 );
nand U15528 ( n4345, n15753, n15754 );
or U15529 ( n15754, n15755, n15730 );
nor U15530 ( n15753, n15756, n15757 );
nor U15531 ( n15757, n19923, g35 );
nor U15532 ( n15756, n10958, n15758 );
nand U15533 ( n15758, n15755, n10795 );
nand U15534 ( n15755, n15759, n15731 );
nor U15535 ( n15731, n19908, n19907 );
nand U15536 ( n4340, n15760, n15761 );
nand U15537 ( n15761, n15762, n10944 );
nor U15538 ( n15760, n15763, n15764 );
nor U15539 ( n15764, n19922, g35 );
nor U15540 ( n15763, n10958, n15765 );
or U15541 ( n15765, n15762, n19923 );
nor U15542 ( n15762, n15766, n19906 );
nand U15543 ( n4335, n15767, n15768 );
nand U15544 ( n15768, n15769, n10943 );
nor U15545 ( n15767, n15770, n15771 );
nor U15546 ( n15771, n19921, g35 );
nor U15547 ( n15770, n10958, n15772 );
or U15548 ( n15772, n15769, n19922 );
nor U15549 ( n15769, n15766, n15773 );
nand U15550 ( n4330, n15774, n15775 );
nand U15551 ( n15775, n15776, n10942 );
nor U15552 ( n15774, n15777, n15778 );
nor U15553 ( n15778, n19920, g35 );
nor U15554 ( n15777, n10958, n15779 );
or U15555 ( n15779, n15776, n19921 );
and U15556 ( n15776, n15780, n15745 );
nand U15557 ( n4325, n15781, n15782 );
nand U15558 ( n15782, n15783, n10944 );
nor U15559 ( n15781, n15784, n15785 );
nor U15560 ( n15785, n19919, g35 );
nor U15561 ( n15784, n10958, n15786 );
or U15562 ( n15786, n15783, n19920 );
nor U15563 ( n15783, n15766, n15787 );
nand U15564 ( n4320, n15788, n15789 );
nand U15565 ( n15789, n15790, n10943 );
nor U15566 ( n15788, n15791, n15792 );
nor U15567 ( n15792, n19918, g35 );
nor U15568 ( n15791, n10958, n15793 );
or U15569 ( n15793, n15790, n19919 );
and U15570 ( n15790, n15780, n15759 );
nand U15571 ( n4315, n15794, n15795 );
nand U15572 ( n15795, n15796, n10942 );
nor U15573 ( n15794, n15797, n15798 );
nor U15574 ( n15798, n19917, g35 );
nor U15575 ( n15797, n10958, n15799 );
or U15576 ( n15799, n15796, n19918 );
nand U15577 ( n4310, n15800, n15801 );
or U15578 ( n15801, n15802, n15730 );
nor U15579 ( n15800, n15803, n15804 );
nor U15580 ( n15804, n19916, g35 );
nor U15581 ( n15803, n10959, n15805 );
nand U15582 ( n15805, n15802, n10839 );
nand U15583 ( n15802, n15806, n15738 );
nand U15584 ( n4305, n15807, n15808 );
nand U15585 ( n15808, n15809, n10944 );
nor U15586 ( n15807, n15810, n15811 );
nor U15587 ( n15811, n19915, g35 );
nor U15588 ( n15810, n10959, n15812 );
or U15589 ( n15812, n15809, n19916 );
and U15590 ( n15809, n15806, n15745 );
nand U15591 ( n4300, n15813, n15814 );
or U15592 ( n15814, n15815, n15730 );
nor U15593 ( n15813, n15816, n15817 );
nor U15594 ( n15817, n19914, g35 );
nor U15595 ( n15816, n10959, n15818 );
nand U15596 ( n15818, n15815, n10840 );
nand U15597 ( n15815, n15806, n15752 );
nand U15598 ( n4295, n15819, n15820 );
or U15599 ( n15820, n15821, n15730 );
nor U15600 ( n15819, n15822, n15823 );
nor U15601 ( n15823, n19913, g35 );
nor U15602 ( n15822, n10959, n15824 );
nand U15603 ( n15824, n15821, n10796 );
nand U15604 ( n15821, n15806, n15759 );
nand U15605 ( n4290, n15825, n15826 );
nand U15606 ( n15826, n15827, n10943 );
nor U15607 ( n15825, n15828, n15829 );
nor U15608 ( n15829, n19912, g35 );
nor U15609 ( n15828, n10959, n15830 );
or U15610 ( n15830, n15827, n19913 );
and U15611 ( n15827, n15831, n10396 );
nand U15612 ( n4285, n15832, n15833 );
nand U15613 ( n15833, n15834, n10942 );
nor U15614 ( n15832, n15835, n15836 );
nor U15615 ( n15836, n19911, g35 );
nor U15616 ( n15835, n10959, n15837 );
or U15617 ( n15837, n15834, n19912 );
and U15618 ( n15834, n15831, n15738 );
nand U15619 ( n4280, n15838, n15839 );
nand U15620 ( n15839, n15840, n10944 );
nor U15621 ( n15838, n15841, n15842 );
nor U15622 ( n15842, n19910, g35 );
nor U15623 ( n15841, n10959, n15843 );
or U15624 ( n15843, n15840, n19911 );
and U15625 ( n15840, n15831, n15745 );
nand U15626 ( n4275, n15844, n15845 );
nand U15627 ( n15845, n15846, n10943 );
nor U15628 ( n15844, n15847, n15848 );
nor U15629 ( n15848, n19909, g35 );
nor U15630 ( n15847, n10959, n15849 );
or U15631 ( n15849, n15846, n19910 );
and U15632 ( n15846, n15831, n15752 );
nand U15633 ( n4270, n15850, n15851 );
nand U15634 ( n15851, n15852, n10942 );
nor U15635 ( n15850, n15853, n15854 );
nor U15636 ( n15854, n19908, g35 );
nor U15637 ( n15853, n10959, n15855 );
or U15638 ( n15855, n15852, n19909 );
and U15639 ( n15852, n15831, n15759 );
and U15640 ( n15759, n15856, n19906 );
nor U15641 ( n15856, n10244, n10463 );
nor U15642 ( n15831, n10595, n10272 );
nand U15643 ( n4265, n15857, n15858 );
nand U15644 ( n15858, n15859, n15860 );
nand U15645 ( n15859, n15861, n15862 );
nand U15646 ( n15862, n4137, n19906 );
nor U15647 ( n15861, n15796, n15863 );
nor U15648 ( n15863, n10959, n15766 );
not U15649 ( n15766, n15780 );
nor U15650 ( n15780, n10272, n19908 );
and U15651 ( n15796, n15806, n10396 );
nor U15652 ( n15806, n10595, n19907 );
nand U15653 ( n15857, n11020, n10272 );
nand U15654 ( n4260, n15864, n15865 );
nand U15655 ( n15865, n15866, n10396 );
nand U15656 ( n15866, g35, n15867 );
nand U15657 ( n15867, n19907, n15860 );
or U15658 ( n15864, n15868, n19907 );
nand U15659 ( n4255, n15869, n15870 );
nand U15660 ( n15870, n15871, n19906 );
nor U15661 ( n15871, n15872, n15773 );
not U15662 ( n15773, n15738 );
nor U15663 ( n15738, n19905, n19904 );
nand U15664 ( n15869, n11020, n10463 );
nand U15665 ( n4250, n15873, n15874 );
nand U15666 ( n15874, n15875, n15860 );
nand U15667 ( n15875, n15787, n15876 );
nand U15668 ( n15876, n15745, g35 );
nor U15669 ( n15745, n10244, n19905 );
not U15670 ( n15787, n15752 );
nor U15671 ( n15752, n10463, n19904 );
nand U15672 ( n15873, n11020, n10244 );
nor U15673 ( n4245, n10244, n15868 );
nand U15674 ( n15868, n15877, n19906 );
nor U15675 ( n15877, n15872, n10988 );
not U15676 ( n15872, n15860 );
nand U15677 ( n15860, n15878, n15879 );
nand U15678 ( n4151, n15880, n15881 );
nand U15679 ( n15881, g35, n10324 );
nand U15680 ( n15880, n11020, n10875 );
nand U15681 ( n4146, n15882, n15883 );
nand U15682 ( n15883, n11020, n10876 );
nand U15683 ( n15882, n15884, g35 );
nor U15684 ( n15884, n15885, g8398 );
nor U15685 ( n15885, n15886, n10875 );
nor U15686 ( n15886, n19903, n10876 );
nor U15687 ( n4137, n10960, n19908 );
nand U15688 ( n4132, n15887, n15888 );
nand U15689 ( n15888, n15889, n15695 );
nor U15690 ( n15887, n15890, n15891 );
nor U15691 ( n15891, n15892, n10988 );
nor U15692 ( n15892, n15893, n15894 );
nor U15693 ( n15894, n15895, n15684 );
nor U15694 ( n15893, n19448, n15643 );
nor U15695 ( n15890, n19902, g35 );
nand U15696 ( n4127, n15896, n15897 );
nand U15697 ( n15897, n15653, n10263 );
nor U15698 ( n15896, n15898, n15899 );
nor U15699 ( n15899, n19901, g35 );
nor U15700 ( n15898, n10960, n15900 );
nand U15701 ( n15900, n15889, n19902 );
nor U15702 ( n15889, n15895, n15637 );
and U15703 ( n15895, n15901, n11120 );
nor U15704 ( n4122, n19900, n15902 );
and U15705 ( n15902, g35, n15903 );
nand U15706 ( n4117, n15904, n15905 );
nand U15707 ( n15905, n11019, n10324 );
nand U15708 ( n15904, n15906, g35 );
nor U15709 ( n15906, n15903, n10692 );
nor U15710 ( n15903, n15907, n19899 );
nand U15711 ( n4112, n15908, n15909 );
or U15712 ( n15909, g35, n19354 );
nand U15713 ( n15908, n15910, g35 );
xnor U15714 ( n15910, n15907, n10324 );
nand U15715 ( n15907, n15911, n15912 );
nor U15716 ( n15912, n19355, n19896 );
nor U15717 ( n15911, n19897, n19898 );
nor U15718 ( n4071, n15913, n15914 );
nand U15719 ( n15914, n15915, n19356 );
nor U15720 ( n15915, n15916, n15917 );
nor U15721 ( n15917, n19897, g13966 );
nor U15722 ( n15916, n19896, g11418 );
nand U15723 ( n15913, n15918, n19357 );
nor U15724 ( n15918, n10960, g16659 );
nor U15725 ( n4066, n19483, n10988 );
nand U15726 ( n4061, n15919, n15920 );
or U15727 ( n15920, n15921, n19535 );
nor U15728 ( n15919, n15922, n15923 );
nor U15729 ( n15923, n10725, n15924 );
nand U15730 ( n15924, n15925, n19894 );
nor U15731 ( n15925, n10960, n11217 );
nor U15732 ( n15922, n19895, n15926 );
nor U15733 ( n15926, n15927, n10988 );
nor U15734 ( n15927, n19894, n11217 );
nand U15735 ( n4056, n15928, n15929 );
nand U15736 ( n15929, n15930, n10725 );
or U15737 ( n15928, n15930, n19894 );
nand U15738 ( n4051, n15931, n15932 );
nand U15739 ( n15932, n11019, n10777 );
nor U15740 ( n15931, n15933, n15934 );
and U15741 ( n15934, n19894, n15935 );
nor U15742 ( n15933, n19894, n15936 );
nand U15743 ( n4046, n15937, n15938 );
nand U15744 ( n15938, n15939, n10777 );
nor U15745 ( n15937, n15940, n15941 );
nor U15746 ( n15941, n10726, n15942 );
nand U15747 ( n15942, n19359, n15935 );
nor U15748 ( n15940, n19358, n15943 );
nor U15749 ( n15943, n15944, n10989 );
nor U15750 ( n15944, n19359, n15945 );
nand U15751 ( n4041, n15946, n15947 );
nand U15752 ( n15947, n15939, n10726 );
nand U15753 ( n15946, n15936, n10565 );
nand U15754 ( n4036, n15948, n15949 );
nand U15755 ( n15949, n15930, n10565 );
nor U15756 ( n15948, n15950, n15951 );
nor U15757 ( n15951, n19519, g35 );
nor U15758 ( n15950, n10961, n15952 );
or U15759 ( n15952, n10565, n11217 );
nand U15760 ( n4031, n15953, n15954 );
nand U15761 ( n15954, n15939, n10640 );
not U15762 ( n15939, n15936 );
nand U15763 ( n15936, g35, n15945 );
nor U15764 ( n15953, n15955, n15956 );
nor U15765 ( n15956, n10485, n15957 );
nand U15766 ( n15957, n15935, n10374 );
nor U15767 ( n15935, n15945, n10989 );
nor U15768 ( n15955, n19893, n15958 );
nor U15769 ( n15958, n15959, n10989 );
nor U15770 ( n15959, n15945, n10374 );
nand U15771 ( n4026, n15960, n15961 );
nand U15772 ( n15961, n11019, n10374 );
nand U15773 ( n15960, n15962, g35 );
nor U15774 ( n15962, n15963, n15964 );
nand U15775 ( n15964, n15965, n15966 );
nand U15776 ( n15966, n15967, n15945 );
nor U15777 ( n15967, n15968, n15969 );
nand U15778 ( n15969, n15970, n10485 );
or U15779 ( n15965, n15970, n15945 );
nand U15780 ( n15945, n15971, n15972 );
nor U15781 ( n15972, n19366, n19863 );
nor U15782 ( n15971, n11110, n15968 );
nor U15783 ( n15963, n15973, n10485 );
and U15784 ( n15973, n15970, n15974 );
nand U15785 ( n4021, n15975, n15976 );
nand U15786 ( n15976, n15930, n10374 );
nand U15787 ( n15975, n15921, n10841 );
nand U15788 ( n4016, n15977, n15978 );
nand U15789 ( n15978, n15979, n15930 );
not U15790 ( n15930, n15921 );
nor U15791 ( n15979, n19360, n15980 );
nand U15792 ( n15977, n10943, n15981 );
nand U15793 ( n15981, n10841, n11217 );
nand U15794 ( n4011, n15982, n15983 );
nand U15795 ( n15983, n15984, n10938 );
nor U15796 ( n15982, n15985, n15986 );
nor U15797 ( n15986, n10961, n15987 );
nand U15798 ( n15987, n15974, n15970 );
nand U15799 ( n15970, n15988, n15989 );
nand U15800 ( n15989, n19863, n15990 );
nand U15801 ( n15990, n15991, n15992 );
nor U15802 ( n15992, n15993, n15994 );
nand U15803 ( n15994, n15995, n15996 );
nand U15804 ( n15996, n15997, n15998 );
nor U15805 ( n15997, n19363, n19885 );
nand U15806 ( n15995, n15999, n16000 );
nor U15807 ( n15999, n19361, n19884 );
nor U15808 ( n15993, n16001, n16002 );
nor U15809 ( n16001, n16003, n16004 );
nor U15810 ( n16004, n19366, n19882 );
nor U15811 ( n16003, n19362, n19886 );
nor U15812 ( n15991, n16005, n16006 );
nand U15813 ( n16006, n16007, n16008 );
nand U15814 ( n16008, n19365, n16009 );
nand U15815 ( n16007, n16010, g11388 );
nand U15816 ( n16010, n16011, n16012 );
nand U15817 ( n16012, n16000, n10797 );
not U15818 ( n16011, n16013 );
nor U15819 ( n16005, n16014, n16015 );
nor U15820 ( n16014, n16016, n16017 );
nor U15821 ( n16017, n19367, n19883 );
nor U15822 ( n16016, n19364, n19887 );
nand U15823 ( n15988, n16018, n10325 );
nand U15824 ( n16018, n16019, n16020 );
nor U15825 ( n16020, n16021, n16022 );
nand U15826 ( n16022, n16023, n16024 );
nand U15827 ( n16024, n16025, n16026 );
nor U15828 ( n16025, n19361, n19874 );
nand U15829 ( n16023, n16027, n16028 );
nor U15830 ( n16027, n19363, n19875 );
nor U15831 ( n16021, n16029, n16030 );
nor U15832 ( n16029, n16031, n16032 );
nor U15833 ( n16032, n19367, n19873 );
nor U15834 ( n16031, n19364, n19877 );
nor U15835 ( n16019, n16033, n16034 );
nand U15836 ( n16034, n16035, n16036 );
nand U15837 ( n16036, n19365, n16013 );
nand U15838 ( n16013, n16037, n16038 );
nand U15839 ( n16038, n16039, n16028 );
nor U15840 ( n16039, n19862, n19891 );
nor U15841 ( n16037, n16040, n16041 );
nor U15842 ( n16041, n16030, n16042 );
nand U15843 ( n16042, n10842, g13926 );
nor U15844 ( n16040, n16002, n16043 );
or U15845 ( n16043, n19890, n19861 );
not U15846 ( n16002, n16026 );
nand U15847 ( n16035, n16044, g11388 );
nand U15848 ( n16044, n16045, n16046 );
nand U15849 ( n16046, n16026, n10798 );
not U15850 ( n16045, n16009 );
nand U15851 ( n16009, n16047, n16048 );
nand U15852 ( n16048, n16049, n16000 );
nor U15853 ( n16049, n19861, n19880 );
nor U15854 ( n16047, n16050, n16051 );
nor U15855 ( n16051, n16015, n16052 );
nand U15856 ( n16052, n10844, g13926 );
nor U15857 ( n16050, n16030, n16053 );
nand U15858 ( n16053, n10843, g16627 );
not U15859 ( n16030, n15998 );
nor U15860 ( n16033, n16054, n11110 );
not U15861 ( n11110, n16000 );
nor U15862 ( n16054, n16055, n16056 );
nor U15863 ( n16056, n19362, n19876 );
nor U15864 ( n16055, n19366, n19892 );
nor U15865 ( n15985, n19892, g35 );
nand U15866 ( n4006, n16057, n16058 );
nand U15867 ( n16058, n11019, n10761 );
nor U15868 ( n16057, n16059, n16060 );
nor U15869 ( n16060, n15730, n11217 );
nor U15870 ( n16059, n19892, n15921 );
nand U15871 ( n15921, g35, n11217 );
nand U15872 ( n11217, n16061, n10397 );
nand U15873 ( n4001, n16062, n16063 );
or U15874 ( n16063, n16064, n15730 );
nor U15875 ( n16062, n16065, n16066 );
nor U15876 ( n16066, n19890, g35 );
nor U15877 ( n16065, n10961, n16067 );
nand U15878 ( n16067, n16064, n10761 );
nand U15879 ( n16064, n16068, n16061 );
nand U15880 ( n3996, n16069, n16070 );
nand U15881 ( n16070, n16071, n10944 );
nor U15882 ( n16069, n16072, n16073 );
nor U15883 ( n16073, n19889, g35 );
nor U15884 ( n16072, n10961, n16074 );
or U15885 ( n16074, n16071, n19890 );
and U15886 ( n16071, n16075, n16061 );
nand U15887 ( n3991, n16076, n16077 );
or U15888 ( n16077, n16078, n15730 );
nor U15889 ( n16076, n16079, n16080 );
nor U15890 ( n16080, n19888, g35 );
nor U15891 ( n16079, n10961, n16081 );
nand U15892 ( n16081, n16078, n10842 );
nand U15893 ( n16078, n16082, n16061 );
nand U15894 ( n3986, n16083, n16084 );
or U15895 ( n16084, n16085, n15730 );
nor U15896 ( n16083, n16086, n16087 );
nor U15897 ( n16087, n19887, g35 );
nor U15898 ( n16086, n10961, n16088 );
nand U15899 ( n16088, n16085, n10797 );
nand U15900 ( n16085, n16089, n16061 );
nor U15901 ( n16061, n19872, n19871 );
nand U15902 ( n3981, n16090, n16091 );
nand U15903 ( n16091, n16092, n10943 );
nor U15904 ( n16090, n16093, n16094 );
nor U15905 ( n16094, n19886, g35 );
nor U15906 ( n16093, n10961, n16095 );
or U15907 ( n16095, n16092, n19887 );
nor U15908 ( n16092, n16096, n19870 );
nand U15909 ( n3976, n16097, n16098 );
nand U15910 ( n16098, n16099, n10942 );
nor U15911 ( n16097, n16100, n16101 );
nor U15912 ( n16101, n19885, g35 );
nor U15913 ( n16100, n10961, n16102 );
or U15914 ( n16102, n16099, n19886 );
nor U15915 ( n16099, n16096, n16103 );
nand U15916 ( n3971, n16104, n16105 );
nand U15917 ( n16105, n16106, n10944 );
nor U15918 ( n16104, n16107, n16108 );
nor U15919 ( n16108, n19884, g35 );
nor U15920 ( n16107, n10962, n16109 );
or U15921 ( n16109, n16106, n19885 );
and U15922 ( n16106, n16110, n16075 );
nand U15923 ( n3966, n16111, n16112 );
nand U15924 ( n16112, n16113, n10943 );
nor U15925 ( n16111, n16114, n16115 );
nor U15926 ( n16115, n19883, g35 );
nor U15927 ( n16114, n10962, n16116 );
or U15928 ( n16116, n16113, n19884 );
nor U15929 ( n16113, n16096, n16117 );
nand U15930 ( n3961, n16118, n16119 );
nand U15931 ( n16119, n16120, n10942 );
nor U15932 ( n16118, n16121, n16122 );
nor U15933 ( n16122, n19882, g35 );
nor U15934 ( n16121, n10962, n16123 );
or U15935 ( n16123, n16120, n19883 );
and U15936 ( n16120, n16110, n16089 );
nand U15937 ( n3956, n16124, n16125 );
nand U15938 ( n16125, n16126, n10944 );
nor U15939 ( n16124, n16127, n16128 );
nor U15940 ( n16128, n19881, g35 );
nor U15941 ( n16127, n10962, n16129 );
or U15942 ( n16129, n16126, n19882 );
nand U15943 ( n3951, n16130, n16131 );
or U15944 ( n16131, n16132, n15730 );
nor U15945 ( n16130, n16133, n16134 );
nor U15946 ( n16134, n19880, g35 );
nor U15947 ( n16133, n10962, n16135 );
nand U15948 ( n16135, n16132, n10843 );
nand U15949 ( n16132, n16136, n16068 );
nand U15950 ( n3946, n16137, n16138 );
nand U15951 ( n16138, n16139, n10943 );
nor U15952 ( n16137, n16140, n16141 );
nor U15953 ( n16141, n19879, g35 );
nor U15954 ( n16140, n10962, n16142 );
or U15955 ( n16142, n16139, n19880 );
and U15956 ( n16139, n16136, n16075 );
nand U15957 ( n3941, n16143, n16144 );
or U15958 ( n16144, n16145, n15730 );
nor U15959 ( n16143, n16146, n16147 );
nor U15960 ( n16147, n19878, g35 );
nor U15961 ( n16146, n10962, n16148 );
nand U15962 ( n16148, n16145, n10844 );
nand U15963 ( n16145, n16136, n16082 );
nand U15964 ( n3936, n16149, n16150 );
or U15965 ( n16150, n16151, n15730 );
nor U15966 ( n16149, n16152, n16153 );
nor U15967 ( n16153, n19877, g35 );
nor U15968 ( n16152, n10962, n16154 );
nand U15969 ( n16154, n16151, n10798 );
nand U15970 ( n16151, n16136, n16089 );
nand U15971 ( n3931, n16155, n16156 );
nand U15972 ( n16156, n16157, n10942 );
nor U15973 ( n16155, n16158, n16159 );
nor U15974 ( n16159, n19876, g35 );
nor U15975 ( n16158, n10962, n16160 );
or U15976 ( n16160, n16157, n19877 );
and U15977 ( n16157, n16161, n10397 );
nand U15978 ( n3926, n16162, n16163 );
nand U15979 ( n16163, n16164, n10944 );
nor U15980 ( n16162, n16165, n16166 );
nor U15981 ( n16166, n19875, g35 );
nor U15982 ( n16165, n10962, n16167 );
or U15983 ( n16167, n16164, n19876 );
and U15984 ( n16164, n16161, n16068 );
nand U15985 ( n3921, n16168, n16169 );
nand U15986 ( n16169, n16170, n10943 );
nor U15987 ( n16168, n16171, n16172 );
nor U15988 ( n16172, n19874, g35 );
nor U15989 ( n16171, n10962, n16173 );
or U15990 ( n16173, n16170, n19875 );
and U15991 ( n16170, n16161, n16075 );
nand U15992 ( n3916, n16174, n16175 );
nand U15993 ( n16175, n16176, n10942 );
nor U15994 ( n16174, n16177, n16178 );
nor U15995 ( n16178, n19873, g35 );
nor U15996 ( n16177, n10962, n16179 );
or U15997 ( n16179, n16176, n19874 );
and U15998 ( n16176, n16161, n16082 );
nand U15999 ( n3911, n16180, n16181 );
nand U16000 ( n16181, n16182, n10944 );
nor U16001 ( n16180, n16183, n16184 );
nor U16002 ( n16184, n19872, g35 );
nor U16003 ( n16183, n10963, n16185 );
or U16004 ( n16185, n16182, n19873 );
and U16005 ( n16182, n16161, n16089 );
and U16006 ( n16089, n16186, n19870 );
nor U16007 ( n16186, n10245, n10464 );
nor U16008 ( n16161, n10596, n10273 );
nand U16009 ( n3906, n16187, n16188 );
nand U16010 ( n16188, n16189, n16190 );
nand U16011 ( n16189, n16191, n16192 );
nand U16012 ( n16192, n3778, n19870 );
nor U16013 ( n16191, n16126, n16193 );
nor U16014 ( n16193, n10963, n16096 );
not U16015 ( n16096, n16110 );
nor U16016 ( n16110, n10273, n19872 );
and U16017 ( n16126, n16136, n10397 );
nor U16018 ( n16136, n10596, n19871 );
nand U16019 ( n16187, n11019, n10273 );
nand U16020 ( n3901, n16194, n16195 );
nand U16021 ( n16195, n16196, n10397 );
nand U16022 ( n16196, g35, n16197 );
nand U16023 ( n16197, n19871, n16190 );
or U16024 ( n16194, n16198, n19871 );
nand U16025 ( n3896, n16199, n16200 );
nand U16026 ( n16200, n16201, n19870 );
nor U16027 ( n16201, n16202, n16103 );
not U16028 ( n16103, n16068 );
nor U16029 ( n16068, n19869, n19868 );
nand U16030 ( n16199, n11019, n10464 );
nand U16031 ( n3891, n16203, n16204 );
nand U16032 ( n16204, n16205, n16190 );
nand U16033 ( n16205, n16117, n16206 );
nand U16034 ( n16206, n16075, g35 );
nor U16035 ( n16075, n10245, n19869 );
not U16036 ( n16117, n16082 );
nor U16037 ( n16082, n10464, n19868 );
nand U16038 ( n16203, n11018, n10245 );
nor U16039 ( n3886, n10245, n16198 );
nand U16040 ( n16198, n16207, n19870 );
nor U16041 ( n16207, n16202, n10990 );
not U16042 ( n16202, n16190 );
nand U16043 ( n16190, n16208, n15879 );
nand U16044 ( n3792, n16209, n16210 );
nand U16045 ( n16210, g35, n10325 );
nand U16046 ( n16209, n11018, n10877 );
nand U16047 ( n3787, n16211, n16212 );
nand U16048 ( n16212, n11018, n10878 );
nand U16049 ( n16211, n16213, g35 );
nor U16050 ( n16213, n16214, g8342 );
nor U16051 ( n16214, n16215, n10877 );
nor U16052 ( n16215, n19867, n10878 );
nor U16053 ( n3778, n10963, n19872 );
nand U16054 ( n3773, n16216, n16217 );
nand U16055 ( n16217, n16218, n16026 );
nor U16056 ( n16216, n16219, n16220 );
nor U16057 ( n16220, n16221, n10990 );
nor U16058 ( n16221, n16222, n16223 );
nor U16059 ( n16223, n16224, n16015 );
nor U16060 ( n16222, n19449, n15974 );
nor U16061 ( n16219, n19866, g35 );
nand U16062 ( n3768, n16225, n16226 );
nand U16063 ( n16226, n15984, n10264 );
nor U16064 ( n16225, n16227, n16228 );
nor U16065 ( n16228, n19865, g35 );
nor U16066 ( n16227, n10949, n16229 );
nand U16067 ( n16229, n16218, n19866 );
nor U16068 ( n16218, n16224, n15968 );
nor U16069 ( n16224, n16230, n11109 );
nor U16070 ( n3763, n19864, n16231 );
and U16071 ( n16231, g35, n16232 );
nand U16072 ( n3758, n16233, n16234 );
nand U16073 ( n16234, n11018, n10325 );
nand U16074 ( n16233, n16235, g35 );
nor U16075 ( n16235, n16232, n10693 );
nor U16076 ( n16232, n16236, n19863 );
nand U16077 ( n3753, n16237, n16238 );
or U16078 ( n16238, g35, n19364 );
nand U16079 ( n16237, n16239, g35 );
xnor U16080 ( n16239, n16236, n10325 );
nand U16081 ( n16236, n16240, n16241 );
nor U16082 ( n16241, n19365, n19860 );
nor U16083 ( n16240, n19861, n19862 );
nor U16084 ( n3712, n16242, n16243 );
nand U16085 ( n16243, n16244, n19366 );
nor U16086 ( n16244, n16245, n16246 );
nor U16087 ( n16246, n19861, g13926 );
nor U16088 ( n16245, n19860, g11388 );
nand U16089 ( n16242, n16247, n19367 );
nor U16090 ( n16247, n10945, g16627 );
nor U16091 ( n3707, n19477, n10990 );
nand U16092 ( n3702, n16248, n16249 );
or U16093 ( n16249, n16250, n19537 );
nor U16094 ( n16248, n16251, n16252 );
nor U16095 ( n16252, n10727, n16253 );
nand U16096 ( n16253, n16254, n19858 );
nor U16097 ( n16254, n11202, n10990 );
nor U16098 ( n16251, n19859, n16255 );
nor U16099 ( n16255, n16256, n10990 );
nor U16100 ( n16256, n19858, n11202 );
nand U16101 ( n3697, n16257, n16258 );
nand U16102 ( n16258, n16259, n10727 );
or U16103 ( n16257, n16259, n19858 );
nand U16104 ( n3692, n16260, n16261 );
nand U16105 ( n16261, n11018, n10778 );
nor U16106 ( n16260, n16262, n16263 );
and U16107 ( n16263, n19858, n16264 );
nor U16108 ( n16262, n19858, n16265 );
nand U16109 ( n3687, n16266, n16267 );
nand U16110 ( n16267, n16268, n10778 );
nor U16111 ( n16266, n16269, n16270 );
nor U16112 ( n16270, n10728, n16271 );
nand U16113 ( n16271, n19369, n16264 );
nor U16114 ( n16269, n19368, n16272 );
nor U16115 ( n16272, n16273, n10990 );
nor U16116 ( n16273, n19369, n16274 );
nand U16117 ( n3682, n16275, n16276 );
nand U16118 ( n16276, n16268, n10728 );
not U16119 ( n16268, n16265 );
nand U16120 ( n16275, n16265, n10566 );
nand U16121 ( n16265, g35, n16274 );
nand U16122 ( n3677, n16277, n16278 );
nand U16123 ( n16278, n16259, n10566 );
nor U16124 ( n16277, n16279, n16280 );
nor U16125 ( n16280, n19518, g35 );
nor U16126 ( n16279, n10945, n16281 );
or U16127 ( n16281, n10566, n11202 );
nand U16128 ( n3672, n16282, n16283 );
nand U16129 ( n16283, n16284, n16274 );
nor U16130 ( n16282, n16285, n16286 );
nor U16131 ( n16286, n10486, n16287 );
nand U16132 ( n16287, n16264, n10375 );
nor U16133 ( n16264, n16274, n10991 );
nor U16134 ( n16285, n19857, n16288 );
nor U16135 ( n16288, n16289, n10991 );
nor U16136 ( n16289, n16274, n10375 );
nand U16137 ( n3667, n16290, n16291 );
nand U16138 ( n16291, n11018, n10375 );
nand U16139 ( n16290, n16292, g35 );
nor U16140 ( n16292, n16293, n16294 );
nand U16141 ( n16294, n16295, n16296 );
nand U16142 ( n16296, n16297, n16274 );
nor U16143 ( n16297, n16298, n16299 );
nand U16144 ( n16299, n16300, n10486 );
or U16145 ( n16295, n16300, n16274 );
nand U16146 ( n16274, n16301, n16302 );
nor U16147 ( n16302, n19376, n19826 );
nor U16148 ( n16301, n11119, n16298 );
nor U16149 ( n16293, n16303, n10486 );
and U16150 ( n16303, n16300, n16304 );
nand U16151 ( n3662, n16305, n16306 );
nand U16152 ( n16306, n16259, n10375 );
nand U16153 ( n16305, n16250, n10845 );
nand U16154 ( n3657, n16307, n16308 );
nand U16155 ( n16308, n16309, n16259 );
not U16156 ( n16259, n16250 );
nor U16157 ( n16309, n19370, n15980 );
nand U16158 ( n16307, n10942, n16310 );
nand U16159 ( n16310, n10845, n11202 );
nand U16160 ( n3652, n16311, n16312 );
nand U16161 ( n16312, n16313, n10894 );
nor U16162 ( n16311, n16314, n16315 );
nor U16163 ( n16315, n10945, n16316 );
nand U16164 ( n16316, n16304, n16300 );
nand U16165 ( n16300, n16317, n16318 );
nand U16166 ( n16318, n19826, n16319 );
nand U16167 ( n16319, n16320, n16321 );
nor U16168 ( n16321, n16322, n16323 );
nand U16169 ( n16323, n16324, n16325 );
nand U16170 ( n16325, n16326, n16327 );
nor U16171 ( n16326, n19373, n19849 );
nand U16172 ( n16324, n16328, n16329 );
nor U16173 ( n16328, n19371, n19848 );
nor U16174 ( n16322, n16330, n16331 );
nor U16175 ( n16330, n16332, n16333 );
nor U16176 ( n16333, n19376, n19846 );
nor U16177 ( n16332, n19372, n19850 );
nor U16178 ( n16320, n16334, n16335 );
nand U16179 ( n16335, n16336, n16337 );
nand U16180 ( n16337, n19375, n16338 );
nand U16181 ( n16336, n16339, g11349 );
nand U16182 ( n16339, n16340, n16341 );
nand U16183 ( n16341, n16329, n10799 );
not U16184 ( n16340, n16342 );
nor U16185 ( n16334, n16343, n16344 );
nor U16186 ( n16343, n16345, n16346 );
nor U16187 ( n16346, n19377, n19847 );
nor U16188 ( n16345, n19374, n19851 );
nand U16189 ( n16317, n16347, n10326 );
nand U16190 ( n16347, n16348, n16349 );
nor U16191 ( n16349, n16350, n16351 );
nand U16192 ( n16351, n16352, n16353 );
nand U16193 ( n16353, n16354, n16355 );
nor U16194 ( n16354, n19371, n19838 );
nand U16195 ( n16352, n16356, n16357 );
nor U16196 ( n16356, n19373, n19839 );
nor U16197 ( n16350, n16358, n16359 );
nor U16198 ( n16358, n16360, n16361 );
nor U16199 ( n16361, n19377, n19837 );
nor U16200 ( n16360, n19374, n19841 );
nor U16201 ( n16348, n16362, n16363 );
nand U16202 ( n16363, n16364, n16365 );
nand U16203 ( n16365, n19375, n16342 );
nand U16204 ( n16342, n16366, n16367 );
nand U16205 ( n16367, n16368, n16357 );
nor U16206 ( n16368, n19825, n19855 );
nor U16207 ( n16366, n16369, n16370 );
nor U16208 ( n16370, n16359, n16371 );
nand U16209 ( n16371, n10846, g13895 );
nor U16210 ( n16369, n16331, n16372 );
or U16211 ( n16372, n19854, n19824 );
nand U16212 ( n16364, n16373, g11349 );
nand U16213 ( n16373, n16374, n16375 );
nand U16214 ( n16375, n16355, n10800 );
not U16215 ( n16374, n16338 );
nand U16216 ( n16338, n16376, n16377 );
nand U16217 ( n16377, n16378, n16329 );
nor U16218 ( n16378, n19824, n19844 );
nor U16219 ( n16376, n16379, n16380 );
nor U16220 ( n16380, n16344, n16381 );
nand U16221 ( n16381, n10848, g13895 );
not U16222 ( n16344, n16357 );
nor U16223 ( n16379, n16359, n16382 );
nand U16224 ( n16382, n10847, g16603 );
nor U16225 ( n16362, n16383, n11119 );
nor U16226 ( n16383, n16384, n16385 );
nor U16227 ( n16385, n19372, n19840 );
nor U16228 ( n16384, n19376, n19856 );
nor U16229 ( n16314, n19856, g35 );
nand U16230 ( n3647, n16386, n16387 );
nand U16231 ( n16387, n11018, n10762 );
nor U16232 ( n16386, n16388, n16389 );
nor U16233 ( n16389, n11202, n15730 );
nor U16234 ( n16388, n19856, n16250 );
nand U16235 ( n16250, g35, n11202 );
nand U16236 ( n11202, n16390, n10336 );
nand U16237 ( n3642, n16391, n16392 );
or U16238 ( n16392, n16393, n15730 );
nor U16239 ( n16391, n16394, n16395 );
nor U16240 ( n16395, n19854, g35 );
nor U16241 ( n16394, n10945, n16396 );
nand U16242 ( n16396, n16393, n10762 );
nand U16243 ( n16393, n16397, n16390 );
nand U16244 ( n3637, n16398, n16399 );
nand U16245 ( n16399, n16400, n10943 );
nor U16246 ( n16398, n16401, n16402 );
nor U16247 ( n16402, n19853, g35 );
nor U16248 ( n16401, n10946, n16403 );
or U16249 ( n16403, n16400, n19854 );
and U16250 ( n16400, n16404, n16390 );
nand U16251 ( n3632, n16405, n16406 );
or U16252 ( n16406, n16407, n15730 );
nor U16253 ( n16405, n16408, n16409 );
nor U16254 ( n16409, n19852, g35 );
nor U16255 ( n16408, n10946, n16410 );
nand U16256 ( n16410, n16407, n10846 );
nand U16257 ( n16407, n16411, n16390 );
nand U16258 ( n3627, n16412, n16413 );
or U16259 ( n16413, n16414, n15730 );
nor U16260 ( n16412, n16415, n16416 );
nor U16261 ( n16416, n19851, g35 );
nor U16262 ( n16415, n10946, n16417 );
nand U16263 ( n16417, n16414, n10799 );
nand U16264 ( n16414, n16418, n16390 );
nor U16265 ( n16390, n19836, n19835 );
nand U16266 ( n3622, n16419, n16420 );
nand U16267 ( n16420, n16421, n10942 );
nor U16268 ( n16419, n16422, n16423 );
nor U16269 ( n16423, n19850, g35 );
nor U16270 ( n16422, n10946, n16424 );
or U16271 ( n16424, n16421, n19851 );
and U16272 ( n16421, n16425, n10336 );
nand U16273 ( n3617, n16426, n16427 );
nand U16274 ( n16427, n16428, n10944 );
nor U16275 ( n16426, n16429, n16430 );
nor U16276 ( n16430, n19849, g35 );
nor U16277 ( n16429, n10946, n16431 );
or U16278 ( n16431, n16428, n19850 );
and U16279 ( n16428, n16425, n16397 );
nand U16280 ( n3612, n16432, n16433 );
nand U16281 ( n16433, n16434, n10943 );
nor U16282 ( n16432, n16435, n16436 );
nor U16283 ( n16436, n19848, g35 );
nor U16284 ( n16435, n10946, n16437 );
or U16285 ( n16437, n16434, n19849 );
and U16286 ( n16434, n16425, n16404 );
nand U16287 ( n3607, n16438, n16439 );
nand U16288 ( n16439, n16440, n10942 );
nor U16289 ( n16438, n16441, n16442 );
nor U16290 ( n16442, n19847, g35 );
nor U16291 ( n16441, n10946, n16443 );
or U16292 ( n16443, n16440, n19848 );
and U16293 ( n16440, n16425, n16411 );
nand U16294 ( n3602, n16444, n16445 );
nand U16295 ( n16445, n16446, n10944 );
nor U16296 ( n16444, n16447, n16448 );
nor U16297 ( n16448, n19846, g35 );
nor U16298 ( n16447, n10946, n16449 );
or U16299 ( n16449, n16446, n19847 );
and U16300 ( n16446, n16425, n16418 );
nand U16301 ( n3597, n16450, n16451 );
nand U16302 ( n16451, n16452, n10943 );
nor U16303 ( n16450, n16453, n16454 );
nor U16304 ( n16454, n19845, g35 );
nor U16305 ( n16453, n10946, n16455 );
or U16306 ( n16455, n16452, n19846 );
nand U16307 ( n3592, n16456, n16457 );
or U16308 ( n16457, n16458, n15730 );
nor U16309 ( n16456, n16459, n16460 );
nor U16310 ( n16460, n19844, g35 );
nor U16311 ( n16459, n10946, n16461 );
nand U16312 ( n16461, n16458, n10847 );
nand U16313 ( n16458, n16462, n16397 );
nand U16314 ( n3587, n16463, n16464 );
nand U16315 ( n16464, n16465, n10942 );
nor U16316 ( n16463, n16466, n16467 );
nor U16317 ( n16467, n19843, g35 );
nor U16318 ( n16466, n10946, n16468 );
or U16319 ( n16468, n16465, n19844 );
and U16320 ( n16465, n16462, n16404 );
nand U16321 ( n3582, n16469, n16470 );
or U16322 ( n16470, n16471, n15730 );
nor U16323 ( n16469, n16472, n16473 );
nor U16324 ( n16473, n19842, g35 );
nor U16325 ( n16472, n10946, n16474 );
nand U16326 ( n16474, n16471, n10848 );
nand U16327 ( n16471, n16462, n16411 );
nand U16328 ( n3577, n16475, n16476 );
or U16329 ( n16476, n16477, n15730 );
nor U16330 ( n16475, n16478, n16479 );
nor U16331 ( n16479, n19841, g35 );
nor U16332 ( n16478, n10947, n16480 );
nand U16333 ( n16480, n16477, n10800 );
nand U16334 ( n16477, n16462, n16418 );
nand U16335 ( n3572, n16481, n16482 );
nand U16336 ( n16482, n16483, n10944 );
nor U16337 ( n16481, n16484, n16485 );
nor U16338 ( n16485, n19840, g35 );
nor U16339 ( n16484, n10947, n16486 );
or U16340 ( n16486, n16483, n19841 );
and U16341 ( n16483, n16487, n10336 );
nand U16342 ( n3567, n16488, n16489 );
nand U16343 ( n16489, n16490, n10943 );
nor U16344 ( n16488, n16491, n16492 );
nor U16345 ( n16492, n19839, g35 );
nor U16346 ( n16491, n10947, n16493 );
or U16347 ( n16493, n16490, n19840 );
and U16348 ( n16490, n16487, n16397 );
nand U16349 ( n3562, n16494, n16495 );
nand U16350 ( n16495, n16496, n10942 );
nor U16351 ( n16494, n16497, n16498 );
nor U16352 ( n16498, n19838, g35 );
nor U16353 ( n16497, n10947, n16499 );
or U16354 ( n16499, n16496, n19839 );
and U16355 ( n16496, n16487, n16404 );
nand U16356 ( n3557, n16500, n16501 );
nand U16357 ( n16501, n16502, n10944 );
nor U16358 ( n16500, n16503, n16504 );
nor U16359 ( n16504, n19837, g35 );
nor U16360 ( n16503, n10947, n16505 );
or U16361 ( n16505, n16502, n19838 );
and U16362 ( n16502, n16487, n16411 );
nand U16363 ( n3552, n16506, n16507 );
nand U16364 ( n16507, n16508, n10943 );
nor U16365 ( n16506, n16509, n16510 );
nor U16366 ( n16510, n19836, g35 );
nor U16367 ( n16509, n10947, n16511 );
or U16368 ( n16511, n16508, n19837 );
and U16369 ( n16508, n16487, n16418 );
and U16370 ( n16418, n16512, n19834 );
nor U16371 ( n16512, n10276, n10465 );
nor U16372 ( n16487, n10266, n10432 );
nand U16373 ( n3547, n16513, n16514 );
nand U16374 ( n16514, n16515, n16516 );
nand U16375 ( n16516, n16517, n16518 );
nand U16376 ( n16518, n19834, n10266 );
nor U16377 ( n16517, n16425, n16452 );
and U16378 ( n16452, n16462, n10336 );
nor U16379 ( n16462, n10266, n19835 );
nor U16380 ( n16425, n10432, n19836 );
nand U16381 ( n16513, n11017, n10432 );
nand U16382 ( n3542, n16519, n16520 );
nand U16383 ( n16520, n16521, n10336 );
nand U16384 ( n16521, g35, n16522 );
nand U16385 ( n16522, n19835, n16523 );
nand U16386 ( n16519, n16524, n19834 );
nor U16387 ( n16524, n19835, n16525 );
nand U16388 ( n3537, n16526, n16527 );
nand U16389 ( n16527, n16528, n19834 );
and U16390 ( n16528, n16523, n16397 );
nor U16391 ( n16397, n19833, n19832 );
nand U16392 ( n16526, n11017, n10465 );
nand U16393 ( n3532, n16529, n16530 );
nand U16394 ( n16530, n11017, n10276 );
nor U16395 ( n16529, n16531, n16532 );
and U16396 ( n16532, n16404, n16515 );
not U16397 ( n16515, n16525 );
nor U16398 ( n16404, n10276, n19833 );
and U16399 ( n16531, n16523, n16411 );
nor U16400 ( n16411, n10465, n19832 );
nor U16401 ( n3527, n16525, n16533 );
nand U16402 ( n16533, n19834, n19832 );
nand U16403 ( n16525, g35, n16523 );
nand U16404 ( n16523, n15879, n11194 );
nand U16405 ( n3433, n16534, n16535 );
nand U16406 ( n16535, g35, n10326 );
nand U16407 ( n16534, n11017, n10879 );
nand U16408 ( n3428, n16536, n16537 );
nand U16409 ( n16537, n11017, n10880 );
nand U16410 ( n16536, n16538, g35 );
nor U16411 ( n16538, n16539, g8277 );
nor U16412 ( n16539, n16540, n10879 );
nor U16413 ( n16540, n19831, n10880 );
nor U16414 ( n3419, n19836, n10991 );
nand U16415 ( n3414, n16541, n16542 );
nand U16416 ( n16542, n11017, n10243 );
nand U16417 ( n16541, n16543, g35 );
nor U16418 ( n16543, n16544, n16545 );
nor U16419 ( n16545, n16357, n16546 );
nand U16420 ( n16546, n16547, n16548 );
nand U16421 ( n16548, n16355, n16304 );
nand U16422 ( n16547, n16298, n10472 );
nand U16423 ( n3409, n16549, n16550 );
nand U16424 ( n16550, n16313, n10243 );
nor U16425 ( n16549, n16551, n16552 );
nor U16426 ( n16552, n19828, g35 );
nor U16427 ( n16551, n10948, n16553 );
nand U16428 ( n16553, n16554, n19829 );
nor U16429 ( n16554, n16544, n16298 );
and U16430 ( n16544, n16555, n16556 );
nor U16431 ( n16556, n19588, n11174 );
nor U16432 ( n16555, n16298, n16557 );
nor U16433 ( n3404, n19827, n16558 );
and U16434 ( n16558, g35, n16559 );
nand U16435 ( n3399, n16560, n16561 );
nand U16436 ( n16561, n11017, n10326 );
nand U16437 ( n16560, n16562, g35 );
nor U16438 ( n16562, n16559, n10740 );
nor U16439 ( n16559, n16563, n19826 );
nand U16440 ( n3394, n16564, n16565 );
or U16441 ( n16565, g35, n19374 );
nand U16442 ( n16564, n16566, g35 );
xnor U16443 ( n16566, n16563, n10326 );
nand U16444 ( n16563, n16567, n16568 );
nor U16445 ( n16568, n19375, n19823 );
nor U16446 ( n16567, n19824, n19825 );
nor U16447 ( n3353, n16569, n16570 );
nand U16448 ( n16570, n16571, n19376 );
nor U16449 ( n16571, n16572, n16573 );
nor U16450 ( n16573, n19824, g13895 );
nor U16451 ( n16572, n19823, g11349 );
nand U16452 ( n16569, n16574, n19377 );
nor U16453 ( n16574, n10948, g16603 );
nor U16454 ( n3348, n19468, n10991 );
nand U16455 ( n3343, n16575, n16576 );
or U16456 ( n16576, n16577, n19533 );
nor U16457 ( n16575, n16578, n16579 );
nor U16458 ( n16579, n10729, n16580 );
nand U16459 ( n16580, n16581, n19821 );
nor U16460 ( n16581, n11200, n10990 );
nor U16461 ( n16578, n19822, n16582 );
nor U16462 ( n16582, n16583, n10992 );
nor U16463 ( n16583, n19821, n11200 );
nand U16464 ( n3338, n16584, n16585 );
nand U16465 ( n16585, n16586, n10729 );
or U16466 ( n16584, n16586, n19821 );
nand U16467 ( n3333, n16587, n16588 );
nand U16468 ( n16588, n11017, n10779 );
nor U16469 ( n16587, n16589, n16590 );
and U16470 ( n16590, n19821, n16591 );
nor U16471 ( n16589, n19821, n16592 );
nand U16472 ( n3328, n16593, n16594 );
nand U16473 ( n16594, n16595, n10779 );
nor U16474 ( n16593, n16596, n16597 );
nor U16475 ( n16597, n10730, n16598 );
nand U16476 ( n16598, n19379, n16591 );
nor U16477 ( n16596, n19378, n16599 );
nor U16478 ( n16599, n16600, n10992 );
nor U16479 ( n16600, n19379, n16601 );
nand U16480 ( n3323, n16602, n16603 );
nand U16481 ( n16603, n16595, n10730 );
not U16482 ( n16595, n16592 );
nand U16483 ( n16602, n16592, n10567 );
nand U16484 ( n16592, g35, n16601 );
nand U16485 ( n3318, n16604, n16605 );
nand U16486 ( n16605, n16586, n10567 );
nor U16487 ( n16604, n16606, n16607 );
nor U16488 ( n16607, n19521, g35 );
nor U16489 ( n16606, n10948, n16608 );
or U16490 ( n16608, n10567, n11200 );
nand U16491 ( n3313, n16609, n16610 );
nand U16492 ( n16610, n16611, n16601 );
nor U16493 ( n16609, n16612, n16613 );
nor U16494 ( n16613, n10487, n16614 );
nand U16495 ( n16614, n16591, n10376 );
nor U16496 ( n16591, n16601, n10992 );
nor U16497 ( n16612, n19820, n16615 );
nor U16498 ( n16615, n16616, n10992 );
nor U16499 ( n16616, n16601, n10376 );
nand U16500 ( n3308, n16617, n16618 );
nand U16501 ( n16618, n11016, n10376 );
nand U16502 ( n16617, n16619, g35 );
nor U16503 ( n16619, n16620, n16621 );
nand U16504 ( n16621, n16622, n16623 );
nand U16505 ( n16623, n16624, n16601 );
nor U16506 ( n16624, n16625, n16626 );
nand U16507 ( n16626, n16627, n10487 );
or U16508 ( n16622, n16627, n16601 );
nand U16509 ( n16601, n16628, n16629 );
nor U16510 ( n16629, n19386, n19789 );
nor U16511 ( n16628, n11123, n16625 );
nor U16512 ( n16620, n16630, n10487 );
and U16513 ( n16630, n16627, n16631 );
nand U16514 ( n3303, n16632, n16633 );
nand U16515 ( n16633, n16586, n10376 );
nand U16516 ( n16632, n16577, n10849 );
nand U16517 ( n3298, n16634, n16635 );
nand U16518 ( n16635, n16636, n16586 );
not U16519 ( n16586, n16577 );
nor U16520 ( n16636, n19380, n15980 );
nand U16521 ( n16634, n10944, n16637 );
nand U16522 ( n16637, n10849, n11200 );
nand U16523 ( n3293, n16638, n16639 );
nand U16524 ( n16639, n16640, n10924 );
nor U16525 ( n16638, n16641, n16642 );
nor U16526 ( n16642, n10948, n16643 );
nand U16527 ( n16643, n16631, n16627 );
nand U16528 ( n16627, n16644, n16645 );
nand U16529 ( n16645, n19789, n16646 );
nand U16530 ( n16646, n16647, n16648 );
nor U16531 ( n16648, n16649, n16650 );
nand U16532 ( n16650, n16651, n16652 );
nand U16533 ( n16652, n16653, n16654 );
nor U16534 ( n16653, n19383, n19811 );
nand U16535 ( n16651, n16655, n16656 );
nor U16536 ( n16655, n19381, n19810 );
nor U16537 ( n16649, n16657, n16658 );
nor U16538 ( n16657, n16659, n16660 );
nor U16539 ( n16660, n19386, n19808 );
nor U16540 ( n16659, n19382, n19812 );
nor U16541 ( n16647, n16661, n16662 );
nand U16542 ( n16662, n16663, n16664 );
nand U16543 ( n16664, n19385, n16665 );
nand U16544 ( n16663, n16666, g12470 );
nand U16545 ( n16666, n16667, n16668 );
nand U16546 ( n16668, n16656, n10801 );
not U16547 ( n16667, n16669 );
nor U16548 ( n16661, n16670, n16671 );
nor U16549 ( n16670, n16672, n16673 );
nor U16550 ( n16673, n19387, n19809 );
nor U16551 ( n16672, n19384, n19813 );
nand U16552 ( n16644, n16674, n10327 );
nand U16553 ( n16674, n16675, n16676 );
nor U16554 ( n16676, n16677, n16678 );
nand U16555 ( n16678, n16679, n16680 );
nand U16556 ( n16680, n16681, n16682 );
nor U16557 ( n16681, n19381, n19800 );
nand U16558 ( n16679, n16683, n16684 );
nor U16559 ( n16683, n19383, n19801 );
nor U16560 ( n16677, n16685, n16686 );
nor U16561 ( n16685, n16687, n16688 );
nor U16562 ( n16688, n19387, n19799 );
nor U16563 ( n16687, n19384, n19803 );
nor U16564 ( n16675, n16689, n16690 );
nand U16565 ( n16690, n16691, n16692 );
nand U16566 ( n16692, n19385, n16669 );
nand U16567 ( n16669, n16693, n16694 );
nand U16568 ( n16694, n16695, n16684 );
nor U16569 ( n16695, n19788, n19817 );
nor U16570 ( n16693, n16696, n16697 );
nor U16571 ( n16697, n16686, n16698 );
nand U16572 ( n16698, n10850, g14828 );
nor U16573 ( n16696, n16658, n16699 );
or U16574 ( n16699, n19816, n19787 );
not U16575 ( n16658, n16682 );
nand U16576 ( n16691, n16700, g12470 );
nand U16577 ( n16700, n16701, n16702 );
nand U16578 ( n16702, n16682, n10802 );
not U16579 ( n16701, n16665 );
nand U16580 ( n16665, n16703, n16704 );
nand U16581 ( n16704, n16705, n16656 );
nor U16582 ( n16705, n19787, n19806 );
nor U16583 ( n16703, n16706, n16707 );
nor U16584 ( n16707, n16671, n16708 );
nand U16585 ( n16708, n10852, g14828 );
nor U16586 ( n16706, n16686, n16709 );
nand U16587 ( n16709, n10851, g17688 );
not U16588 ( n16686, n16654 );
nor U16589 ( n16689, n16710, n11123 );
not U16590 ( n11123, n16656 );
nor U16591 ( n16710, n16711, n16712 );
nor U16592 ( n16712, n19382, n19802 );
nor U16593 ( n16711, n19386, n19818 );
nor U16594 ( n16641, n19818, g35 );
nand U16595 ( n3288, n16713, n16714 );
nand U16596 ( n16714, n11016, n10763 );
nor U16597 ( n16713, n16715, n16716 );
nor U16598 ( n16716, n11200, n15730 );
nor U16599 ( n16715, n19818, n16577 );
nand U16600 ( n16577, g35, n11200 );
nand U16601 ( n11200, n16717, n10304 );
nand U16602 ( n3283, n16718, n16719 );
or U16603 ( n16719, n16720, n15730 );
nor U16604 ( n16718, n16721, n16722 );
nor U16605 ( n16722, n19816, g35 );
nor U16606 ( n16721, n10948, n16723 );
nand U16607 ( n16723, n16720, n10763 );
nand U16608 ( n16720, n16724, n16717 );
nand U16609 ( n3278, n16725, n16726 );
nand U16610 ( n16726, n16727, n10942 );
nor U16611 ( n16725, n16728, n16729 );
nor U16612 ( n16729, n19815, g35 );
nor U16613 ( n16728, n10949, n16730 );
or U16614 ( n16730, n16727, n19816 );
and U16615 ( n16727, n16731, n16717 );
nand U16616 ( n3273, n16732, n16733 );
or U16617 ( n16733, n16734, n15730 );
nor U16618 ( n16732, n16735, n16736 );
nor U16619 ( n16736, n19814, g35 );
nor U16620 ( n16735, n10949, n16737 );
nand U16621 ( n16737, n16734, n10850 );
nand U16622 ( n16734, n16738, n16717 );
nand U16623 ( n3268, n16739, n16740 );
or U16624 ( n16740, n16741, n15730 );
nor U16625 ( n16739, n16742, n16743 );
nor U16626 ( n16743, n19813, g35 );
nor U16627 ( n16742, n10949, n16744 );
nand U16628 ( n16744, n16741, n10801 );
nand U16629 ( n16741, n16745, n16717 );
nor U16630 ( n16717, n19798, n19797 );
nand U16631 ( n3263, n16746, n16747 );
nand U16632 ( n16747, n16748, n10944 );
nor U16633 ( n16746, n16749, n16750 );
nor U16634 ( n16750, n19812, g35 );
nor U16635 ( n16749, n10949, n16751 );
or U16636 ( n16751, n16748, n19813 );
and U16637 ( n16748, n16752, n10304 );
nand U16638 ( n3258, n16753, n16754 );
nand U16639 ( n16754, n16755, n10943 );
nor U16640 ( n16753, n16756, n16757 );
nor U16641 ( n16757, n19811, g35 );
nor U16642 ( n16756, n10949, n16758 );
or U16643 ( n16758, n16755, n19812 );
and U16644 ( n16755, n16752, n16724 );
nand U16645 ( n3253, n16759, n16760 );
nand U16646 ( n16760, n16761, n10942 );
nor U16647 ( n16759, n16762, n16763 );
nor U16648 ( n16763, n19810, g35 );
nor U16649 ( n16762, n10949, n16764 );
or U16650 ( n16764, n16761, n19811 );
and U16651 ( n16761, n16752, n16731 );
nand U16652 ( n3248, n16765, n16766 );
nand U16653 ( n16766, n16767, n10944 );
nor U16654 ( n16765, n16768, n16769 );
nor U16655 ( n16769, n19809, g35 );
nor U16656 ( n16768, n10949, n16770 );
or U16657 ( n16770, n16767, n19810 );
and U16658 ( n16767, n16752, n16738 );
nand U16659 ( n3243, n16771, n16772 );
nand U16660 ( n16772, n16773, n10943 );
nor U16661 ( n16771, n16774, n16775 );
nor U16662 ( n16775, n19808, g35 );
nor U16663 ( n16774, n10949, n16776 );
or U16664 ( n16776, n16773, n19809 );
and U16665 ( n16773, n16752, n16745 );
nand U16666 ( n3238, n16777, n16778 );
nand U16667 ( n16778, n16779, n10942 );
nor U16668 ( n16777, n16780, n16781 );
nor U16669 ( n16781, n19807, g35 );
nor U16670 ( n16780, n10949, n16782 );
or U16671 ( n16782, n16779, n19808 );
and U16672 ( n16779, n16783, n10304 );
nand U16673 ( n3233, n16784, n16785 );
or U16674 ( n16785, n16786, n15730 );
nor U16675 ( n16784, n16787, n16788 );
nor U16676 ( n16788, n19806, g35 );
nor U16677 ( n16787, n10949, n16789 );
nand U16678 ( n16789, n16786, n10851 );
nand U16679 ( n16786, n16783, n16724 );
nand U16680 ( n3228, n16790, n16791 );
nand U16681 ( n16791, n16792, n10944 );
nor U16682 ( n16790, n16793, n16794 );
nor U16683 ( n16794, n19805, g35 );
nor U16684 ( n16793, n10949, n16795 );
or U16685 ( n16795, n16792, n19806 );
and U16686 ( n16792, n16783, n16731 );
nand U16687 ( n3223, n16796, n16797 );
or U16688 ( n16797, n16798, n15730 );
nor U16689 ( n16796, n16799, n16800 );
nor U16690 ( n16800, n19804, g35 );
nor U16691 ( n16799, n10950, n16801 );
nand U16692 ( n16801, n16798, n10852 );
nand U16693 ( n16798, n16783, n16738 );
nand U16694 ( n3218, n16802, n16803 );
or U16695 ( n16803, n16804, n15730 );
nor U16696 ( n16802, n16805, n16806 );
nor U16697 ( n16806, n19803, g35 );
nor U16698 ( n16805, n10950, n16807 );
nand U16699 ( n16807, n16804, n10802 );
nand U16700 ( n16804, n16783, n16745 );
nand U16701 ( n3213, n16808, n16809 );
nand U16702 ( n16809, n16810, n10943 );
nor U16703 ( n16808, n16811, n16812 );
nor U16704 ( n16812, n19802, g35 );
nor U16705 ( n16811, n10950, n16813 );
or U16706 ( n16813, n16810, n19803 );
and U16707 ( n16810, n16814, n10304 );
nand U16708 ( n3208, n16815, n16816 );
nand U16709 ( n16816, n16817, n10942 );
nor U16710 ( n16815, n16818, n16819 );
nor U16711 ( n16819, n19801, g35 );
nor U16712 ( n16818, n10950, n16820 );
or U16713 ( n16820, n16817, n19802 );
and U16714 ( n16817, n16814, n16724 );
nand U16715 ( n3203, n16821, n16822 );
nand U16716 ( n16822, n16823, n10944 );
nor U16717 ( n16821, n16824, n16825 );
nor U16718 ( n16825, n19800, g35 );
nor U16719 ( n16824, n10950, n16826 );
or U16720 ( n16826, n16823, n19801 );
and U16721 ( n16823, n16814, n16731 );
nand U16722 ( n3198, n16827, n16828 );
nand U16723 ( n16828, n16829, n10943 );
nor U16724 ( n16827, n16830, n16831 );
nor U16725 ( n16831, n19799, g35 );
nor U16726 ( n16830, n10950, n16832 );
or U16727 ( n16832, n16829, n19800 );
and U16728 ( n16829, n16814, n16738 );
nand U16729 ( n3193, n16833, n16834 );
nand U16730 ( n16834, n16835, n10942 );
nor U16731 ( n16833, n16836, n16837 );
nor U16732 ( n16837, n19798, g35 );
nor U16733 ( n16836, n10950, n16838 );
or U16734 ( n16838, n16835, n19799 );
and U16735 ( n16835, n16814, n16745 );
and U16736 ( n16745, n16839, n19796 );
nor U16737 ( n16839, n10246, n10466 );
nor U16738 ( n16814, n10267, n10434 );
nand U16739 ( n3188, n16840, n16841 );
nand U16740 ( n16841, n11016, n10434 );
nand U16741 ( n16840, n16842, g35 );
nor U16742 ( n16842, n16843, n16844 );
nor U16743 ( n16844, n16752, n16845 );
nand U16744 ( n16845, n16846, n16847 );
nand U16745 ( n16847, n19796, n10267 );
nand U16746 ( n16846, n16783, n10304 );
nor U16747 ( n16783, n10267, n19797 );
nor U16748 ( n16752, n10434, n19798 );
nand U16749 ( n3183, n16848, n16849 );
nand U16750 ( n16849, n16850, n10304 );
nand U16751 ( n16850, g35, n16851 );
nand U16752 ( n16851, n19797, n16852 );
or U16753 ( n16848, n16853, n19797 );
nand U16754 ( n3178, n16854, n16855 );
nand U16755 ( n16855, n16856, n19796 );
and U16756 ( n16856, n16852, n16724 );
nor U16757 ( n16724, n19795, n19794 );
nand U16758 ( n16854, n11016, n10466 );
nand U16759 ( n3173, n16857, n16858 );
nand U16760 ( n16858, n16859, n16852 );
nand U16761 ( n16859, n16860, n16861 );
nand U16762 ( n16861, n16731, g35 );
nor U16763 ( n16731, n10246, n19795 );
not U16764 ( n16860, n16738 );
nor U16765 ( n16738, n10466, n19794 );
nand U16766 ( n16857, n11016, n10246 );
nor U16767 ( n3168, n10246, n16853 );
nand U16768 ( n16853, n16862, n19796 );
nor U16769 ( n16862, n16843, n10992 );
not U16770 ( n16843, n16852 );
nand U16771 ( n16852, n15879, n15513 );
and U16772 ( n15879, n16863, n16864 );
nor U16773 ( n16864, n19425, n19939 );
nand U16774 ( n3074, n16865, n16866 );
nand U16775 ( n16866, g35, n10327 );
nand U16776 ( n16865, n11016, n10881 );
nand U16777 ( n3069, n16867, n16868 );
nand U16778 ( n16868, n11016, n10882 );
nand U16779 ( n16867, n16869, g35 );
nor U16780 ( n16869, n16870, g9817 );
nor U16781 ( n16870, n16871, n10881 );
nor U16782 ( n16871, n19793, n10882 );
nor U16783 ( n3060, n19798, n10991 );
nand U16784 ( n3055, n16872, n16873 );
nand U16785 ( n16873, n16874, n16682 );
nor U16786 ( n16872, n16875, n16876 );
nor U16787 ( n16876, n16877, n10992 );
nor U16788 ( n16877, n16878, n16879 );
nor U16789 ( n16879, n16880, n16671 );
nor U16790 ( n16878, n19452, n16631 );
nor U16791 ( n16875, n19792, g35 );
nand U16792 ( n3050, n16881, n16882 );
nand U16793 ( n16882, n16640, n10265 );
nor U16794 ( n16881, n16883, n16884 );
nor U16795 ( n16884, n19791, g35 );
nor U16796 ( n16883, n10951, n16885 );
nand U16797 ( n16885, n16874, n19792 );
nor U16798 ( n16874, n16880, n16625 );
nor U16799 ( n16880, n16557, n11109 );
nand U16800 ( n11109, n19588, n11120 );
not U16801 ( n11120, n11174 );
nor U16802 ( n3045, n19790, n16886 );
and U16803 ( n16886, g35, n16887 );
nand U16804 ( n3040, n16888, n16889 );
nand U16805 ( n16889, n11016, n10327 );
nand U16806 ( n16888, n16890, g35 );
nor U16807 ( n16890, n16887, n10694 );
nor U16808 ( n16887, n16891, n19789 );
nand U16809 ( n3035, n16892, n16893 );
or U16810 ( n16893, g35, n19384 );
nand U16811 ( n16892, n16894, g35 );
xnor U16812 ( n16894, n16891, n10327 );
nand U16813 ( n16891, n16895, n16896 );
nor U16814 ( n16896, n19385, n19786 );
nor U16815 ( n16895, n19787, n19788 );
nor U16816 ( n2994, n16897, n16898 );
nand U16817 ( n16898, n16899, n19386 );
nor U16818 ( n16899, n16900, n16901 );
nor U16819 ( n16901, n19787, g14828 );
nor U16820 ( n16900, n19786, g12470 );
nand U16821 ( n16897, n16902, n19387 );
nor U16822 ( n16902, n10951, g17688 );
nor U16823 ( n2989, n19491, n10993 );
nand U16824 ( n2984, n16903, n16904 );
nand U16825 ( n16904, n16905, n10896 );
nor U16826 ( n16903, n16906, n16907 );
nor U16827 ( n16907, n10731, n16908 );
nand U16828 ( n16908, n16909, n19784 );
nor U16829 ( n16909, n10951, n11211 );
nor U16830 ( n16906, n19785, n16910 );
nor U16831 ( n16910, n16911, n10991 );
nor U16832 ( n16911, n19784, n11211 );
nand U16833 ( n2979, n16912, n16913 );
nand U16834 ( n16913, n16905, n10731 );
or U16835 ( n16912, n16905, n19784 );
nand U16836 ( n2974, n16914, n16915 );
nand U16837 ( n16915, n11015, n10279 );
nor U16838 ( n16914, n16916, n16917 );
and U16839 ( n16917, n19784, n16918 );
nor U16840 ( n16916, n19784, n16919 );
nand U16841 ( n2969, n16920, n16921 );
nand U16842 ( n16921, n16922, n10279 );
nor U16843 ( n16920, n16923, n16924 );
nor U16844 ( n16924, n10732, n16925 );
nand U16845 ( n16925, n19389, n16918 );
nor U16846 ( n16923, n19388, n16926 );
nor U16847 ( n16926, n16927, n10993 );
nor U16848 ( n16927, n19389, n16928 );
nand U16849 ( n2964, n16929, n16930 );
nand U16850 ( n16930, n16922, n10732 );
not U16851 ( n16922, n16919 );
nand U16852 ( n16929, n16919, n10568 );
nand U16853 ( n16919, g35, n16928 );
nand U16854 ( n2959, n16931, n16932 );
nand U16855 ( n16932, n16905, n10568 );
nor U16856 ( n16931, n16933, n16934 );
nor U16857 ( n16934, n19522, g35 );
nor U16858 ( n16933, n10951, n16935 );
or U16859 ( n16935, n10568, n11211 );
nand U16860 ( n2954, n16936, n16937 );
nand U16861 ( n16937, n16938, n16928 );
nor U16862 ( n16936, n16939, n16940 );
nor U16863 ( n16940, n10488, n16941 );
nand U16864 ( n16941, n16918, n10377 );
nor U16865 ( n16918, n16928, n10990 );
nor U16866 ( n16939, n19783, n16942 );
nor U16867 ( n16942, n16943, n10993 );
nor U16868 ( n16943, n16928, n10377 );
nand U16869 ( n2949, n16944, n16945 );
nand U16870 ( n16945, n11015, n10377 );
nand U16871 ( n16944, n16946, g35 );
nor U16872 ( n16946, n16947, n16948 );
nand U16873 ( n16948, n16949, n16950 );
nand U16874 ( n16950, n16951, n16928 );
nor U16875 ( n16951, n16952, n16953 );
nand U16876 ( n16953, n16954, n10488 );
or U16877 ( n16949, n16954, n16928 );
nand U16878 ( n16928, n16955, n16956 );
nor U16879 ( n16956, n19396, n19753 );
nor U16880 ( n16955, n11104, n16952 );
nor U16881 ( n16947, n16957, n10488 );
and U16882 ( n16957, n16954, n16958 );
nand U16883 ( n2944, n16959, n16960 );
nand U16884 ( n16960, n16905, n10377 );
nand U16885 ( n16959, n16961, n10853 );
nand U16886 ( n2939, n16962, n16963 );
nand U16887 ( n16963, n16964, n16905 );
not U16888 ( n16905, n16961 );
nor U16889 ( n16964, n19390, n15980 );
nand U16890 ( n16962, n10943, n16965 );
nand U16891 ( n16965, n10853, n11211 );
nand U16892 ( n2934, n16966, n16967 );
nand U16893 ( n16967, n16968, n10929 );
nor U16894 ( n16966, n16969, n16970 );
nor U16895 ( n16970, n10952, n16971 );
nand U16896 ( n16971, n16958, n16954 );
nand U16897 ( n16954, n16972, n16973 );
nand U16898 ( n16973, n19753, n16974 );
nand U16899 ( n16974, n16975, n16976 );
nor U16900 ( n16976, n16977, n16978 );
nand U16901 ( n16978, n16979, n16980 );
nand U16902 ( n16980, n16981, n16982 );
nor U16903 ( n16981, n19393, n19775 );
nand U16904 ( n16979, n16983, n16984 );
nor U16905 ( n16983, n19391, n19774 );
nor U16906 ( n16977, n16985, n16986 );
nor U16907 ( n16985, n16987, n16988 );
nor U16908 ( n16988, n19396, n19772 );
nor U16909 ( n16987, n19392, n19776 );
nor U16910 ( n16975, n16989, n16990 );
nand U16911 ( n16990, n16991, n16992 );
nand U16912 ( n16992, n19395, n16993 );
nand U16913 ( n16991, n16994, g12422 );
nand U16914 ( n16994, n16995, n16996 );
nand U16915 ( n16996, n16984, n10803 );
not U16916 ( n16995, n16997 );
nor U16917 ( n16989, n16998, n16999 );
nor U16918 ( n16998, n17000, n17001 );
nor U16919 ( n17001, n19397, n19773 );
nor U16920 ( n17000, n19394, n19777 );
nand U16921 ( n16972, n17002, n10328 );
nand U16922 ( n17002, n17003, n17004 );
nor U16923 ( n17004, n17005, n17006 );
nand U16924 ( n17006, n17007, n17008 );
nand U16925 ( n17008, n17009, n17010 );
nor U16926 ( n17009, n19391, n19764 );
nand U16927 ( n17007, n17011, n17012 );
nor U16928 ( n17011, n19393, n19765 );
nor U16929 ( n17005, n17013, n17014 );
nor U16930 ( n17013, n17015, n17016 );
nor U16931 ( n17016, n19397, n19763 );
nor U16932 ( n17015, n19394, n19767 );
nor U16933 ( n17003, n17017, n17018 );
nand U16934 ( n17018, n17019, n17020 );
nand U16935 ( n17020, n19395, n16997 );
nand U16936 ( n16997, n17021, n17022 );
nand U16937 ( n17022, n17023, n17012 );
nor U16938 ( n17023, n19752, n19781 );
nor U16939 ( n17021, n17024, n17025 );
nor U16940 ( n17025, n17014, n17026 );
nand U16941 ( n17026, n10854, g14779 );
nor U16942 ( n17024, n16986, n17027 );
or U16943 ( n17027, n19780, n19751 );
not U16944 ( n16986, n17010 );
nand U16945 ( n17019, n17028, g12422 );
nand U16946 ( n17028, n17029, n17030 );
nand U16947 ( n17030, n17010, n10804 );
not U16948 ( n17029, n16993 );
nand U16949 ( n16993, n17031, n17032 );
nand U16950 ( n17032, n17033, n16984 );
nor U16951 ( n17033, n19751, n19770 );
nor U16952 ( n17031, n17034, n17035 );
nor U16953 ( n17035, n16999, n17036 );
nand U16954 ( n17036, n10856, g14779 );
nor U16955 ( n17034, n17014, n17037 );
nand U16956 ( n17037, n10855, g17649 );
not U16957 ( n17014, n16982 );
nor U16958 ( n17017, n17038, n11104 );
not U16959 ( n11104, n16984 );
nor U16960 ( n17038, n17039, n17040 );
nor U16961 ( n17040, n19392, n19766 );
nor U16962 ( n17039, n19396, n19782 );
nor U16963 ( n16969, n19782, g35 );
nand U16964 ( n2929, n17041, n17042 );
nand U16965 ( n17042, n11019, n10764 );
nor U16966 ( n17041, n17043, n17044 );
nor U16967 ( n17044, n15730, n11211 );
nor U16968 ( n17043, n19782, n16961 );
nand U16969 ( n16961, g35, n11211 );
nand U16970 ( n11211, n17045, n10398 );
nand U16971 ( n2924, n17046, n17047 );
or U16972 ( n17047, n17048, n15730 );
nor U16973 ( n17046, n17049, n17050 );
nor U16974 ( n17050, n19780, g35 );
nor U16975 ( n17049, n10952, n17051 );
nand U16976 ( n17051, n17048, n10764 );
nand U16977 ( n17048, n17052, n17045 );
nand U16978 ( n2919, n17053, n17054 );
nand U16979 ( n17054, n17055, n10944 );
nor U16980 ( n17053, n17056, n17057 );
nor U16981 ( n17057, n19779, g35 );
nor U16982 ( n17056, n10952, n17058 );
or U16983 ( n17058, n17055, n19780 );
and U16984 ( n17055, n17059, n17045 );
nand U16985 ( n2914, n17060, n17061 );
or U16986 ( n17061, n17062, n15730 );
nor U16987 ( n17060, n17063, n17064 );
nor U16988 ( n17064, n19778, g35 );
nor U16989 ( n17063, n10952, n17065 );
nand U16990 ( n17065, n17062, n10854 );
nand U16991 ( n17062, n17066, n17045 );
nand U16992 ( n2909, n17067, n17068 );
or U16993 ( n17068, n17069, n15730 );
nor U16994 ( n17067, n17070, n17071 );
nor U16995 ( n17071, n19777, g35 );
nor U16996 ( n17070, n10952, n17072 );
nand U16997 ( n17072, n17069, n10803 );
nand U16998 ( n17069, n17073, n17045 );
nor U16999 ( n17045, n19762, n19761 );
nand U17000 ( n2904, n17074, n17075 );
nand U17001 ( n17075, n17076, n10943 );
nor U17002 ( n17074, n17077, n17078 );
nor U17003 ( n17078, n19776, g35 );
nor U17004 ( n17077, n10952, n17079 );
or U17005 ( n17079, n17076, n19777 );
nor U17006 ( n17076, n17080, n19760 );
nand U17007 ( n2899, n17081, n17082 );
nand U17008 ( n17082, n17083, n10942 );
nor U17009 ( n17081, n17084, n17085 );
nor U17010 ( n17085, n19775, g35 );
nor U17011 ( n17084, n10952, n17086 );
or U17012 ( n17086, n17083, n19776 );
nor U17013 ( n17083, n17080, n17087 );
nand U17014 ( n2894, n17088, n17089 );
nand U17015 ( n17089, n17090, n10944 );
nor U17016 ( n17088, n17091, n17092 );
nor U17017 ( n17092, n19774, g35 );
nor U17018 ( n17091, n10952, n17093 );
or U17019 ( n17093, n17090, n19775 );
and U17020 ( n17090, n17094, n17059 );
nand U17021 ( n2889, n17095, n17096 );
nand U17022 ( n17096, n17097, n10943 );
nor U17023 ( n17095, n17098, n17099 );
nor U17024 ( n17099, n19773, g35 );
nor U17025 ( n17098, n10972, n17100 );
or U17026 ( n17100, n17097, n19774 );
nor U17027 ( n17097, n17080, n17101 );
nand U17028 ( n2884, n17102, n17103 );
nand U17029 ( n17103, n17104, n10942 );
nor U17030 ( n17102, n17105, n17106 );
nor U17031 ( n17106, n19772, g35 );
nor U17032 ( n17105, n10952, n17107 );
or U17033 ( n17107, n17104, n19773 );
and U17034 ( n17104, n17094, n17073 );
nand U17035 ( n2879, n17108, n17109 );
nand U17036 ( n17109, n17110, n10944 );
nor U17037 ( n17108, n17111, n17112 );
nor U17038 ( n17112, n19771, g35 );
nor U17039 ( n17111, n10952, n17113 );
or U17040 ( n17113, n17110, n19772 );
nand U17041 ( n2874, n17114, n17115 );
or U17042 ( n17115, n17116, n15730 );
nor U17043 ( n17114, n17117, n17118 );
nor U17044 ( n17118, n19770, g35 );
nor U17045 ( n17117, n10953, n17119 );
nand U17046 ( n17119, n17116, n10855 );
nand U17047 ( n17116, n17120, n17052 );
nand U17048 ( n2869, n17121, n17122 );
nand U17049 ( n17122, n17123, n10943 );
nor U17050 ( n17121, n17124, n17125 );
nor U17051 ( n17125, n19769, g35 );
nor U17052 ( n17124, n10953, n17126 );
or U17053 ( n17126, n17123, n19770 );
and U17054 ( n17123, n17120, n17059 );
nand U17055 ( n2864, n17127, n17128 );
or U17056 ( n17128, n17129, n15730 );
nor U17057 ( n17127, n17130, n17131 );
nor U17058 ( n17131, n19768, g35 );
nor U17059 ( n17130, n10953, n17132 );
nand U17060 ( n17132, n17129, n10856 );
nand U17061 ( n17129, n17120, n17066 );
nand U17062 ( n2859, n17133, n17134 );
or U17063 ( n17134, n17135, n15730 );
nor U17064 ( n17133, n17136, n17137 );
nor U17065 ( n17137, n19767, g35 );
nor U17066 ( n17136, n10953, n17138 );
nand U17067 ( n17138, n17135, n10804 );
nand U17068 ( n17135, n17120, n17073 );
nand U17069 ( n2854, n17139, n17140 );
nand U17070 ( n17140, n17141, n10942 );
nor U17071 ( n17139, n17142, n17143 );
nor U17072 ( n17143, n19766, g35 );
nor U17073 ( n17142, n10953, n17144 );
or U17074 ( n17144, n17141, n19767 );
and U17075 ( n17141, n17145, n10398 );
nand U17076 ( n2849, n17146, n17147 );
nand U17077 ( n17147, n17148, n10944 );
nor U17078 ( n17146, n17149, n17150 );
nor U17079 ( n17150, n19765, g35 );
nor U17080 ( n17149, n10953, n17151 );
or U17081 ( n17151, n17148, n19766 );
and U17082 ( n17148, n17145, n17052 );
nand U17083 ( n2844, n17152, n17153 );
nand U17084 ( n17153, n17154, n10943 );
nor U17085 ( n17152, n17155, n17156 );
nor U17086 ( n17156, n19764, g35 );
nor U17087 ( n17155, n10953, n17157 );
or U17088 ( n17157, n17154, n19765 );
and U17089 ( n17154, n17145, n17059 );
nand U17090 ( n2839, n17158, n17159 );
nand U17091 ( n17159, n17160, n10942 );
nor U17092 ( n17158, n17161, n17162 );
nor U17093 ( n17162, n19763, g35 );
nor U17094 ( n17161, n10953, n17163 );
or U17095 ( n17163, n17160, n19764 );
and U17096 ( n17160, n17145, n17066 );
nand U17097 ( n2834, n17164, n17165 );
nand U17098 ( n17165, n17166, n10944 );
nor U17099 ( n17164, n17167, n17168 );
nor U17100 ( n17168, n19762, g35 );
nor U17101 ( n17167, n10953, n17169 );
or U17102 ( n17169, n17166, n19763 );
and U17103 ( n17166, n17145, n17073 );
and U17104 ( n17073, n17170, n19760 );
nor U17105 ( n17170, n10247, n10467 );
nor U17106 ( n17145, n10597, n10274 );
nand U17107 ( n2829, n17171, n17172 );
nand U17108 ( n17172, n17173, n17174 );
nand U17109 ( n17173, n17175, n17176 );
nand U17110 ( n17176, n2701, n19760 );
nor U17111 ( n17175, n17110, n17177 );
nor U17112 ( n17177, n10953, n17080 );
not U17113 ( n17080, n17094 );
nor U17114 ( n17094, n10274, n19762 );
and U17115 ( n17110, n17120, n10398 );
nor U17116 ( n17120, n10597, n19761 );
nand U17117 ( n17171, n10997, n10274 );
nand U17118 ( n2824, n17178, n17179 );
nand U17119 ( n17179, n17180, n10398 );
nand U17120 ( n17180, g35, n17181 );
nand U17121 ( n17181, n19761, n17174 );
or U17122 ( n17178, n17182, n19761 );
nand U17123 ( n2819, n17183, n17184 );
nand U17124 ( n17184, n17185, n19760 );
nor U17125 ( n17185, n17186, n17087 );
not U17126 ( n17087, n17052 );
nor U17127 ( n17052, n19759, n19758 );
nand U17128 ( n17183, n10997, n10467 );
nand U17129 ( n2814, n17187, n17188 );
nand U17130 ( n17188, n17189, n17174 );
nand U17131 ( n17189, n17101, n17190 );
nand U17132 ( n17190, n17059, g35 );
nor U17133 ( n17059, n10247, n19759 );
not U17134 ( n17101, n17066 );
nor U17135 ( n17066, n10467, n19758 );
nand U17136 ( n17187, n10996, n10247 );
nor U17137 ( n2809, n10247, n17182 );
nand U17138 ( n17182, n17191, n19760 );
nor U17139 ( n17191, n17186, n10992 );
not U17140 ( n17186, n17174 );
nand U17141 ( n17174, n15878, n17192 );
nor U17142 ( n15878, n19937, n19938 );
nand U17143 ( n2715, n17193, n17194 );
nand U17144 ( n17194, g35, n10328 );
nand U17145 ( n17193, n10996, n10883 );
nand U17146 ( n2710, n17195, n17196 );
nand U17147 ( n17196, n10995, n10884 );
nand U17148 ( n17195, n17197, g35 );
nor U17149 ( n17197, n17198, g9741 );
nor U17150 ( n17198, n17199, n10883 );
nor U17151 ( n17199, n19757, n10884 );
nor U17152 ( n2701, n10954, n19762 );
nand U17153 ( n2696, n17200, n17201 );
nand U17154 ( n17201, n17202, n17010 );
nor U17155 ( n17200, n17203, n17204 );
nor U17156 ( n17204, n17205, n10991 );
nor U17157 ( n17205, n17206, n17207 );
nor U17158 ( n17207, n17208, n16999 );
nor U17159 ( n17206, n19436, n16958 );
nor U17160 ( n17203, n19756, g35 );
nand U17161 ( n2691, n17209, n17210 );
nand U17162 ( n17210, n16968, n10261 );
nor U17163 ( n17209, n17211, n17212 );
nor U17164 ( n17212, n19755, g35 );
nor U17165 ( n17211, n10978, n17213 );
nand U17166 ( n17213, n17202, n19756 );
nor U17167 ( n17202, n17208, n16952 );
and U17168 ( n17208, n15901, n17214 );
nor U17169 ( n15901, n16230, n19588 );
nor U17170 ( n2686, n19754, n17215 );
and U17171 ( n17215, g35, n17216 );
nand U17172 ( n2681, n17217, n17218 );
nand U17173 ( n17218, n10996, n10328 );
nand U17174 ( n17217, n17219, g35 );
nor U17175 ( n17219, n17216, n10689 );
nor U17176 ( n17216, n17220, n19753 );
nand U17177 ( n2676, n17221, n17222 );
or U17178 ( n17222, g35, n19394 );
nand U17179 ( n17221, n17223, g35 );
xnor U17180 ( n17223, n17220, n10328 );
nand U17181 ( n17220, n17224, n17225 );
nor U17182 ( n17225, n19395, n19750 );
nor U17183 ( n17224, n19751, n19752 );
nor U17184 ( n2635, n17226, n17227 );
nand U17185 ( n17227, n17228, n19396 );
nor U17186 ( n17228, n17229, n17230 );
nor U17187 ( n17230, n19751, g14779 );
nor U17188 ( n17229, n19750, g12422 );
nand U17189 ( n17226, n17231, n19397 );
nor U17190 ( n17231, n10978, g17649 );
nor U17191 ( n2630, n19485, n10992 );
nand U17192 ( n2625, n17232, n17233 );
nand U17193 ( n17233, n17234, n10759 );
nor U17194 ( n17232, n17235, n17236 );
nor U17195 ( n17236, n10733, n17237 );
nand U17196 ( n17237, n17238, n19748 );
nor U17197 ( n17238, n10978, n11216 );
nor U17198 ( n17235, n19749, n17239 );
nor U17199 ( n17239, n17240, n10992 );
nor U17200 ( n17240, n19748, n11216 );
nand U17201 ( n2620, n17241, n17242 );
nand U17202 ( n17242, n17234, n10733 );
or U17203 ( n17241, n17234, n19748 );
nand U17204 ( n2615, n17243, n17244 );
nand U17205 ( n17244, n10996, n10282 );
nor U17206 ( n17243, n17245, n17246 );
and U17207 ( n17246, n19748, n17247 );
nor U17208 ( n17245, n19748, n17248 );
nand U17209 ( n2610, n17249, n17250 );
nand U17210 ( n17250, n17251, n10282 );
nor U17211 ( n17249, n17252, n17253 );
nor U17212 ( n17253, n10734, n17254 );
nand U17213 ( n17254, n19399, n17247 );
nor U17214 ( n17252, n19398, n17255 );
nor U17215 ( n17255, n17256, n10992 );
nor U17216 ( n17256, n19399, n17257 );
nand U17217 ( n2605, n17258, n17259 );
nand U17218 ( n17259, n17251, n10734 );
not U17219 ( n17251, n17248 );
nand U17220 ( n17258, n17248, n10569 );
nand U17221 ( n2600, n17260, n17261 );
nand U17222 ( n17261, n17234, n10569 );
nor U17223 ( n17260, n17262, n17263 );
nor U17224 ( n17263, n19516, g35 );
nor U17225 ( n17262, n10975, n17264 );
or U17226 ( n17264, n10569, n11216 );
nand U17227 ( n2595, n17265, n17266 );
or U17228 ( n17266, n17248, n19516 );
nand U17229 ( n17248, g35, n17257 );
nor U17230 ( n17265, n17267, n17268 );
nor U17231 ( n17268, n10489, n17269 );
nand U17232 ( n17269, n17247, n10378 );
nor U17233 ( n17247, n17257, n10992 );
nor U17234 ( n17267, n19747, n17270 );
nor U17235 ( n17270, n17271, n10991 );
nor U17236 ( n17271, n17257, n10378 );
nand U17237 ( n2590, n17272, n17273 );
nand U17238 ( n17273, n10994, n10378 );
nand U17239 ( n17272, n17274, g35 );
nor U17240 ( n17274, n17275, n17276 );
nand U17241 ( n17276, n17277, n17278 );
nand U17242 ( n17278, n17279, n17257 );
nor U17243 ( n17279, n17280, n17281 );
nand U17244 ( n17281, n17282, n10489 );
or U17245 ( n17277, n17282, n17257 );
nand U17246 ( n17257, n17283, n17284 );
nor U17247 ( n17284, n19406, n19716 );
nor U17248 ( n17283, n11112, n17280 );
nor U17249 ( n17275, n17285, n10489 );
and U17250 ( n17285, n17282, n17286 );
nand U17251 ( n2585, n17287, n17288 );
nand U17252 ( n17288, n17234, n10378 );
nand U17253 ( n17287, n17289, n10857 );
nand U17254 ( n2580, n17290, n17291 );
nand U17255 ( n17291, n17292, n17234 );
not U17256 ( n17234, n17289 );
nor U17257 ( n17292, n19400, n15980 );
nand U17258 ( n17290, n10942, n17293 );
nand U17259 ( n17293, n10857, n11216 );
nand U17260 ( n2575, n17294, n17295 );
nand U17261 ( n17295, n17296, n10925 );
nor U17262 ( n17294, n17297, n17298 );
nor U17263 ( n17298, n10974, n17299 );
nand U17264 ( n17299, n17286, n17282 );
nand U17265 ( n17282, n17300, n17301 );
nand U17266 ( n17301, n19716, n17302 );
nand U17267 ( n17302, n17303, n17304 );
nor U17268 ( n17304, n17305, n17306 );
nand U17269 ( n17306, n17307, n17308 );
nand U17270 ( n17308, n17309, n17310 );
nor U17271 ( n17309, n19403, n19738 );
nand U17272 ( n17307, n17311, n17312 );
nor U17273 ( n17311, n19401, n19737 );
nor U17274 ( n17305, n17313, n17314 );
nor U17275 ( n17313, n17315, n17316 );
nor U17276 ( n17316, n19406, n19735 );
nor U17277 ( n17315, n19402, n19739 );
nor U17278 ( n17303, n17317, n17318 );
nand U17279 ( n17318, n17319, n17320 );
nand U17280 ( n17320, n19405, n17321 );
nand U17281 ( n17319, n17322, g12350 );
nand U17282 ( n17322, n17323, n17324 );
nand U17283 ( n17324, n17312, n10805 );
not U17284 ( n17323, n17325 );
nor U17285 ( n17317, n17326, n17327 );
nor U17286 ( n17326, n17328, n17329 );
nor U17287 ( n17329, n19407, n19736 );
nor U17288 ( n17328, n19404, n19740 );
nand U17289 ( n17300, n17330, n10329 );
nand U17290 ( n17330, n17331, n17332 );
nor U17291 ( n17332, n17333, n17334 );
nand U17292 ( n17334, n17335, n17336 );
nand U17293 ( n17336, n17337, n17338 );
nor U17294 ( n17337, n19401, n19727 );
nand U17295 ( n17335, n17339, n17340 );
nor U17296 ( n17339, n19403, n19728 );
nor U17297 ( n17333, n17341, n17342 );
nor U17298 ( n17341, n17343, n17344 );
nor U17299 ( n17344, n19407, n19726 );
nor U17300 ( n17343, n19404, n19730 );
nor U17301 ( n17331, n17345, n17346 );
nand U17302 ( n17346, n17347, n17348 );
nand U17303 ( n17348, n19405, n17325 );
nand U17304 ( n17325, n17349, n17350 );
nand U17305 ( n17350, n17351, n17340 );
nor U17306 ( n17351, n19715, n19744 );
nor U17307 ( n17349, n17352, n17353 );
nor U17308 ( n17353, n17342, n17354 );
nand U17309 ( n17354, n10858, g14738 );
nor U17310 ( n17352, n17314, n17355 );
or U17311 ( n17355, n19743, n19714 );
not U17312 ( n17314, n17338 );
nand U17313 ( n17347, n17356, g12350 );
nand U17314 ( n17356, n17357, n17358 );
nand U17315 ( n17358, n17338, n10806 );
not U17316 ( n17357, n17321 );
nand U17317 ( n17321, n17359, n17360 );
nand U17318 ( n17360, n17361, n17312 );
nor U17319 ( n17361, n19714, n19733 );
nor U17320 ( n17359, n17362, n17363 );
nor U17321 ( n17363, n17327, n17364 );
nand U17322 ( n17364, n10860, g14738 );
nor U17323 ( n17362, n17342, n17365 );
nand U17324 ( n17365, n10859, g17607 );
not U17325 ( n17342, n17310 );
nor U17326 ( n17345, n17366, n11112 );
not U17327 ( n11112, n17312 );
nor U17328 ( n17366, n17367, n17368 );
nor U17329 ( n17368, n19402, n19729 );
nor U17330 ( n17367, n19406, n19745 );
nor U17331 ( n17297, n19745, g35 );
nand U17332 ( n2570, n17369, n17370 );
nand U17333 ( n17370, n10994, n10765 );
nor U17334 ( n17369, n17371, n17372 );
nor U17335 ( n17372, n15730, n11216 );
nor U17336 ( n17371, n19745, n17289 );
nand U17337 ( n17289, g35, n11216 );
nand U17338 ( n11216, n17373, n10399 );
nand U17339 ( n2565, n17374, n17375 );
or U17340 ( n17375, n17376, n15730 );
nor U17341 ( n17374, n17377, n17378 );
nor U17342 ( n17378, n19743, g35 );
nor U17343 ( n17377, n10973, n17379 );
nand U17344 ( n17379, n17376, n10765 );
nand U17345 ( n17376, n17380, n17373 );
nand U17346 ( n2560, n17381, n17382 );
nand U17347 ( n17382, n17383, n10943 );
nor U17348 ( n17381, n17384, n17385 );
nor U17349 ( n17385, n19742, g35 );
nor U17350 ( n17384, n10973, n17386 );
or U17351 ( n17386, n17383, n19743 );
and U17352 ( n17383, n17387, n17373 );
nand U17353 ( n2555, n17388, n17389 );
or U17354 ( n17389, n17390, n15730 );
nor U17355 ( n17388, n17391, n17392 );
nor U17356 ( n17392, n19741, g35 );
nor U17357 ( n17391, n10973, n17393 );
nand U17358 ( n17393, n17390, n10858 );
nand U17359 ( n17390, n17394, n17373 );
nand U17360 ( n2550, n17395, n17396 );
or U17361 ( n17396, n17397, n15730 );
nor U17362 ( n17395, n17398, n17399 );
nor U17363 ( n17399, n19740, g35 );
nor U17364 ( n17398, n10973, n17400 );
nand U17365 ( n17400, n17397, n10805 );
nand U17366 ( n17397, n17401, n17373 );
nor U17367 ( n17373, n19725, n19724 );
nand U17368 ( n2545, n17402, n17403 );
nand U17369 ( n17403, n17404, n10942 );
nor U17370 ( n17402, n17405, n17406 );
nor U17371 ( n17406, n19739, g35 );
nor U17372 ( n17405, n10972, n17407 );
or U17373 ( n17407, n17404, n19740 );
nor U17374 ( n17404, n17408, n19723 );
nand U17375 ( n2540, n17409, n17410 );
nand U17376 ( n17410, n17411, n10944 );
nor U17377 ( n17409, n17412, n17413 );
nor U17378 ( n17413, n19738, g35 );
nor U17379 ( n17412, n10972, n17414 );
or U17380 ( n17414, n17411, n19739 );
nor U17381 ( n17411, n17408, n17415 );
nand U17382 ( n2535, n17416, n17417 );
nand U17383 ( n17417, n17418, n10943 );
nor U17384 ( n17416, n17419, n17420 );
nor U17385 ( n17420, n19737, g35 );
nor U17386 ( n17419, n10972, n17421 );
or U17387 ( n17421, n17418, n19738 );
and U17388 ( n17418, n17422, n17387 );
nand U17389 ( n2530, n17423, n17424 );
nand U17390 ( n17424, n17425, n10942 );
nor U17391 ( n17423, n17426, n17427 );
nor U17392 ( n17427, n19736, g35 );
nor U17393 ( n17426, n10972, n17428 );
or U17394 ( n17428, n17425, n19737 );
nor U17395 ( n17425, n17408, n17429 );
nand U17396 ( n2525, n17430, n17431 );
nand U17397 ( n17431, n17432, n10944 );
nor U17398 ( n17430, n17433, n17434 );
nor U17399 ( n17434, n19735, g35 );
nor U17400 ( n17433, n10973, n17435 );
or U17401 ( n17435, n17432, n19736 );
and U17402 ( n17432, n17422, n17401 );
nand U17403 ( n2520, n17436, n17437 );
nand U17404 ( n17437, n17438, n10943 );
nor U17405 ( n17436, n17439, n17440 );
nor U17406 ( n17440, n19734, g35 );
nor U17407 ( n17439, n10973, n17441 );
or U17408 ( n17441, n17438, n19735 );
nand U17409 ( n2515, n17442, n17443 );
or U17410 ( n17443, n17444, n15730 );
nor U17411 ( n17442, n17445, n17446 );
nor U17412 ( n17446, n19733, g35 );
nor U17413 ( n17445, n10973, n17447 );
nand U17414 ( n17447, n17444, n10859 );
nand U17415 ( n17444, n17448, n17380 );
nand U17416 ( n2510, n17449, n17450 );
nand U17417 ( n17450, n17451, n10942 );
nor U17418 ( n17449, n17452, n17453 );
nor U17419 ( n17453, n19732, g35 );
nor U17420 ( n17452, n10973, n17454 );
or U17421 ( n17454, n17451, n19733 );
and U17422 ( n17451, n17448, n17387 );
nand U17423 ( n2505, n17455, n17456 );
or U17424 ( n17456, n17457, n15730 );
nor U17425 ( n17455, n17458, n17459 );
nor U17426 ( n17459, n19731, g35 );
nor U17427 ( n17458, n10973, n17460 );
nand U17428 ( n17460, n17457, n10860 );
nand U17429 ( n17457, n17448, n17394 );
nand U17430 ( n2500, n17461, n17462 );
or U17431 ( n17462, n17463, n15730 );
nor U17432 ( n17461, n17464, n17465 );
nor U17433 ( n17465, n19730, g35 );
nor U17434 ( n17464, n10973, n17466 );
nand U17435 ( n17466, n17463, n10806 );
nand U17436 ( n17463, n17448, n17401 );
nand U17437 ( n2495, n17467, n17468 );
nand U17438 ( n17468, n17469, n10944 );
nor U17439 ( n17467, n17470, n17471 );
nor U17440 ( n17471, n19729, g35 );
nor U17441 ( n17470, n10973, n17472 );
or U17442 ( n17472, n17469, n19730 );
and U17443 ( n17469, n17473, n10399 );
nand U17444 ( n2490, n17474, n17475 );
nand U17445 ( n17475, n17476, n10943 );
nor U17446 ( n17474, n17477, n17478 );
nor U17447 ( n17478, n19728, g35 );
nor U17448 ( n17477, n10973, n17479 );
or U17449 ( n17479, n17476, n19729 );
and U17450 ( n17476, n17473, n17380 );
nand U17451 ( n2485, n17480, n17481 );
nand U17452 ( n17481, n17482, n10942 );
nor U17453 ( n17480, n17483, n17484 );
nor U17454 ( n17484, n19727, g35 );
nor U17455 ( n17483, n10974, n17485 );
or U17456 ( n17485, n17482, n19728 );
and U17457 ( n17482, n17473, n17387 );
nand U17458 ( n2480, n17486, n17487 );
nand U17459 ( n17487, n17488, n10944 );
nor U17460 ( n17486, n17489, n17490 );
nor U17461 ( n17490, n19726, g35 );
nor U17462 ( n17489, n10974, n17491 );
or U17463 ( n17491, n17488, n19727 );
and U17464 ( n17488, n17473, n17394 );
nand U17465 ( n2475, n17492, n17493 );
nand U17466 ( n17493, n17494, n10943 );
nor U17467 ( n17492, n17495, n17496 );
nor U17468 ( n17496, n19725, g35 );
nor U17469 ( n17495, n10974, n17497 );
or U17470 ( n17497, n17494, n19726 );
and U17471 ( n17494, n17473, n17401 );
and U17472 ( n17401, n17498, n19723 );
nor U17473 ( n17498, n10248, n10468 );
nor U17474 ( n17473, n10598, n10275 );
nand U17475 ( n2470, n17499, n17500 );
nand U17476 ( n17500, n17501, n17502 );
nand U17477 ( n17501, n17503, n17504 );
nand U17478 ( n17504, n2342, n19723 );
nor U17479 ( n17503, n17438, n17505 );
nor U17480 ( n17505, n10976, n17408 );
not U17481 ( n17408, n17422 );
nor U17482 ( n17422, n10275, n19725 );
and U17483 ( n17438, n17448, n10399 );
nor U17484 ( n17448, n10598, n19724 );
nand U17485 ( n17499, n10993, n10275 );
nand U17486 ( n2465, n17506, n17507 );
nand U17487 ( n17507, n17508, n10399 );
nand U17488 ( n17508, g35, n17509 );
nand U17489 ( n17509, n19724, n17502 );
or U17490 ( n17506, n17510, n19724 );
nand U17491 ( n2460, n17511, n17512 );
nand U17492 ( n17512, n17513, n19723 );
nor U17493 ( n17513, n17514, n17415 );
not U17494 ( n17415, n17380 );
nor U17495 ( n17380, n19722, n19721 );
nand U17496 ( n17511, n10995, n10468 );
nand U17497 ( n2455, n17515, n17516 );
nand U17498 ( n17516, n17517, n17502 );
nand U17499 ( n17517, n17429, n17518 );
nand U17500 ( n17518, n17387, g35 );
nor U17501 ( n17387, n10248, n19722 );
not U17502 ( n17429, n17394 );
nor U17503 ( n17394, n10468, n19721 );
nand U17504 ( n17515, n10994, n10248 );
nor U17505 ( n2450, n10248, n17510 );
nand U17506 ( n17510, n17519, n19723 );
nor U17507 ( n17519, n17514, n10991 );
not U17508 ( n17514, n17502 );
nand U17509 ( n17502, n16208, n17192 );
nor U17510 ( n16208, n19938, n10232 );
nand U17511 ( n2356, n17520, n17521 );
nand U17512 ( n17521, g35, n10329 );
nand U17513 ( n17520, n10994, n10885 );
nand U17514 ( n2351, n17522, n17523 );
nand U17515 ( n17523, n10993, n10886 );
nand U17516 ( n17522, n17524, g35 );
nor U17517 ( n17524, n17525, g9680 );
nor U17518 ( n17525, n17526, n10885 );
nor U17519 ( n17526, n19720, n10886 );
nor U17520 ( n2342, n10974, n19725 );
nand U17521 ( n2337, n17527, n17528 );
nand U17522 ( n17528, n17529, n17338 );
nor U17523 ( n17527, n17530, n17531 );
nor U17524 ( n17531, n17532, n10991 );
nor U17525 ( n17532, n17533, n17534 );
nor U17526 ( n17534, n17535, n17327 );
nor U17527 ( n17533, n19437, n17286 );
nor U17528 ( n17530, n19719, g35 );
nand U17529 ( n2332, n17536, n17537 );
nand U17530 ( n17537, n17296, n10262 );
nor U17531 ( n17536, n17538, n17539 );
nor U17532 ( n17539, n19718, g35 );
nor U17533 ( n17538, n10974, n17540 );
nand U17534 ( n17540, n17529, n19719 );
nor U17535 ( n17529, n17535, n17280 );
nor U17536 ( n17535, n16230, n11111 );
nand U17537 ( n16230, n17541, n13438 );
nor U17538 ( n17541, n19430, n19589 );
nor U17539 ( n2327, n19717, n17542 );
and U17540 ( n17542, g35, n17543 );
nand U17541 ( n2322, n17544, n17545 );
nand U17542 ( n17545, n10995, n10329 );
nand U17543 ( n17544, n17546, g35 );
nor U17544 ( n17546, n17543, n10690 );
nor U17545 ( n17543, n17547, n19716 );
nand U17546 ( n2317, n17548, n17549 );
or U17547 ( n17549, g35, n19404 );
nand U17548 ( n17548, n17550, g35 );
xnor U17549 ( n17550, n17547, n10329 );
nand U17550 ( n17547, n17551, n17552 );
nor U17551 ( n17552, n19405, n19713 );
nor U17552 ( n17551, n19714, n19715 );
nor U17553 ( n2276, n17553, n17554 );
nand U17554 ( n17554, n17555, n19406 );
nor U17555 ( n17555, n17556, n17557 );
nor U17556 ( n17557, n19714, g14738 );
nor U17557 ( n17556, n19713, g12350 );
nand U17558 ( n17553, n17558, n19407 );
nor U17559 ( n17558, n10975, g17607 );
nor U17560 ( n2271, n19481, n10990 );
nand U17561 ( n2266, n17559, n17560 );
or U17562 ( n17560, n17561, n19529 );
nor U17563 ( n17559, n17562, n17563 );
nor U17564 ( n17563, n10735, n17564 );
nand U17565 ( n17564, n17565, n19711 );
nor U17566 ( n17565, n17566, n10990 );
nor U17567 ( n17562, n19712, n17567 );
nor U17568 ( n17567, n17568, n10989 );
nor U17569 ( n17568, n19711, n17566 );
nand U17570 ( n2261, n17569, n17570 );
nand U17571 ( n17570, n17571, n10735 );
or U17572 ( n17569, n17571, n19711 );
nand U17573 ( n2256, n17572, n17573 );
nand U17574 ( n17573, n10993, n10780 );
nor U17575 ( n17572, n17574, n17575 );
and U17576 ( n17575, n19711, n17576 );
nor U17577 ( n17574, n19711, n17577 );
nand U17578 ( n2251, n17578, n17579 );
nand U17579 ( n17579, n17580, n10780 );
nor U17580 ( n17578, n17581, n17582 );
nor U17581 ( n17582, n10736, n17583 );
nand U17582 ( n17583, n19409, n17576 );
nor U17583 ( n17581, n19408, n17584 );
nor U17584 ( n17584, n17585, n10989 );
nor U17585 ( n17585, n19409, n17586 );
nand U17586 ( n2246, n17587, n17588 );
nand U17587 ( n17588, n17580, n10736 );
nand U17588 ( n17587, n17577, n10623 );
nand U17589 ( n2241, n17589, n17590 );
nand U17590 ( n17590, n17571, n10623 );
nor U17591 ( n17589, n17591, n17592 );
nor U17592 ( n17592, n19514, g35 );
nor U17593 ( n17591, n10975, n17593 );
nand U17594 ( n17593, n19409, n11195 );
nand U17595 ( n2236, n17594, n17595 );
nand U17596 ( n17595, n17580, n10625 );
not U17597 ( n17580, n17577 );
nand U17598 ( n17577, g35, n17586 );
nor U17599 ( n17594, n17596, n17597 );
nor U17600 ( n17597, n10490, n17598 );
nand U17601 ( n17598, n17576, n10379 );
nor U17602 ( n17576, n17586, n10989 );
nor U17603 ( n17596, n19710, n17599 );
nor U17604 ( n17599, n17600, n10989 );
nor U17605 ( n17600, n17586, n10379 );
nand U17606 ( n2231, n17601, n17602 );
nand U17607 ( n17602, n10993, n10379 );
nand U17608 ( n17601, n17603, g35 );
nor U17609 ( n17603, n17604, n17605 );
nand U17610 ( n17605, n17606, n17607 );
nand U17611 ( n17607, n17608, n17586 );
nor U17612 ( n17608, n17609, n17610 );
nand U17613 ( n17610, n17611, n10490 );
or U17614 ( n17606, n17611, n17586 );
nand U17615 ( n17586, n17612, n17613 );
nor U17616 ( n17613, n19416, n19680 );
nor U17617 ( n17612, n11118, n17609 );
nor U17618 ( n17604, n17614, n10490 );
and U17619 ( n17614, n17611, n17615 );
nand U17620 ( n2226, n17616, n17617 );
nand U17621 ( n17617, n17571, n10379 );
nand U17622 ( n17616, n17561, n10861 );
nand U17623 ( n2221, n17618, n17619 );
nand U17624 ( n17619, n17620, n17571 );
nor U17625 ( n17620, n19410, n15980 );
nand U17626 ( n17618, n10944, n17621 );
nand U17627 ( n17621, n10861, n17566 );
nand U17628 ( n2216, n17622, n17623 );
nand U17629 ( n17623, n17624, n10892 );
nor U17630 ( n17622, n17625, n17626 );
nor U17631 ( n17626, n10975, n17627 );
nand U17632 ( n17627, n17615, n17611 );
nand U17633 ( n17611, n17628, n17629 );
nand U17634 ( n17629, n19680, n17630 );
nand U17635 ( n17630, n17631, n17632 );
nor U17636 ( n17632, n17633, n17634 );
nand U17637 ( n17634, n17635, n17636 );
nand U17638 ( n17636, n17637, n17638 );
nor U17639 ( n17637, n19413, n19702 );
nand U17640 ( n17635, n17639, n17640 );
nor U17641 ( n17639, n19411, n19701 );
nor U17642 ( n17633, n17641, n17642 );
nor U17643 ( n17641, n17643, n17644 );
nor U17644 ( n17644, n19416, n19699 );
nor U17645 ( n17643, n19412, n19703 );
nor U17646 ( n17631, n17645, n17646 );
nand U17647 ( n17646, n17647, n17648 );
nand U17648 ( n17648, n19415, n17649 );
nand U17649 ( n17647, n17650, g12300 );
nand U17650 ( n17650, n17651, n17652 );
nand U17651 ( n17652, n17640, n10807 );
not U17652 ( n17651, n17653 );
nor U17653 ( n17645, n17654, n17655 );
nor U17654 ( n17654, n17656, n17657 );
nor U17655 ( n17657, n19417, n19700 );
nor U17656 ( n17656, n19414, n19704 );
nand U17657 ( n17628, n17658, n10330 );
nand U17658 ( n17658, n17659, n17660 );
nor U17659 ( n17660, n17661, n17662 );
nand U17660 ( n17662, n17663, n17664 );
nand U17661 ( n17664, n17665, n17666 );
nor U17662 ( n17665, n19411, n19691 );
nand U17663 ( n17663, n17667, n17668 );
nor U17664 ( n17667, n19413, n19692 );
nor U17665 ( n17661, n17669, n17670 );
nor U17666 ( n17669, n17671, n17672 );
nor U17667 ( n17672, n19417, n19690 );
nor U17668 ( n17671, n19414, n19694 );
nor U17669 ( n17659, n17673, n17674 );
nand U17670 ( n17674, n17675, n17676 );
nand U17671 ( n17676, n19415, n17653 );
nand U17672 ( n17653, n17677, n17678 );
nand U17673 ( n17678, n17679, n17668 );
nor U17674 ( n17679, n19679, n19708 );
nor U17675 ( n17677, n17680, n17681 );
nor U17676 ( n17681, n17670, n17682 );
nand U17677 ( n17682, n10862, g14694 );
nor U17678 ( n17680, n17642, n17683 );
or U17679 ( n17683, n19707, n19678 );
nand U17680 ( n17675, n17684, g12300 );
nand U17681 ( n17684, n17685, n17686 );
nand U17682 ( n17686, n17666, n10808 );
not U17683 ( n17685, n17649 );
nand U17684 ( n17649, n17687, n17688 );
nand U17685 ( n17688, n17689, n17640 );
nor U17686 ( n17689, n19678, n19697 );
nor U17687 ( n17687, n17690, n17691 );
nor U17688 ( n17691, n17655, n17692 );
nand U17689 ( n17692, n10864, g14694 );
nor U17690 ( n17690, n17670, n17693 );
nand U17691 ( n17693, n10863, g17580 );
nor U17692 ( n17673, n17694, n11118 );
nor U17693 ( n17694, n17695, n17696 );
nor U17694 ( n17696, n19412, n19693 );
nor U17695 ( n17695, n19416, n19709 );
nor U17696 ( n17625, n19709, g35 );
nand U17697 ( n2211, n17697, n17698 );
nand U17698 ( n17698, n10994, n10766 );
nor U17699 ( n17697, n17699, n17700 );
nor U17700 ( n17700, n17566, n15730 );
nor U17701 ( n17699, n19709, n17561 );
not U17702 ( n17561, n17571 );
nor U17703 ( n17571, n10976, n11195 );
not U17704 ( n11195, n17566 );
nand U17705 ( n17566, n17701, n10305 );
nand U17706 ( n2206, n17702, n17703 );
or U17707 ( n17703, n17704, n15730 );
nor U17708 ( n17702, n17705, n17706 );
nor U17709 ( n17706, n19707, g35 );
nor U17710 ( n17705, n10976, n17707 );
nand U17711 ( n17707, n17704, n10766 );
nand U17712 ( n17704, n17708, n17701 );
nand U17713 ( n2201, n17709, n17710 );
nand U17714 ( n17710, n17711, n10942 );
nor U17715 ( n17709, n17712, n17713 );
nor U17716 ( n17713, n19706, g35 );
nor U17717 ( n17712, n10976, n17714 );
or U17718 ( n17714, n17711, n19707 );
and U17719 ( n17711, n17715, n17701 );
nand U17720 ( n2196, n17716, n17717 );
or U17721 ( n17717, n17718, n15730 );
nor U17722 ( n17716, n17719, n17720 );
nor U17723 ( n17720, n19705, g35 );
nor U17724 ( n17719, n10976, n17721 );
nand U17725 ( n17721, n17718, n10862 );
nand U17726 ( n17718, n17722, n17701 );
nand U17727 ( n2191, n17723, n17724 );
or U17728 ( n17724, n17725, n15730 );
nor U17729 ( n17723, n17726, n17727 );
nor U17730 ( n17727, n19704, g35 );
nor U17731 ( n17726, n10976, n17728 );
nand U17732 ( n17728, n17725, n10807 );
nand U17733 ( n17725, n17729, n17701 );
nor U17734 ( n17701, n19689, n19688 );
nand U17735 ( n2186, n17730, n17731 );
nand U17736 ( n17731, n17732, n10944 );
nor U17737 ( n17730, n17733, n17734 );
nor U17738 ( n17734, n19703, g35 );
nor U17739 ( n17733, n10976, n17735 );
or U17740 ( n17735, n17732, n19704 );
and U17741 ( n17732, n17736, n10305 );
nand U17742 ( n2181, n17737, n17738 );
nand U17743 ( n17738, n17739, n10943 );
nor U17744 ( n17737, n17740, n17741 );
nor U17745 ( n17741, n19702, g35 );
nor U17746 ( n17740, n10976, n17742 );
or U17747 ( n17742, n17739, n19703 );
and U17748 ( n17739, n17736, n17708 );
nand U17749 ( n2176, n17743, n17744 );
nand U17750 ( n17744, n17745, n10942 );
nor U17751 ( n17743, n17746, n17747 );
nor U17752 ( n17747, n19701, g35 );
nor U17753 ( n17746, n10976, n17748 );
or U17754 ( n17748, n17745, n19702 );
and U17755 ( n17745, n17736, n17715 );
nand U17756 ( n2171, n17749, n17750 );
nand U17757 ( n17750, n17751, n10944 );
nor U17758 ( n17749, n17752, n17753 );
nor U17759 ( n17753, n19700, g35 );
nor U17760 ( n17752, n10977, n17754 );
or U17761 ( n17754, n17751, n19701 );
and U17762 ( n17751, n17736, n17722 );
nand U17763 ( n2166, n17755, n17756 );
nand U17764 ( n17756, n17757, n10943 );
nor U17765 ( n17755, n17758, n17759 );
nor U17766 ( n17759, n19699, g35 );
nor U17767 ( n17758, n10977, n17760 );
or U17768 ( n17760, n17757, n19700 );
and U17769 ( n17757, n17736, n17729 );
nand U17770 ( n2161, n17761, n17762 );
nand U17771 ( n17762, n17763, n10942 );
nor U17772 ( n17761, n17764, n17765 );
nor U17773 ( n17765, n19698, g35 );
nor U17774 ( n17764, n10977, n17766 );
or U17775 ( n17766, n17763, n19699 );
and U17776 ( n17763, n17767, n10305 );
nand U17777 ( n2156, n17768, n17769 );
or U17778 ( n17769, n17770, n15730 );
nor U17779 ( n17768, n17771, n17772 );
nor U17780 ( n17772, n19697, g35 );
nor U17781 ( n17771, n10977, n17773 );
nand U17782 ( n17773, n17770, n10863 );
nand U17783 ( n17770, n17767, n17708 );
nand U17784 ( n2151, n17774, n17775 );
nand U17785 ( n17775, n17776, n10944 );
nor U17786 ( n17774, n17777, n17778 );
nor U17787 ( n17778, n19696, g35 );
nor U17788 ( n17777, n10977, n17779 );
or U17789 ( n17779, n17776, n19697 );
and U17790 ( n17776, n17767, n17715 );
nand U17791 ( n2146, n17780, n17781 );
or U17792 ( n17781, n17782, n15730 );
nor U17793 ( n17780, n17783, n17784 );
nor U17794 ( n17784, n19695, g35 );
nor U17795 ( n17783, n10977, n17785 );
nand U17796 ( n17785, n17782, n10864 );
nand U17797 ( n17782, n17767, n17722 );
nand U17798 ( n2141, n17786, n17787 );
or U17799 ( n17787, n17788, n15730 );
nor U17800 ( n17786, n17789, n17790 );
nor U17801 ( n17790, n19694, g35 );
nor U17802 ( n17789, n10977, n17791 );
nand U17803 ( n17791, n17788, n10808 );
nand U17804 ( n17788, n17767, n17729 );
nand U17805 ( n2136, n17792, n17793 );
nand U17806 ( n17793, n17794, n10943 );
nor U17807 ( n17792, n17795, n17796 );
nor U17808 ( n17796, n19693, g35 );
nor U17809 ( n17795, n10977, n17797 );
or U17810 ( n17797, n17794, n19694 );
and U17811 ( n17794, n17798, n10305 );
nand U17812 ( n2131, n17799, n17800 );
nand U17813 ( n17800, n17801, n10942 );
nor U17814 ( n17799, n17802, n17803 );
nor U17815 ( n17803, n19692, g35 );
nor U17816 ( n17802, n10977, n17804 );
or U17817 ( n17804, n17801, n19693 );
and U17818 ( n17801, n17798, n17708 );
nand U17819 ( n2126, n17805, n17806 );
nand U17820 ( n17806, n17807, n10944 );
nor U17821 ( n17805, n17808, n17809 );
nor U17822 ( n17809, n19691, g35 );
nor U17823 ( n17808, n10978, n17810 );
or U17824 ( n17810, n17807, n19692 );
and U17825 ( n17807, n17798, n17715 );
nand U17826 ( n2121, n17811, n17812 );
nand U17827 ( n17812, n17813, n10943 );
nor U17828 ( n17811, n17814, n17815 );
nor U17829 ( n17815, n19690, g35 );
nor U17830 ( n17814, n10977, n17816 );
or U17831 ( n17816, n17813, n19691 );
and U17832 ( n17813, n17798, n17722 );
nand U17833 ( n2116, n17817, n17818 );
nand U17834 ( n17818, n17819, n10942 );
nor U17835 ( n17817, n17820, n17821 );
nor U17836 ( n17821, n19689, g35 );
nor U17837 ( n17820, n10978, n17822 );
or U17838 ( n17822, n17819, n19690 );
and U17839 ( n17819, n17798, n17729 );
and U17840 ( n17729, n17823, n19687 );
nor U17841 ( n17823, n10249, n10469 );
nor U17842 ( n17798, n10268, n10435 );
nand U17843 ( n2111, n17824, n17825 );
nand U17844 ( n17825, n10993, n10435 );
nand U17845 ( n17824, n17826, g35 );
nor U17846 ( n17826, n17827, n17828 );
nor U17847 ( n17828, n17736, n17829 );
nand U17848 ( n17829, n17830, n17831 );
nand U17849 ( n17831, n19687, n10268 );
nand U17850 ( n17830, n17767, n10305 );
nor U17851 ( n17767, n10268, n19688 );
nor U17852 ( n17736, n10435, n19689 );
nand U17853 ( n2106, n17832, n17833 );
nand U17854 ( n17833, n17834, n10305 );
nand U17855 ( n17834, g35, n17835 );
nand U17856 ( n17835, n19688, n17836 );
or U17857 ( n17832, n17837, n19688 );
nand U17858 ( n2101, n17838, n17839 );
nand U17859 ( n17839, n17840, n19687 );
and U17860 ( n17840, n17836, n17708 );
nor U17861 ( n17708, n19686, n19685 );
nand U17862 ( n17838, n10994, n10469 );
not U17863 ( n210, n17841 );
nand U17864 ( n2096, n17842, n17843 );
nand U17865 ( n17843, n17844, n17836 );
nand U17866 ( n17844, n17845, n17846 );
nand U17867 ( n17846, n17715, g35 );
nor U17868 ( n17715, n10249, n19686 );
not U17869 ( n17845, n17722 );
nor U17870 ( n17722, n10469, n19685 );
nand U17871 ( n17842, n10994, n10249 );
nor U17872 ( n2091, n10249, n17837 );
nand U17873 ( n17837, n17847, n19687 );
nor U17874 ( n17847, n17827, n10988 );
not U17875 ( n17827, n17836 );
nand U17876 ( n17836, n17192, n11194 );
nor U17877 ( n11194, n10421, n19937 );
nand U17878 ( n1997, n17848, n17849 );
nand U17879 ( n17849, g35, n10330 );
nand U17880 ( n17848, n10995, n10887 );
nand U17881 ( n1992, n17850, n17851 );
nand U17882 ( n17851, n10995, n10888 );
nand U17883 ( n17850, n17852, g35 );
nor U17884 ( n17852, n17853, g9615 );
nor U17885 ( n17853, n17854, n10887 );
nor U17886 ( n17854, n19684, n10888 );
nor U17887 ( n1983, n19689, n10988 );
nand U17888 ( n1978, n17855, n17856 );
nand U17889 ( n17856, n17857, n17858 );
nand U17890 ( n17857, n17859, n17860 );
nand U17891 ( n17860, g35, n17861 );
nand U17892 ( n17861, n17655, n17862 );
nand U17893 ( n17862, n17609, n10471 );
not U17894 ( n17655, n17668 );
nand U17895 ( n17859, n17666, n17615 );
nand U17896 ( n17855, n10997, n10242 );
nand U17897 ( n1973, n17863, n17864 );
nand U17898 ( n17864, n17624, n10242 );
nor U17899 ( n17863, n17865, n17866 );
nor U17900 ( n17866, n19682, g35 );
nor U17901 ( n17865, n10979, n17867 );
nand U17902 ( n17867, n17868, n19683 );
and U17903 ( n17868, n17858, n17615 );
nand U17904 ( n17858, n17869, n17615 );
nor U17905 ( n17869, n11103, n16557 );
nand U17906 ( n11103, n17214, n10223 );
nor U17907 ( n1968, n19681, n17870 );
and U17908 ( n17870, g35, n17871 );
nand U17909 ( n1963, n17872, n17873 );
nand U17910 ( n17873, n10995, n10330 );
nand U17911 ( n17872, n17874, g35 );
nor U17912 ( n17874, n17871, n10739 );
nor U17913 ( n17871, n17875, n19680 );
nand U17914 ( n1958, n17876, n17877 );
or U17915 ( n17877, g35, n19414 );
nand U17916 ( n17876, n17878, g35 );
xnor U17917 ( n17878, n17875, n10330 );
nand U17918 ( n17875, n17879, n17880 );
nor U17919 ( n17880, n19415, n19677 );
nor U17920 ( n17879, n19678, n19679 );
nor U17921 ( n1917, n17881, n17882 );
nand U17922 ( n17882, n17883, n19416 );
nor U17923 ( n17883, n17884, n17885 );
nor U17924 ( n17885, n19678, g14694 );
nor U17925 ( n17884, n19677, g12300 );
nand U17926 ( n17881, n17886, n19417 );
nor U17927 ( n17886, n10979, g17580 );
nor U17928 ( n1912, n19472, n10987 );
nand U17929 ( n1907, n17887, n17888 );
or U17930 ( n17888, n17889, n19527 );
nor U17931 ( n17887, n17890, n17891 );
nor U17932 ( n17891, n10737, n17892 );
nand U17933 ( n17892, n17893, n19675 );
nor U17934 ( n17893, n11219, n10987 );
nor U17935 ( n17890, n19676, n17894 );
nor U17936 ( n17894, n17895, n10987 );
nor U17937 ( n17895, n19675, n11219 );
nand U17938 ( n1902, n17896, n17897 );
nand U17939 ( n17897, n17898, n10737 );
or U17940 ( n17896, n17898, n19675 );
nand U17941 ( n1897, n17899, n17900 );
nand U17942 ( n17900, n10995, n10781 );
nor U17943 ( n17899, n17901, n17902 );
and U17944 ( n17902, n19675, n17903 );
nor U17945 ( n17901, n19675, n17904 );
nand U17946 ( n1892, n17905, n17906 );
nand U17947 ( n17906, n17907, n10781 );
nor U17948 ( n17905, n17908, n17909 );
nor U17949 ( n17909, n10738, n17910 );
nand U17950 ( n17910, n19419, n17903 );
nor U17951 ( n17908, n19418, n17911 );
nor U17952 ( n17911, n17912, n10987 );
nor U17953 ( n17912, n19419, n17913 );
nand U17954 ( n1887, n17914, n17915 );
nand U17955 ( n17915, n17907, n10738 );
not U17956 ( n17907, n17904 );
nand U17957 ( n17914, n17904, n10624 );
nand U17958 ( n17904, g35, n17913 );
nand U17959 ( n1882, n17916, n17917 );
nand U17960 ( n17917, n17898, n10624 );
nor U17961 ( n17916, n17918, n17919 );
nor U17962 ( n17919, n19515, g35 );
nor U17963 ( n17918, n10979, n17920 );
nand U17964 ( n17920, n19419, g26801 );
nand U17965 ( n1877, n17921, n17922 );
nand U17966 ( n17922, n17923, n17913 );
nor U17967 ( n17921, n17924, n17925 );
nor U17968 ( n17925, n10491, n17926 );
nand U17969 ( n17926, n17903, n10380 );
nor U17970 ( n17903, n17913, n10986 );
nor U17971 ( n17924, n19674, n17927 );
nor U17972 ( n17927, n17928, n10986 );
nor U17973 ( n17928, n17913, n10380 );
nand U17974 ( n1872, n17929, n17930 );
nand U17975 ( n17930, n10996, n10380 );
nand U17976 ( n17929, n17931, g35 );
nor U17977 ( n17931, n17932, n17933 );
nand U17978 ( n17933, n17934, n17935 );
nand U17979 ( n17935, n17936, n17913 );
nor U17980 ( n17936, n17937, n17938 );
nand U17981 ( n17938, n17939, n10491 );
or U17982 ( n17934, n17939, n17913 );
nand U17983 ( n17913, n17940, n17941 );
nor U17984 ( n17941, n19434, n19629 );
nor U17985 ( n17940, n11124, n17937 );
nor U17986 ( n17932, n17942, n10491 );
and U17987 ( n17942, n17939, g33959 );
nand U17988 ( n1867, n17943, n17944 );
nand U17989 ( n17944, n17898, n10380 );
nand U17990 ( n17943, n17889, n10865 );
nand U17991 ( n1862, n17945, n17946 );
nand U17992 ( n17946, n17947, n17898 );
nor U17993 ( n17947, n19420, n15980 );
nand U17994 ( n17945, n10943, n17948 );
nand U17995 ( n17948, n10865, n11219 );
nand U17996 ( n1857, n17949, n17950 );
nand U17997 ( n17950, n17951, g21245 );
nor U17998 ( n17949, n17952, n17953 );
nor U17999 ( n17953, n10979, n17954 );
nand U18000 ( n17954, g33959, n17939 );
nand U18001 ( n17939, n17955, n17956 );
nand U18002 ( n17956, n19629, n17957 );
nand U18003 ( n17957, n17958, n17959 );
nor U18004 ( n17959, n17960, n17961 );
nand U18005 ( n17961, n17962, n17963 );
nand U18006 ( n17963, n17964, n17965 );
nor U18007 ( n17964, n19423, n19667 );
nand U18008 ( n17962, n17966, g31860 );
nor U18009 ( n17966, n19422, n19666 );
nor U18010 ( n17960, n17967, n17968 );
nor U18011 ( n17967, n17969, n17970 );
nor U18012 ( n17970, n19435, n19665 );
nor U18013 ( n17969, n19431, n19669 );
nor U18014 ( n17958, n17971, n17972 );
nand U18015 ( n17972, n17973, n17974 );
nand U18016 ( n17974, n19433, n17975 );
nand U18017 ( n17973, n17976, g12238 );
nand U18018 ( n17976, n17977, n17978 );
nand U18019 ( n17978, g31860, n10809 );
not U18020 ( n17977, n17979 );
nor U18021 ( n17971, n17980, n17981 );
not U18022 ( n17981, n17982 );
nor U18023 ( n17980, n17983, n17984 );
nor U18024 ( n17984, n19434, n19664 );
nor U18025 ( n17983, n19421, n19668 );
nand U18026 ( n17955, n17985, g25219 );
nand U18027 ( n17985, n17986, n17987 );
nor U18028 ( n17987, n17988, n17989 );
nand U18029 ( n17989, n17990, n17991 );
nand U18030 ( n17991, n17992, n17993 );
nor U18031 ( n17992, n19423, n19657 );
nand U18032 ( n17990, n17994, n17982 );
nor U18033 ( n17994, n19422, n19656 );
nor U18034 ( n17988, n17995, n17996 );
nor U18035 ( n17995, n17997, n17998 );
nor U18036 ( n17998, n19435, n19655 );
nor U18037 ( n17997, n19431, n19659 );
nor U18038 ( n17986, n17999, n18000 );
nand U18039 ( n18000, n18001, n18002 );
nand U18040 ( n18002, n19433, n17979 );
nand U18041 ( n17979, n18003, n18004 );
nand U18042 ( n18004, n18005, n17982 );
nor U18043 ( n18005, n19432, n19672 );
nor U18044 ( n18003, n18006, n18007 );
nor U18045 ( n18007, n17968, n18008 );
nand U18046 ( n18008, n10563, g17519 );
nor U18047 ( n18006, n17996, n18009 );
nand U18048 ( n18009, n10866, g14662 );
nand U18049 ( n18001, n18010, g12238 );
nand U18050 ( n18010, n18011, n18012 );
nand U18051 ( n18012, n17982, n10810 );
not U18052 ( n18011, n17975 );
nand U18053 ( n17975, n18013, n18014 );
nand U18054 ( n18014, n18015, g31860 );
nor U18055 ( n18015, n19432, n19662 );
nor U18056 ( n18013, n18016, n18017 );
nor U18057 ( n18017, n17968, n18018 );
nand U18058 ( n18018, n10868, g14662 );
nor U18059 ( n18016, n17996, n18019 );
nand U18060 ( n18019, n10867, g17519 );
not U18061 ( n17996, n17965 );
nor U18062 ( n17999, n18020, n11124 );
not U18063 ( n11124, g31860 );
nor U18064 ( n18020, n18021, n18022 );
nor U18065 ( n18022, n19421, n19658 );
nor U18066 ( n18021, n19434, n19673 );
nor U18067 ( n17952, n19673, g35 );
nand U18068 ( n1852, n18023, n18024 );
nand U18069 ( n18024, n10996, n10563 );
nor U18070 ( n18023, n18025, n18026 );
nor U18071 ( n18026, n11219, n15730 );
nor U18072 ( n18025, n19673, n17889 );
not U18073 ( n17889, n17898 );
nor U18074 ( n17898, n10968, g26801 );
not U18075 ( g26801, n11219 );
nand U18076 ( n11219, n18027, n10306 );
nand U18077 ( n1847, n18028, n18029 );
or U18078 ( n18029, n18030, n15730 );
nor U18079 ( n18028, n18031, n18032 );
nor U18080 ( n18032, n19672, g35 );
nor U18081 ( n18031, n10963, n18033 );
nand U18082 ( n18033, n18030, n10563 );
nand U18083 ( n18030, n18034, n18027 );
nand U18084 ( n1842, n18035, n18036 );
nand U18085 ( n18036, n18037, n10944 );
nor U18086 ( n18035, n18038, n18039 );
nor U18087 ( n18039, n19671, g35 );
nor U18088 ( n18038, n10963, n18040 );
or U18089 ( n18040, n18037, n19672 );
and U18090 ( n18037, n18041, n18027 );
nand U18091 ( n1837, n18042, n18043 );
or U18092 ( n18043, n18044, n15730 );
nor U18093 ( n18042, n18045, n18046 );
nor U18094 ( n18046, n19670, g35 );
nor U18095 ( n18045, n10963, n18047 );
nand U18096 ( n18047, n18044, n10866 );
nand U18097 ( n18044, n18048, n18027 );
nand U18098 ( n1832, n18049, n18050 );
or U18099 ( n18050, n18051, n15730 );
nor U18100 ( n18049, n18052, n18053 );
nor U18101 ( n18053, n19669, g35 );
nor U18102 ( n18052, n10964, n18054 );
nand U18103 ( n18054, n18051, n10809 );
nand U18104 ( n18051, n18055, n18027 );
nor U18105 ( n18027, n19654, n19653 );
nand U18106 ( n1827, n18056, n18057 );
nand U18107 ( n18057, n18058, n10943 );
nor U18108 ( n18056, n18059, n18060 );
nor U18109 ( n18060, n19668, g35 );
nor U18110 ( n18059, n10964, n18061 );
or U18111 ( n18061, n18058, n19669 );
and U18112 ( n18058, n18062, n10306 );
nand U18113 ( n1822, n18063, n18064 );
nand U18114 ( n18064, n18065, n10942 );
nor U18115 ( n18063, n18066, n18067 );
nor U18116 ( n18067, n19667, g35 );
nor U18117 ( n18066, n10964, n18068 );
or U18118 ( n18068, n18065, n19668 );
and U18119 ( n18065, n18062, n18034 );
nand U18120 ( n1817, n18069, n18070 );
nand U18121 ( n18070, n18071, n10944 );
nor U18122 ( n18069, n18072, n18073 );
nor U18123 ( n18073, n19666, g35 );
nor U18124 ( n18072, n10964, n18074 );
or U18125 ( n18074, n18071, n19667 );
and U18126 ( n18071, n18062, n18041 );
nand U18127 ( n1812, n18075, n18076 );
nand U18128 ( n18076, n18077, n10943 );
nor U18129 ( n18075, n18078, n18079 );
nor U18130 ( n18079, n19665, g35 );
nor U18131 ( n18078, n10964, n18080 );
or U18132 ( n18080, n18077, n19666 );
and U18133 ( n18077, n18062, n18048 );
nand U18134 ( n1807, n18081, n18082 );
nand U18135 ( n18082, n18083, n10942 );
nor U18136 ( n18081, n18084, n18085 );
nor U18137 ( n18085, n19664, g35 );
nor U18138 ( n18084, n10964, n18086 );
or U18139 ( n18086, n18083, n19665 );
and U18140 ( n18083, n18062, n18055 );
nand U18141 ( n1802, n18087, n18088 );
nand U18142 ( n18088, n18089, n10944 );
nor U18143 ( n18087, n18090, n18091 );
nor U18144 ( n18091, n19663, g35 );
nor U18145 ( n18090, n10964, n18092 );
or U18146 ( n18092, n18089, n19664 );
and U18147 ( n18089, n18093, n10306 );
nand U18148 ( n1797, n18094, n18095 );
or U18149 ( n18095, n18096, n15730 );
nor U18150 ( n18094, n18097, n18098 );
nor U18151 ( n18098, n19662, g35 );
nor U18152 ( n18097, n10964, n18099 );
nand U18153 ( n18099, n18096, n10867 );
nand U18154 ( n18096, n18093, n18034 );
nand U18155 ( n1792, n18100, n18101 );
nand U18156 ( n18101, n18102, n10943 );
nor U18157 ( n18100, n18103, n18104 );
nor U18158 ( n18104, n19661, g35 );
nor U18159 ( n18103, n10964, n18105 );
or U18160 ( n18105, n18102, n19662 );
and U18161 ( n18102, n18093, n18041 );
nand U18162 ( n1787, n18106, n18107 );
or U18163 ( n18107, n18108, n15730 );
nor U18164 ( n18106, n18109, n18110 );
nor U18165 ( n18110, n19660, g35 );
nor U18166 ( n18109, n10964, n18111 );
nand U18167 ( n18111, n18108, n10868 );
nand U18168 ( n18108, n18093, n18048 );
nand U18169 ( n1782, n18112, n18113 );
or U18170 ( n18113, n18114, n15730 );
nor U18171 ( n18112, n18115, n18116 );
nor U18172 ( n18116, n19659, g35 );
nor U18173 ( n18115, n10964, n18117 );
nand U18174 ( n18117, n18114, n10810 );
nand U18175 ( n18114, n18093, n18055 );
nand U18176 ( n1777, n18118, n18119 );
nand U18177 ( n18119, n18120, n10942 );
nor U18178 ( n18118, n18121, n18122 );
nor U18179 ( n18122, n19658, g35 );
nor U18180 ( n18121, n10964, n18123 );
or U18181 ( n18123, n18120, n19659 );
and U18182 ( n18120, n18124, n10306 );
nand U18183 ( n1772, n18125, n18126 );
nand U18184 ( n18126, n18127, n10944 );
nor U18185 ( n18125, n18128, n18129 );
nor U18186 ( n18129, n19657, g35 );
nor U18187 ( n18128, n10965, n18130 );
or U18188 ( n18130, n18127, n19658 );
and U18189 ( n18127, n18124, n18034 );
not U18190 ( n177, n18131 );
nand U18191 ( n1767, n18132, n18133 );
nand U18192 ( n18133, n18134, n10943 );
nor U18193 ( n18132, n18135, n18136 );
nor U18194 ( n18136, n19656, g35 );
nor U18195 ( n18135, n10965, n18137 );
or U18196 ( n18137, n18134, n19657 );
and U18197 ( n18134, n18124, n18041 );
nand U18198 ( n1762, n18138, n18139 );
nand U18199 ( n18139, n18140, n10944 );
nor U18200 ( n18138, n18141, n18142 );
nor U18201 ( n18142, n19655, g35 );
nor U18202 ( n18141, n10965, n18143 );
or U18203 ( n18143, n18140, n19656 );
and U18204 ( n18140, n18124, n18048 );
nand U18205 ( n1757, n18144, n18145 );
nand U18206 ( n18145, n18146, n10943 );
not U18207 ( n15649, n15980 );
nand U18208 ( n15980, n19424, n10457 );
nor U18209 ( n18144, n18147, n18148 );
nor U18210 ( n18148, n19654, g35 );
nor U18211 ( n18147, n10965, n18149 );
or U18212 ( n18149, n18146, n19655 );
and U18213 ( n18146, n18124, n18055 );
and U18214 ( n18055, n18150, n19652 );
nor U18215 ( n18150, n10250, n10470 );
nor U18216 ( n18124, n10269, n10436 );
nand U18217 ( n1752, n18151, n18152 );
nand U18218 ( n18152, n10997, n10436 );
nand U18219 ( n18151, n18153, g35 );
nor U18220 ( n18153, n18154, n18155 );
nor U18221 ( n18155, n18062, n18156 );
nand U18222 ( n18156, n18157, n18158 );
nand U18223 ( n18158, n19652, n10269 );
nand U18224 ( n18157, n18093, n10306 );
nor U18225 ( n18093, n10269, n19653 );
nor U18226 ( n18062, n10436, n19654 );
nand U18227 ( n1747, n18159, n18160 );
nand U18228 ( n18160, n18161, n10306 );
nand U18229 ( n18161, g35, n18162 );
nand U18230 ( n18162, n19653, n18163 );
or U18231 ( n18159, n18164, n19653 );
nand U18232 ( n1742, n18165, n18166 );
nand U18233 ( n18166, n18167, n19652 );
and U18234 ( n18167, n18163, n18034 );
nor U18235 ( n18034, n19651, n19650 );
nand U18236 ( n18165, n10997, n10470 );
nand U18237 ( n1737, n18168, n18169 );
nand U18238 ( n18169, n18170, n18163 );
nand U18239 ( n18170, n18171, n18172 );
nand U18240 ( n18172, n18041, g35 );
nor U18241 ( n18041, n10250, n19651 );
not U18242 ( n18171, n18048 );
nor U18243 ( n18048, n10470, n19650 );
nand U18244 ( n18168, n10997, n10250 );
nor U18245 ( n1732, n10250, n18164 );
nand U18246 ( n18164, n18173, n19652 );
nor U18247 ( n18173, n18154, n10990 );
not U18248 ( n18154, n18163 );
nand U18249 ( n18163, n17192, n15513 );
nor U18250 ( n15513, n10232, n10421 );
and U18251 ( n17192, n16863, n18174 );
nor U18252 ( n18174, n19425, n10293 );
nor U18253 ( n16863, n11187, n13560 );
nand U18254 ( n11187, n18175, n18176 );
xnor U18255 ( n18176, n19940, n19562 );
xnor U18256 ( n18175, n19426, n19563 );
nand U18257 ( n1727, n18177, n18178 );
nand U18258 ( n18178, n19649, n18179 );
nor U18259 ( n18177, n18180, n18181 );
nor U18260 ( n18181, n19648, g35 );
nor U18261 ( n18180, n10965, n18182 );
or U18262 ( n18182, n18179, n19649 );
nor U18263 ( n18179, n18183, n19648 );
not U18264 ( n18183, n18184 );
nand U18265 ( n1722, n18185, n18186 );
nand U18266 ( n18186, n19648, n18184 );
nor U18267 ( n18185, n18187, n18188 );
nor U18268 ( n18188, n19427, g35 );
nor U18269 ( n18187, n10965, n18189 );
or U18270 ( n18189, n18184, n19648 );
nor U18271 ( n18184, n19427, n19647 );
xnor U18272 ( n1717, n18190, n10402 );
or U18273 ( n18190, n11024, n19427 );
nand U18274 ( n1712, n18191, n18192 );
nand U18275 ( n18192, n18193, n19644 );
nor U18276 ( n18193, n19645, n10985 );
nor U18277 ( n18191, n18194, n18195 );
nor U18278 ( n18195, n10923, n18196 );
nand U18279 ( n18196, n18197, n18198 );
or U18280 ( n18198, n10579, n19645 );
nor U18281 ( n18194, n19646, n18197 );
nor U18282 ( n18197, n10402, n10986 );
nor U18283 ( n1707, n19645, n18199 );
nor U18284 ( n18199, n10966, n18200 );
nand U18285 ( n18200, n18201, n18202 );
nand U18286 ( n18202, n19643, n10402 );
nand U18287 ( n18201, n19644, n19647 );
nor U18288 ( n1702, n19644, n18203 );
nor U18289 ( n18203, n10966, n10579 );
nand U18290 ( n1697, n18204, n18205 );
nand U18291 ( n18205, n11006, n10579 );
nand U18292 ( n18204, g35, n18206 );
nand U18293 ( n1692, n18207, n18208 );
nand U18294 ( n18208, n11006, n10445 );
nand U18295 ( n18207, g35, n18209 );
nand U18296 ( n1687, n18210, n18211 );
nand U18297 ( n18211, n18212, n19642 );
nor U18298 ( n18210, n18213, n18214 );
nor U18299 ( n18214, n19429, n18215 );
nor U18300 ( n18215, n10966, n18216 );
nand U18301 ( n18216, n18217, n18218 );
nand U18302 ( n18218, n18219, n10445 );
nor U18303 ( n18219, n18220, n18221 );
nand U18304 ( n18217, n18220, n19642 );
nor U18305 ( n18213, n10447, n18222 );
nand U18306 ( n18222, n18223, n10445 );
nand U18307 ( n1682, n18224, n18225 );
nor U18308 ( n18225, n18226, n18227 );
nor U18309 ( n18227, n10447, n18228 );
nor U18310 ( n18226, n19429, n18229 );
nand U18311 ( n18229, n18230, n18223 );
nor U18312 ( n18230, n18231, n18220 );
not U18313 ( n18220, n18228 );
nand U18314 ( n18228, n18232, n18233 );
nor U18315 ( n18232, n19640, n19641 );
nor U18316 ( n18224, n18212, n18234 );
nor U18317 ( n18234, n19641, g35 );
and U18318 ( n18212, n18235, n18231 );
and U18319 ( n18231, n18236, n18237 );
and U18320 ( n18236, n19640, n19641 );
nor U18321 ( n18235, n10966, n10447 );
nand U18322 ( n1677, n18238, n18239 );
nand U18323 ( n18239, n18240, n18241 );
not U18324 ( n18241, n18242 );
nor U18325 ( n18240, n19641, n18221 );
nor U18326 ( n18238, n18243, n18244 );
nor U18327 ( n18244, n19640, g35 );
nor U18328 ( n18243, n10966, n18245 );
nand U18329 ( n18245, n19641, n18242 );
nand U18330 ( n18242, n18246, n18247 );
nand U18331 ( n18247, n18233, n10583 );
nand U18332 ( n18246, n18237, n19640 );
nand U18333 ( n1672, n18248, n18249 );
nand U18334 ( n18249, n18250, n18251 );
nor U18335 ( n18250, n19640, n18221 );
nor U18336 ( n18248, n18252, n18253 );
nor U18337 ( n18253, n19639, g35 );
nor U18338 ( n18252, n10966, n18254 );
or U18339 ( n18254, n10583, n18251 );
nor U18340 ( n18251, n18237, n18233 );
and U18341 ( n18233, n18255, n18256 );
nor U18342 ( n18255, n19638, n19639 );
and U18343 ( n18237, n18257, n19638 );
nor U18344 ( n18257, n18258, n10591 );
nand U18345 ( n1667, n18259, n18260 );
nand U18346 ( n18260, n18261, n19639 );
nor U18347 ( n18259, n18262, n18263 );
nor U18348 ( n18263, n19638, n18264 );
nor U18349 ( n18264, n10966, n18265 );
nand U18350 ( n18265, n18266, n18267 );
nand U18351 ( n18267, n18268, n10591 );
nor U18352 ( n18268, n18256, n18221 );
nand U18353 ( n18266, n19639, n18256 );
nor U18354 ( n18262, n10594, n18269 );
nand U18355 ( n18269, n18270, n18223 );
nor U18356 ( n18270, n19639, n18271 );
nand U18357 ( n1662, n18272, n18273 );
nor U18358 ( n18273, n18274, n18275 );
nor U18359 ( n18275, n18276, n10594 );
nor U18360 ( n18274, n19638, n18277 );
nand U18361 ( n18277, n18278, n18223 );
nor U18362 ( n18278, n18271, n18256 );
not U18363 ( n18256, n18276 );
nand U18364 ( n18276, n18279, n10362 );
nor U18365 ( n18279, n19428, n19634 );
nor U18366 ( n18272, n18261, n18280 );
nor U18367 ( n18280, n19428, g35 );
and U18368 ( n18261, n18281, n19638 );
nor U18369 ( n18281, n10966, n18258 );
nand U18370 ( n1657, n18282, n18283 );
nand U18371 ( n18283, n18271, g35 );
not U18372 ( n18271, n18258 );
nand U18373 ( n18258, n18284, n19428 );
nor U18374 ( n18284, n19636, n10362 );
nor U18375 ( n18282, n18285, n18286 );
nor U18376 ( n18286, n10362, n18287 );
nand U18377 ( n18287, n18288, n19636 );
nor U18378 ( n18288, n19428, n18221 );
nor U18379 ( n18285, n19637, n18289 );
nor U18380 ( n18289, n10966, n18290 );
nand U18381 ( n18290, n18291, n18292 );
nand U18382 ( n18292, n18293, n10901 );
nor U18383 ( n18293, n18294, n10236 );
nand U18384 ( n18291, n19428, n10236 );
nand U18385 ( n1652, n18295, n18296 );
nand U18386 ( n18296, n18297, n19637 );
nor U18387 ( n18297, n18298, n18221 );
not U18388 ( n18221, n18223 );
nor U18389 ( n18223, n18294, n10986 );
nand U18390 ( n18294, n18209, n18206 );
nand U18391 ( n18206, n18299, n18300 );
and U18392 ( n18300, n18301, n19642 );
nor U18393 ( n18301, n19634, n19641 );
not U18394 ( n18299, n18302 );
nand U18395 ( n18209, n18302, n18303 );
and U18396 ( n18303, n18304, n19641 );
nor U18397 ( n18304, n19636, n19642 );
nand U18398 ( n18302, n18305, n18306 );
or U18399 ( n18306, n10583, n19564 );
nand U18400 ( n18305, n19564, n19429 );
nor U18401 ( n18295, n18307, n18308 );
nor U18402 ( n18308, n19636, g35 );
nor U18403 ( n18307, n10967, n18309 );
nand U18404 ( n18309, n18298, n10362 );
nor U18405 ( n18298, n10236, n10603 );
nand U18406 ( n1647, n18310, n18311 );
nand U18407 ( n18311, n11006, n10889 );
nand U18408 ( n18310, n18312, g35 );
nor U18409 ( n18312, n18313, g9497 );
nor U18410 ( n18313, n18314, n10603 );
nor U18411 ( n18314, n19635, n10889 );
nand U18412 ( n1638, n18315, n18316 );
nand U18413 ( n18316, g35, g25219 );
nand U18414 ( n18315, n11006, n10236 );
nand U18415 ( n1633, n18317, n18318 );
nand U18416 ( n18318, n11006, n10890 );
nand U18417 ( n18317, n18319, g35 );
nor U18418 ( n18319, n18320, g9553 );
nor U18419 ( n18320, n18321, n10236 );
nor U18420 ( n18321, n19633, n10890 );
nor U18421 ( n1624, n19654, n10986 );
nand U18422 ( n1619, n18322, n18323 );
nand U18423 ( n18323, n18324, n17982 );
nor U18424 ( n18322, n18325, n18326 );
nor U18425 ( n18326, n18327, n10986 );
nor U18426 ( n18327, n18328, n18329 );
nor U18427 ( n18329, n18330, n17968 );
nor U18428 ( n18328, n19441, g33959 );
nor U18429 ( n18325, n19632, g35 );
nand U18430 ( n1614, n18331, n18332 );
nand U18431 ( n18332, n17951, n10270 );
nor U18432 ( n18331, n18333, n18334 );
nor U18433 ( n18334, n19631, g35 );
nor U18434 ( n18333, n10967, n18335 );
nand U18435 ( n18335, n18324, n19632 );
nor U18436 ( n18324, n18330, n17937 );
nor U18437 ( n18330, n16557, n11111 );
nand U18438 ( n11111, n19588, n17214 );
not U18439 ( n17214, n11178 );
nand U18440 ( n16557, n18336, n13438 );
nor U18441 ( n18336, n19430, n10292 );
nor U18442 ( n1609, n19630, n18337 );
and U18443 ( n18337, g35, n18338 );
nand U18444 ( n1604, n18339, n18340 );
nand U18445 ( n18340, n11005, g25219 );
nand U18446 ( n18339, n18341, g35 );
nor U18447 ( n18341, n18338, n10691 );
nor U18448 ( n18338, n18342, n19629 );
nand U18449 ( n1599, n18343, n18344 );
or U18450 ( n18344, g35, n19431 );
nand U18451 ( n18343, n18345, g35 );
xnor U18452 ( n18345, n18342, g25219 );
nand U18453 ( n18342, n18346, n18347 );
nor U18454 ( n18347, n19432, n19433 );
nor U18455 ( n18346, n19627, n19628 );
nor U18456 ( n1558, n18348, n18349 );
nand U18457 ( n18349, n18350, n19434 );
nor U18458 ( n18350, n18351, n18352 );
nor U18459 ( n18352, n19627, g12238 );
nor U18460 ( n18351, n19432, g14662 );
nand U18461 ( n18348, n18353, n19435 );
nor U18462 ( n18353, n10967, g17519 );
nand U18463 ( n1553, n18354, n18355 );
nand U18464 ( n18355, n18356, n10550 );
nand U18465 ( n18356, g35, n18357 );
nand U18466 ( n18357, n18358, n18359 );
nor U18467 ( n18354, n18360, n18361 );
nor U18468 ( n18361, n18362, n18363 );
or U18469 ( n18363, n18358, n19626 );
nand U18470 ( n1548, n18364, n18365 );
nand U18471 ( n18365, n18366, n18358 );
nor U18472 ( n18358, n18367, n18368 );
nor U18473 ( n18366, n18369, n10986 );
nor U18474 ( n18369, n18370, n10550 );
nor U18475 ( n18370, n18371, n16952 );
nor U18476 ( n18371, n18372, n18373 );
nand U18477 ( n18373, n18374, n18375 );
or U18478 ( n18375, n16999, n19754 );
not U18479 ( n16999, n17012 );
nor U18480 ( n17012, n10261, n19436 );
nand U18481 ( n18374, n19754, n16982 );
nor U18482 ( n16982, n10261, n10612 );
nand U18483 ( n18372, n18376, n18377 );
nand U18484 ( n18377, n16984, n10689 );
nor U18485 ( n16984, n19436, n19756 );
nand U18486 ( n18376, n19755, n17010 );
nor U18487 ( n17010, n10612, n19756 );
nand U18488 ( n18364, n16968, n10550 );
nor U18489 ( n16968, n10967, n16958 );
not U18490 ( n16958, n16952 );
nand U18491 ( n16952, n10459, n18378 );
nand U18492 ( n18378, n18379, n18380 );
nand U18493 ( n1543, n18381, n18382 );
nand U18494 ( n18382, n18383, n10551 );
nand U18495 ( n18383, g35, n18384 );
nand U18496 ( n18384, n18385, n18359 );
nor U18497 ( n18381, n18360, n18386 );
nor U18498 ( n18386, n18362, n18387 );
or U18499 ( n18387, n18385, n19625 );
nand U18500 ( n1538, n18388, n18389 );
nand U18501 ( n18389, n18390, n18385 );
nor U18502 ( n18385, n18391, n18368 );
nor U18503 ( n18390, n18392, n10986 );
nor U18504 ( n18392, n18393, n10551 );
nor U18505 ( n18393, n18394, n17280 );
nor U18506 ( n18394, n18395, n18396 );
nand U18507 ( n18396, n18397, n18398 );
or U18508 ( n18398, n17327, n19717 );
not U18509 ( n17327, n17340 );
nor U18510 ( n17340, n10262, n19437 );
nand U18511 ( n18397, n19717, n17310 );
nor U18512 ( n17310, n10262, n10613 );
nand U18513 ( n18395, n18399, n18400 );
nand U18514 ( n18400, n17312, n10690 );
nor U18515 ( n17312, n19437, n19719 );
nand U18516 ( n18399, n19718, n17338 );
nor U18517 ( n17338, n10613, n19719 );
nand U18518 ( n18388, n17296, n10551 );
nor U18519 ( n17296, n10967, n17286 );
not U18520 ( n17286, n17280 );
nand U18521 ( n17280, n10290, n18401 );
nand U18522 ( n18401, n18402, n18380 );
nand U18523 ( n1533, n18403, n18404 );
nand U18524 ( n18404, n18405, n10552 );
nand U18525 ( n18405, g35, n18406 );
nand U18526 ( n18406, n18407, n18359 );
nor U18527 ( n18403, n18360, n18408 );
nor U18528 ( n18408, n18362, n18409 );
or U18529 ( n18409, n18407, n19624 );
nand U18530 ( n1528, n18410, n18411 );
nand U18531 ( n18411, n18412, n18407 );
and U18532 ( n18407, n18413, n19622 );
nor U18533 ( n18413, n18368, n10444 );
nor U18534 ( n18412, n18414, n10987 );
nor U18535 ( n18414, n18415, n10552 );
nor U18536 ( n18415, n18416, n18417 );
nand U18537 ( n18417, n18418, n17615 );
nor U18538 ( n18418, n18419, n18420 );
nor U18539 ( n18420, n11118, n10739 );
not U18540 ( n11118, n17640 );
nor U18541 ( n17640, n19438, n19683 );
nor U18542 ( n18419, n19682, n17642 );
not U18543 ( n17642, n17666 );
nor U18544 ( n17666, n10471, n19683 );
nand U18545 ( n18416, n18421, n18422 );
or U18546 ( n18422, n17670, n19681 );
not U18547 ( n17670, n17638 );
nor U18548 ( n17638, n10242, n10471 );
nand U18549 ( n18421, n19681, n17668 );
nor U18550 ( n17668, n10242, n19438 );
nand U18551 ( n18410, n17624, n10552 );
nor U18552 ( n17624, n10968, n17615 );
not U18553 ( n17615, n17609 );
nand U18554 ( n17609, n10811, n18423 );
nand U18555 ( n18423, n18424, n18380 );
nand U18556 ( n1523, n18425, n18426 );
nand U18557 ( n18426, n18427, n10553 );
nand U18558 ( n18427, g35, n18428 );
nand U18559 ( n18428, n18429, n18359 );
nor U18560 ( n18425, n18360, n18430 );
nor U18561 ( n18430, n18362, n18431 );
or U18562 ( n18431, n18429, n19444 );
nand U18563 ( n18362, g35, n18359 );
nor U18564 ( n18360, n18432, n18359 );
nand U18565 ( n18359, n18433, n19440 );
nor U18566 ( n18433, n11183, n10891 );
or U18567 ( n18432, n19439, n11024 );
nand U18568 ( n1518, n18434, n18435 );
nand U18569 ( n18435, n17951, n10553 );
nor U18570 ( n17951, n10968, g33959 );
nand U18571 ( n18434, n18436, g35 );
nor U18572 ( n18436, n18437, n11179 );
not U18573 ( n11179, n18429 );
nor U18574 ( n18429, n18368, n18438 );
nor U18575 ( n18437, n18439, n10553 );
nor U18576 ( n18439, n18440, n17937 );
not U18577 ( n17937, g33959 );
nor U18578 ( n18440, n18441, n18442 );
nand U18579 ( n18442, n18443, n18444 );
nand U18580 ( n18444, g31860, n10691 );
nand U18581 ( n18443, n19631, n17982 );
nor U18582 ( n17982, n10604, n19632 );
nand U18583 ( n18441, n18445, n18446 );
or U18584 ( n18446, n17968, n19630 );
not U18585 ( n17968, n17993 );
nor U18586 ( n17993, n10270, n19441 );
nand U18587 ( n18445, n19630, n17965 );
nor U18588 ( n17965, n10604, n10270 );
nand U18589 ( n1513, n18447, n18448 );
nor U18590 ( n18448, n18449, n18450 );
nor U18591 ( n18450, n10968, n18451 );
nand U18592 ( n18451, n18452, n18453 );
nor U18593 ( n18449, n19622, g35 );
nor U18594 ( n18447, n18454, n18455 );
nor U18595 ( n18455, n19623, n18456 );
nor U18596 ( n18454, n18391, n18457 );
nand U18597 ( n1508, n18458, n18459 );
nand U18598 ( n18459, n11005, n10309 );
nor U18599 ( n18458, n18460, n18461 );
nor U18600 ( n18461, n10406, n18457 );
nand U18601 ( n18457, n18462, n18463 );
nor U18602 ( n18462, n19621, n18464 );
nor U18603 ( n18460, n19622, n18456 );
nand U18604 ( n1503, n18465, n18466 );
nand U18605 ( n18466, n18467, n10450 );
nand U18606 ( n18467, g35, n18468 );
nand U18607 ( n18465, n18469, n10309 );
nand U18608 ( n1498, n18470, n18471 );
nand U18609 ( n18471, n11005, n10392 );
nor U18610 ( n18470, n18472, n18473 );
nor U18611 ( n18473, n10450, n18468 );
nand U18612 ( n18468, n18474, n18463 );
nor U18613 ( n18472, n19620, n18475 );
or U18614 ( n18475, n18456, n18463 );
nand U18615 ( n1493, n18476, n18477 );
nand U18616 ( n18477, n18478, n18469 );
not U18617 ( n18469, n18456 );
nand U18618 ( n18456, n18474, g35 );
and U18619 ( n18474, n18453, n18479 );
nand U18620 ( n18479, n18463, n10309 );
and U18621 ( n18463, n11177, n10392 );
xnor U18622 ( n18478, n19445, n11177 );
nand U18623 ( n18476, n11005, n10891 );
nor U18624 ( n1476, n19566, n10987 );
nand U18625 ( n1471, n17841, n18480 );
or U18626 ( n18480, g35, n19442 );
nand U18627 ( n17841, g35, n18481 );
nand U18628 ( n18481, n18482, n18483 );
nor U18629 ( n18483, n18484, n18485 );
nor U18630 ( n18485, n19613, n10892 );
nor U18631 ( n18484, n19614, n19746 );
nor U18632 ( n18482, n18486, n18487 );
nand U18633 ( n18487, n18488, n18489 );
nand U18634 ( n18489, n19446, n10459 );
nand U18635 ( n18488, n18490, n19615 );
nor U18636 ( n18490, n18491, n18492 );
nor U18637 ( n18491, n18493, n18494 );
nand U18638 ( n18494, n18495, n18496 );
nand U18639 ( n18496, n18497, n10392 );
and U18640 ( n18497, new_g34657_, n19621 );
nand U18641 ( n18495, n18498, n19445 );
nor U18642 ( n18498, n18499, n10450 );
nand U18643 ( n18499, n18500, n18501 );
nand U18644 ( n18501, n18502, n10309 );
xor U18645 ( n18502, new_g34657_, n18503 );
nor U18646 ( n18503, n18504, n18505 );
nand U18647 ( n18505, n18506, n18507 );
nand U18648 ( n18507, n18452, n10367 );
or U18649 ( n18506, n18391, n19479 );
nand U18650 ( n18504, n18508, n18509 );
nand U18651 ( n18509, n18510, n19622 );
nor U18652 ( n18510, n19470, n10444 );
nand U18653 ( n18508, n18511, n10511 );
nand U18654 ( new_g34657_, n18512, n18513 );
nor U18655 ( n18513, n18514, n18379 );
nor U18656 ( n18379, n19626, n18438 );
nor U18657 ( n18512, n18402, n18424 );
nor U18658 ( n18424, n19624, n18391 );
nor U18659 ( n18402, n19625, n18367 );
nand U18660 ( n18500, n18515, n19621 );
nor U18661 ( n18515, n18516, n18517 );
nand U18662 ( n18517, n18367, n18391 );
nand U18663 ( n18391, n19623, n10406 );
not U18664 ( n18367, n18452 );
nor U18665 ( n18452, n10406, n19623 );
nor U18666 ( n18516, n10702, n18438 );
not U18667 ( n18438, n18511 );
nor U18668 ( n18511, n19623, n19622 );
not U18669 ( n18493, n18368 );
nand U18670 ( n18368, n18518, n19620 );
nor U18671 ( n18518, n19445, n19621 );
nor U18672 ( n18486, n19443, n19612 );
nand U18673 ( n1451, n18519, n18520 );
nand U18674 ( n18520, g35, n10702 );
nand U18675 ( n18519, n11005, n10510 );
nand U18676 ( n1446, n18521, n18522 );
nand U18677 ( n18522, g35, n10510 );
nand U18678 ( n18521, n11005, n10515 );
nand U18679 ( n1441, n18523, n18524 );
nand U18680 ( n18524, g35, n10515 );
nand U18681 ( n18523, n11005, n10367 );
nand U18682 ( n1436, n18525, n18526 );
nand U18683 ( n18526, g35, n10367 );
nand U18684 ( n18525, n11004, n10511 );
nor U18685 ( n1431, n19490, n10987 );
nand U18686 ( n1426, n18527, n18528 );
nand U18687 ( n18528, n18529, n10919 );
nand U18688 ( n18529, g35, n18530 );
nand U18689 ( n18530, n18531, n18532 );
nand U18690 ( n18527, n18533, n10768 );
nand U18691 ( n1421, n18534, n18535 );
nand U18692 ( n18535, n18536, n18533 );
xnor U18693 ( n18536, n18532, n19618 );
nand U18694 ( n18534, n11004, n10609 );
nand U18695 ( n1416, n18537, n18538 );
nand U18696 ( n18538, n11004, n10288 );
nor U18697 ( n18537, n18539, n18540 );
nor U18698 ( n18540, n10609, n18541 );
nand U18699 ( n18541, n18531, n18542 );
nor U18700 ( n18539, n19617, n18543 );
nand U18701 ( n18543, n18533, n18544 );
not U18702 ( n18533, n18545 );
nand U18703 ( n1411, n18546, n18547 );
nand U18704 ( n18547, n18548, n10459 );
nand U18705 ( n18548, g35, n18549 );
nand U18706 ( n18549, n19616, n18531 );
nand U18707 ( n18546, n18550, n19615 );
nor U18708 ( n18550, n19616, n18545 );
nor U18709 ( n1406, n19614, n18551 );
nor U18710 ( n1401, n19613, n18551 );
nor U18711 ( n1396, n19612, n18551 );
nor U18712 ( n18551, n18453, n10988 );
nor U18713 ( n1391, n18492, n18545 );
nand U18714 ( n18545, n18531, g35 );
nor U18715 ( n18531, n18464, n11177 );
nor U18716 ( n11177, n18552, n19447 );
not U18717 ( n18552, n18532 );
nor U18718 ( n18532, n18544, n19617 );
not U18719 ( n18544, n18542 );
nor U18720 ( n18542, n19615, n19616 );
not U18721 ( n18464, n18453 );
nand U18722 ( n18453, n18553, n13438 );
nor U18723 ( n18553, n19499, n11178 );
nand U18724 ( n18492, n18554, n19612 );
nor U18725 ( n18554, n10290, n10811 );
not U18726 ( n139, n14483 );
nand U18727 ( n14483, g35, g64 );
nand U18728 ( n1386, n18555, n18556 );
nand U18729 ( n18556, n18557, n10554 );
nand U18730 ( n18557, g35, n18558 );
nand U18731 ( n18558, n18559, n18560 );
nor U18732 ( n18555, n18561, n18562 );
nor U18733 ( n18562, n18563, n18564 );
or U18734 ( n18564, n18559, n19611 );
nand U18735 ( n1381, n18565, n18566 );
nand U18736 ( n18566, n18567, n18559 );
nor U18737 ( n18559, n18568, n18569 );
nor U18738 ( n18567, n18570, n10988 );
nor U18739 ( n18570, n18571, n10554 );
nor U18740 ( n18571, n18572, n15637 );
nor U18741 ( n18572, n18573, n18574 );
nand U18742 ( n18574, n18575, n18576 );
or U18743 ( n18576, n15684, n19900 );
not U18744 ( n15684, n15697 );
nor U18745 ( n15697, n10263, n19448 );
nand U18746 ( n18575, n19900, n15667 );
nor U18747 ( n15667, n10263, n10614 );
nand U18748 ( n18573, n18577, n18578 );
nand U18749 ( n18578, n15669, n10692 );
nor U18750 ( n15669, n19448, n19902 );
nand U18751 ( n18577, n19901, n15695 );
nor U18752 ( n15695, n10614, n19902 );
nand U18753 ( n18565, n15653, n10554 );
nor U18754 ( n15653, n10969, n15643 );
not U18755 ( n15643, n15637 );
nand U18756 ( n15637, n10460, n18579 );
nand U18757 ( n18579, n18580, n18581 );
nand U18758 ( n1376, n18582, n18583 );
nand U18759 ( n18583, n18584, n10555 );
nand U18760 ( n18584, g35, n18585 );
nand U18761 ( n18585, n18586, n18560 );
nor U18762 ( n18582, n18561, n18587 );
nor U18763 ( n18587, n18563, n18588 );
or U18764 ( n18588, n18586, n19610 );
nand U18765 ( n1371, n18589, n18590 );
nand U18766 ( n18590, n18591, n18586 );
nor U18767 ( n18586, n18592, n18569 );
nor U18768 ( n18591, n18593, n10988 );
nor U18769 ( n18593, n18594, n10555 );
nor U18770 ( n18594, n18595, n15968 );
nor U18771 ( n18595, n18596, n18597 );
nand U18772 ( n18597, n18598, n18599 );
or U18773 ( n18599, n16015, n19864 );
not U18774 ( n16015, n16028 );
nor U18775 ( n16028, n10264, n19449 );
nand U18776 ( n18598, n19864, n15998 );
nor U18777 ( n15998, n10264, n10615 );
nand U18778 ( n18596, n18600, n18601 );
nand U18779 ( n18601, n16000, n10693 );
nor U18780 ( n16000, n19449, n19866 );
nand U18781 ( n18600, n19865, n16026 );
nor U18782 ( n16026, n10615, n19866 );
nand U18783 ( n18589, n15984, n10555 );
nor U18784 ( n15984, n10969, n15974 );
not U18785 ( n15974, n15968 );
nand U18786 ( n15968, n10289, n18602 );
nand U18787 ( n18602, n18603, n18581 );
not U18788 ( n137, n15049 );
nand U18789 ( n15049, n18604, n18605 );
nor U18790 ( n18605, n15053, n10939 );
nand U18791 ( n15053, n19569, g54 );
nor U18792 ( n18604, g57, g53 );
nand U18793 ( n1366, n18606, n18607 );
nand U18794 ( n18607, n18608, n10556 );
nand U18795 ( n18608, g35, n18609 );
nand U18796 ( n18609, n18610, n18560 );
nor U18797 ( n18606, n18561, n18611 );
nor U18798 ( n18611, n18563, n18612 );
or U18799 ( n18612, n18610, n19609 );
nand U18800 ( n1361, n18613, n18614 );
nand U18801 ( n18614, n18615, n18610 );
and U18802 ( n18610, n18616, n19607 );
nor U18803 ( n18616, n18569, n10443 );
nor U18804 ( n18615, n18617, n10988 );
nor U18805 ( n18617, n18618, n10556 );
nor U18806 ( n18618, n18619, n18620 );
nand U18807 ( n18620, n18621, n16304 );
nor U18808 ( n18621, n18622, n18623 );
nor U18809 ( n18623, n11119, n10740 );
not U18810 ( n11119, n16329 );
nor U18811 ( n16329, n19830, n19829 );
nor U18812 ( n18622, n19828, n16331 );
not U18813 ( n16331, n16355 );
nor U18814 ( n16355, n10472, n19829 );
nand U18815 ( n18619, n18624, n18625 );
or U18816 ( n18625, n16359, n19827 );
not U18817 ( n16359, n16327 );
nor U18818 ( n16327, n10243, n10472 );
nand U18819 ( n18624, n19827, n16357 );
nor U18820 ( n16357, n10243, n19830 );
nand U18821 ( n18613, n16313, n10556 );
nor U18822 ( n16313, n10969, n16304 );
not U18823 ( n16304, n16298 );
nand U18824 ( n16298, n10812, n18626 );
nand U18825 ( n18626, n18627, n18581 );
nand U18826 ( n1356, n18628, n18629 );
nand U18827 ( n18629, n18630, n10557 );
nand U18828 ( n18630, g35, n18631 );
nand U18829 ( n18631, n18632, n18560 );
nor U18830 ( n18628, n18561, n18633 );
nor U18831 ( n18633, n18563, n18634 );
or U18832 ( n18634, n18632, n19456 );
nand U18833 ( n18563, g35, n18560 );
nor U18834 ( n18561, n18635, n18560 );
nand U18835 ( n18560, n18636, n19451 );
nor U18836 ( n18636, n11183, n10893 );
or U18837 ( n18635, n19450, n11024 );
nand U18838 ( n1351, n18637, n18638 );
nand U18839 ( n18638, n16640, n10557 );
nor U18840 ( n16640, n10969, n16631 );
nand U18841 ( n18637, n18639, g35 );
nor U18842 ( n18639, n18640, n11175 );
not U18843 ( n11175, n18632 );
nor U18844 ( n18632, n18569, n18641 );
nor U18845 ( n18640, n18642, n10557 );
nor U18846 ( n18642, n18643, n16625 );
not U18847 ( n16625, n16631 );
nor U18848 ( n16631, n19597, n18644 );
and U18849 ( n18644, n18645, n18581 );
and U18850 ( n18581, n18646, n18647 );
nor U18851 ( n18647, n19602, n18648 );
nand U18852 ( n18648, n10287, n10767 );
nor U18853 ( n18646, n10391, n18649 );
nand U18854 ( n18649, n19605, n10308 );
nor U18855 ( n18643, n18650, n18651 );
nand U18856 ( n18651, n18652, n18653 );
nand U18857 ( n18653, n16656, n10694 );
nor U18858 ( n16656, n19452, n19792 );
nand U18859 ( n18652, n19791, n16682 );
nor U18860 ( n16682, n10616, n19792 );
nand U18861 ( n18650, n18654, n18655 );
or U18862 ( n18655, n16671, n19790 );
not U18863 ( n16671, n16684 );
nor U18864 ( n16684, n10265, n19452 );
nand U18865 ( n18654, n19790, n16654 );
nor U18866 ( n16654, n10265, n10616 );
nand U18867 ( n1346, n18656, n18657 );
nor U18868 ( n18657, n18658, n18659 );
nor U18869 ( n18659, n10969, n18660 );
nand U18870 ( n18660, n18661, n18662 );
nor U18871 ( n18658, n19607, g35 );
nor U18872 ( n18656, n18663, n18664 );
nor U18873 ( n18664, n19608, n18665 );
nor U18874 ( n18663, n18592, n18666 );
nand U18875 ( n1341, n18667, n18668 );
nand U18876 ( n18668, n11004, n10308 );
nor U18877 ( n18667, n18669, n18670 );
nor U18878 ( n18670, n10407, n18666 );
nand U18879 ( n18666, n18671, n18672 );
nor U18880 ( n18671, n19606, n18673 );
nor U18881 ( n18669, n19607, n18665 );
nand U18882 ( n1336, n18674, n18675 );
nand U18883 ( n18675, n18676, n10451 );
nand U18884 ( n18676, g35, n18677 );
nand U18885 ( n18674, n18678, n10308 );
nand U18886 ( n1331, n18679, n18680 );
nand U18887 ( n18680, n11004, n10391 );
nor U18888 ( n18679, n18681, n18682 );
nor U18889 ( n18682, n10451, n18677 );
nand U18890 ( n18677, n18683, n18672 );
nor U18891 ( n18681, n19605, n18684 );
or U18892 ( n18684, n18665, n18672 );
nand U18893 ( n1326, n18685, n18686 );
nand U18894 ( n18686, n18687, n18678 );
not U18895 ( n18678, n18665 );
nand U18896 ( n18665, n18683, g35 );
and U18897 ( n18683, n18662, n18688 );
nand U18898 ( n18688, n18672, n10308 );
and U18899 ( n18672, n11173, n10391 );
xnor U18900 ( n18687, n19457, n11173 );
nand U18901 ( n18685, n11004, n10893 );
nand U18902 ( n1304, n18131, n18689 );
or U18903 ( n18689, g35, n19453 );
nand U18904 ( n18131, g35, n18690 );
nand U18905 ( n18690, n18691, n18692 );
nor U18906 ( n18692, n18693, n18694 );
nor U18907 ( n18694, n19597, n19819 );
nor U18908 ( n18693, n19598, n10894 );
nor U18909 ( n18691, n18695, n18696 );
nand U18910 ( n18696, n18697, n18698 );
nand U18911 ( n18698, n19455, n10460 );
nand U18912 ( n18697, n18699, n19600 );
nor U18913 ( n18699, n18700, n18701 );
nor U18914 ( n18700, n18702, n18703 );
nand U18915 ( n18703, n18704, n18705 );
nand U18916 ( n18705, n18706, n10391 );
and U18917 ( n18706, new_g34649_, n19606 );
nand U18918 ( n18704, n18707, n19457 );
nor U18919 ( n18707, n18708, n10451 );
nand U18920 ( n18708, n18709, n18710 );
nand U18921 ( n18710, n18711, n10308 );
xor U18922 ( n18711, new_g34649_, n18712 );
nor U18923 ( n18712, n18713, n18714 );
nand U18924 ( n18714, n18715, n18716 );
nand U18925 ( n18716, n18661, n10368 );
or U18926 ( n18715, n18592, n19480 );
nand U18927 ( n18713, n18717, n18718 );
nand U18928 ( n18718, n18719, n19607 );
nor U18929 ( n18719, n19471, n10443 );
nand U18930 ( n18717, n18720, n10513 );
nand U18931 ( new_g34649_, n18721, n18722 );
nor U18932 ( n18722, n18645, n18580 );
nor U18933 ( n18580, n19611, n18641 );
and U18934 ( n18645, n18723, n19607 );
nor U18935 ( n18723, n19456, n10443 );
nor U18936 ( n18721, n18603, n18627 );
nor U18937 ( n18627, n19609, n18592 );
nor U18938 ( n18603, n19610, n18568 );
nand U18939 ( n18709, n18724, n19606 );
nor U18940 ( n18724, n18725, n18726 );
nand U18941 ( n18726, n18568, n18592 );
nand U18942 ( n18592, n19608, n10407 );
not U18943 ( n18568, n18661 );
nor U18944 ( n18661, n10407, n19608 );
nor U18945 ( n18725, n10703, n18641 );
not U18946 ( n18641, n18720 );
nor U18947 ( n18720, n19608, n19607 );
not U18948 ( n18702, n18569 );
nand U18949 ( n18569, n18727, n19605 );
nor U18950 ( n18727, n19457, n19606 );
nor U18951 ( n18695, n19454, n19599 );
nand U18952 ( n1284, n18728, n18729 );
nand U18953 ( n18729, g35, n10703 );
nand U18954 ( n18728, n11004, n10512 );
nand U18955 ( n1279, n18730, n18731 );
nand U18956 ( n18731, g35, n10512 );
nand U18957 ( n18730, n11004, n10516 );
nand U18958 ( n1274, n18732, n18733 );
nand U18959 ( n18733, g35, n10516 );
nand U18960 ( n18732, n11003, n10368 );
nand U18961 ( n1269, n18734, n18735 );
nand U18962 ( n18735, g35, n10368 );
nand U18963 ( n18734, n11003, n10513 );
nor U18964 ( n1264, n19494, n10988 );
nand U18965 ( n1259, n18736, n18737 );
nand U18966 ( n18737, n18738, n10920 );
nand U18967 ( n18738, g35, n18739 );
nand U18968 ( n18739, n18740, n18741 );
nand U18969 ( n18736, n18742, n10767 );
nand U18970 ( n1254, n18743, n18744 );
nand U18971 ( n18744, n18745, n18742 );
xnor U18972 ( n18745, n18741, n19603 );
nand U18973 ( n18743, n11003, n10610 );
nand U18974 ( n1249, n18746, n18747 );
nand U18975 ( n18747, n11003, n10287 );
nor U18976 ( n18746, n18748, n18749 );
nor U18977 ( n18749, n10610, n18750 );
nand U18978 ( n18750, n18740, n18751 );
nor U18979 ( n18748, n19602, n18752 );
nand U18980 ( n18752, n18742, n18753 );
not U18981 ( n18742, n18754 );
nand U18982 ( n1244, n18755, n18756 );
nand U18983 ( n18756, n18757, n10460 );
nand U18984 ( n18757, g35, n18758 );
nand U18985 ( n18758, n19601, n18740 );
nand U18986 ( n18755, n18759, n19600 );
nor U18987 ( n18759, n19601, n18754 );
nor U18988 ( n1239, n19599, n18760 );
nor U18989 ( n1234, n19598, n18760 );
nor U18990 ( n1229, n19597, n18760 );
nor U18991 ( n18760, n18662, n10989 );
nor U18992 ( n1224, n18701, n18754 );
nand U18993 ( n18754, n18740, g35 );
nor U18994 ( n18740, n18673, n11173 );
nor U18995 ( n11173, n18761, n19500 );
not U18996 ( n18761, n18741 );
nor U18997 ( n18741, n18753, n19602 );
not U18998 ( n18753, n18751 );
nor U18999 ( n18751, n19600, n19601 );
not U19000 ( n18673, n18662 );
nand U19001 ( n18662, n18762, n13438 );
nor U19002 ( n18762, n19499, n11174 );
nand U19003 ( n11174, n18763, n18764 );
nor U19004 ( n18763, n19590, n18765 );
nand U19005 ( n18701, n18766, n19597 );
nor U19006 ( n18766, n10289, n10812 );
nand U19007 ( n1219, n18767, n18768 );
nand U19008 ( n18768, n11003, n10895 );
nand U19009 ( n18767, n18769, g35 );
nand U19010 ( n18769, n18770, n18771 );
nand U19011 ( n18771, n18772, n10292 );
nand U19012 ( n18772, n18773, n18774 );
nand U19013 ( n18774, n10223, n10302 );
nand U19014 ( n18773, n19587, n18775 );
nand U19015 ( n18770, n18776, n19589 );
nand U19016 ( n18776, n18777, n18778 );
nand U19017 ( n18778, n19588, n18779 );
nand U19018 ( n18779, n18780, n19587 );
nor U19019 ( n18780, n18781, n18782 );
nor U19020 ( n18782, n19592, n18783 );
nand U19021 ( n18783, n19591, n10346 );
nor U19022 ( n18781, n18784, n10351 );
nor U19023 ( n18784, n11304, n18785 );
nand U19024 ( n18785, n18786, n18787 );
nand U19025 ( n18787, n19501, n10227 );
nand U19026 ( n18786, n18788, n19591 );
nor U19027 ( n18788, n19502, n10517 );
not U19028 ( n11304, n11266 );
nand U19029 ( n18777, n18789, n10223 );
nor U19030 ( n18789, n11327, n10302 );
nor U19031 ( n1214, n18790, n10989 );
nor U19032 ( n18790, n18791, n18792 );
nand U19033 ( n18792, n18793, n18775 );
not U19034 ( n18775, n11327 );
nand U19035 ( n11327, n19503, n18794 );
nand U19036 ( n18794, n18795, n18796 );
nand U19037 ( n18796, n18797, n18798 );
xnor U19038 ( n18798, n19595, n19593 );
nor U19039 ( n18797, n10478, n18799 );
xnor U19040 ( n18799, n10334, n19594 );
nor U19041 ( n18795, n18800, n18801 );
nor U19042 ( n18801, n10585, n18802 );
nand U19043 ( n18802, n19594, n10430 );
nor U19044 ( n18800, n19593, n18803 );
nand U19045 ( n18803, n18804, n19595 );
nor U19046 ( n18804, n19594, n10334 );
nand U19047 ( n18791, n18805, n10292 );
nor U19048 ( n18805, n19587, n19588 );
nand U19049 ( n1209, n18806, n18807 );
nand U19050 ( n18807, n18808, n10430 );
nand U19051 ( n18808, g35, n18809 );
nand U19052 ( n18806, n18810, n10478 );
nand U19053 ( n1204, n18811, n18812 );
nand U19054 ( n18812, n11003, n10334 );
nor U19055 ( n18811, n18813, n18814 );
nor U19056 ( n18814, n10430, n18809 );
nand U19057 ( n18809, n18815, n18816 );
not U19058 ( n18816, n18817 );
nor U19059 ( n18813, n19595, n18818 );
nand U19060 ( n18818, n18810, n18817 );
nand U19061 ( n18817, n18819, n10334 );
nand U19062 ( n1199, n18820, n18821 );
nand U19063 ( n18821, n18822, n18810 );
xnor U19064 ( n18822, n19504, n18819 );
nor U19065 ( n18819, n18823, n19594 );
nand U19066 ( n18820, n11003, n10584 );
nand U19067 ( n1194, n18824, n18825 );
nand U19068 ( n18825, n11003, n10585 );
nor U19069 ( n18824, n18826, n18827 );
nor U19070 ( n18827, n10584, n18828 );
nand U19071 ( n18828, n18815, n18829 );
nor U19072 ( n18826, n19594, n18830 );
nand U19073 ( n18830, n18810, n18823 );
not U19074 ( n18823, n18829 );
nand U19075 ( n1189, n18831, n18832 );
nand U19076 ( n18832, n18833, n18810 );
and U19077 ( n18810, n18815, g35 );
and U19078 ( n18815, n18834, n18835 );
nand U19079 ( n18835, n18829, n10478 );
nor U19080 ( n18829, n18836, n19593 );
xnor U19081 ( n18833, n19593, n18837 );
nand U19082 ( n18831, n11002, n10351 );
nand U19083 ( n1184, n18838, n18839 );
nand U19084 ( n18839, n18840, n18841 );
nand U19085 ( n18841, n18842, n18843 );
nand U19086 ( n18843, n18844, n10227 );
nand U19087 ( n18842, g35, n10351 );
nand U19088 ( n18838, n11002, n10227 );
nand U19089 ( n1179, n18845, n18846 );
nand U19090 ( n18846, n18840, n18847 );
nor U19091 ( n18847, n18848, n18849 );
nor U19092 ( n18849, n18844, n18850 );
nor U19093 ( n18850, n19591, n10989 );
and U19094 ( n18848, n10227, n18844 );
nor U19095 ( n18844, n18851, n19590 );
nor U19096 ( n18840, n18852, n18837 );
nand U19097 ( n18845, n11002, n10346 );
nor U19098 ( n1174, n18853, n18854 );
nand U19099 ( n18854, n18855, n18836 );
not U19100 ( n18836, n18837 );
nor U19101 ( n18837, n18856, n18851 );
nand U19102 ( n18856, n10227, n10351 );
xnor U19103 ( n18853, n19590, n18851 );
nand U19104 ( n18851, n18857, n10292 );
nand U19105 ( n1169, n18858, n18859 );
nand U19106 ( n18859, n18860, n18861 );
nor U19107 ( n18860, n19586, n10302 );
nand U19108 ( n18858, g29218, n10979 );
nand U19109 ( n1164, n18862, n18863 );
nand U19110 ( n18863, n18864, n18865 );
nor U19111 ( n18865, n18866, n18867 );
nand U19112 ( n18867, n19593, n19594 );
nand U19113 ( n18866, n19504, n10302 );
nor U19114 ( n18864, n18868, n18869 );
nand U19115 ( n18869, n18861, n18793 );
and U19116 ( n18861, n18870, n18871 );
nor U19117 ( n18871, n10346, n18872 );
nand U19118 ( n18872, n19591, n19592 );
nor U19119 ( n18870, n10971, n18873 );
nand U19120 ( n18873, n19589, n19588 );
nand U19121 ( n18868, n19596, n19595 );
nand U19122 ( n18862, n11002, n10292 );
nand U19123 ( n1159, n18874, n18875 );
nand U19124 ( n18875, n11002, n10223 );
nor U19125 ( n18874, n18876, n18877 );
nor U19126 ( n18877, n10292, n18878 );
nand U19127 ( n18878, n18857, n18834 );
nor U19128 ( n18876, n19589, n18879 );
nand U19129 ( n18879, n18855, n18880 );
not U19130 ( n18880, n18857 );
nor U19131 ( n18857, n18881, n19588 );
nand U19132 ( n1154, n18882, n18883 );
nand U19133 ( n18883, n18884, n18855 );
xnor U19134 ( n18884, n18881, n10223 );
nand U19135 ( n18881, n18885, n18886 );
nor U19136 ( n18885, n19587, n10593 );
nand U19137 ( n18882, n11002, n10302 );
nand U19138 ( n1149, n18887, n18888 );
or U19139 ( n18888, g35, n19586 );
nand U19140 ( n18887, g35, n18889 );
nand U19141 ( n18889, n18890, n18834 );
xnor U19142 ( n18890, n19587, n18891 );
nand U19143 ( n18891, n18886, n19582 );
nand U19144 ( n1144, n18892, n18893 );
nand U19145 ( n18893, n18894, n18793 );
and U19146 ( n18793, n18895, n19582 );
nor U19147 ( n18895, n19583, n19585 );
nand U19148 ( n18892, n11002, n10658 );
nand U19149 ( n1139, n18896, n18897 );
nand U19150 ( n18897, n11001, n10666 );
nor U19151 ( n18896, n18898, n18899 );
nor U19152 ( n18899, n10658, n18900 );
nand U19153 ( n18900, n18901, n18894 );
nor U19154 ( n18901, n19582, n18902 );
nor U19155 ( n18898, n19585, n18903 );
nor U19156 ( n18903, n18904, n40 );
nor U19157 ( n18904, n18905, n18906 );
nand U19158 ( n18906, g35, n18902 );
not U19159 ( n18902, n18886 );
nor U19160 ( n18886, n19583, n19584 );
nand U19161 ( n1134, n18907, n18908 );
nand U19162 ( n18908, n18909, n10666 );
nand U19163 ( n18909, n18910, n18911 );
nand U19164 ( n18911, n18912, n19583 );
nor U19165 ( n18912, n10971, n18905 );
nand U19166 ( n18907, n18913, n10601 );
nand U19167 ( n18913, g35, n18914 );
nand U19168 ( n18914, n18915, n19584 );
nor U19169 ( n18915, n19582, n18905 );
nand U19170 ( n1129, n18916, n18917 );
nand U19171 ( n18917, n18918, n10593 );
nand U19172 ( n18918, g35, n18919 );
nand U19173 ( n18919, n19583, n18894 );
not U19174 ( n18894, n18905 );
nand U19175 ( n18905, n19586, n18834 );
nand U19176 ( n18916, n40, n10601 );
not U19177 ( n40, n18910 );
nand U19178 ( n18910, n18920, n19582 );
and U19179 ( n18920, n18855, n19586 );
nor U19180 ( n18855, n10971, n18852 );
not U19181 ( n18852, n18834 );
nand U19182 ( n18834, g65, n18921 );
nand U19183 ( n18921, n11266, n13560 );
nor U19184 ( n11266, g72, g73 );
nand U19185 ( n1119, n18922, n18923 );
or U19186 ( n18923, g35, n19506 );
nand U19187 ( n18922, n18924, g35 );
nor U19188 ( n1110, n18925, n10991 );
xnor U19189 ( n18925, n19505, n18924 );
xor U19190 ( n18924, n19506, n19505 );
nand U19191 ( n1105, n18926, n18927 );
nand U19192 ( n18927, n10998, g4455 );
nand U19193 ( n1090, n18926, n18928 );
nand U19194 ( n18928, n10998, n10704 );
nand U19195 ( n18926, n18929, n18930 );
nand U19196 ( n18930, n19580, n18931 );
nand U19197 ( n18931, n19507, n18932 );
nand U19198 ( n1085, n13422, n18933 );
or U19199 ( n18933, g35, n19579 );
not U19200 ( n13422, n11572 );
nor U19201 ( n11572, n13560, n10993 );
not U19202 ( n13560, n13438 );
nor U19203 ( n13438, g113, n11183 );
not U19204 ( n11183, n11221 );
nand U19205 ( n11221, n19567, n18934 );
nand U19206 ( n18934, n10386, g99 );
nand U19207 ( n1080, n18935, n18936 );
nand U19208 ( n18936, n10997, n10514 );
nand U19209 ( n18935, n18937, g35 );
nand U19210 ( n18937, n18938, n18939 );
nand U19211 ( n18939, n18940, n18941 );
xnor U19212 ( n18940, n10592, n19579 );
nand U19213 ( n18938, n18942, n18932 );
nor U19214 ( n18942, n10704, n10251 );
nand U19215 ( n1075, n18943, n18944 );
or U19216 ( n18944, n18929, n19508 );
and U19217 ( n18929, g35, n18945 );
nand U19218 ( n18945, n18932, n10251 );
nand U19219 ( n18943, g35, n10558 );
nand U19220 ( n1070, n19578, n18946 );
nand U19221 ( n18946, n18947, n18948 );
nor U19222 ( n18947, n19509, n18941 );
nand U19223 ( n1061, n18949, n18950 );
nand U19224 ( n18950, n10997, n10558 );
nor U19225 ( n18949, n18951, n18952 );
nor U19226 ( n18952, n19577, n18953 );
nor U19227 ( n18951, n18941, n18954 );
nand U19228 ( n1052, n18955, n18956 );
nand U19229 ( n18956, n18957, n18932 );
not U19230 ( n18932, n18941 );
nand U19231 ( n18941, n18958, n18959 );
nor U19232 ( n18959, g7243, n18960 );
nand U19233 ( n18960, n19577, n19578 );
nor U19234 ( n18958, g7257, n10558 );
nand U19235 ( n18955, n18953, n10592 );
nand U19236 ( n1047, n18961, n18962 );
or U19237 ( n18962, g35, n19517 );
not U19238 ( n18961, n145 );
nor U19239 ( n145, n10972, n19512 );
nand U19240 ( n1042, n18963, n18964 );
nand U19241 ( n18964, n18965, n10906 );
nand U19242 ( n18965, g35, n10514 );
nand U19243 ( n18963, g35, n18966 );
nand U19244 ( n18966, n18967, n18968 );
nand U19245 ( n18968, n19511, n10514 );
xnor U19246 ( n18967, n19510, n19508 );
nand U19247 ( n1037, n18969, n18970 );
nand U19248 ( n18970, n18971, n10921 );
nand U19249 ( n18971, g35, n18972 );
nand U19250 ( n18972, n18973, n10251 );
nand U19251 ( n18969, g35, n10493 );
nand U19252 ( n1032, n19576, n18974 );
nand U19253 ( n18974, n18975, n18973 );
nor U19254 ( n18975, n19511, n18954 );
nand U19255 ( n1023, n18976, n18977 );
nand U19256 ( n18977, n10997, n10493 );
nor U19257 ( n18976, n18978, n18979 );
nor U19258 ( n18979, n19575, n18953 );
nor U19259 ( n18978, n18954, n18980 );
not U19260 ( n18954, n18948 );
nor U19261 ( n18948, n10251, n10992 );
nand U19262 ( n1014, n18981, n18982 );
nand U19263 ( n18982, n18957, n18973 );
not U19264 ( n18973, n18980 );
nand U19265 ( n18980, n18983, n18984 );
nor U19266 ( n18984, n10493, n18985 );
nand U19267 ( n18985, n19575, n19576 );
nor U19268 ( n18983, g7245, g7260 );
nor U19269 ( n18957, n19580, n10990 );
nand U19270 ( n18981, n18953, n10907 );
nand U19271 ( n18953, n19579, g35 );
xor U19272 ( n1004, n18986, n19513 );
nand U19273 ( n18986, g35, g10306 );
nor U19274 ( g34839, n19571, n18987 );
nor U19275 ( n18987, n11178, n10895 );
nand U19276 ( n11178, n18988, n18764 );
xnor U19277 ( n18764, n19592, n19563 );
nor U19278 ( n18988, n10346, n18765 );
xnor U19279 ( n18765, n10227, n19562 );
nor U19280 ( g33959, n19612, n18989 );
and U19281 ( n18989, n18514, n18380 );
and U19282 ( n18380, n18990, n18991 );
nor U19283 ( n18991, n19617, n18992 );
nand U19284 ( n18992, n10288, n10768 );
nor U19285 ( n18990, n10392, n18993 );
nand U19286 ( n18993, n19620, n10309 );
and U19287 ( n18514, n18994, n19622 );
nor U19288 ( n18994, n19444, n10444 );
nor U19289 ( g32185, n18995, n18996 );
nand U19290 ( n18996, n18997, n18998 );
nand U19291 ( n18998, n10562, n10281 );
nor U19292 ( n18997, n18999, n19000 );
nor U19293 ( n19000, n20226, n20232 );
nor U19294 ( n18999, n20227, n20233 );
nand U19295 ( n18995, n19001, n19002 );
nor U19296 ( n19002, n19003, n19004 );
nor U19297 ( n19004, n20223, n20230 );
nor U19298 ( n19003, n20224, n20231 );
nor U19299 ( n19001, n19005, n19006 );
nor U19300 ( n19006, n20221, n20228 );
nor U19301 ( n19005, n20222, n20229 );
nor U19302 ( g31860, n19441, n19632 );
nand U19303 ( g31793, n19007, n19008 );
nand U19304 ( n19008, n19009, n19010 );
nor U19305 ( n19009, n19011, n11475 );
and U19306 ( n19011, n16611, n16938 );
nand U19307 ( n19007, n11474, n19012 );
nand U19308 ( n19012, n19013, n19014 );
nand U19309 ( n19014, n19015, n19016 );
nand U19310 ( n19016, n19017, n19018 );
nand U19311 ( n19018, n19019, n19517 );
nor U19312 ( n19019, n19020, n10897 );
nor U19313 ( n19020, n19021, n19022 );
nor U19314 ( n19022, n16284, n10640 );
nor U19315 ( n19021, n19023, n10698 );
nor U19316 ( n19023, n19519, n19024 );
not U19317 ( n19015, n11475 );
nand U19318 ( n11475, n19025, n19026 );
nand U19319 ( n19026, g35, n19027 );
nand U19320 ( n19027, n19514, n19516 );
nand U19321 ( n19013, n19010, n19028 );
nand U19322 ( n19028, n19029, n19030 );
nand U19323 ( n19030, n19516, n19031 );
nand U19324 ( n19031, n17923, n10625 );
nand U19325 ( n19029, n19514, n19025 );
not U19326 ( n19025, n17923 );
nor U19327 ( n17923, n10972, n19515 );
not U19328 ( n19010, n11476 );
nand U19329 ( n11476, n19032, n19517 );
nor U19330 ( n19032, n19017, n10897 );
nand U19331 ( n19017, n19024, n19033 );
nand U19332 ( n19033, g35, n19034 );
nand U19333 ( n19034, n19519, n19520 );
not U19334 ( n19024, n16284 );
nor U19335 ( n16284, n10972, n19518 );
nor U19336 ( n11474, n16938, n16611 );
nor U19337 ( n16611, n10972, n19521 );
nor U19338 ( n16938, n10972, n19522 );
nand U19339 ( g28042, n19035, n19523 );
nor U19340 ( n19035, n10963, n10381 );
nand U19341 ( g28041, n19036, g35 );
nor U19342 ( n19036, n11419, n11418 );
nor U19343 ( n11418, n20033, n14165 );
not U19344 ( n14165, n14152 );
nand U19345 ( n14152, n20036, n20037 );
nor U19346 ( n11419, n20071, n13817 );
not U19347 ( n13817, n13804 );
nand U19348 ( n13804, n20074, n20075 );
nand U19349 ( g28030, n19037, n19038 );
nand U19350 ( n19038, n19039, n19040 );
nor U19351 ( n19040, n19041, n19042 );
nor U19352 ( n19041, n19043, n19044 );
nor U19353 ( n19044, n19045, n19046 );
nor U19354 ( n19045, n19047, n19048 );
nor U19355 ( n19048, n19049, n19050 );
not U19356 ( n19050, n19051 );
nor U19357 ( n19049, n19052, n19053 );
nor U19358 ( n19053, n19054, n19055 );
nor U19359 ( n19055, n19056, n10982 );
not U19360 ( n11226, g35 );
nor U19361 ( n19054, n19057, n19058 );
nor U19362 ( n19057, n10759, n10282 );
nand U19363 ( n19037, n19059, n19043 );
not U19364 ( n19043, n11469 );
nand U19365 ( n11469, n19047, n19051 );
nand U19366 ( n19051, g35, n19060 );
nand U19367 ( n19060, n19532, n19533 );
and U19368 ( n19047, n19052, n19056 );
nor U19369 ( n19056, n10279, n10896 );
and U19370 ( n19052, n19061, n19530 );
and U19371 ( n19061, n19058, n19531 );
nand U19372 ( n19058, g35, n19062 );
nand U19373 ( n19062, n19528, n19529 );
nor U19374 ( n19059, n19046, n19063 );
nor U19375 ( n19063, n19064, n19039 );
nor U19376 ( n19039, n11464, n11468 );
not U19377 ( n11468, n19065 );
not U19378 ( n11464, n19066 );
nor U19379 ( n19064, n19042, n19067 );
nor U19380 ( n19067, n19065, n19066 );
nand U19381 ( n19066, g35, n19068 );
nand U19382 ( n19068, n19526, n19527 );
nand U19383 ( n19065, g35, n19069 );
nand U19384 ( n19069, n19524, n19525 );
not U19385 ( n19042, n11467 );
nand U19386 ( n11467, g35, n19070 );
nand U19387 ( n19070, n19536, n19537 );
not U19388 ( n19046, n11466 );
nand U19389 ( n11466, g35, n19071 );
nand U19390 ( n19071, n19534, n19535 );
nand U19391 ( g26877, n11458, n11457 );
nand U19392 ( n11457, n19072, n19073 );
nor U19393 ( n19073, n19074, n19075 );
nand U19394 ( n19075, n20170, n20179 );
nand U19395 ( n19074, n20183, n20192 );
nor U19396 ( n19072, n19076, n19077 );
nand U19397 ( n19077, n20143, n20152 );
nand U19398 ( n19076, n20157, n20166 );
and U19399 ( n11458, g35, n19078 );
nand U19400 ( n19078, n19079, n19080 );
nor U19401 ( n19080, n19081, n19082 );
nand U19402 ( n19082, n20115, n20124 );
nand U19403 ( n19081, n20128, n20137 );
nor U19404 ( n19079, n19083, n19084 );
nand U19405 ( n19084, n20090, n20097 );
nand U19406 ( n19083, n20102, n20111 );
nand U19407 ( g26876, n19085, g35 );
and U19408 ( n19085, n11405, n11399 );
nand U19409 ( n11399, n19086, n19087 );
nor U19410 ( n19087, n19088, n19089 );
nand U19411 ( n19089, n19542, n19543 );
nand U19412 ( n19088, n19544, n19545 );
nor U19413 ( n19086, n19090, n19091 );
nand U19414 ( n19091, n19538, n19539 );
nand U19415 ( n19090, n19540, n19541 );
nand U19416 ( n11405, n19092, n19093 );
nor U19417 ( n19093, n19094, n19095 );
nand U19418 ( n19095, n19550, n19551 );
nand U19419 ( n19094, n19552, n19553 );
nor U19420 ( n19092, n19096, n19097 );
nand U19421 ( n19097, n19546, n19547 );
nand U19422 ( n19096, n19548, n19549 );
nand U19423 ( g26875, n11485, n11404 );
nand U19424 ( n11404, n19098, n19099 );
and U19425 ( n19099, n19557, n19556 );
and U19426 ( n19098, n19555, n19554 );
not U19427 ( n11485, n11401 );
nand U19428 ( n11401, g35, n19100 );
nand U19429 ( n19100, n19101, n19102 );
and U19430 ( n19102, n19561, n19560 );
and U19431 ( n19101, n19559, n19558 );
endmodule

