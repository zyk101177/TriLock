
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule


module s35932_ori ( clk, reset, DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27,
DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22, DATA_0_21,
DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15,
DATA_0_14, DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9,
DATA_0_8, DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2,
DATA_0_1, DATA_0_0, RESET, TM1, TM0, DATA_9_31, DATA_9_30, DATA_9_29,
DATA_9_28, DATA_9_27, DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23,
DATA_9_22, DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17,
DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12, DATA_9_11,
DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4,
DATA_9_3, DATA_9_2, DATA_9_1, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1,
CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11,
CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21,
CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26,
CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31,
CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4,
CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9,
CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14,
CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19,
CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24,
CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29,
CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2,
CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7,
CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12,
CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17,
CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22,
CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27,
CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0,
CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5,
CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10,
CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15,
CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20,
CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25,
CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30,
CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3,
CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8,
CRC_OUT_5_9, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13,
CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18,
CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
CRC_OUT_5_29, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1,
CRC_OUT_4_2, CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11,
CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21,
CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26,
CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31,
CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4,
CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9,
CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14,
CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19,
CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24,
CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29,
CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2,
CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7,
CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12,
CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17,
CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22,
CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27,
CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0,
CRC_OUT_1_1, CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5,
CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10,
CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15,
CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20,
CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25,
CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30,
CRC_OUT_1_31 );
input clk, reset, DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27, DATA_0_26,
DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20,
DATA_0_19, DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14,
DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8,
DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2, DATA_0_1,
DATA_0_0, RESET, TM1, TM0;
output DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27, DATA_9_26,
DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22, DATA_9_21, DATA_9_20,
DATA_9_19, DATA_9_18, DATA_9_17, DATA_9_16, DATA_9_15, DATA_9_14,
DATA_9_13, DATA_9_12, DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8,
DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2, DATA_9_1,
DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3,
CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8,
CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13,
CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18,
CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23,
CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28,
CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1,
CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6,
CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10, CRC_OUT_8_11,
CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16,
CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21,
CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26,
CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30, CRC_OUT_8_31,
CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3, CRC_OUT_7_4,
CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9,
CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14,
CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19,
CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2,
CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22,
CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27,
CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0,
CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5,
CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10,
CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15,
CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_20,
CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25,
CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30,
CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2, CRC_OUT_4_3,
CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8,
CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13,
CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18,
CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23,
CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28,
CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0, CRC_OUT_3_1,
CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6,
CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10, CRC_OUT_3_11,
CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16,
CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21,
CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26,
CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30, CRC_OUT_3_31,
CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4,
CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9,
CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14,
CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19,
CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2,
CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22,
CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27,
CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31;
wire WX485, WX837, WX839, WX841, WX843, WX845, WX847, WX849, WX851, WX853,
WX855, WX857, WX859, WX861, WX863, WX865, WX867, WX869, WX871, WX873,
WX875, WX877, WX879, WX881, WX883, WX885, WX887, WX889, WX891, WX893,
WX895, WX897, WX899, WX1778, WX2130, WX2132, WX2134, WX2136, WX2138,
WX2140, WX2142, WX2144, WX2146, WX2148, WX2150, WX2152, WX2154,
WX2156, WX2158, WX2160, WX2162, WX2164, WX2166, WX2168, WX2170,
WX2172, WX2174, WX2176, WX2178, WX2180, WX2182, WX2184, WX2186,
WX2188, WX2190, WX2192, WX3071, WX3423, WX3425, WX3427, WX3429,
WX3431, WX3433, WX3435, WX3437, WX3439, WX3441, WX3443, WX3445,
WX3447, WX3449, WX3451, WX3453, WX3455, WX3457, WX3459, WX3461,
WX3463, WX3465, WX3467, WX3469, WX3471, WX3473, WX3475, WX3477,
WX3479, WX3481, WX3483, WX3485, WX4364, WX4716, WX4718, WX4720,
WX4722, WX4724, WX4726, WX4728, WX4730, WX4732, WX4734, WX4736,
WX4738, WX4740, WX4742, WX4744, WX4746, WX4748, WX4750, WX4752,
WX4754, WX4756, WX4758, WX4760, WX4762, WX4764, WX4766, WX4768,
WX4770, WX4772, WX4774, WX4776, WX4778, WX5657, WX6009, WX6011,
WX6013, WX6015, WX6017, WX6019, WX6021, WX6023, WX6025, WX6027,
WX6029, WX6031, WX6033, WX6035, WX6037, WX6039, WX6041, WX6043,
WX6045, WX6047, WX6049, WX6051, WX6053, WX6055, WX6057, WX6059,
WX6061, WX6063, WX6065, WX6067, WX6069, WX6071, WX6950, WX7302,
WX7304, WX7306, WX7308, WX7310, WX7312, WX7314, WX7316, WX7318,
WX7320, WX7322, WX7324, WX7326, WX7328, WX7330, WX7332, WX7334,
WX7336, WX7338, WX7340, WX7342, WX7344, WX7346, WX7348, WX7350,
WX7352, WX7354, WX7356, WX7358, WX7360, WX7362, WX7364, WX8243,
WX8595, WX8597, WX8599, WX8601, WX8603, WX8605, WX8607, WX8609,
WX8611, WX8613, WX8615, WX8617, WX8619, WX8621, WX8623, WX8625,
WX8627, WX8629, WX8631, WX8633, WX8635, WX8637, WX8639, WX8641,
WX8643, WX8645, WX8647, WX8649, WX8651, WX8653, WX8655, WX8657,
WX9536, WX9888, WX9890, WX9892, WX9894, WX9896, WX9898, WX9900,
WX9902, WX9904, WX9906, WX9908, WX9910, WX9912, WX9914, WX9916,
WX9918, WX9920, WX9922, WX9924, WX9926, WX9928, WX9930, WX9932,
WX9934, WX9936, WX9938, WX9940, WX9942, WX9944, WX9946, WX9948,
WX9950, WX10829, WX11181, WX11183, WX11185, WX11187, WX11189, WX11191,
WX11193, WX11195, WX11197, WX11199, WX11201, WX11203, WX11205,
WX11207, WX11209, WX11211, WX11213, WX11215, WX11217, WX11219,
WX11221, WX11223, WX11225, WX11227, WX11229, WX11231, WX11233,
WX11235, WX11237, WX11239, WX11241, WX11243, WX487, WX489, WX491,
WX493, WX495, WX497, WX499, WX501, WX503, WX505, WX507, WX509, WX511,
WX513, WX515, WX517, WX519, WX521, WX523, WX525, WX527, WX529, WX531,
WX533, WX535, WX537, WX539, WX541, WX543, WX545, WX547, n867, n872,
n877, n882, n887, n892, n897, n902, n907, n912, n917, n922, n927,
n932, n937, n942, n947, n952, n957, n962, n967, n972, n977, n982,
n987, n992, n997, n1002, n1007, n1012, n1017, n1022, n1027, WX645,
n1032, WX647, n1037, WX649, n1042, WX651, n1047, WX653, n1052, WX655,
n1057, WX657, n1062, WX659, n1067, WX661, n1072, WX663, n1077, WX665,
n1082, WX667, n1087, WX669, n1092, WX671, n1097, WX673, n1102, WX675,
n1107, WX677, n1112, WX679, n1117, WX681, n1122, WX683, n1127, WX685,
n1132, WX687, n1137, WX689, n1142, WX691, n1147, WX693, n1152, WX695,
n1157, WX697, n1162, WX699, n1167, WX701, n1172, WX703, n1177, WX705,
n1182, WX707, n1187, WX709, n1192, WX711, n1197, WX713, n1202, WX715,
n1207, WX717, n1212, WX719, n1217, WX721, n1222, WX723, n1227, WX725,
n1232, WX727, n1237, WX729, n1242, WX731, n1247, WX733, n1252, WX735,
n1257, WX737, n1262, WX739, n1267, WX741, n1272, WX743, n1277, WX745,
n1282, WX747, n1287, WX749, n1292, WX751, n1297, WX753, n1302, WX755,
n1307, WX757, n1312, WX759, n1317, WX761, n1322, WX763, n1327, WX765,
n1332, WX767, n1337, WX769, n1342, WX771, n1347, WX773, n1352, WX775,
n1357, WX777, n1362, WX779, n1367, WX781, n1372, WX783, n1377, WX785,
n1382, WX787, n1387, WX789, n1392, WX791, n1397, WX793, n1402, WX795,
n1407, WX797, n1412, WX799, n1417, WX801, n1422, WX803, n1427, WX805,
n1432, WX807, n1437, WX809, n1442, WX811, n1447, WX813, n1452, WX815,
n1457, WX817, n1462, WX819, n1467, WX821, n1472, WX823, n1477, WX825,
n1482, WX827, n1487, WX829, n1492, WX831, n1497, WX833, n1502, WX835,
n1507, n1512, n1516, n1520, n1524, n1528, n1532, n1536, n1540, n1544,
n1548, n1552, n1556, n1560, n1564, n1568, n1572, n1576, n1580, n1584,
n1588, n1592, n1596, n1600, n1604, n1608, n1612, n1616, n1620, n1624,
n1628, n1632, n1636, WX1780, WX1782, WX1784, WX1786, WX1788, WX1790,
WX1792, WX1794, WX1796, WX1798, WX1800, WX1802, WX1804, WX1806,
WX1808, WX1810, WX1812, WX1814, WX1816, WX1818, WX1820, WX1822,
WX1824, WX1826, WX1828, WX1830, WX1832, WX1834, WX1836, WX1838,
WX1840, n1795, n1800, n1805, n1810, n1815, n1820, n1825, n1830, n1835,
n1840, n1845, n1850, n1855, n1860, n1865, n1870, n1875, n1880, n1885,
n1890, n1895, n1900, n1905, n1910, n1915, n1920, n1925, n1930, n1935,
n1940, n1945, n1950, n1955, WX1938, n1960, WX1940, n1965, WX1942,
n1970, WX1944, n1975, WX1946, n1980, WX1948, n1985, WX1950, n1990,
WX1952, n1995, WX1954, n2000, WX1956, n2005, WX1958, n2010, WX1960,
n2015, WX1962, n2020, WX1964, n2025, WX1966, n2030, WX1968, n2035,
WX1970, n2040, WX1972, n2045, WX1974, n2050, WX1976, n2055, WX1978,
n2060, WX1980, n2065, WX1982, n2070, WX1984, n2075, WX1986, n2080,
WX1988, n2085, WX1990, n2090, WX1992, n2095, WX1994, n2100, WX1996,
n2105, WX1998, n2110, WX2000, n2115, WX2002, n2120, WX2004, n2125,
WX2006, n2130, WX2008, n2135, WX2010, n2140, WX2012, n2145, WX2014,
n2150, WX2016, n2155, WX2018, n2160, WX2020, n2165, WX2022, n2170,
WX2024, n2175, WX2026, n2180, WX2028, n2185, WX2030, n2190, WX2032,
n2195, WX2034, n2200, WX2036, n2205, WX2038, n2210, WX2040, n2215,
WX2042, n2220, WX2044, n2225, WX2046, n2230, WX2048, n2235, WX2050,
n2240, WX2052, n2245, WX2054, n2250, WX2056, n2255, WX2058, n2260,
WX2060, n2265, WX2062, n2270, WX2064, n2275, WX2066, n2280, WX2068,
n2285, WX2070, n2290, WX2072, n2295, WX2074, n2300, WX2076, n2305,
WX2078, n2310, WX2080, n2315, WX2082, n2320, WX2084, n2325, WX2086,
n2330, WX2088, n2335, WX2090, n2340, WX2092, n2345, WX2094, n2350,
WX2096, n2355, WX2098, n2360, WX2100, n2365, WX2102, n2370, WX2104,
n2375, WX2106, n2380, WX2108, n2385, WX2110, n2390, WX2112, n2395,
WX2114, n2400, WX2116, n2405, WX2118, n2410, WX2120, n2415, WX2122,
n2420, WX2124, n2425, WX2126, n2430, WX2128, n2435, n2440, n2444,
n2448, n2452, n2456, n2460, n2464, n2468, n2472, n2476, n2480, n2484,
n2488, n2492, n2496, n2500, n2504, n2508, n2512, n2516, n2520, n2524,
n2528, n2532, n2536, n2540, n2544, n2548, n2552, n2556, n2560, n2564,
WX3073, WX3075, WX3077, WX3079, WX3081, WX3083, WX3085, WX3087,
WX3089, WX3091, WX3093, WX3095, WX3097, WX3099, WX3101, WX3103,
WX3105, WX3107, WX3109, WX3111, WX3113, WX3115, WX3117, WX3119,
WX3121, WX3123, WX3125, WX3127, WX3129, WX3131, WX3133, n2723, n2728,
n2733, n2738, n2743, n2748, n2753, n2758, n2763, n2768, n2773, n2778,
n2783, n2788, n2793, n2798, n2803, n2808, n2813, n2818, n2823, n2828,
n2833, n2838, n2843, n2848, n2853, n2858, n2863, n2868, n2873, n2878,
n2883, WX3231, n2888, WX3233, n2893, WX3235, n2898, WX3237, n2903,
WX3239, n2908, WX3241, n2913, WX3243, n2918, WX3245, n2923, WX3247,
n2928, WX3249, n2933, WX3251, n2938, WX3253, n2943, WX3255, n2948,
WX3257, n2953, WX3259, n2958, WX3261, n2963, WX3263, n2968, WX3265,
n2973, WX3267, n2978, WX3269, n2983, WX3271, n2988, WX3273, n2993,
WX3275, n2998, WX3277, n3003, WX3279, n3008, WX3281, n3013, WX3283,
n3018, WX3285, n3023, WX3287, n3028, WX3289, n3033, WX3291, n3038,
WX3293, n3043, WX3295, n3048, WX3297, n3053, WX3299, n3058, WX3301,
n3063, WX3303, n3068, WX3305, n3073, WX3307, n3078, WX3309, n3083,
WX3311, n3088, WX3313, n3093, WX3315, n3098, WX3317, n3103, WX3319,
n3108, WX3321, n3113, WX3323, n3118, WX3325, n3123, WX3327, n3128,
WX3329, n3133, WX3331, n3138, WX3333, n3143, WX3335, n3148, WX3337,
n3153, WX3339, n3158, WX3341, n3163, WX3343, n3168, WX3345, n3173,
WX3347, n3178, WX3349, n3183, WX3351, n3188, WX3353, n3193, WX3355,
n3198, WX3357, n3203, WX3359, n3208, WX3361, n3213, WX3363, n3218,
WX3365, n3223, WX3367, n3228, WX3369, n3233, WX3371, n3238, WX3373,
n3243, WX3375, n3248, WX3377, n3253, WX3379, n3258, WX3381, n3263,
WX3383, n3268, WX3385, n3273, WX3387, n3278, WX3389, n3283, WX3391,
n3288, WX3393, n3293, WX3395, n3298, WX3397, n3303, WX3399, n3308,
WX3401, n3313, WX3403, n3318, WX3405, n3323, WX3407, n3328, WX3409,
n3333, WX3411, n3338, WX3413, n3343, WX3415, n3348, WX3417, n3353,
WX3419, n3358, WX3421, n3363, n3368, n3372, n3376, n3380, n3384,
n3388, n3392, n3396, n3400, n3404, n3408, n3412, n3416, n3420, n3424,
n3428, n3432, n3436, n3440, n3444, n3448, n3452, n3456, n3460, n3464,
n3468, n3472, n3476, n3480, n3484, n3488, n3492, WX4366, WX4368,
WX4370, WX4372, WX4374, WX4376, WX4378, WX4380, WX4382, WX4384,
WX4386, WX4388, WX4390, WX4392, WX4394, WX4396, WX4398, WX4400,
WX4402, WX4404, WX4406, WX4408, WX4410, WX4412, WX4414, WX4416,
WX4418, WX4420, WX4422, WX4424, WX4426, n3651, n3656, n3661, n3666,
n3671, n3676, n3681, n3686, n3691, n3696, n3701, n3706, n3711, n3716,
n3721, n3726, n3731, n3736, n3741, n3746, n3751, n3756, n3761, n3766,
n3771, n3776, n3781, n3786, n3791, n3796, n3801, n3806, n3811, WX4524,
n3816, WX4526, n3821, WX4528, n3826, WX4530, n3831, WX4532, n3836,
WX4534, n3841, WX4536, n3846, WX4538, n3851, WX4540, n3856, WX4542,
n3861, WX4544, n3866, WX4546, n3871, WX4548, n3876, WX4550, n3881,
WX4552, n3886, WX4554, n3891, WX4556, n3896, WX4558, n3901, WX4560,
n3906, WX4562, n3911, WX4564, n3916, WX4566, n3921, WX4568, n3926,
WX4570, n3931, WX4572, n3936, WX4574, n3941, WX4576, n3946, WX4578,
n3951, WX4580, n3956, WX4582, n3961, WX4584, n3966, WX4586, n3971,
WX4588, n3976, WX4590, n3981, WX4592, n3986, WX4594, n3991, WX4596,
n3996, WX4598, n4001, WX4600, n4006, WX4602, n4011, WX4604, n4016,
WX4606, n4021, WX4608, n4026, WX4610, n4031, WX4612, n4036, WX4614,
n4041, WX4616, n4046, WX4618, n4051, WX4620, n4056, WX4622, n4061,
WX4624, n4066, WX4626, n4071, WX4628, n4076, WX4630, n4081, WX4632,
n4086, WX4634, n4091, WX4636, n4096, WX4638, n4101, WX4640, n4106,
WX4642, n4111, WX4644, n4116, WX4646, n4121, WX4648, n4126, WX4650,
n4131, WX4652, n4136, WX4654, n4141, WX4656, n4146, WX4658, n4151,
WX4660, n4156, WX4662, n4161, WX4664, n4166, WX4666, n4171, WX4668,
n4176, WX4670, n4181, WX4672, n4186, WX4674, n4191, WX4676, n4196,
WX4678, n4201, WX4680, n4206, WX4682, n4211, WX4684, n4216, WX4686,
n4221, WX4688, n4226, WX4690, n4231, WX4692, n4236, WX4694, n4241,
WX4696, n4246, WX4698, n4251, WX4700, n4256, WX4702, n4261, WX4704,
n4266, WX4706, n4271, WX4708, n4276, WX4710, n4281, WX4712, n4286,
WX4714, n4291, n4296, n4300, n4304, n4308, n4312, n4316, n4320, n4324,
n4328, n4332, n4336, n4340, n4344, n4348, n4352, n4356, n4360, n4364,
n4368, n4372, n4376, n4380, n4384, n4388, n4392, n4396, n4400, n4404,
n4408, n4412, n4416, n4420, WX5659, WX5661, WX5663, WX5665, WX5667,
WX5669, WX5671, WX5673, WX5675, WX5677, WX5679, WX5681, WX5683,
WX5685, WX5687, WX5689, WX5691, WX5693, WX5695, WX5697, WX5699,
WX5701, WX5703, WX5705, WX5707, WX5709, WX5711, WX5713, WX5715,
WX5717, WX5719, n4579, n4584, n4589, n4594, n4599, n4604, n4609,
n4614, n4619, n4624, n4629, n4634, n4639, n4644, n4649, n4654, n4659,
n4664, n4669, n4674, n4679, n4684, n4689, n4694, n4699, n4704, n4709,
n4714, n4719, n4724, n4729, n4734, n4739, WX5817, n4744, WX5819,
n4749, WX5821, n4754, WX5823, n4759, WX5825, n4764, WX5827, n4769,
WX5829, n4774, WX5831, n4779, WX5833, n4784, WX5835, n4789, WX5837,
n4794, WX5839, n4799, WX5841, n4804, WX5843, n4809, WX5845, n4814,
WX5847, n4819, WX5849, n4824, WX5851, n4829, WX5853, n4834, WX5855,
n4839, WX5857, n4844, WX5859, n4849, WX5861, n4854, WX5863, n4859,
WX5865, n4864, WX5867, n4869, WX5869, n4874, WX5871, n4879, WX5873,
n4884, WX5875, n4889, WX5877, n4894, WX5879, n4899, WX5881, n4904,
WX5883, n4909, WX5885, n4914, WX5887, n4919, WX5889, n4924, WX5891,
n4929, WX5893, n4934, WX5895, n4939, WX5897, n4944, WX5899, n4949,
WX5901, n4954, WX5903, n4959, WX5905, n4964, WX5907, n4969, WX5909,
n4974, WX5911, n4979, WX5913, n4984, WX5915, n4989, WX5917, n4994,
WX5919, n4999, WX5921, n5004, WX5923, n5009, WX5925, n5014, WX5927,
n5019, WX5929, n5024, WX5931, n5029, WX5933, n5034, WX5935, n5039,
WX5937, n5044, WX5939, n5049, WX5941, n5054, WX5943, n5059, WX5945,
n5064, WX5947, n5069, WX5949, n5074, WX5951, n5079, WX5953, n5084,
WX5955, n5089, WX5957, n5094, WX5959, n5099, WX5961, n5104, WX5963,
n5109, WX5965, n5114, WX5967, n5119, WX5969, n5124, WX5971, n5129,
WX5973, n5134, WX5975, n5139, WX5977, n5144, WX5979, n5149, WX5981,
n5154, WX5983, n5159, WX5985, n5164, WX5987, n5169, WX5989, n5174,
WX5991, n5179, WX5993, n5184, WX5995, n5189, WX5997, n5194, WX5999,
n5199, WX6001, n5204, WX6003, n5209, WX6005, n5214, WX6007, n5219,
n5224, n5228, n5232, n5236, n5240, n5244, n5248, n5252, n5256, n5260,
n5264, n5268, n5272, n5276, n5280, n5284, n5288, n5292, n5296, n5300,
n5304, n5308, n5312, n5316, n5320, n5324, n5328, n5332, n5336, n5340,
n5344, n5348, WX6952, WX6954, WX6956, WX6958, WX6960, WX6962, WX6964,
WX6966, WX6968, WX6970, WX6972, WX6974, WX6976, WX6978, WX6980,
WX6982, WX6984, WX6986, WX6988, WX6990, WX6992, WX6994, WX6996,
WX6998, WX7000, WX7002, WX7004, WX7006, WX7008, WX7010, WX7012, n5507,
n5512, n5517, n5522, n5527, n5532, n5537, n5542, n5547, n5552, n5557,
n5562, n5567, n5572, n5577, n5582, n5587, n5592, n5597, n5602, n5607,
n5612, n5617, n5622, n5627, n5632, n5637, n5642, n5647, n5652, n5657,
n5662, n5667, WX7110, n5672, WX7112, n5677, WX7114, n5682, WX7116,
n5687, WX7118, n5692, WX7120, n5697, WX7122, n5702, WX7124, n5707,
WX7126, n5712, WX7128, n5717, WX7130, n5722, WX7132, n5727, WX7134,
n5732, WX7136, n5737, WX7138, n5742, WX7140, n5747, WX7142, n5752,
WX7144, n5757, WX7146, n5762, WX7148, n5767, WX7150, n5772, WX7152,
n5777, WX7154, n5782, WX7156, n5787, WX7158, n5792, WX7160, n5797,
WX7162, n5802, WX7164, n5807, WX7166, n5812, WX7168, n5817, WX7170,
n5822, WX7172, n5827, WX7174, n5832, WX7176, n5837, WX7178, n5842,
WX7180, n5847, WX7182, n5852, WX7184, n5857, WX7186, n5862, WX7188,
n5867, WX7190, n5872, WX7192, n5877, WX7194, n5882, WX7196, n5887,
WX7198, n5892, WX7200, n5897, WX7202, n5902, WX7204, n5907, WX7206,
n5912, WX7208, n5917, WX7210, n5922, WX7212, n5927, WX7214, n5932,
WX7216, n5937, WX7218, n5942, WX7220, n5947, WX7222, n5952, WX7224,
n5957, WX7226, n5962, WX7228, n5967, WX7230, n5972, WX7232, n5977,
WX7234, n5982, WX7236, n5987, WX7238, n5992, WX7240, n5997, WX7242,
n6002, WX7244, n6007, WX7246, n6012, WX7248, n6017, WX7250, n6022,
WX7252, n6027, WX7254, n6032, WX7256, n6037, WX7258, n6042, WX7260,
n6047, WX7262, n6052, WX7264, n6057, WX7266, n6062, WX7268, n6067,
WX7270, n6072, WX7272, n6077, WX7274, n6082, WX7276, n6087, WX7278,
n6092, WX7280, n6097, WX7282, n6102, WX7284, n6107, WX7286, n6112,
WX7288, n6117, WX7290, n6122, WX7292, n6127, WX7294, n6132, WX7296,
n6137, WX7298, n6142, WX7300, n6147, n6152, n6156, n6160, n6164,
n6168, n6172, n6176, n6180, n6184, n6188, n6192, n6196, n6200, n6204,
n6208, n6212, n6216, n6220, n6224, n6228, n6232, n6236, n6240, n6244,
n6248, n6252, n6256, n6260, n6264, n6268, n6272, n6276, WX8245,
WX8247, WX8249, WX8251, WX8253, WX8255, WX8257, WX8259, WX8261,
WX8263, WX8265, WX8267, WX8269, WX8271, WX8273, WX8275, WX8277,
WX8279, WX8281, WX8283, WX8285, WX8287, WX8289, WX8291, WX8293,
WX8295, WX8297, WX8299, WX8301, WX8303, WX8305, n6435, n6440, n6445,
n6450, n6455, n6460, n6465, n6470, n6475, n6480, n6485, n6490, n6495,
n6500, n6505, n6510, n6515, n6520, n6525, n6530, n6535, n6540, n6545,
n6550, n6555, n6560, n6565, n6570, n6575, n6580, n6585, n6590, n6595,
WX8403, n6600, WX8405, n6605, WX8407, n6610, WX8409, n6615, WX8411,
n6620, WX8413, n6625, WX8415, n6630, WX8417, n6635, WX8419, n6640,
WX8421, n6645, WX8423, n6650, WX8425, n6655, WX8427, n6660, WX8429,
n6665, WX8431, n6670, WX8433, n6675, WX8435, n6680, WX8437, n6685,
WX8439, n6690, WX8441, n6695, WX8443, n6700, WX8445, n6705, WX8447,
n6710, WX8449, n6715, WX8451, n6720, WX8453, n6725, WX8455, n6730,
WX8457, n6735, WX8459, n6740, WX8461, n6745, WX8463, n6750, WX8465,
n6755, WX8467, n6760, WX8469, n6765, WX8471, n6770, WX8473, n6775,
WX8475, n6780, WX8477, n6785, WX8479, n6790, WX8481, n6795, WX8483,
n6800, WX8485, n6805, WX8487, n6810, WX8489, n6815, WX8491, n6820,
WX8493, n6825, WX8495, n6830, WX8497, n6835, WX8499, n6840, WX8501,
n6845, WX8503, n6850, WX8505, n6855, WX8507, n6860, WX8509, n6865,
WX8511, n6870, WX8513, n6875, WX8515, n6880, WX8517, n6885, WX8519,
n6890, WX8521, n6895, WX8523, n6900, WX8525, n6905, WX8527, n6910,
WX8529, n6915, WX8531, n6920, WX8533, n6925, WX8535, n6930, WX8537,
n6935, WX8539, n6940, WX8541, n6945, WX8543, n6950, WX8545, n6955,
WX8547, n6960, WX8549, n6965, WX8551, n6970, WX8553, n6975, WX8555,
n6980, WX8557, n6985, WX8559, n6990, WX8561, n6995, WX8563, n7000,
WX8565, n7005, WX8567, n7010, WX8569, n7015, WX8571, n7020, WX8573,
n7025, WX8575, n7030, WX8577, n7035, WX8579, n7040, WX8581, n7045,
WX8583, n7050, WX8585, n7055, WX8587, n7060, WX8589, n7065, WX8591,
n7070, WX8593, n7075, n7080, n7084, n7088, n7092, n7096, n7100, n7104,
n7108, n7112, n7116, n7120, n7124, n7128, n7132, n7136, n7140, n7144,
n7148, n7152, n7156, n7160, n7164, n7168, n7172, n7176, n7180, n7184,
n7188, n7192, n7196, n7200, n7204, WX9538, WX9540, WX9542, WX9544,
WX9546, WX9548, WX9550, WX9552, WX9554, WX9556, WX9558, WX9560,
WX9562, WX9564, WX9566, WX9568, WX9570, WX9572, WX9574, WX9576,
WX9578, WX9580, WX9582, WX9584, WX9586, WX9588, WX9590, WX9592,
WX9594, WX9596, WX9598, n7363, n7368, n7373, n7378, n7383, n7388,
n7393, n7398, n7403, n7408, n7413, n7418, n7423, n7428, n7433, n7438,
n7443, n7448, n7453, n7458, n7463, n7468, n7473, n7478, n7483, n7488,
n7493, n7498, n7503, n7508, n7513, n7518, n7523, WX9696, n7528,
WX9698, n7533, WX9700, n7538, WX9702, n7543, WX9704, n7548, WX9706,
n7553, WX9708, n7558, WX9710, n7563, WX9712, n7568, WX9714, n7573,
WX9716, n7578, WX9718, n7583, WX9720, n7588, WX9722, n7593, WX9724,
n7598, WX9726, n7603, WX9728, n7608, WX9730, n7613, WX9732, n7618,
WX9734, n7623, WX9736, n7628, WX9738, n7633, WX9740, n7638, WX9742,
n7643, WX9744, n7648, WX9746, n7653, WX9748, n7658, WX9750, n7663,
WX9752, n7668, WX9754, n7673, WX9756, n7678, WX9758, n7683, WX9760,
n7688, WX9762, n7693, WX9764, n7698, WX9766, n7703, WX9768, n7708,
WX9770, n7713, WX9772, n7718, WX9774, n7723, WX9776, n7728, WX9778,
n7733, WX9780, n7738, WX9782, n7743, WX9784, n7748, WX9786, n7753,
WX9788, n7758, WX9790, n7763, WX9792, n7768, WX9794, n7773, WX9796,
n7778, WX9798, n7783, WX9800, n7788, WX9802, n7793, WX9804, n7798,
WX9806, n7803, WX9808, n7808, WX9810, n7813, WX9812, n7818, WX9814,
n7823, WX9816, n7828, WX9818, n7833, WX9820, n7838, WX9822, n7843,
WX9824, n7848, WX9826, n7853, WX9828, n7858, WX9830, n7863, WX9832,
n7868, WX9834, n7873, WX9836, n7878, WX9838, n7883, WX9840, n7888,
WX9842, n7893, WX9844, n7898, WX9846, n7903, WX9848, n7908, WX9850,
n7913, WX9852, n7918, WX9854, n7923, WX9856, n7928, WX9858, n7933,
WX9860, n7938, WX9862, n7943, WX9864, n7948, WX9866, n7953, WX9868,
n7958, WX9870, n7963, WX9872, n7968, WX9874, n7973, WX9876, n7978,
WX9878, n7983, WX9880, n7988, WX9882, n7993, WX9884, n7998, WX9886,
n8003, n8008, n8012, n8016, n8020, n8024, n8028, n8032, n8036, n8040,
n8044, n8048, n8052, n8056, n8060, n8064, n8068, n8072, n8076, n8080,
n8084, n8088, n8092, n8096, n8100, n8104, n8108, n8112, n8116, n8120,
n8124, n8128, n8132, WX10831, WX10833, WX10835, WX10837, WX10839,
WX10841, WX10843, WX10845, WX10847, WX10849, WX10851, WX10853,
WX10855, WX10857, WX10859, WX10861, WX10863, WX10865, WX10867,
WX10869, WX10871, WX10873, WX10875, WX10877, WX10879, WX10881,
WX10883, WX10885, WX10887, WX10889, WX10891, n8291, n8296, n8301,
n8306, n8311, n8316, n8321, n8326, n8331, n8336, n8341, n8346, n8351,
n8356, n8361, n8366, n8371, n8376, n8381, n8386, n8391, n8396, n8401,
n8406, n8411, n8416, n8421, n8426, n8431, n8436, n8441, n8446, n8451,
WX10989, n8456, WX10991, n8461, WX10993, n8466, WX10995, n8471,
WX10997, n8476, WX10999, n8481, WX11001, n8486, WX11003, n8491,
WX11005, n8496, WX11007, n8501, WX11009, n8506, WX11011, n8511,
WX11013, n8516, WX11015, n8521, WX11017, n8526, WX11019, n8531,
WX11021, n8536, WX11023, n8541, WX11025, n8546, WX11027, n8551,
WX11029, n8556, WX11031, n8561, WX11033, n8566, WX11035, n8571,
WX11037, n8576, WX11039, n8581, WX11041, n8586, WX11043, n8591,
WX11045, n8596, WX11047, n8601, WX11049, n8606, WX11051, n8611,
WX11053, n8616, WX11055, n8621, WX11057, n8626, WX11059, n8631,
WX11061, n8636, WX11063, n8641, WX11065, n8646, WX11067, n8651,
WX11069, n8656, WX11071, n8661, WX11073, n8666, WX11075, n8671,
WX11077, n8676, WX11079, n8681, WX11081, n8686, WX11083, n8691,
WX11085, n8696, WX11087, n8701, WX11089, n8706, WX11091, n8711,
WX11093, n8716, WX11095, n8721, WX11097, n8726, WX11099, n8731,
WX11101, n8736, WX11103, n8741, WX11105, n8746, WX11107, n8751,
WX11109, n8756, WX11111, n8761, WX11113, n8766, WX11115, n8771,
WX11117, n8776, WX11119, n8781, WX11121, n8786, WX11123, n8791,
WX11125, n8796, WX11127, n8801, WX11129, n8806, WX11131, n8811,
WX11133, n8816, WX11135, n8821, WX11137, n8826, WX11139, n8831,
WX11141, n8836, WX11143, n8841, WX11145, n8846, WX11147, n8851,
WX11149, n8856, WX11151, n8861, WX11153, n8866, WX11155, n8871,
WX11157, n8876, WX11159, n8881, WX11161, n8886, WX11163, n8891,
WX11165, n8896, WX11167, n8901, WX11169, n8906, WX11171, n8911,
WX11173, n8916, WX11175, n8921, WX11177, n8926, WX11179, n8931, n8936,
n8940, n8944, n8948, n8952, n8956, n8960, n8964, n8968, n8972, n8976,
n8980, n8984, n8988, n8992, n8996, n9000, n9004, n9008, n9012, n9016,
n9020, n9024, n9028, n9032, n9036, n9040, n9044, n9048, n9052, n9056,
n9060, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
n276, n277, n278, n279, n285, n287, n289, n291, n293, n295, n297,
n299, n301, n303, n305, n307, n309, n311, n313, n315, n317, n319,
n321, n323, n325, n327, n329, n331, n333, n335, n337, n339, n341,
n343, n345, n347, n348, n349, n350, n351, n352, n353, n354, n355,
n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
n862, n863, n864, n865, n866, n868, n869, n870, n871, n873, n874,
n875, n876, n878, n879, n880, n881, n883, n884, n885, n886, n888,
n889, n890, n891, n893, n894, n895, n896, n898, n899, n900, n901,
n903, n904, n905, n906, n908, n909, n910, n911, n913, n914, n915,
n916, n918, n919, n920, n921, n923, n924, n925, n926, n928, n929,
n930, n931, n933, n934, n935, n936, n938, n939, n940, n941, n943,
n944, n945, n946, n948, n949, n950, n951, n953, n954, n955, n956,
n958, n959, n960, n961, n963, n964, n965, n966, n968, n969, n970,
n971, n973, n974, n975, n976, n978, n979, n980, n981, n983, n984,
n985, n986, n988, n989, n990, n991, n993, n994, n995, n996, n998,
n999, n1000, n1001, n1003, n1004, n1005, n1006, n1008, n1009, n1010,
n1011, n1013, n1014, n1015, n1016, n1018, n1019, n1020, n1021, n1023,
n1024, n1025, n1026, n1028, n1029, n1030, n1031, n1033, n1034, n1035,
n1036, n1038, n1039, n1040, n1041, n1043, n1044, n1045, n1046, n1048,
n1049, n1050, n1051, n1053, n1054, n1055, n1056, n1058, n1059, n1060,
n1061, n1063, n1064, n1065, n1066, n1068, n1069, n1070, n1071, n1073,
n1074, n1075, n1076, n1078, n1079, n1080, n1081, n1083, n1084, n1085,
n1086, n1088, n1089, n1090, n1091, n1093, n1094, n1095, n1096, n1098,
n1099, n1100, n1101, n1103, n1104, n1105, n1106, n1108, n1109, n1110,
n1111, n1113, n1114, n1115, n1116, n1118, n1119, n1120, n1121, n1123,
n1124, n1125, n1126, n1128, n1129, n1130, n1131, n1133, n1134, n1135,
n1136, n1138, n1139, n1140, n1141, n1143, n1144, n1145, n1146, n1148,
n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1158, n1159, n1160,
n1161, n1163, n1164, n1165, n1166, n1168, n1169, n1170, n1171, n1173,
n1174, n1175, n1176, n1178, n1179, n1180, n1181, n1183, n1184, n1185,
n1186, n1188, n1189, n1190, n1191, n1193, n1194, n1195, n1196, n1198,
n1199, n1200, n1201, n1203, n1204, n1205, n1206, n1208, n1209, n1210,
n1211, n1213, n1214, n1215, n1216, n1218, n1219, n1220, n1221, n1223,
n1224, n1225, n1226, n1228, n1229, n1230, n1231, n1233, n1234, n1235,
n1236, n1238, n1239, n1240, n1241, n1243, n1244, n1245, n1246, n1248,
n1249, n1250, n1251, n1253, n1254, n1255, n1256, n1258, n1259, n1260,
n1261, n1263, n1264, n1265, n1266, n1268, n1269, n1270, n1271, n1273,
n1274, n1275, n1276, n1278, n1279, n1280, n1281, n1283, n1284, n1285,
n1286, n1288, n1289, n1290, n1291, n1293, n1294, n1295, n1296, n1298,
n1299, n1300, n1301, n1303, n1304, n1305, n1306, n1308, n1309, n1310,
n1311, n1313, n1314, n1315, n1316, n1318, n1319, n1320, n1321, n1323,
n1324, n1325, n1326, n1328, n1329, n1330, n1331, n1333, n1334, n1335,
n1336, n1338, n1339, n1340, n1341, n1343, n1344, n1345, n1346, n1348,
n1349, n1350, n1351, n1353, n1354, n1355, n1356, n1358, n1359, n1360,
n1361, n1363, n1364, n1365, n1366, n1368, n1369, n1370, n1371, n1373,
n1374, n1375, n1376, n1378, n1379, n1380, n1381, n1383, n1384, n1385,
n1386, n1388, n1389, n1390, n1391, n1393, n1394, n1395, n1396, n1398,
n1399, n1400, n1401, n1403, n1404, n1405, n1406, n1408, n1409, n1410,
n1411, n1413, n1414, n1415, n1416, n1418, n1419, n1420, n1421, n1423,
n1424, n1425, n1426, n1428, n1429, n1430, n1431, n1433, n1434, n1435,
n1436, n1438, n1439, n1440, n1441, n1443, n1444, n1445, n1446, n1448,
n1449, n1450, n1451, n1453, n1454, n1455, n1456, n1458, n1459, n1460,
n1461, n1463, n1464, n1465, n1466, n1468, n1469, n1470, n1471, n1473,
n1474, n1475, n1476, n1478, n1479, n1480, n1481, n1483, n1484, n1485,
n1486, n1488, n1489, n1490, n1491, n1493, n1494, n1495, n1496, n1498,
n1499, n1500, n1501, n1503, n1504, n1505, n1506, n1508, n1509, n1510,
n1511, n1513, n1514, n1515, n1517, n1518, n1519, n1521, n1522, n1523,
n1525, n1526, n1527, n1529, n1530, n1531, n1533, n1534, n1535, n1537,
n1538, n1539, n1541, n1542, n1543, n1545, n1546, n1547, n1549, n1550,
n1551, n1553, n1554, n1555, n1557, n1558, n1559, n1561, n1562, n1563,
n1565, n1566, n1567, n1569, n1570, n1571, n1573, n1574, n1575, n1577,
n1578, n1579, n1581, n1582, n1583, n1585, n1586, n1587, n1589, n1590,
n1591, n1593, n1594, n1595, n1597, n1598, n1599, n1601, n1602, n1603,
n1605, n1606, n1607, n1609, n1610, n1611, n1613, n1614, n1615, n1617,
n1618, n1619, n1621, n1622, n1623, n1625, n1626, n1627, n1629, n1630,
n1631, n1633, n1634, n1635, n1637, n1638, n1639, n1640, n1641, n1642,
n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
n1793, n1794, n1796, n1797, n1798, n1799, n1801, n1802, n1803, n1804,
n1806, n1807, n1808, n1809, n1811, n1812, n1813, n1814, n1816, n1817,
n1818, n1819, n1821, n1822, n1823, n1824, n1826, n1827, n1828, n1829,
n1831, n1832, n1833, n1834, n1836, n1837, n1838, n1839, n1841, n1842,
n1843, n1844, n1846, n1847, n1848, n1849, n1851, n1852, n1853, n1854,
n1856, n1857, n1858, n1859, n1861, n1862, n1863, n1864, n1866, n1867,
n1868, n1869, n1871, n1872, n1873, n1874, n1876, n1877, n1878, n1879,
n1881, n1882, n1883, n1884, n1886, n1887, n1888, n1889, n1891, n1892,
n1893, n1894, n1896, n1897, n1898, n1899, n1901, n1902, n1903, n1904,
n1906, n1907, n1908, n1909, n1911, n1912, n1913, n1914, n1916, n1917,
n1918, n1919, n1921, n1922, n1923, n1924, n1926, n1927, n1928, n1929,
n1931, n1932, n1933, n1934, n1936, n1937, n1938, n1939, n1941, n1942,
n1943, n1944, n1946, n1947, n1948, n1949, n1951, n1952, n1953, n1954,
n1956, n1957, n1958, n1959, n1961, n1962, n1963, n1964, n1966, n1967,
n1968, n1969, n1971, n1972, n1973, n1974, n1976, n1977, n1978, n1979,
n1981, n1982, n1983, n1984, n1986, n1987, n1988, n1989, n1991, n1992,
n1993, n1994, n1996, n1997, n1998, n1999, n2001, n2002, n2003, n2004,
n2006, n2007, n2008, n2009, n2011, n2012, n2013, n2014, n2016, n2017,
n2018, n2019, n2021, n2022, n2023, n2024, n2026, n2027, n2028, n2029,
n2031, n2032, n2033, n2034, n2036, n2037, n2038, n2039, n2041, n2042,
n2043, n2044, n2046, n2047, n2048, n2049, n2051, n2052, n2053, n2054,
n2056, n2057, n2058, n2059, n2061, n2062, n2063, n2064, n2066, n2067,
n2068, n2069, n2071, n2072, n2073, n2074, n2076, n2077, n2078, n2079,
n2081, n2082, n2083, n2084, n2086, n2087, n2088, n2089, n2091, n2092,
n2093, n2094, n2096, n2097, n2098, n2099, n2101, n2102, n2103, n2104,
n2106, n2107, n2108, n2109, n2111, n2112, n2113, n2114, n2116, n2117,
n2118, n2119, n2121, n2122, n2123, n2124, n2126, n2127, n2128, n2129,
n2131, n2132, n2133, n2134, n2136, n2137, n2138, n2139, n2141, n2142,
n2143, n2144, n2146, n2147, n2148, n2149, n2151, n2152, n2153, n2154,
n2156, n2157, n2158, n2159, n2161, n2162, n2163, n2164, n2166, n2167,
n2168, n2169, n2171, n2172, n2173, n2174, n2176, n2177, n2178, n2179,
n2181, n2182, n2183, n2184, n2186, n2187, n2188, n2189, n2191, n2192,
n2193, n2194, n2196, n2197, n2198, n2199, n2201, n2202, n2203, n2204,
n2206, n2207, n2208, n2209, n2211, n2212, n2213, n2214, n2216, n2217,
n2218, n2219, n2221, n2222, n2223, n2224, n2226, n2227, n2228, n2229,
n2231, n2232, n2233, n2234, n2236, n2237, n2238, n2239, n2241, n2242,
n2243, n2244, n2246, n2247, n2248, n2249, n2251, n2252, n2253, n2254,
n2256, n2257, n2258, n2259, n2261, n2262, n2263, n2264, n2266, n2267,
n2268, n2269, n2271, n2272, n2273, n2274, n2276, n2277, n2278, n2279,
n2281, n2282, n2283, n2284, n2286, n2287, n2288, n2289, n2291, n2292,
n2293, n2294, n2296, n2297, n2298, n2299, n2301, n2302, n2303, n2304,
n2306, n2307, n2308, n2309, n2311, n2312, n2313, n2314, n2316, n2317,
n2318, n2319, n2321, n2322, n2323, n2324, n2326, n2327, n2328, n2329,
n2331, n2332, n2333, n2334, n2336, n2337, n2338, n2339, n2341, n2342,
n2343, n2344, n2346, n2347, n2348, n2349, n2351, n2352, n2353, n2354,
n2356, n2357, n2358, n2359, n2361, n2362, n2363, n2364, n2366, n2367,
n2368, n2369, n2371, n2372, n2373, n2374, n2376, n2377, n2378, n2379,
n2381, n2382, n2383, n2384, n2386, n2387, n2388, n2389, n2391, n2392,
n2393, n2394, n2396, n2397, n2398, n2399, n2401, n2402, n2403, n2404,
n2406, n2407, n2408, n2409, n2411, n2412, n2413, n2414, n2416, n2417,
n2418, n2419, n2421, n2422, n2423, n2424, n2426, n2427, n2428, n2429,
n2431, n2432, n2433, n2434, n2436, n2437, n2438, n2439, n2441, n2442,
n2443, n2445, n2446, n2447, n2449, n2450, n2451, n2453, n2454, n2455,
n2457, n2458, n2459, n2461, n2462, n2463, n2465, n2466, n2467, n2469,
n2470, n2471, n2473, n2474, n2475, n2477, n2478, n2479, n2481, n2482,
n2483, n2485, n2486, n2487, n2489, n2490, n2491, n2493, n2494, n2495,
n2497, n2498, n2499, n2501, n2502, n2503, n2505, n2506, n2507, n2509,
n2510, n2511, n2513, n2514, n2515, n2517, n2518, n2519, n2521, n2522,
n2523, n2525, n2526, n2527, n2529, n2530, n2531, n2533, n2534, n2535,
n2537, n2538, n2539, n2541, n2542, n2543, n2545, n2546, n2547, n2549,
n2550, n2551, n2553, n2554, n2555, n2557, n2558, n2559, n2561, n2562,
n2563, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2724,
n2725, n2726, n2727, n2729, n2730, n2731, n2732, n2734, n2735, n2736,
n2737, n2739, n2740, n2741, n2742, n2744, n2745, n2746, n2747, n2749,
n2750, n2751, n2752, n2754, n2755, n2756, n2757, n2759, n2760, n2761,
n2762, n2764, n2765, n2766, n2767, n2769, n2770, n2771, n2772, n2774,
n2775, n2776, n2777, n2779, n2780, n2781, n2782, n2784, n2785, n2786,
n2787, n2789, n2790, n2791, n2792, n2794, n2795, n2796, n2797, n2799,
n2800, n2801, n2802, n2804, n2805, n2806, n2807, n2809, n2810, n2811,
n2812, n2814, n2815, n2816, n2817, n2819, n2820, n2821, n2822, n2824,
n2825, n2826, n2827, n2829, n2830, n2831, n2832, n2834, n2835, n2836,
n2837, n2839, n2840, n2841, n2842, n2844, n2845, n2846, n2847, n2849,
n2850, n2851, n2852, n2854, n2855, n2856, n2857, n2859, n2860, n2861,
n2862, n2864, n2865, n2866, n2867, n2869, n2870, n2871, n2872, n2874,
n2875, n2876, n2877, n2879, n2880, n2881, n2882, n2884, n2885, n2886,
n2887, n2889, n2890, n2891, n2892, n2894, n2895, n2896, n2897, n2899,
n2900, n2901, n2902, n2904, n2905, n2906, n2907, n2909, n2910, n2911,
n2912, n2914, n2915, n2916, n2917, n2919, n2920, n2921, n2922, n2924,
n2925, n2926, n2927, n2929, n2930, n2931, n2932, n2934, n2935, n2936,
n2937, n2939, n2940, n2941, n2942, n2944, n2945, n2946, n2947, n2949,
n2950, n2951, n2952, n2954, n2955, n2956, n2957, n2959, n2960, n2961,
n2962, n2964, n2965, n2966, n2967, n2969, n2970, n2971, n2972, n2974,
n2975, n2976, n2977, n2979, n2980, n2981, n2982, n2984, n2985, n2986,
n2987, n2989, n2990, n2991, n2992, n2994, n2995, n2996, n2997, n2999,
n3000, n3001, n3002, n3004, n3005, n3006, n3007, n3009, n3010, n3011,
n3012, n3014, n3015, n3016, n3017, n3019, n3020, n3021, n3022, n3024,
n3025, n3026, n3027, n3029, n3030, n3031, n3032, n3034, n3035, n3036,
n3037, n3039, n3040, n3041, n3042, n3044, n3045, n3046, n3047, n3049,
n3050, n3051, n3052, n3054, n3055, n3056, n3057, n3059, n3060, n3061,
n3062, n3064, n3065, n3066, n3067, n3069, n3070, n3071, n3072, n3074,
n3075, n3076, n3077, n3079, n3080, n3081, n3082, n3084, n3085, n3086,
n3087, n3089, n3090, n3091, n3092, n3094, n3095, n3096, n3097, n3099,
n3100, n3101, n3102, n3104, n3105, n3106, n3107, n3109, n3110, n3111,
n3112, n3114, n3115, n3116, n3117, n3119, n3120, n3121, n3122, n3124,
n3125, n3126, n3127, n3129, n3130, n3131, n3132, n3134, n3135, n3136,
n3137, n3139, n3140, n3141, n3142, n3144, n3145, n3146, n3147, n3149,
n3150, n3151, n3152, n3154, n3155, n3156, n3157, n3159, n3160, n3161,
n3162, n3164, n3165, n3166, n3167, n3169, n3170, n3171, n3172, n3174,
n3175, n3176, n3177, n3179, n3180, n3181, n3182, n3184, n3185, n3186,
n3187, n3189, n3190, n3191, n3192, n3194, n3195, n3196, n3197, n3199,
n3200, n3201, n3202, n3204, n3205, n3206, n3207, n3209, n3210, n3211,
n3212, n3214, n3215, n3216, n3217, n3219, n3220, n3221, n3222, n3224,
n3225, n3226, n3227, n3229, n3230, n3231, n3232, n3234, n3235, n3236,
n3237, n3239, n3240, n3241, n3242, n3244, n3245, n3246, n3247, n3249,
n3250, n3251, n3252, n3254, n3255, n3256, n3257, n3259, n3260, n3261,
n3262, n3264, n3265, n3266, n3267, n3269, n3270, n3271, n3272, n3274,
n3275, n3276, n3277, n3279, n3280, n3281, n3282, n3284, n3285, n3286,
n3287, n3289, n3290, n3291, n3292, n3294, n3295, n3296, n3297, n3299,
n3300, n3301, n3302, n3304, n3305, n3306, n3307, n3309, n3310, n3311,
n3312, n3314, n3315, n3316, n3317, n3319, n3320, n3321, n3322, n3324,
n3325, n3326, n3327, n3329, n3330, n3331, n3332, n3334, n3335, n3336,
n3337, n3339, n3340, n3341, n3342, n3344, n3345, n3346, n3347, n3349,
n3350, n3351, n3352, n3354, n3355, n3356, n3357, n3359, n3360, n3361,
n3362, n3364, n3365, n3366, n3367, n3369, n3370, n3371, n3373, n3374,
n3375, n3377, n3378, n3379, n3381, n3382, n3383, n3385, n3386, n3387,
n3389, n3390, n3391, n3393, n3394, n3395, n3397, n3398, n3399, n3401,
n3402, n3403, n3405, n3406, n3407, n3409, n3410, n3411, n3413, n3414,
n3415, n3417, n3418, n3419, n3421, n3422, n3423, n3425, n3426, n3427,
n3429, n3430, n3431, n3433, n3434, n3435, n3437, n3438, n3439, n3441,
n3442, n3443, n3445, n3446, n3447, n3449, n3450, n3451, n3453, n3454,
n3455, n3457, n3458, n3459, n3461, n3462, n3463, n3465, n3466, n3467,
n3469, n3470, n3471, n3473, n3474, n3475, n3477, n3478, n3479, n3481,
n3482, n3483, n3485, n3486, n3487, n3489, n3490, n3491, n3493, n3494,
n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
n3645, n3646, n3647, n3648, n3649, n3650, n3652, n3653, n3654, n3655,
n3657, n3658, n3659, n3660, n3662, n3663, n3664, n3665, n3667, n3668,
n3669, n3670, n3672, n3673, n3674, n3675, n3677, n3678, n3679, n3680,
n3682, n3683, n3684, n3685, n3687, n3688, n3689, n3690, n3692, n3693,
n3694, n3695, n3697, n3698, n3699, n3700, n3702, n3703, n3704, n3705,
n3707, n3708, n3709, n3710, n3712, n3713, n3714, n3715, n3717, n3718,
n3719, n3720, n3722, n3723, n3724, n3725, n3727, n3728, n3729, n3730,
n3732, n3733, n3734, n3735, n3737, n3738, n3739, n3740, n3742, n3743,
n3744, n3745, n3747, n3748, n3749, n3750, n3752, n3753, n3754, n3755,
n3757, n3758, n3759, n3760, n3762, n3763, n3764, n3765, n3767, n3768,
n3769, n3770, n3772, n3773, n3774, n3775, n3777, n3778, n3779, n3780,
n3782, n3783, n3784, n3785, n3787, n3788, n3789, n3790, n3792, n3793,
n3794, n3795, n3797, n3798, n3799, n3800, n3802, n3803, n3804, n3805,
n3807, n3808, n3809, n3810, n3812, n3813, n3814, n3815, n3817, n3818,
n3819, n3820, n3822, n3823, n3824, n3825, n3827, n3828, n3829, n3830,
n3832, n3833, n3834, n3835, n3837, n3838, n3839, n3840, n3842, n3843,
n3844, n3845, n3847, n3848, n3849, n3850, n3852, n3853, n3854, n3855,
n3857, n3858, n3859, n3860, n3862, n3863, n3864, n3865, n3867, n3868,
n3869, n3870, n3872, n3873, n3874, n3875, n3877, n3878, n3879, n3880,
n3882, n3883, n3884, n3885, n3887, n3888, n3889, n3890, n3892, n3893,
n3894, n3895, n3897, n3898, n3899, n3900, n3902, n3903, n3904, n3905,
n3907, n3908, n3909, n3910, n3912, n3913, n3914, n3915, n3917, n3918,
n3919, n3920, n3922, n3923, n3924, n3925, n3927, n3928, n3929, n3930,
n3932, n3933, n3934, n3935, n3937, n3938, n3939, n3940, n3942, n3943,
n3944, n3945, n3947, n3948, n3949, n3950, n3952, n3953, n3954, n3955,
n3957, n3958, n3959, n3960, n3962, n3963, n3964, n3965, n3967, n3968,
n3969, n3970, n3972, n3973, n3974, n3975, n3977, n3978, n3979, n3980,
n3982, n3983, n3984, n3985, n3987, n3988, n3989, n3990, n3992, n3993,
n3994, n3995, n3997, n3998, n3999, n4000, n4002, n4003, n4004, n4005,
n4007, n4008, n4009, n4010, n4012, n4013, n4014, n4015, n4017, n4018,
n4019, n4020, n4022, n4023, n4024, n4025, n4027, n4028, n4029, n4030,
n4032, n4033, n4034, n4035, n4037, n4038, n4039, n4040, n4042, n4043,
n4044, n4045, n4047, n4048, n4049, n4050, n4052, n4053, n4054, n4055,
n4057, n4058, n4059, n4060, n4062, n4063, n4064, n4065, n4067, n4068,
n4069, n4070, n4072, n4073, n4074, n4075, n4077, n4078, n4079, n4080,
n4082, n4083, n4084, n4085, n4087, n4088, n4089, n4090, n4092, n4093,
n4094, n4095, n4097, n4098, n4099, n4100, n4102, n4103, n4104, n4105,
n4107, n4108, n4109, n4110, n4112, n4113, n4114, n4115, n4117, n4118,
n4119, n4120, n4122, n4123, n4124, n4125, n4127, n4128, n4129, n4130,
n4132, n4133, n4134, n4135, n4137, n4138, n4139, n4140, n4142, n4143,
n4144, n4145, n4147, n4148, n4149, n4150, n4152, n4153, n4154, n4155,
n4157, n4158, n4159, n4160, n4162, n4163, n4164, n4165, n4167, n4168,
n4169, n4170, n4172, n4173, n4174, n4175, n4177, n4178, n4179, n4180,
n4182, n4183, n4184, n4185, n4187, n4188, n4189, n4190, n4192, n4193,
n4194, n4195, n4197, n4198, n4199, n4200, n4202, n4203, n4204, n4205,
n4207, n4208, n4209, n4210, n4212, n4213, n4214, n4215, n4217, n4218,
n4219, n4220, n4222, n4223, n4224, n4225, n4227, n4228, n4229, n4230,
n4232, n4233, n4234, n4235, n4237, n4238, n4239, n4240, n4242, n4243,
n4244, n4245, n4247, n4248, n4249, n4250, n4252, n4253, n4254, n4255,
n4257, n4258, n4259, n4260, n4262, n4263, n4264, n4265, n4267, n4268,
n4269, n4270, n4272, n4273, n4274, n4275, n4277, n4278, n4279, n4280,
n4282, n4283, n4284, n4285, n4287, n4288, n4289, n4290, n4292, n4293,
n4294, n4295, n4297, n4298, n4299, n4301, n4302, n4303, n4305, n4306,
n4307, n4309, n4310, n4311, n4313, n4314, n4315, n4317, n4318, n4319,
n4321, n4322, n4323, n4325, n4326, n4327, n4329, n4330, n4331, n4333,
n4334, n4335, n4337, n4338, n4339, n4341, n4342, n4343, n4345, n4346,
n4347, n4349, n4350, n4351, n4353, n4354, n4355, n4357, n4358, n4359,
n4361, n4362, n4363, n4365, n4366, n4367, n4369, n4370, n4371, n4373,
n4374, n4375, n4377, n4378, n4379, n4381, n4382, n4383, n4385, n4386,
n4387, n4389, n4390, n4391, n4393, n4394, n4395, n4397, n4398, n4399,
n4401, n4402, n4403, n4405, n4406, n4407, n4409, n4410, n4411, n4413,
n4414, n4415, n4417, n4418, n4419, n4421, n4422, n4423, n4424, n4425,
n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
n4576, n4577, n4578, n4580, n4581, n4582, n4583, n4585, n4586, n4587,
n4588, n4590, n4591, n4592, n4593, n4595, n4596, n4597, n4598, n4600,
n4601, n4602, n4603, n4605, n4606, n4607, n4608, n4610, n4611, n4612,
n4613, n4615, n4616, n4617, n4618, n4620, n4621, n4622, n4623, n4625,
n4626, n4627, n4628, n4630, n4631, n4632, n4633, n4635, n4636, n4637,
n4638, n4640, n4641, n4642, n4643, n4645, n4646, n4647, n4648, n4650,
n4651, n4652, n4653, n4655, n4656, n4657, n4658, n4660, n4661, n4662,
n4663, n4665, n4666, n4667, n4668, n4670, n4671, n4672, n4673, n4675;

dff WX547_reg ( clk, reset, WX547, n867 );
dff WX545_reg ( clk, reset, WX545, n31 );
dff WX543_reg ( clk, reset, WX543, n30 );
dff WX541_reg ( clk, reset, WX541, n29 );
dff WX539_reg ( clk, reset, WX539, n28 );
dff WX537_reg ( clk, reset, WX537, n27 );
dff WX535_reg ( clk, reset, WX535, n26 );
dff WX533_reg ( clk, reset, WX533, n25 );
dff WX531_reg ( clk, reset, WX531, n24 );
dff WX529_reg ( clk, reset, WX529, n23 );
dff WX527_reg ( clk, reset, WX527, n22 );
dff WX525_reg ( clk, reset, WX525, n21 );
dff WX523_reg ( clk, reset, WX523, n20 );
dff WX521_reg ( clk, reset, WX521, n19 );
dff WX519_reg ( clk, reset, WX519, n18 );
dff WX517_reg ( clk, reset, WX517, n17 );
dff WX515_reg ( clk, reset, WX515, n16 );
dff WX513_reg ( clk, reset, WX513, n15 );
dff WX511_reg ( clk, reset, WX511, n14 );
dff WX509_reg ( clk, reset, WX509, n13 );
dff WX507_reg ( clk, reset, WX507, n12 );
dff WX505_reg ( clk, reset, WX505, n11 );
dff WX503_reg ( clk, reset, WX503, n10 );
dff WX501_reg ( clk, reset, WX501, n9 );
dff WX499_reg ( clk, reset, WX499, n8 );
dff WX497_reg ( clk, reset, WX497, n7 );
dff WX495_reg ( clk, reset, WX495, n6 );
dff WX493_reg ( clk, reset, WX493, n5 );
dff WX491_reg ( clk, reset, WX491, n4 );
dff WX489_reg ( clk, reset, WX489, n3 );
dff WX487_reg ( clk, reset, WX487, n2 );
dff WX485_reg ( clk, reset, WX485, n1 );
dff WX1840_reg ( clk, reset, WX1840, n1795 );
dff WX1838_reg ( clk, reset, WX1838, n62 );
dff WX1836_reg ( clk, reset, WX1836, n61 );
dff WX1834_reg ( clk, reset, WX1834, n60 );
dff WX1832_reg ( clk, reset, WX1832, n59 );
dff WX1830_reg ( clk, reset, WX1830, n58 );
dff WX1828_reg ( clk, reset, WX1828, n57 );
dff WX1826_reg ( clk, reset, WX1826, n56 );
dff WX1824_reg ( clk, reset, WX1824, n55 );
dff WX1822_reg ( clk, reset, WX1822, n54 );
dff WX1820_reg ( clk, reset, WX1820, n53 );
dff WX1818_reg ( clk, reset, WX1818, n52 );
dff WX1816_reg ( clk, reset, WX1816, n51 );
dff WX1814_reg ( clk, reset, WX1814, n50 );
dff WX1812_reg ( clk, reset, WX1812, n49 );
dff WX1810_reg ( clk, reset, WX1810, n48 );
dff WX1808_reg ( clk, reset, WX1808, n47 );
dff WX1806_reg ( clk, reset, WX1806, n46 );
dff WX1804_reg ( clk, reset, WX1804, n45 );
dff WX1802_reg ( clk, reset, WX1802, n44 );
dff WX1800_reg ( clk, reset, WX1800, n43 );
dff WX1798_reg ( clk, reset, WX1798, n42 );
dff WX1796_reg ( clk, reset, WX1796, n41 );
dff WX1794_reg ( clk, reset, WX1794, n40 );
dff WX1792_reg ( clk, reset, WX1792, n39 );
dff WX1790_reg ( clk, reset, WX1790, n38 );
dff WX1788_reg ( clk, reset, WX1788, n37 );
dff WX1786_reg ( clk, reset, WX1786, n36 );
dff WX1784_reg ( clk, reset, WX1784, n35 );
dff WX1782_reg ( clk, reset, WX1782, n34 );
dff WX1780_reg ( clk, reset, WX1780, n33 );
dff WX1778_reg ( clk, reset, WX1778, n32 );
dff WX3133_reg ( clk, reset, WX3133, n2723 );
dff WX3131_reg ( clk, reset, WX3131, n93 );
dff WX3129_reg ( clk, reset, WX3129, n92 );
dff WX3127_reg ( clk, reset, WX3127, n91 );
dff WX3125_reg ( clk, reset, WX3125, n90 );
dff WX3123_reg ( clk, reset, WX3123, n89 );
dff WX3121_reg ( clk, reset, WX3121, n88 );
dff WX3119_reg ( clk, reset, WX3119, n87 );
dff WX3117_reg ( clk, reset, WX3117, n86 );
dff WX3115_reg ( clk, reset, WX3115, n85 );
dff WX3113_reg ( clk, reset, WX3113, n84 );
dff WX3111_reg ( clk, reset, WX3111, n83 );
dff WX3109_reg ( clk, reset, WX3109, n82 );
dff WX3107_reg ( clk, reset, WX3107, n81 );
dff WX3105_reg ( clk, reset, WX3105, n80 );
dff WX3103_reg ( clk, reset, WX3103, n79 );
dff WX3101_reg ( clk, reset, WX3101, n78 );
dff WX3099_reg ( clk, reset, WX3099, n77 );
dff WX3097_reg ( clk, reset, WX3097, n76 );
dff WX3095_reg ( clk, reset, WX3095, n75 );
dff WX3093_reg ( clk, reset, WX3093, n74 );
dff WX3091_reg ( clk, reset, WX3091, n73 );
dff WX3089_reg ( clk, reset, WX3089, n72 );
dff WX3087_reg ( clk, reset, WX3087, n71 );
dff WX3085_reg ( clk, reset, WX3085, n70 );
dff WX3083_reg ( clk, reset, WX3083, n69 );
dff WX3081_reg ( clk, reset, WX3081, n68 );
dff WX3079_reg ( clk, reset, WX3079, n67 );
dff WX3077_reg ( clk, reset, WX3077, n66 );
dff WX3075_reg ( clk, reset, WX3075, n65 );
dff WX3073_reg ( clk, reset, WX3073, n64 );
dff WX3071_reg ( clk, reset, WX3071, n63 );
dff WX4426_reg ( clk, reset, WX4426, n3651 );
dff WX4424_reg ( clk, reset, WX4424, n124 );
dff WX4422_reg ( clk, reset, WX4422, n123 );
dff WX4420_reg ( clk, reset, WX4420, n122 );
dff WX4418_reg ( clk, reset, WX4418, n121 );
dff WX4416_reg ( clk, reset, WX4416, n120 );
dff WX4414_reg ( clk, reset, WX4414, n119 );
dff WX4412_reg ( clk, reset, WX4412, n118 );
dff WX4410_reg ( clk, reset, WX4410, n117 );
dff WX4408_reg ( clk, reset, WX4408, n116 );
dff WX4406_reg ( clk, reset, WX4406, n115 );
dff WX4404_reg ( clk, reset, WX4404, n114 );
dff WX4402_reg ( clk, reset, WX4402, n113 );
dff WX4400_reg ( clk, reset, WX4400, n112 );
dff WX4398_reg ( clk, reset, WX4398, n111 );
dff WX4396_reg ( clk, reset, WX4396, n110 );
dff WX4394_reg ( clk, reset, WX4394, n109 );
dff WX4392_reg ( clk, reset, WX4392, n108 );
dff WX4390_reg ( clk, reset, WX4390, n107 );
dff WX4388_reg ( clk, reset, WX4388, n106 );
dff WX4386_reg ( clk, reset, WX4386, n105 );
dff WX4384_reg ( clk, reset, WX4384, n104 );
dff WX4382_reg ( clk, reset, WX4382, n103 );
dff WX4380_reg ( clk, reset, WX4380, n102 );
dff WX4378_reg ( clk, reset, WX4378, n101 );
dff WX4376_reg ( clk, reset, WX4376, n100 );
dff WX4374_reg ( clk, reset, WX4374, n99 );
dff WX4372_reg ( clk, reset, WX4372, n98 );
dff WX4370_reg ( clk, reset, WX4370, n97 );
dff WX4368_reg ( clk, reset, WX4368, n96 );
dff WX4366_reg ( clk, reset, WX4366, n95 );
dff WX4364_reg ( clk, reset, WX4364, n94 );
dff WX5719_reg ( clk, reset, WX5719, n4579 );
dff WX5717_reg ( clk, reset, WX5717, n155 );
dff WX5715_reg ( clk, reset, WX5715, n154 );
dff WX5713_reg ( clk, reset, WX5713, n153 );
dff WX5711_reg ( clk, reset, WX5711, n152 );
dff WX5709_reg ( clk, reset, WX5709, n151 );
dff WX5707_reg ( clk, reset, WX5707, n150 );
dff WX5705_reg ( clk, reset, WX5705, n149 );
dff WX5703_reg ( clk, reset, WX5703, n148 );
dff WX5701_reg ( clk, reset, WX5701, n147 );
dff WX5699_reg ( clk, reset, WX5699, n146 );
dff WX5697_reg ( clk, reset, WX5697, n145 );
dff WX5695_reg ( clk, reset, WX5695, n144 );
dff WX5693_reg ( clk, reset, WX5693, n143 );
dff WX5691_reg ( clk, reset, WX5691, n142 );
dff WX5689_reg ( clk, reset, WX5689, n141 );
dff WX5687_reg ( clk, reset, WX5687, n140 );
dff WX5685_reg ( clk, reset, WX5685, n139 );
dff WX5683_reg ( clk, reset, WX5683, n138 );
dff WX5681_reg ( clk, reset, WX5681, n137 );
dff WX5679_reg ( clk, reset, WX5679, n136 );
dff WX5677_reg ( clk, reset, WX5677, n135 );
dff WX5675_reg ( clk, reset, WX5675, n134 );
dff WX5673_reg ( clk, reset, WX5673, n133 );
dff WX5671_reg ( clk, reset, WX5671, n132 );
dff WX5669_reg ( clk, reset, WX5669, n131 );
dff WX5667_reg ( clk, reset, WX5667, n130 );
dff WX5665_reg ( clk, reset, WX5665, n129 );
dff WX5663_reg ( clk, reset, WX5663, n128 );
dff WX5661_reg ( clk, reset, WX5661, n127 );
dff WX5659_reg ( clk, reset, WX5659, n126 );
dff WX5657_reg ( clk, reset, WX5657, n125 );
dff WX7012_reg ( clk, reset, WX7012, n5507 );
dff WX7010_reg ( clk, reset, WX7010, n186 );
dff WX7008_reg ( clk, reset, WX7008, n185 );
dff WX7006_reg ( clk, reset, WX7006, n184 );
dff WX7004_reg ( clk, reset, WX7004, n183 );
dff WX7002_reg ( clk, reset, WX7002, n182 );
dff WX7000_reg ( clk, reset, WX7000, n181 );
dff WX6998_reg ( clk, reset, WX6998, n180 );
dff WX6996_reg ( clk, reset, WX6996, n179 );
dff WX6994_reg ( clk, reset, WX6994, n178 );
dff WX6992_reg ( clk, reset, WX6992, n177 );
dff WX6990_reg ( clk, reset, WX6990, n176 );
dff WX6988_reg ( clk, reset, WX6988, n175 );
dff WX6986_reg ( clk, reset, WX6986, n174 );
dff WX6984_reg ( clk, reset, WX6984, n173 );
dff WX6982_reg ( clk, reset, WX6982, n172 );
dff WX6980_reg ( clk, reset, WX6980, n171 );
dff WX6978_reg ( clk, reset, WX6978, n170 );
dff WX6976_reg ( clk, reset, WX6976, n169 );
dff WX6974_reg ( clk, reset, WX6974, n168 );
dff WX6972_reg ( clk, reset, WX6972, n167 );
dff WX6970_reg ( clk, reset, WX6970, n166 );
dff WX6968_reg ( clk, reset, WX6968, n165 );
dff WX6966_reg ( clk, reset, WX6966, n164 );
dff WX6964_reg ( clk, reset, WX6964, n163 );
dff WX6962_reg ( clk, reset, WX6962, n162 );
dff WX6960_reg ( clk, reset, WX6960, n161 );
dff WX6958_reg ( clk, reset, WX6958, n160 );
dff WX6956_reg ( clk, reset, WX6956, n159 );
dff WX6954_reg ( clk, reset, WX6954, n158 );
dff WX6952_reg ( clk, reset, WX6952, n157 );
dff WX6950_reg ( clk, reset, WX6950, n156 );
dff WX8305_reg ( clk, reset, WX8305, n6435 );
dff WX8303_reg ( clk, reset, WX8303, n217 );
dff WX8301_reg ( clk, reset, WX8301, n216 );
dff WX8299_reg ( clk, reset, WX8299, n215 );
dff WX8297_reg ( clk, reset, WX8297, n214 );
dff WX8295_reg ( clk, reset, WX8295, n213 );
dff WX8293_reg ( clk, reset, WX8293, n212 );
dff WX8291_reg ( clk, reset, WX8291, n211 );
dff WX8289_reg ( clk, reset, WX8289, n210 );
dff WX8287_reg ( clk, reset, WX8287, n209 );
dff WX8285_reg ( clk, reset, WX8285, n208 );
dff WX8283_reg ( clk, reset, WX8283, n207 );
dff WX8281_reg ( clk, reset, WX8281, n206 );
dff WX8279_reg ( clk, reset, WX8279, n205 );
dff WX8277_reg ( clk, reset, WX8277, n204 );
dff WX8275_reg ( clk, reset, WX8275, n203 );
dff WX8273_reg ( clk, reset, WX8273, n202 );
dff WX8271_reg ( clk, reset, WX8271, n201 );
dff WX8269_reg ( clk, reset, WX8269, n200 );
dff WX8267_reg ( clk, reset, WX8267, n199 );
dff WX8265_reg ( clk, reset, WX8265, n198 );
dff WX8263_reg ( clk, reset, WX8263, n197 );
dff WX8261_reg ( clk, reset, WX8261, n196 );
dff WX8259_reg ( clk, reset, WX8259, n195 );
dff WX8257_reg ( clk, reset, WX8257, n194 );
dff WX8255_reg ( clk, reset, WX8255, n193 );
dff WX8253_reg ( clk, reset, WX8253, n192 );
dff WX8251_reg ( clk, reset, WX8251, n191 );
dff WX8249_reg ( clk, reset, WX8249, n190 );
dff WX8247_reg ( clk, reset, WX8247, n189 );
dff WX8245_reg ( clk, reset, WX8245, n188 );
dff WX8243_reg ( clk, reset, WX8243, n187 );
dff WX9598_reg ( clk, reset, WX9598, n7363 );
dff WX9596_reg ( clk, reset, WX9596, n248 );
dff WX9594_reg ( clk, reset, WX9594, n247 );
dff WX9592_reg ( clk, reset, WX9592, n246 );
dff WX9590_reg ( clk, reset, WX9590, n245 );
dff WX9588_reg ( clk, reset, WX9588, n244 );
dff WX9586_reg ( clk, reset, WX9586, n243 );
dff WX9584_reg ( clk, reset, WX9584, n242 );
dff WX9582_reg ( clk, reset, WX9582, n241 );
dff WX9580_reg ( clk, reset, WX9580, n240 );
dff WX9578_reg ( clk, reset, WX9578, n239 );
dff WX9576_reg ( clk, reset, WX9576, n238 );
dff WX9574_reg ( clk, reset, WX9574, n237 );
dff WX9572_reg ( clk, reset, WX9572, n236 );
dff WX9570_reg ( clk, reset, WX9570, n235 );
dff WX9568_reg ( clk, reset, WX9568, n234 );
dff WX9566_reg ( clk, reset, WX9566, n233 );
dff WX9564_reg ( clk, reset, WX9564, n232 );
dff WX9562_reg ( clk, reset, WX9562, n231 );
dff WX9560_reg ( clk, reset, WX9560, n230 );
dff WX9558_reg ( clk, reset, WX9558, n229 );
dff WX9556_reg ( clk, reset, WX9556, n228 );
dff WX9554_reg ( clk, reset, WX9554, n227 );
dff WX9552_reg ( clk, reset, WX9552, n226 );
dff WX9550_reg ( clk, reset, WX9550, n225 );
dff WX9548_reg ( clk, reset, WX9548, n224 );
dff WX9546_reg ( clk, reset, WX9546, n223 );
dff WX9544_reg ( clk, reset, WX9544, n222 );
dff WX9542_reg ( clk, reset, WX9542, n221 );
dff WX9540_reg ( clk, reset, WX9540, n220 );
dff WX9538_reg ( clk, reset, WX9538, n219 );
dff WX9536_reg ( clk, reset, WX9536, n218 );
dff WX10891_reg ( clk, reset, WX10891, n8291 );
dff WX10889_reg ( clk, reset, WX10889, n279 );
dff WX10887_reg ( clk, reset, WX10887, n278 );
dff WX10885_reg ( clk, reset, WX10885, n277 );
dff WX10883_reg ( clk, reset, WX10883, n276 );
dff WX10881_reg ( clk, reset, WX10881, n275 );
dff WX10879_reg ( clk, reset, WX10879, n274 );
dff WX10877_reg ( clk, reset, WX10877, n273 );
dff WX10875_reg ( clk, reset, WX10875, n272 );
dff WX10873_reg ( clk, reset, WX10873, n271 );
dff WX10871_reg ( clk, reset, WX10871, n270 );
dff WX10869_reg ( clk, reset, WX10869, n269 );
dff WX10867_reg ( clk, reset, WX10867, n268 );
dff WX10865_reg ( clk, reset, WX10865, n267 );
dff WX10863_reg ( clk, reset, WX10863, n266 );
dff WX10861_reg ( clk, reset, WX10861, n265 );
dff WX10859_reg ( clk, reset, WX10859, n264 );
dff WX10857_reg ( clk, reset, WX10857, n263 );
dff WX10855_reg ( clk, reset, WX10855, n262 );
dff WX10853_reg ( clk, reset, WX10853, n261 );
dff WX10851_reg ( clk, reset, WX10851, n260 );
dff WX10849_reg ( clk, reset, WX10849, n259 );
dff WX10847_reg ( clk, reset, WX10847, n258 );
dff WX10845_reg ( clk, reset, WX10845, n257 );
dff WX10843_reg ( clk, reset, WX10843, n256 );
dff WX10841_reg ( clk, reset, WX10841, n255 );
dff WX10839_reg ( clk, reset, WX10839, n254 );
dff WX10837_reg ( clk, reset, WX10837, n253 );
dff WX10835_reg ( clk, reset, WX10835, n252 );
dff WX10833_reg ( clk, reset, WX10833, n251 );
dff WX10831_reg ( clk, reset, WX10831, n250 );
dff WX10829_reg ( clk, reset, WX10829, n249 );
dff CRC_OUT_1_31_reg ( clk, reset, CRC_OUT_1_31, n9060 );
dff CRC_OUT_1_0_reg ( clk, reset, CRC_OUT_1_0, n8936 );
dff CRC_OUT_1_1_reg ( clk, reset, CRC_OUT_1_1, n8940 );
dff CRC_OUT_1_2_reg ( clk, reset, CRC_OUT_1_2, n8944 );
dff CRC_OUT_1_3_reg ( clk, reset, CRC_OUT_1_3, n8948 );
dff CRC_OUT_1_4_reg ( clk, reset, CRC_OUT_1_4, n8952 );
dff CRC_OUT_1_5_reg ( clk, reset, CRC_OUT_1_5, n8956 );
dff CRC_OUT_1_6_reg ( clk, reset, CRC_OUT_1_6, n8960 );
dff CRC_OUT_1_7_reg ( clk, reset, CRC_OUT_1_7, n8964 );
dff CRC_OUT_1_8_reg ( clk, reset, CRC_OUT_1_8, n8968 );
dff CRC_OUT_1_9_reg ( clk, reset, CRC_OUT_1_9, n8972 );
dff CRC_OUT_1_10_reg ( clk, reset, CRC_OUT_1_10, n8976 );
dff CRC_OUT_1_11_reg ( clk, reset, CRC_OUT_1_11, n8980 );
dff CRC_OUT_1_12_reg ( clk, reset, CRC_OUT_1_12, n8984 );
dff CRC_OUT_1_13_reg ( clk, reset, CRC_OUT_1_13, n8988 );
dff CRC_OUT_1_14_reg ( clk, reset, CRC_OUT_1_14, n8992 );
dff CRC_OUT_1_15_reg ( clk, reset, CRC_OUT_1_15, n8996 );
dff CRC_OUT_1_16_reg ( clk, reset, CRC_OUT_1_16, n9000 );
dff CRC_OUT_1_17_reg ( clk, reset, CRC_OUT_1_17, n9004 );
dff CRC_OUT_1_18_reg ( clk, reset, CRC_OUT_1_18, n9008 );
dff CRC_OUT_1_19_reg ( clk, reset, CRC_OUT_1_19, n9012 );
dff CRC_OUT_1_20_reg ( clk, reset, CRC_OUT_1_20, n9016 );
dff CRC_OUT_1_21_reg ( clk, reset, CRC_OUT_1_21, n9020 );
dff CRC_OUT_1_22_reg ( clk, reset, CRC_OUT_1_22, n9024 );
dff CRC_OUT_1_23_reg ( clk, reset, CRC_OUT_1_23, n9028 );
dff CRC_OUT_1_24_reg ( clk, reset, CRC_OUT_1_24, n9032 );
dff CRC_OUT_1_25_reg ( clk, reset, CRC_OUT_1_25, n9036 );
dff CRC_OUT_1_26_reg ( clk, reset, CRC_OUT_1_26, n9040 );
dff CRC_OUT_1_27_reg ( clk, reset, CRC_OUT_1_27, n9044 );
dff CRC_OUT_1_28_reg ( clk, reset, CRC_OUT_1_28, n9048 );
dff CRC_OUT_1_29_reg ( clk, reset, CRC_OUT_1_29, n9052 );
dff CRC_OUT_1_30_reg ( clk, reset, CRC_OUT_1_30, n9056 );
dff WX10991_reg ( clk, reset, WX10991, n8301 );
dff WX11055_reg ( clk, reset, WX11055, n8461 );
dff WX11119_reg ( clk, reset, WX11119, n8621 );
dff WX11183_reg ( clk, reset, WX11183, n8781 );
dff WX10993_reg ( clk, reset, WX10993, n8306 );
dff WX11057_reg ( clk, reset, WX11057, n8466 );
dff WX11121_reg ( clk, reset, WX11121, n8626 );
dff WX11185_reg ( clk, reset, WX11185, n8786 );
dff WX10995_reg ( clk, reset, WX10995, n8311 );
dff WX11059_reg ( clk, reset, WX11059, n8471 );
dff WX11123_reg ( clk, reset, WX11123, n8631 );
dff WX11187_reg ( clk, reset, WX11187, n8791 );
dff WX10997_reg ( clk, reset, WX10997, n8316 );
dff WX11061_reg ( clk, reset, WX11061, n8476 );
dff WX11125_reg ( clk, reset, WX11125, n8636 );
dff WX11189_reg ( clk, reset, WX11189, n8796 );
dff WX10999_reg ( clk, reset, WX10999, n8321 );
dff WX11063_reg ( clk, reset, WX11063, n8481 );
dff WX11127_reg ( clk, reset, WX11127, n8641 );
dff WX11191_reg ( clk, reset, WX11191, n8801 );
dff WX11001_reg ( clk, reset, WX11001, n8326 );
dff WX11065_reg ( clk, reset, WX11065, n8486 );
dff WX11129_reg ( clk, reset, WX11129, n8646 );
dff WX11193_reg ( clk, reset, WX11193, n8806 );
dff WX11003_reg ( clk, reset, WX11003, n8331 );
dff WX11067_reg ( clk, reset, WX11067, n8491 );
dff WX11131_reg ( clk, reset, WX11131, n8651 );
dff WX11195_reg ( clk, reset, WX11195, n8811 );
dff WX11005_reg ( clk, reset, WX11005, n8336 );
dff WX11069_reg ( clk, reset, WX11069, n8496 );
dff WX11133_reg ( clk, reset, WX11133, n8656 );
dff WX11197_reg ( clk, reset, WX11197, n8816 );
dff WX11007_reg ( clk, reset, WX11007, n8341 );
dff WX11071_reg ( clk, reset, WX11071, n8501 );
dff WX11135_reg ( clk, reset, WX11135, n8661 );
dff WX11199_reg ( clk, reset, WX11199, n8821 );
dff WX11009_reg ( clk, reset, WX11009, n8346 );
dff WX11073_reg ( clk, reset, WX11073, n8506 );
dff WX11137_reg ( clk, reset, WX11137, n8666 );
dff WX11201_reg ( clk, reset, WX11201, n8826 );
dff WX11011_reg ( clk, reset, WX11011, n8351 );
dff WX11075_reg ( clk, reset, WX11075, n8511 );
dff WX11139_reg ( clk, reset, WX11139, n8671 );
dff WX11203_reg ( clk, reset, WX11203, n8831 );
dff WX11013_reg ( clk, reset, WX11013, n8356 );
dff WX11077_reg ( clk, reset, WX11077, n8516 );
dff WX11141_reg ( clk, reset, WX11141, n8676 );
dff WX11205_reg ( clk, reset, WX11205, n8836 );
dff WX11015_reg ( clk, reset, WX11015, n8361 );
dff WX11079_reg ( clk, reset, WX11079, n8521 );
dff WX11143_reg ( clk, reset, WX11143, n8681 );
dff WX11207_reg ( clk, reset, WX11207, n8841 );
dff WX11017_reg ( clk, reset, WX11017, n8366 );
dff WX11081_reg ( clk, reset, WX11081, n8526 );
dff WX11145_reg ( clk, reset, WX11145, n8686 );
dff WX11209_reg ( clk, reset, WX11209, n8846 );
dff WX11019_reg ( clk, reset, WX11019, n8371 );
dff WX11083_reg ( clk, reset, WX11083, n8531 );
dff WX11147_reg ( clk, reset, WX11147, n8691 );
dff WX11211_reg ( clk, reset, WX11211, n8851 );
dff WX11021_reg ( clk, reset, WX11021, n8376 );
dff WX11085_reg ( clk, reset, WX11085, n8536 );
dff WX11149_reg ( clk, reset, WX11149, n8696 );
dff WX11213_reg ( clk, reset, WX11213, n8856 );
dff WX11023_reg ( clk, reset, WX11023, n8381 );
dff WX11087_reg ( clk, reset, WX11087, n8541 );
dff WX11151_reg ( clk, reset, WX11151, n8701 );
dff WX11215_reg ( clk, reset, WX11215, n8861 );
dff WX11025_reg ( clk, reset, WX11025, n8386 );
dff WX11089_reg ( clk, reset, WX11089, n8546 );
dff WX11153_reg ( clk, reset, WX11153, n8706 );
dff WX11217_reg ( clk, reset, WX11217, n8866 );
dff WX11027_reg ( clk, reset, WX11027, n8391 );
dff WX11091_reg ( clk, reset, WX11091, n8551 );
dff WX11155_reg ( clk, reset, WX11155, n8711 );
dff WX11219_reg ( clk, reset, WX11219, n8871 );
dff WX11029_reg ( clk, reset, WX11029, n8396 );
dff WX11093_reg ( clk, reset, WX11093, n8556 );
dff WX11157_reg ( clk, reset, WX11157, n8716 );
dff WX11221_reg ( clk, reset, WX11221, n8876 );
dff WX11031_reg ( clk, reset, WX11031, n8401 );
dff WX11095_reg ( clk, reset, WX11095, n8561 );
dff WX11159_reg ( clk, reset, WX11159, n8721 );
dff WX11223_reg ( clk, reset, WX11223, n8881 );
dff WX11033_reg ( clk, reset, WX11033, n8406 );
dff WX11097_reg ( clk, reset, WX11097, n8566 );
dff WX11161_reg ( clk, reset, WX11161, n8726 );
dff WX11225_reg ( clk, reset, WX11225, n8886 );
dff WX11035_reg ( clk, reset, WX11035, n8411 );
dff WX11099_reg ( clk, reset, WX11099, n8571 );
dff WX11163_reg ( clk, reset, WX11163, n8731 );
dff WX11227_reg ( clk, reset, WX11227, n8891 );
dff WX11037_reg ( clk, reset, WX11037, n8416 );
dff WX11101_reg ( clk, reset, WX11101, n8576 );
dff WX11165_reg ( clk, reset, WX11165, n8736 );
dff WX11229_reg ( clk, reset, WX11229, n8896 );
dff WX11039_reg ( clk, reset, WX11039, n8421 );
dff WX11103_reg ( clk, reset, WX11103, n8581 );
dff WX11167_reg ( clk, reset, WX11167, n8741 );
dff WX11231_reg ( clk, reset, WX11231, n8901 );
dff WX11041_reg ( clk, reset, WX11041, n8426 );
dff WX11105_reg ( clk, reset, WX11105, n8586 );
dff WX11169_reg ( clk, reset, WX11169, n8746 );
dff WX11233_reg ( clk, reset, WX11233, n8906 );
dff WX11043_reg ( clk, reset, WX11043, n8431 );
dff WX11107_reg ( clk, reset, WX11107, n8591 );
dff WX11171_reg ( clk, reset, WX11171, n8751 );
dff WX11235_reg ( clk, reset, WX11235, n8911 );
dff WX11045_reg ( clk, reset, WX11045, n8436 );
dff WX11109_reg ( clk, reset, WX11109, n8596 );
dff WX11173_reg ( clk, reset, WX11173, n8756 );
dff WX11237_reg ( clk, reset, WX11237, n8916 );
dff WX11047_reg ( clk, reset, WX11047, n8441 );
dff WX11111_reg ( clk, reset, WX11111, n8601 );
dff WX11175_reg ( clk, reset, WX11175, n8761 );
dff WX11239_reg ( clk, reset, WX11239, n8921 );
dff WX11049_reg ( clk, reset, WX11049, n8446 );
dff WX11113_reg ( clk, reset, WX11113, n8606 );
dff WX11177_reg ( clk, reset, WX11177, n8766 );
dff WX11241_reg ( clk, reset, WX11241, n8926 );
dff WX11051_reg ( clk, reset, WX11051, n8451 );
dff WX11115_reg ( clk, reset, WX11115, n8611 );
dff WX11179_reg ( clk, reset, WX11179, n8771 );
dff WX11243_reg ( clk, reset, WX11243, n8931 );
dff WX10989_reg ( clk, reset, WX10989, n8296 );
dff WX11053_reg ( clk, reset, WX11053, n8456 );
dff WX11117_reg ( clk, reset, WX11117, n8616 );
dff WX11181_reg ( clk, reset, WX11181, n8776 );
dff WX9696_reg ( clk, reset, WX9696, n7368 );
dff WX9760_reg ( clk, reset, WX9760, n7528 );
dff WX9824_reg ( clk, reset, WX9824, n7688 );
dff WX9888_reg ( clk, reset, WX9888, n7848 );
dff CRC_OUT_2_31_reg ( clk, reset, CRC_OUT_2_31, n8132 );
dff CRC_OUT_2_0_reg ( clk, reset, CRC_OUT_2_0, n8008 );
dff CRC_OUT_2_1_reg ( clk, reset, CRC_OUT_2_1, n8012 );
dff CRC_OUT_2_2_reg ( clk, reset, CRC_OUT_2_2, n8016 );
dff CRC_OUT_2_3_reg ( clk, reset, CRC_OUT_2_3, n8020 );
dff CRC_OUT_2_4_reg ( clk, reset, CRC_OUT_2_4, n8024 );
dff CRC_OUT_2_5_reg ( clk, reset, CRC_OUT_2_5, n8028 );
dff CRC_OUT_2_6_reg ( clk, reset, CRC_OUT_2_6, n8032 );
dff CRC_OUT_2_7_reg ( clk, reset, CRC_OUT_2_7, n8036 );
dff CRC_OUT_2_8_reg ( clk, reset, CRC_OUT_2_8, n8040 );
dff CRC_OUT_2_9_reg ( clk, reset, CRC_OUT_2_9, n8044 );
dff CRC_OUT_2_10_reg ( clk, reset, CRC_OUT_2_10, n8048 );
dff CRC_OUT_2_11_reg ( clk, reset, CRC_OUT_2_11, n8052 );
dff CRC_OUT_2_12_reg ( clk, reset, CRC_OUT_2_12, n8056 );
dff CRC_OUT_2_13_reg ( clk, reset, CRC_OUT_2_13, n8060 );
dff CRC_OUT_2_14_reg ( clk, reset, CRC_OUT_2_14, n8064 );
dff CRC_OUT_2_15_reg ( clk, reset, CRC_OUT_2_15, n8068 );
dff CRC_OUT_2_16_reg ( clk, reset, CRC_OUT_2_16, n8072 );
dff CRC_OUT_2_17_reg ( clk, reset, CRC_OUT_2_17, n8076 );
dff CRC_OUT_2_18_reg ( clk, reset, CRC_OUT_2_18, n8080 );
dff CRC_OUT_2_19_reg ( clk, reset, CRC_OUT_2_19, n8084 );
dff CRC_OUT_2_20_reg ( clk, reset, CRC_OUT_2_20, n8088 );
dff CRC_OUT_2_21_reg ( clk, reset, CRC_OUT_2_21, n8092 );
dff CRC_OUT_2_22_reg ( clk, reset, CRC_OUT_2_22, n8096 );
dff CRC_OUT_2_23_reg ( clk, reset, CRC_OUT_2_23, n8100 );
dff CRC_OUT_2_24_reg ( clk, reset, CRC_OUT_2_24, n8104 );
dff CRC_OUT_2_25_reg ( clk, reset, CRC_OUT_2_25, n8108 );
dff CRC_OUT_2_26_reg ( clk, reset, CRC_OUT_2_26, n8112 );
dff CRC_OUT_2_27_reg ( clk, reset, CRC_OUT_2_27, n8116 );
dff CRC_OUT_2_28_reg ( clk, reset, CRC_OUT_2_28, n8120 );
dff CRC_OUT_2_29_reg ( clk, reset, CRC_OUT_2_29, n8124 );
dff CRC_OUT_2_30_reg ( clk, reset, CRC_OUT_2_30, n8128 );
dff WX9698_reg ( clk, reset, WX9698, n7373 );
dff WX9762_reg ( clk, reset, WX9762, n7533 );
dff WX9826_reg ( clk, reset, WX9826, n7693 );
dff WX9890_reg ( clk, reset, WX9890, n7853 );
dff WX9700_reg ( clk, reset, WX9700, n7378 );
dff WX9764_reg ( clk, reset, WX9764, n7538 );
dff WX9828_reg ( clk, reset, WX9828, n7698 );
dff WX9892_reg ( clk, reset, WX9892, n7858 );
dff WX9702_reg ( clk, reset, WX9702, n7383 );
dff WX9766_reg ( clk, reset, WX9766, n7543 );
dff WX9830_reg ( clk, reset, WX9830, n7703 );
dff WX9894_reg ( clk, reset, WX9894, n7863 );
dff WX9704_reg ( clk, reset, WX9704, n7388 );
dff WX9768_reg ( clk, reset, WX9768, n7548 );
dff WX9832_reg ( clk, reset, WX9832, n7708 );
dff WX9896_reg ( clk, reset, WX9896, n7868 );
dff WX9706_reg ( clk, reset, WX9706, n7393 );
dff WX9770_reg ( clk, reset, WX9770, n7553 );
dff WX9834_reg ( clk, reset, WX9834, n7713 );
dff WX9898_reg ( clk, reset, WX9898, n7873 );
dff WX9708_reg ( clk, reset, WX9708, n7398 );
dff WX9772_reg ( clk, reset, WX9772, n7558 );
dff WX9836_reg ( clk, reset, WX9836, n7718 );
dff WX9900_reg ( clk, reset, WX9900, n7878 );
dff WX9710_reg ( clk, reset, WX9710, n7403 );
dff WX9774_reg ( clk, reset, WX9774, n7563 );
dff WX9838_reg ( clk, reset, WX9838, n7723 );
dff WX9902_reg ( clk, reset, WX9902, n7883 );
dff WX9712_reg ( clk, reset, WX9712, n7408 );
dff WX9776_reg ( clk, reset, WX9776, n7568 );
dff WX9840_reg ( clk, reset, WX9840, n7728 );
dff WX9904_reg ( clk, reset, WX9904, n7888 );
dff WX9714_reg ( clk, reset, WX9714, n7413 );
dff WX9778_reg ( clk, reset, WX9778, n7573 );
dff WX9842_reg ( clk, reset, WX9842, n7733 );
dff WX9906_reg ( clk, reset, WX9906, n7893 );
dff WX9716_reg ( clk, reset, WX9716, n7418 );
dff WX9780_reg ( clk, reset, WX9780, n7578 );
dff WX9844_reg ( clk, reset, WX9844, n7738 );
dff WX9908_reg ( clk, reset, WX9908, n7898 );
dff WX9718_reg ( clk, reset, WX9718, n7423 );
dff WX9782_reg ( clk, reset, WX9782, n7583 );
dff WX9846_reg ( clk, reset, WX9846, n7743 );
dff WX9910_reg ( clk, reset, WX9910, n7903 );
dff WX9720_reg ( clk, reset, WX9720, n7428 );
dff WX9784_reg ( clk, reset, WX9784, n7588 );
dff WX9848_reg ( clk, reset, WX9848, n7748 );
dff WX9912_reg ( clk, reset, WX9912, n7908 );
dff WX9722_reg ( clk, reset, WX9722, n7433 );
dff WX9786_reg ( clk, reset, WX9786, n7593 );
dff WX9850_reg ( clk, reset, WX9850, n7753 );
dff WX9914_reg ( clk, reset, WX9914, n7913 );
dff WX9724_reg ( clk, reset, WX9724, n7438 );
dff WX9788_reg ( clk, reset, WX9788, n7598 );
dff WX9852_reg ( clk, reset, WX9852, n7758 );
dff WX9916_reg ( clk, reset, WX9916, n7918 );
dff WX9726_reg ( clk, reset, WX9726, n7443 );
dff WX9790_reg ( clk, reset, WX9790, n7603 );
dff WX9854_reg ( clk, reset, WX9854, n7763 );
dff WX9918_reg ( clk, reset, WX9918, n7923 );
dff WX9728_reg ( clk, reset, WX9728, n7448 );
dff WX9792_reg ( clk, reset, WX9792, n7608 );
dff WX9856_reg ( clk, reset, WX9856, n7768 );
dff WX9920_reg ( clk, reset, WX9920, n7928 );
dff WX9730_reg ( clk, reset, WX9730, n7453 );
dff WX9794_reg ( clk, reset, WX9794, n7613 );
dff WX9858_reg ( clk, reset, WX9858, n7773 );
dff WX9922_reg ( clk, reset, WX9922, n7933 );
dff WX9732_reg ( clk, reset, WX9732, n7458 );
dff WX9796_reg ( clk, reset, WX9796, n7618 );
dff WX9860_reg ( clk, reset, WX9860, n7778 );
dff WX9924_reg ( clk, reset, WX9924, n7938 );
dff WX9734_reg ( clk, reset, WX9734, n7463 );
dff WX9798_reg ( clk, reset, WX9798, n7623 );
dff WX9862_reg ( clk, reset, WX9862, n7783 );
dff WX9926_reg ( clk, reset, WX9926, n7943 );
dff WX9736_reg ( clk, reset, WX9736, n7468 );
dff WX9800_reg ( clk, reset, WX9800, n7628 );
dff WX9864_reg ( clk, reset, WX9864, n7788 );
dff WX9928_reg ( clk, reset, WX9928, n7948 );
dff WX9738_reg ( clk, reset, WX9738, n7473 );
dff WX9802_reg ( clk, reset, WX9802, n7633 );
dff WX9866_reg ( clk, reset, WX9866, n7793 );
dff WX9930_reg ( clk, reset, WX9930, n7953 );
dff WX9740_reg ( clk, reset, WX9740, n7478 );
dff WX9804_reg ( clk, reset, WX9804, n7638 );
dff WX9868_reg ( clk, reset, WX9868, n7798 );
dff WX9932_reg ( clk, reset, WX9932, n7958 );
dff WX9742_reg ( clk, reset, WX9742, n7483 );
dff WX9806_reg ( clk, reset, WX9806, n7643 );
dff WX9870_reg ( clk, reset, WX9870, n7803 );
dff WX9934_reg ( clk, reset, WX9934, n7963 );
dff WX9744_reg ( clk, reset, WX9744, n7488 );
dff WX9808_reg ( clk, reset, WX9808, n7648 );
dff WX9872_reg ( clk, reset, WX9872, n7808 );
dff WX9936_reg ( clk, reset, WX9936, n7968 );
dff WX9746_reg ( clk, reset, WX9746, n7493 );
dff WX9810_reg ( clk, reset, WX9810, n7653 );
dff WX9874_reg ( clk, reset, WX9874, n7813 );
dff WX9938_reg ( clk, reset, WX9938, n7973 );
dff WX9748_reg ( clk, reset, WX9748, n7498 );
dff WX9812_reg ( clk, reset, WX9812, n7658 );
dff WX9876_reg ( clk, reset, WX9876, n7818 );
dff WX9940_reg ( clk, reset, WX9940, n7978 );
dff WX9750_reg ( clk, reset, WX9750, n7503 );
dff WX9814_reg ( clk, reset, WX9814, n7663 );
dff WX9878_reg ( clk, reset, WX9878, n7823 );
dff WX9942_reg ( clk, reset, WX9942, n7983 );
dff WX9752_reg ( clk, reset, WX9752, n7508 );
dff WX9816_reg ( clk, reset, WX9816, n7668 );
dff WX9880_reg ( clk, reset, WX9880, n7828 );
dff WX9944_reg ( clk, reset, WX9944, n7988 );
dff WX9754_reg ( clk, reset, WX9754, n7513 );
dff WX9818_reg ( clk, reset, WX9818, n7673 );
dff WX9882_reg ( clk, reset, WX9882, n7833 );
dff WX9946_reg ( clk, reset, WX9946, n7993 );
dff WX9756_reg ( clk, reset, WX9756, n7518 );
dff WX9820_reg ( clk, reset, WX9820, n7678 );
dff WX9884_reg ( clk, reset, WX9884, n7838 );
dff WX9948_reg ( clk, reset, WX9948, n7998 );
dff WX9758_reg ( clk, reset, WX9758, n7523 );
dff WX9822_reg ( clk, reset, WX9822, n7683 );
dff WX9886_reg ( clk, reset, WX9886, n7843 );
dff WX9950_reg ( clk, reset, WX9950, n8003 );
dff WX8403_reg ( clk, reset, WX8403, n6440 );
dff WX8467_reg ( clk, reset, WX8467, n6600 );
dff WX8531_reg ( clk, reset, WX8531, n6760 );
dff WX8595_reg ( clk, reset, WX8595, n6920 );
dff CRC_OUT_3_31_reg ( clk, reset, CRC_OUT_3_31, n7204 );
dff CRC_OUT_3_0_reg ( clk, reset, CRC_OUT_3_0, n7080 );
dff CRC_OUT_3_1_reg ( clk, reset, CRC_OUT_3_1, n7084 );
dff CRC_OUT_3_2_reg ( clk, reset, CRC_OUT_3_2, n7088 );
dff CRC_OUT_3_3_reg ( clk, reset, CRC_OUT_3_3, n7092 );
dff CRC_OUT_3_4_reg ( clk, reset, CRC_OUT_3_4, n7096 );
dff CRC_OUT_3_5_reg ( clk, reset, CRC_OUT_3_5, n7100 );
dff CRC_OUT_3_6_reg ( clk, reset, CRC_OUT_3_6, n7104 );
dff CRC_OUT_3_7_reg ( clk, reset, CRC_OUT_3_7, n7108 );
dff CRC_OUT_3_8_reg ( clk, reset, CRC_OUT_3_8, n7112 );
dff CRC_OUT_3_9_reg ( clk, reset, CRC_OUT_3_9, n7116 );
dff CRC_OUT_3_10_reg ( clk, reset, CRC_OUT_3_10, n7120 );
dff CRC_OUT_3_11_reg ( clk, reset, CRC_OUT_3_11, n7124 );
dff CRC_OUT_3_12_reg ( clk, reset, CRC_OUT_3_12, n7128 );
dff CRC_OUT_3_13_reg ( clk, reset, CRC_OUT_3_13, n7132 );
dff CRC_OUT_3_14_reg ( clk, reset, CRC_OUT_3_14, n7136 );
dff CRC_OUT_3_15_reg ( clk, reset, CRC_OUT_3_15, n7140 );
dff CRC_OUT_3_16_reg ( clk, reset, CRC_OUT_3_16, n7144 );
dff CRC_OUT_3_17_reg ( clk, reset, CRC_OUT_3_17, n7148 );
dff CRC_OUT_3_18_reg ( clk, reset, CRC_OUT_3_18, n7152 );
dff CRC_OUT_3_19_reg ( clk, reset, CRC_OUT_3_19, n7156 );
dff CRC_OUT_3_20_reg ( clk, reset, CRC_OUT_3_20, n7160 );
dff CRC_OUT_3_21_reg ( clk, reset, CRC_OUT_3_21, n7164 );
dff CRC_OUT_3_22_reg ( clk, reset, CRC_OUT_3_22, n7168 );
dff CRC_OUT_3_23_reg ( clk, reset, CRC_OUT_3_23, n7172 );
dff CRC_OUT_3_24_reg ( clk, reset, CRC_OUT_3_24, n7176 );
dff CRC_OUT_3_25_reg ( clk, reset, CRC_OUT_3_25, n7180 );
dff CRC_OUT_3_26_reg ( clk, reset, CRC_OUT_3_26, n7184 );
dff CRC_OUT_3_27_reg ( clk, reset, CRC_OUT_3_27, n7188 );
dff CRC_OUT_3_28_reg ( clk, reset, CRC_OUT_3_28, n7192 );
dff CRC_OUT_3_29_reg ( clk, reset, CRC_OUT_3_29, n7196 );
dff CRC_OUT_3_30_reg ( clk, reset, CRC_OUT_3_30, n7200 );
dff WX8405_reg ( clk, reset, WX8405, n6445 );
dff WX8469_reg ( clk, reset, WX8469, n6605 );
dff WX8533_reg ( clk, reset, WX8533, n6765 );
dff WX8597_reg ( clk, reset, WX8597, n6925 );
dff WX8407_reg ( clk, reset, WX8407, n6450 );
dff WX8471_reg ( clk, reset, WX8471, n6610 );
dff WX8535_reg ( clk, reset, WX8535, n6770 );
dff WX8599_reg ( clk, reset, WX8599, n6930 );
dff WX8409_reg ( clk, reset, WX8409, n6455 );
dff WX8473_reg ( clk, reset, WX8473, n6615 );
dff WX8537_reg ( clk, reset, WX8537, n6775 );
dff WX8601_reg ( clk, reset, WX8601, n6935 );
dff WX8411_reg ( clk, reset, WX8411, n6460 );
dff WX8475_reg ( clk, reset, WX8475, n6620 );
dff WX8539_reg ( clk, reset, WX8539, n6780 );
dff WX8603_reg ( clk, reset, WX8603, n6940 );
dff WX8413_reg ( clk, reset, WX8413, n6465 );
dff WX8477_reg ( clk, reset, WX8477, n6625 );
dff WX8541_reg ( clk, reset, WX8541, n6785 );
dff WX8605_reg ( clk, reset, WX8605, n6945 );
dff WX8415_reg ( clk, reset, WX8415, n6470 );
dff WX8479_reg ( clk, reset, WX8479, n6630 );
dff WX8543_reg ( clk, reset, WX8543, n6790 );
dff WX8607_reg ( clk, reset, WX8607, n6950 );
dff WX8417_reg ( clk, reset, WX8417, n6475 );
dff WX8481_reg ( clk, reset, WX8481, n6635 );
dff WX8545_reg ( clk, reset, WX8545, n6795 );
dff WX8609_reg ( clk, reset, WX8609, n6955 );
dff WX8419_reg ( clk, reset, WX8419, n6480 );
dff WX8483_reg ( clk, reset, WX8483, n6640 );
dff WX8547_reg ( clk, reset, WX8547, n6800 );
dff WX8611_reg ( clk, reset, WX8611, n6960 );
dff WX8421_reg ( clk, reset, WX8421, n6485 );
dff WX8485_reg ( clk, reset, WX8485, n6645 );
dff WX8549_reg ( clk, reset, WX8549, n6805 );
dff WX8613_reg ( clk, reset, WX8613, n6965 );
dff WX8423_reg ( clk, reset, WX8423, n6490 );
dff WX8487_reg ( clk, reset, WX8487, n6650 );
dff WX8551_reg ( clk, reset, WX8551, n6810 );
dff WX8615_reg ( clk, reset, WX8615, n6970 );
dff WX8425_reg ( clk, reset, WX8425, n6495 );
dff WX8489_reg ( clk, reset, WX8489, n6655 );
dff WX8553_reg ( clk, reset, WX8553, n6815 );
dff WX8617_reg ( clk, reset, WX8617, n6975 );
dff WX8427_reg ( clk, reset, WX8427, n6500 );
dff WX8491_reg ( clk, reset, WX8491, n6660 );
dff WX8555_reg ( clk, reset, WX8555, n6820 );
dff WX8619_reg ( clk, reset, WX8619, n6980 );
dff WX8429_reg ( clk, reset, WX8429, n6505 );
dff WX8493_reg ( clk, reset, WX8493, n6665 );
dff WX8557_reg ( clk, reset, WX8557, n6825 );
dff WX8621_reg ( clk, reset, WX8621, n6985 );
dff WX8431_reg ( clk, reset, WX8431, n6510 );
dff WX8495_reg ( clk, reset, WX8495, n6670 );
dff WX8559_reg ( clk, reset, WX8559, n6830 );
dff WX8623_reg ( clk, reset, WX8623, n6990 );
dff WX8433_reg ( clk, reset, WX8433, n6515 );
dff WX8497_reg ( clk, reset, WX8497, n6675 );
dff WX8561_reg ( clk, reset, WX8561, n6835 );
dff WX8625_reg ( clk, reset, WX8625, n6995 );
dff WX8435_reg ( clk, reset, WX8435, n6520 );
dff WX8499_reg ( clk, reset, WX8499, n6680 );
dff WX8563_reg ( clk, reset, WX8563, n6840 );
dff WX8627_reg ( clk, reset, WX8627, n7000 );
dff WX8437_reg ( clk, reset, WX8437, n6525 );
dff WX8501_reg ( clk, reset, WX8501, n6685 );
dff WX8565_reg ( clk, reset, WX8565, n6845 );
dff WX8629_reg ( clk, reset, WX8629, n7005 );
dff WX8439_reg ( clk, reset, WX8439, n6530 );
dff WX8503_reg ( clk, reset, WX8503, n6690 );
dff WX8567_reg ( clk, reset, WX8567, n6850 );
dff WX8631_reg ( clk, reset, WX8631, n7010 );
dff WX8441_reg ( clk, reset, WX8441, n6535 );
dff WX8505_reg ( clk, reset, WX8505, n6695 );
dff WX8569_reg ( clk, reset, WX8569, n6855 );
dff WX8633_reg ( clk, reset, WX8633, n7015 );
dff WX8443_reg ( clk, reset, WX8443, n6540 );
dff WX8507_reg ( clk, reset, WX8507, n6700 );
dff WX8571_reg ( clk, reset, WX8571, n6860 );
dff WX8635_reg ( clk, reset, WX8635, n7020 );
dff WX8445_reg ( clk, reset, WX8445, n6545 );
dff WX8509_reg ( clk, reset, WX8509, n6705 );
dff WX8573_reg ( clk, reset, WX8573, n6865 );
dff WX8637_reg ( clk, reset, WX8637, n7025 );
dff WX8447_reg ( clk, reset, WX8447, n6550 );
dff WX8511_reg ( clk, reset, WX8511, n6710 );
dff WX8575_reg ( clk, reset, WX8575, n6870 );
dff WX8639_reg ( clk, reset, WX8639, n7030 );
dff WX8449_reg ( clk, reset, WX8449, n6555 );
dff WX8513_reg ( clk, reset, WX8513, n6715 );
dff WX8577_reg ( clk, reset, WX8577, n6875 );
dff WX8641_reg ( clk, reset, WX8641, n7035 );
dff WX8451_reg ( clk, reset, WX8451, n6560 );
dff WX8515_reg ( clk, reset, WX8515, n6720 );
dff WX8579_reg ( clk, reset, WX8579, n6880 );
dff WX8643_reg ( clk, reset, WX8643, n7040 );
dff WX8453_reg ( clk, reset, WX8453, n6565 );
dff WX8517_reg ( clk, reset, WX8517, n6725 );
dff WX8581_reg ( clk, reset, WX8581, n6885 );
dff WX8645_reg ( clk, reset, WX8645, n7045 );
dff WX8455_reg ( clk, reset, WX8455, n6570 );
dff WX8519_reg ( clk, reset, WX8519, n6730 );
dff WX8583_reg ( clk, reset, WX8583, n6890 );
dff WX8647_reg ( clk, reset, WX8647, n7050 );
dff WX8457_reg ( clk, reset, WX8457, n6575 );
dff WX8521_reg ( clk, reset, WX8521, n6735 );
dff WX8585_reg ( clk, reset, WX8585, n6895 );
dff WX8649_reg ( clk, reset, WX8649, n7055 );
dff WX8459_reg ( clk, reset, WX8459, n6580 );
dff WX8523_reg ( clk, reset, WX8523, n6740 );
dff WX8587_reg ( clk, reset, WX8587, n6900 );
dff WX8651_reg ( clk, reset, WX8651, n7060 );
dff WX8461_reg ( clk, reset, WX8461, n6585 );
dff WX8525_reg ( clk, reset, WX8525, n6745 );
dff WX8589_reg ( clk, reset, WX8589, n6905 );
dff WX8653_reg ( clk, reset, WX8653, n7065 );
dff WX8463_reg ( clk, reset, WX8463, n6590 );
dff WX8527_reg ( clk, reset, WX8527, n6750 );
dff WX8591_reg ( clk, reset, WX8591, n6910 );
dff WX8655_reg ( clk, reset, WX8655, n7070 );
dff WX8465_reg ( clk, reset, WX8465, n6595 );
dff WX8529_reg ( clk, reset, WX8529, n6755 );
dff WX8593_reg ( clk, reset, WX8593, n6915 );
dff WX8657_reg ( clk, reset, WX8657, n7075 );
dff WX7110_reg ( clk, reset, WX7110, n5512 );
dff WX7174_reg ( clk, reset, WX7174, n5672 );
dff WX7238_reg ( clk, reset, WX7238, n5832 );
dff WX7302_reg ( clk, reset, WX7302, n5992 );
dff CRC_OUT_4_31_reg ( clk, reset, CRC_OUT_4_31, n6276 );
dff CRC_OUT_4_0_reg ( clk, reset, CRC_OUT_4_0, n6152 );
dff CRC_OUT_4_1_reg ( clk, reset, CRC_OUT_4_1, n6156 );
dff CRC_OUT_4_2_reg ( clk, reset, CRC_OUT_4_2, n6160 );
dff CRC_OUT_4_3_reg ( clk, reset, CRC_OUT_4_3, n6164 );
dff CRC_OUT_4_4_reg ( clk, reset, CRC_OUT_4_4, n6168 );
dff CRC_OUT_4_5_reg ( clk, reset, CRC_OUT_4_5, n6172 );
dff CRC_OUT_4_6_reg ( clk, reset, CRC_OUT_4_6, n6176 );
dff CRC_OUT_4_7_reg ( clk, reset, CRC_OUT_4_7, n6180 );
dff CRC_OUT_4_8_reg ( clk, reset, CRC_OUT_4_8, n6184 );
dff CRC_OUT_4_9_reg ( clk, reset, CRC_OUT_4_9, n6188 );
dff CRC_OUT_4_10_reg ( clk, reset, CRC_OUT_4_10, n6192 );
dff CRC_OUT_4_11_reg ( clk, reset, CRC_OUT_4_11, n6196 );
dff CRC_OUT_4_12_reg ( clk, reset, CRC_OUT_4_12, n6200 );
dff CRC_OUT_4_13_reg ( clk, reset, CRC_OUT_4_13, n6204 );
dff CRC_OUT_4_14_reg ( clk, reset, CRC_OUT_4_14, n6208 );
dff CRC_OUT_4_15_reg ( clk, reset, CRC_OUT_4_15, n6212 );
dff CRC_OUT_4_16_reg ( clk, reset, CRC_OUT_4_16, n6216 );
dff CRC_OUT_4_17_reg ( clk, reset, CRC_OUT_4_17, n6220 );
dff CRC_OUT_4_18_reg ( clk, reset, CRC_OUT_4_18, n6224 );
dff CRC_OUT_4_19_reg ( clk, reset, CRC_OUT_4_19, n6228 );
dff CRC_OUT_4_20_reg ( clk, reset, CRC_OUT_4_20, n6232 );
dff CRC_OUT_4_21_reg ( clk, reset, CRC_OUT_4_21, n6236 );
dff CRC_OUT_4_22_reg ( clk, reset, CRC_OUT_4_22, n6240 );
dff CRC_OUT_4_23_reg ( clk, reset, CRC_OUT_4_23, n6244 );
dff CRC_OUT_4_24_reg ( clk, reset, CRC_OUT_4_24, n6248 );
dff CRC_OUT_4_25_reg ( clk, reset, CRC_OUT_4_25, n6252 );
dff CRC_OUT_4_26_reg ( clk, reset, CRC_OUT_4_26, n6256 );
dff CRC_OUT_4_27_reg ( clk, reset, CRC_OUT_4_27, n6260 );
dff CRC_OUT_4_28_reg ( clk, reset, CRC_OUT_4_28, n6264 );
dff CRC_OUT_4_29_reg ( clk, reset, CRC_OUT_4_29, n6268 );
dff CRC_OUT_4_30_reg ( clk, reset, CRC_OUT_4_30, n6272 );
dff WX7112_reg ( clk, reset, WX7112, n5517 );
dff WX7176_reg ( clk, reset, WX7176, n5677 );
dff WX7240_reg ( clk, reset, WX7240, n5837 );
dff WX7304_reg ( clk, reset, WX7304, n5997 );
dff WX7114_reg ( clk, reset, WX7114, n5522 );
dff WX7178_reg ( clk, reset, WX7178, n5682 );
dff WX7242_reg ( clk, reset, WX7242, n5842 );
dff WX7306_reg ( clk, reset, WX7306, n6002 );
dff WX7116_reg ( clk, reset, WX7116, n5527 );
dff WX7180_reg ( clk, reset, WX7180, n5687 );
dff WX7244_reg ( clk, reset, WX7244, n5847 );
dff WX7308_reg ( clk, reset, WX7308, n6007 );
dff WX7118_reg ( clk, reset, WX7118, n5532 );
dff WX7182_reg ( clk, reset, WX7182, n5692 );
dff WX7246_reg ( clk, reset, WX7246, n5852 );
dff WX7310_reg ( clk, reset, WX7310, n6012 );
dff WX7120_reg ( clk, reset, WX7120, n5537 );
dff WX7184_reg ( clk, reset, WX7184, n5697 );
dff WX7248_reg ( clk, reset, WX7248, n5857 );
dff WX7312_reg ( clk, reset, WX7312, n6017 );
dff WX7122_reg ( clk, reset, WX7122, n5542 );
dff WX7186_reg ( clk, reset, WX7186, n5702 );
dff WX7250_reg ( clk, reset, WX7250, n5862 );
dff WX7314_reg ( clk, reset, WX7314, n6022 );
dff WX7124_reg ( clk, reset, WX7124, n5547 );
dff WX7188_reg ( clk, reset, WX7188, n5707 );
dff WX7252_reg ( clk, reset, WX7252, n5867 );
dff WX7316_reg ( clk, reset, WX7316, n6027 );
dff WX7126_reg ( clk, reset, WX7126, n5552 );
dff WX7190_reg ( clk, reset, WX7190, n5712 );
dff WX7254_reg ( clk, reset, WX7254, n5872 );
dff WX7318_reg ( clk, reset, WX7318, n6032 );
dff WX7128_reg ( clk, reset, WX7128, n5557 );
dff WX7192_reg ( clk, reset, WX7192, n5717 );
dff WX7256_reg ( clk, reset, WX7256, n5877 );
dff WX7320_reg ( clk, reset, WX7320, n6037 );
dff WX7130_reg ( clk, reset, WX7130, n5562 );
dff WX7194_reg ( clk, reset, WX7194, n5722 );
dff WX7258_reg ( clk, reset, WX7258, n5882 );
dff WX7322_reg ( clk, reset, WX7322, n6042 );
dff WX7132_reg ( clk, reset, WX7132, n5567 );
dff WX7196_reg ( clk, reset, WX7196, n5727 );
dff WX7260_reg ( clk, reset, WX7260, n5887 );
dff WX7324_reg ( clk, reset, WX7324, n6047 );
dff WX7134_reg ( clk, reset, WX7134, n5572 );
dff WX7198_reg ( clk, reset, WX7198, n5732 );
dff WX7262_reg ( clk, reset, WX7262, n5892 );
dff WX7326_reg ( clk, reset, WX7326, n6052 );
dff WX7136_reg ( clk, reset, WX7136, n5577 );
dff WX7200_reg ( clk, reset, WX7200, n5737 );
dff WX7264_reg ( clk, reset, WX7264, n5897 );
dff WX7328_reg ( clk, reset, WX7328, n6057 );
dff WX7138_reg ( clk, reset, WX7138, n5582 );
dff WX7202_reg ( clk, reset, WX7202, n5742 );
dff WX7266_reg ( clk, reset, WX7266, n5902 );
dff WX7330_reg ( clk, reset, WX7330, n6062 );
dff WX7140_reg ( clk, reset, WX7140, n5587 );
dff WX7204_reg ( clk, reset, WX7204, n5747 );
dff WX7268_reg ( clk, reset, WX7268, n5907 );
dff WX7332_reg ( clk, reset, WX7332, n6067 );
dff WX7142_reg ( clk, reset, WX7142, n5592 );
dff WX7206_reg ( clk, reset, WX7206, n5752 );
dff WX7270_reg ( clk, reset, WX7270, n5912 );
dff WX7334_reg ( clk, reset, WX7334, n6072 );
dff WX7144_reg ( clk, reset, WX7144, n5597 );
dff WX7208_reg ( clk, reset, WX7208, n5757 );
dff WX7272_reg ( clk, reset, WX7272, n5917 );
dff WX7336_reg ( clk, reset, WX7336, n6077 );
dff WX7146_reg ( clk, reset, WX7146, n5602 );
dff WX7210_reg ( clk, reset, WX7210, n5762 );
dff WX7274_reg ( clk, reset, WX7274, n5922 );
dff WX7338_reg ( clk, reset, WX7338, n6082 );
dff WX7148_reg ( clk, reset, WX7148, n5607 );
dff WX7212_reg ( clk, reset, WX7212, n5767 );
dff WX7276_reg ( clk, reset, WX7276, n5927 );
dff WX7340_reg ( clk, reset, WX7340, n6087 );
dff WX7150_reg ( clk, reset, WX7150, n5612 );
dff WX7214_reg ( clk, reset, WX7214, n5772 );
dff WX7278_reg ( clk, reset, WX7278, n5932 );
dff WX7342_reg ( clk, reset, WX7342, n6092 );
dff WX7152_reg ( clk, reset, WX7152, n5617 );
dff WX7216_reg ( clk, reset, WX7216, n5777 );
dff WX7280_reg ( clk, reset, WX7280, n5937 );
dff WX7344_reg ( clk, reset, WX7344, n6097 );
dff WX7154_reg ( clk, reset, WX7154, n5622 );
dff WX7218_reg ( clk, reset, WX7218, n5782 );
dff WX7282_reg ( clk, reset, WX7282, n5942 );
dff WX7346_reg ( clk, reset, WX7346, n6102 );
dff WX7156_reg ( clk, reset, WX7156, n5627 );
dff WX7220_reg ( clk, reset, WX7220, n5787 );
dff WX7284_reg ( clk, reset, WX7284, n5947 );
dff WX7348_reg ( clk, reset, WX7348, n6107 );
dff WX7158_reg ( clk, reset, WX7158, n5632 );
dff WX7222_reg ( clk, reset, WX7222, n5792 );
dff WX7286_reg ( clk, reset, WX7286, n5952 );
dff WX7350_reg ( clk, reset, WX7350, n6112 );
dff WX7160_reg ( clk, reset, WX7160, n5637 );
dff WX7224_reg ( clk, reset, WX7224, n5797 );
dff WX7288_reg ( clk, reset, WX7288, n5957 );
dff WX7352_reg ( clk, reset, WX7352, n6117 );
dff WX7162_reg ( clk, reset, WX7162, n5642 );
dff WX7226_reg ( clk, reset, WX7226, n5802 );
dff WX7290_reg ( clk, reset, WX7290, n5962 );
dff WX7354_reg ( clk, reset, WX7354, n6122 );
dff WX7164_reg ( clk, reset, WX7164, n5647 );
dff WX7228_reg ( clk, reset, WX7228, n5807 );
dff WX7292_reg ( clk, reset, WX7292, n5967 );
dff WX7356_reg ( clk, reset, WX7356, n6127 );
dff WX7166_reg ( clk, reset, WX7166, n5652 );
dff WX7230_reg ( clk, reset, WX7230, n5812 );
dff WX7294_reg ( clk, reset, WX7294, n5972 );
dff WX7358_reg ( clk, reset, WX7358, n6132 );
dff WX7168_reg ( clk, reset, WX7168, n5657 );
dff WX7232_reg ( clk, reset, WX7232, n5817 );
dff WX7296_reg ( clk, reset, WX7296, n5977 );
dff WX7360_reg ( clk, reset, WX7360, n6137 );
dff WX7170_reg ( clk, reset, WX7170, n5662 );
dff WX7234_reg ( clk, reset, WX7234, n5822 );
dff WX7298_reg ( clk, reset, WX7298, n5982 );
dff WX7362_reg ( clk, reset, WX7362, n6142 );
dff WX7172_reg ( clk, reset, WX7172, n5667 );
dff WX7236_reg ( clk, reset, WX7236, n5827 );
dff WX7300_reg ( clk, reset, WX7300, n5987 );
dff WX7364_reg ( clk, reset, WX7364, n6147 );
dff WX5817_reg ( clk, reset, WX5817, n4584 );
dff WX5881_reg ( clk, reset, WX5881, n4744 );
dff WX5945_reg ( clk, reset, WX5945, n4904 );
dff WX6009_reg ( clk, reset, WX6009, n5064 );
dff CRC_OUT_5_31_reg ( clk, reset, CRC_OUT_5_31, n5348 );
dff CRC_OUT_5_0_reg ( clk, reset, CRC_OUT_5_0, n5224 );
dff CRC_OUT_5_1_reg ( clk, reset, CRC_OUT_5_1, n5228 );
dff CRC_OUT_5_2_reg ( clk, reset, CRC_OUT_5_2, n5232 );
dff CRC_OUT_5_3_reg ( clk, reset, CRC_OUT_5_3, n5236 );
dff CRC_OUT_5_4_reg ( clk, reset, CRC_OUT_5_4, n5240 );
dff CRC_OUT_5_5_reg ( clk, reset, CRC_OUT_5_5, n5244 );
dff CRC_OUT_5_6_reg ( clk, reset, CRC_OUT_5_6, n5248 );
dff CRC_OUT_5_7_reg ( clk, reset, CRC_OUT_5_7, n5252 );
dff CRC_OUT_5_8_reg ( clk, reset, CRC_OUT_5_8, n5256 );
dff CRC_OUT_5_9_reg ( clk, reset, CRC_OUT_5_9, n5260 );
dff CRC_OUT_5_10_reg ( clk, reset, CRC_OUT_5_10, n5264 );
dff CRC_OUT_5_11_reg ( clk, reset, CRC_OUT_5_11, n5268 );
dff CRC_OUT_5_12_reg ( clk, reset, CRC_OUT_5_12, n5272 );
dff CRC_OUT_5_13_reg ( clk, reset, CRC_OUT_5_13, n5276 );
dff CRC_OUT_5_14_reg ( clk, reset, CRC_OUT_5_14, n5280 );
dff CRC_OUT_5_15_reg ( clk, reset, CRC_OUT_5_15, n5284 );
dff CRC_OUT_5_16_reg ( clk, reset, CRC_OUT_5_16, n5288 );
dff CRC_OUT_5_17_reg ( clk, reset, CRC_OUT_5_17, n5292 );
dff CRC_OUT_5_18_reg ( clk, reset, CRC_OUT_5_18, n5296 );
dff CRC_OUT_5_19_reg ( clk, reset, CRC_OUT_5_19, n5300 );
dff CRC_OUT_5_20_reg ( clk, reset, CRC_OUT_5_20, n5304 );
dff CRC_OUT_5_21_reg ( clk, reset, CRC_OUT_5_21, n5308 );
dff CRC_OUT_5_22_reg ( clk, reset, CRC_OUT_5_22, n5312 );
dff CRC_OUT_5_23_reg ( clk, reset, CRC_OUT_5_23, n5316 );
dff CRC_OUT_5_24_reg ( clk, reset, CRC_OUT_5_24, n5320 );
dff CRC_OUT_5_25_reg ( clk, reset, CRC_OUT_5_25, n5324 );
dff CRC_OUT_5_26_reg ( clk, reset, CRC_OUT_5_26, n5328 );
dff CRC_OUT_5_27_reg ( clk, reset, CRC_OUT_5_27, n5332 );
dff CRC_OUT_5_28_reg ( clk, reset, CRC_OUT_5_28, n5336 );
dff CRC_OUT_5_29_reg ( clk, reset, CRC_OUT_5_29, n5340 );
dff CRC_OUT_5_30_reg ( clk, reset, CRC_OUT_5_30, n5344 );
dff WX5819_reg ( clk, reset, WX5819, n4589 );
dff WX5883_reg ( clk, reset, WX5883, n4749 );
dff WX5947_reg ( clk, reset, WX5947, n4909 );
dff WX6011_reg ( clk, reset, WX6011, n5069 );
dff WX5821_reg ( clk, reset, WX5821, n4594 );
dff WX5885_reg ( clk, reset, WX5885, n4754 );
dff WX5949_reg ( clk, reset, WX5949, n4914 );
dff WX6013_reg ( clk, reset, WX6013, n5074 );
dff WX5823_reg ( clk, reset, WX5823, n4599 );
dff WX5887_reg ( clk, reset, WX5887, n4759 );
dff WX5951_reg ( clk, reset, WX5951, n4919 );
dff WX6015_reg ( clk, reset, WX6015, n5079 );
dff WX5825_reg ( clk, reset, WX5825, n4604 );
dff WX5889_reg ( clk, reset, WX5889, n4764 );
dff WX5953_reg ( clk, reset, WX5953, n4924 );
dff WX6017_reg ( clk, reset, WX6017, n5084 );
dff WX5827_reg ( clk, reset, WX5827, n4609 );
dff WX5891_reg ( clk, reset, WX5891, n4769 );
dff WX5955_reg ( clk, reset, WX5955, n4929 );
dff WX6019_reg ( clk, reset, WX6019, n5089 );
dff WX5829_reg ( clk, reset, WX5829, n4614 );
dff WX5893_reg ( clk, reset, WX5893, n4774 );
dff WX5957_reg ( clk, reset, WX5957, n4934 );
dff WX6021_reg ( clk, reset, WX6021, n5094 );
dff WX5831_reg ( clk, reset, WX5831, n4619 );
dff WX5895_reg ( clk, reset, WX5895, n4779 );
dff WX5959_reg ( clk, reset, WX5959, n4939 );
dff WX6023_reg ( clk, reset, WX6023, n5099 );
dff WX5833_reg ( clk, reset, WX5833, n4624 );
dff WX5897_reg ( clk, reset, WX5897, n4784 );
dff WX5961_reg ( clk, reset, WX5961, n4944 );
dff WX6025_reg ( clk, reset, WX6025, n5104 );
dff WX5835_reg ( clk, reset, WX5835, n4629 );
dff WX5899_reg ( clk, reset, WX5899, n4789 );
dff WX5963_reg ( clk, reset, WX5963, n4949 );
dff WX6027_reg ( clk, reset, WX6027, n5109 );
dff WX5837_reg ( clk, reset, WX5837, n4634 );
dff WX5901_reg ( clk, reset, WX5901, n4794 );
dff WX5965_reg ( clk, reset, WX5965, n4954 );
dff WX6029_reg ( clk, reset, WX6029, n5114 );
dff WX5839_reg ( clk, reset, WX5839, n4639 );
dff WX5903_reg ( clk, reset, WX5903, n4799 );
dff WX5967_reg ( clk, reset, WX5967, n4959 );
dff WX6031_reg ( clk, reset, WX6031, n5119 );
dff WX5841_reg ( clk, reset, WX5841, n4644 );
dff WX5905_reg ( clk, reset, WX5905, n4804 );
dff WX5969_reg ( clk, reset, WX5969, n4964 );
dff WX6033_reg ( clk, reset, WX6033, n5124 );
dff WX5843_reg ( clk, reset, WX5843, n4649 );
dff WX5907_reg ( clk, reset, WX5907, n4809 );
dff WX5971_reg ( clk, reset, WX5971, n4969 );
dff WX6035_reg ( clk, reset, WX6035, n5129 );
dff WX5845_reg ( clk, reset, WX5845, n4654 );
dff WX5909_reg ( clk, reset, WX5909, n4814 );
dff WX5973_reg ( clk, reset, WX5973, n4974 );
dff WX6037_reg ( clk, reset, WX6037, n5134 );
dff WX5847_reg ( clk, reset, WX5847, n4659 );
dff WX5911_reg ( clk, reset, WX5911, n4819 );
dff WX5975_reg ( clk, reset, WX5975, n4979 );
dff WX6039_reg ( clk, reset, WX6039, n5139 );
dff WX5849_reg ( clk, reset, WX5849, n4664 );
dff WX5913_reg ( clk, reset, WX5913, n4824 );
dff WX5977_reg ( clk, reset, WX5977, n4984 );
dff WX6041_reg ( clk, reset, WX6041, n5144 );
dff WX5851_reg ( clk, reset, WX5851, n4669 );
dff WX5915_reg ( clk, reset, WX5915, n4829 );
dff WX5979_reg ( clk, reset, WX5979, n4989 );
dff WX6043_reg ( clk, reset, WX6043, n5149 );
dff WX5853_reg ( clk, reset, WX5853, n4674 );
dff WX5917_reg ( clk, reset, WX5917, n4834 );
dff WX5981_reg ( clk, reset, WX5981, n4994 );
dff WX6045_reg ( clk, reset, WX6045, n5154 );
dff WX5855_reg ( clk, reset, WX5855, n4679 );
dff WX5919_reg ( clk, reset, WX5919, n4839 );
dff WX5983_reg ( clk, reset, WX5983, n4999 );
dff WX6047_reg ( clk, reset, WX6047, n5159 );
dff WX5857_reg ( clk, reset, WX5857, n4684 );
dff WX5921_reg ( clk, reset, WX5921, n4844 );
dff WX5985_reg ( clk, reset, WX5985, n5004 );
dff WX6049_reg ( clk, reset, WX6049, n5164 );
dff WX5859_reg ( clk, reset, WX5859, n4689 );
dff WX5923_reg ( clk, reset, WX5923, n4849 );
dff WX5987_reg ( clk, reset, WX5987, n5009 );
dff WX6051_reg ( clk, reset, WX6051, n5169 );
dff WX5861_reg ( clk, reset, WX5861, n4694 );
dff WX5925_reg ( clk, reset, WX5925, n4854 );
dff WX5989_reg ( clk, reset, WX5989, n5014 );
dff WX6053_reg ( clk, reset, WX6053, n5174 );
dff WX5863_reg ( clk, reset, WX5863, n4699 );
dff WX5927_reg ( clk, reset, WX5927, n4859 );
dff WX5991_reg ( clk, reset, WX5991, n5019 );
dff WX6055_reg ( clk, reset, WX6055, n5179 );
dff WX5865_reg ( clk, reset, WX5865, n4704 );
dff WX5929_reg ( clk, reset, WX5929, n4864 );
dff WX5993_reg ( clk, reset, WX5993, n5024 );
dff WX6057_reg ( clk, reset, WX6057, n5184 );
dff WX5867_reg ( clk, reset, WX5867, n4709 );
dff WX5931_reg ( clk, reset, WX5931, n4869 );
dff WX5995_reg ( clk, reset, WX5995, n5029 );
dff WX6059_reg ( clk, reset, WX6059, n5189 );
dff WX5869_reg ( clk, reset, WX5869, n4714 );
dff WX5933_reg ( clk, reset, WX5933, n4874 );
dff WX5997_reg ( clk, reset, WX5997, n5034 );
dff WX6061_reg ( clk, reset, WX6061, n5194 );
dff WX5871_reg ( clk, reset, WX5871, n4719 );
dff WX5935_reg ( clk, reset, WX5935, n4879 );
dff WX5999_reg ( clk, reset, WX5999, n5039 );
dff WX6063_reg ( clk, reset, WX6063, n5199 );
dff WX5873_reg ( clk, reset, WX5873, n4724 );
dff WX5937_reg ( clk, reset, WX5937, n4884 );
dff WX6001_reg ( clk, reset, WX6001, n5044 );
dff WX6065_reg ( clk, reset, WX6065, n5204 );
dff WX5875_reg ( clk, reset, WX5875, n4729 );
dff WX5939_reg ( clk, reset, WX5939, n4889 );
dff WX6003_reg ( clk, reset, WX6003, n5049 );
dff WX6067_reg ( clk, reset, WX6067, n5209 );
dff WX5877_reg ( clk, reset, WX5877, n4734 );
dff WX5941_reg ( clk, reset, WX5941, n4894 );
dff WX6005_reg ( clk, reset, WX6005, n5054 );
dff WX6069_reg ( clk, reset, WX6069, n5214 );
dff WX5879_reg ( clk, reset, WX5879, n4739 );
dff WX5943_reg ( clk, reset, WX5943, n4899 );
dff WX6007_reg ( clk, reset, WX6007, n5059 );
dff WX6071_reg ( clk, reset, WX6071, n5219 );
dff WX4524_reg ( clk, reset, WX4524, n3656 );
dff WX4588_reg ( clk, reset, WX4588, n3816 );
dff WX4652_reg ( clk, reset, WX4652, n3976 );
dff WX4716_reg ( clk, reset, WX4716, n4136 );
dff CRC_OUT_6_31_reg ( clk, reset, CRC_OUT_6_31, n4420 );
dff CRC_OUT_6_0_reg ( clk, reset, CRC_OUT_6_0, n4296 );
dff CRC_OUT_6_1_reg ( clk, reset, CRC_OUT_6_1, n4300 );
dff CRC_OUT_6_2_reg ( clk, reset, CRC_OUT_6_2, n4304 );
dff CRC_OUT_6_3_reg ( clk, reset, CRC_OUT_6_3, n4308 );
dff CRC_OUT_6_4_reg ( clk, reset, CRC_OUT_6_4, n4312 );
dff CRC_OUT_6_5_reg ( clk, reset, CRC_OUT_6_5, n4316 );
dff CRC_OUT_6_6_reg ( clk, reset, CRC_OUT_6_6, n4320 );
dff CRC_OUT_6_7_reg ( clk, reset, CRC_OUT_6_7, n4324 );
dff CRC_OUT_6_8_reg ( clk, reset, CRC_OUT_6_8, n4328 );
dff CRC_OUT_6_9_reg ( clk, reset, CRC_OUT_6_9, n4332 );
dff CRC_OUT_6_10_reg ( clk, reset, CRC_OUT_6_10, n4336 );
dff CRC_OUT_6_11_reg ( clk, reset, CRC_OUT_6_11, n4340 );
dff CRC_OUT_6_12_reg ( clk, reset, CRC_OUT_6_12, n4344 );
dff CRC_OUT_6_13_reg ( clk, reset, CRC_OUT_6_13, n4348 );
dff CRC_OUT_6_14_reg ( clk, reset, CRC_OUT_6_14, n4352 );
dff CRC_OUT_6_15_reg ( clk, reset, CRC_OUT_6_15, n4356 );
dff CRC_OUT_6_16_reg ( clk, reset, CRC_OUT_6_16, n4360 );
dff CRC_OUT_6_17_reg ( clk, reset, CRC_OUT_6_17, n4364 );
dff CRC_OUT_6_18_reg ( clk, reset, CRC_OUT_6_18, n4368 );
dff CRC_OUT_6_19_reg ( clk, reset, CRC_OUT_6_19, n4372 );
dff CRC_OUT_6_20_reg ( clk, reset, CRC_OUT_6_20, n4376 );
dff CRC_OUT_6_21_reg ( clk, reset, CRC_OUT_6_21, n4380 );
dff CRC_OUT_6_22_reg ( clk, reset, CRC_OUT_6_22, n4384 );
dff CRC_OUT_6_23_reg ( clk, reset, CRC_OUT_6_23, n4388 );
dff CRC_OUT_6_24_reg ( clk, reset, CRC_OUT_6_24, n4392 );
dff CRC_OUT_6_25_reg ( clk, reset, CRC_OUT_6_25, n4396 );
dff CRC_OUT_6_26_reg ( clk, reset, CRC_OUT_6_26, n4400 );
dff CRC_OUT_6_27_reg ( clk, reset, CRC_OUT_6_27, n4404 );
dff CRC_OUT_6_28_reg ( clk, reset, CRC_OUT_6_28, n4408 );
dff CRC_OUT_6_29_reg ( clk, reset, CRC_OUT_6_29, n4412 );
dff CRC_OUT_6_30_reg ( clk, reset, CRC_OUT_6_30, n4416 );
dff WX4526_reg ( clk, reset, WX4526, n3661 );
dff WX4590_reg ( clk, reset, WX4590, n3821 );
dff WX4654_reg ( clk, reset, WX4654, n3981 );
dff WX4718_reg ( clk, reset, WX4718, n4141 );
dff WX4528_reg ( clk, reset, WX4528, n3666 );
dff WX4592_reg ( clk, reset, WX4592, n3826 );
dff WX4656_reg ( clk, reset, WX4656, n3986 );
dff WX4720_reg ( clk, reset, WX4720, n4146 );
dff WX4530_reg ( clk, reset, WX4530, n3671 );
dff WX4594_reg ( clk, reset, WX4594, n3831 );
dff WX4658_reg ( clk, reset, WX4658, n3991 );
dff WX4722_reg ( clk, reset, WX4722, n4151 );
dff WX4532_reg ( clk, reset, WX4532, n3676 );
dff WX4596_reg ( clk, reset, WX4596, n3836 );
dff WX4660_reg ( clk, reset, WX4660, n3996 );
dff WX4724_reg ( clk, reset, WX4724, n4156 );
dff WX4534_reg ( clk, reset, WX4534, n3681 );
dff WX4598_reg ( clk, reset, WX4598, n3841 );
dff WX4662_reg ( clk, reset, WX4662, n4001 );
dff WX4726_reg ( clk, reset, WX4726, n4161 );
dff WX4536_reg ( clk, reset, WX4536, n3686 );
dff WX4600_reg ( clk, reset, WX4600, n3846 );
dff WX4664_reg ( clk, reset, WX4664, n4006 );
dff WX4728_reg ( clk, reset, WX4728, n4166 );
dff WX4538_reg ( clk, reset, WX4538, n3691 );
dff WX4602_reg ( clk, reset, WX4602, n3851 );
dff WX4666_reg ( clk, reset, WX4666, n4011 );
dff WX4730_reg ( clk, reset, WX4730, n4171 );
dff WX4540_reg ( clk, reset, WX4540, n3696 );
dff WX4604_reg ( clk, reset, WX4604, n3856 );
dff WX4668_reg ( clk, reset, WX4668, n4016 );
dff WX4732_reg ( clk, reset, WX4732, n4176 );
dff WX4542_reg ( clk, reset, WX4542, n3701 );
dff WX4606_reg ( clk, reset, WX4606, n3861 );
dff WX4670_reg ( clk, reset, WX4670, n4021 );
dff WX4734_reg ( clk, reset, WX4734, n4181 );
dff WX4544_reg ( clk, reset, WX4544, n3706 );
dff WX4608_reg ( clk, reset, WX4608, n3866 );
dff WX4672_reg ( clk, reset, WX4672, n4026 );
dff WX4736_reg ( clk, reset, WX4736, n4186 );
dff WX4546_reg ( clk, reset, WX4546, n3711 );
dff WX4610_reg ( clk, reset, WX4610, n3871 );
dff WX4674_reg ( clk, reset, WX4674, n4031 );
dff WX4738_reg ( clk, reset, WX4738, n4191 );
dff WX4548_reg ( clk, reset, WX4548, n3716 );
dff WX4612_reg ( clk, reset, WX4612, n3876 );
dff WX4676_reg ( clk, reset, WX4676, n4036 );
dff WX4740_reg ( clk, reset, WX4740, n4196 );
dff WX4550_reg ( clk, reset, WX4550, n3721 );
dff WX4614_reg ( clk, reset, WX4614, n3881 );
dff WX4678_reg ( clk, reset, WX4678, n4041 );
dff WX4742_reg ( clk, reset, WX4742, n4201 );
dff WX4552_reg ( clk, reset, WX4552, n3726 );
dff WX4616_reg ( clk, reset, WX4616, n3886 );
dff WX4680_reg ( clk, reset, WX4680, n4046 );
dff WX4744_reg ( clk, reset, WX4744, n4206 );
dff WX4554_reg ( clk, reset, WX4554, n3731 );
dff WX4618_reg ( clk, reset, WX4618, n3891 );
dff WX4682_reg ( clk, reset, WX4682, n4051 );
dff WX4746_reg ( clk, reset, WX4746, n4211 );
dff WX4556_reg ( clk, reset, WX4556, n3736 );
dff WX4620_reg ( clk, reset, WX4620, n3896 );
dff WX4684_reg ( clk, reset, WX4684, n4056 );
dff WX4748_reg ( clk, reset, WX4748, n4216 );
dff WX4558_reg ( clk, reset, WX4558, n3741 );
dff WX4622_reg ( clk, reset, WX4622, n3901 );
dff WX4686_reg ( clk, reset, WX4686, n4061 );
dff WX4750_reg ( clk, reset, WX4750, n4221 );
dff WX4560_reg ( clk, reset, WX4560, n3746 );
dff WX4624_reg ( clk, reset, WX4624, n3906 );
dff WX4688_reg ( clk, reset, WX4688, n4066 );
dff WX4752_reg ( clk, reset, WX4752, n4226 );
dff WX4562_reg ( clk, reset, WX4562, n3751 );
dff WX4626_reg ( clk, reset, WX4626, n3911 );
dff WX4690_reg ( clk, reset, WX4690, n4071 );
dff WX4754_reg ( clk, reset, WX4754, n4231 );
dff WX4564_reg ( clk, reset, WX4564, n3756 );
dff WX4628_reg ( clk, reset, WX4628, n3916 );
dff WX4692_reg ( clk, reset, WX4692, n4076 );
dff WX4756_reg ( clk, reset, WX4756, n4236 );
dff WX4566_reg ( clk, reset, WX4566, n3761 );
dff WX4630_reg ( clk, reset, WX4630, n3921 );
dff WX4694_reg ( clk, reset, WX4694, n4081 );
dff WX4758_reg ( clk, reset, WX4758, n4241 );
dff WX4568_reg ( clk, reset, WX4568, n3766 );
dff WX4632_reg ( clk, reset, WX4632, n3926 );
dff WX4696_reg ( clk, reset, WX4696, n4086 );
dff WX4760_reg ( clk, reset, WX4760, n4246 );
dff WX4570_reg ( clk, reset, WX4570, n3771 );
dff WX4634_reg ( clk, reset, WX4634, n3931 );
dff WX4698_reg ( clk, reset, WX4698, n4091 );
dff WX4762_reg ( clk, reset, WX4762, n4251 );
dff WX4572_reg ( clk, reset, WX4572, n3776 );
dff WX4636_reg ( clk, reset, WX4636, n3936 );
dff WX4700_reg ( clk, reset, WX4700, n4096 );
dff WX4764_reg ( clk, reset, WX4764, n4256 );
dff WX4574_reg ( clk, reset, WX4574, n3781 );
dff WX4638_reg ( clk, reset, WX4638, n3941 );
dff WX4702_reg ( clk, reset, WX4702, n4101 );
dff WX4766_reg ( clk, reset, WX4766, n4261 );
dff WX4576_reg ( clk, reset, WX4576, n3786 );
dff WX4640_reg ( clk, reset, WX4640, n3946 );
dff WX4704_reg ( clk, reset, WX4704, n4106 );
dff WX4768_reg ( clk, reset, WX4768, n4266 );
dff WX4578_reg ( clk, reset, WX4578, n3791 );
dff WX4642_reg ( clk, reset, WX4642, n3951 );
dff WX4706_reg ( clk, reset, WX4706, n4111 );
dff WX4770_reg ( clk, reset, WX4770, n4271 );
dff WX4580_reg ( clk, reset, WX4580, n3796 );
dff WX4644_reg ( clk, reset, WX4644, n3956 );
dff WX4708_reg ( clk, reset, WX4708, n4116 );
dff WX4772_reg ( clk, reset, WX4772, n4276 );
dff WX4582_reg ( clk, reset, WX4582, n3801 );
dff WX4646_reg ( clk, reset, WX4646, n3961 );
dff WX4710_reg ( clk, reset, WX4710, n4121 );
dff WX4774_reg ( clk, reset, WX4774, n4281 );
dff WX4584_reg ( clk, reset, WX4584, n3806 );
dff WX4648_reg ( clk, reset, WX4648, n3966 );
dff WX4712_reg ( clk, reset, WX4712, n4126 );
dff WX4776_reg ( clk, reset, WX4776, n4286 );
dff WX4586_reg ( clk, reset, WX4586, n3811 );
dff WX4650_reg ( clk, reset, WX4650, n3971 );
dff WX4714_reg ( clk, reset, WX4714, n4131 );
dff WX4778_reg ( clk, reset, WX4778, n4291 );
dff WX3231_reg ( clk, reset, WX3231, n2728 );
dff WX3295_reg ( clk, reset, WX3295, n2888 );
dff WX3359_reg ( clk, reset, WX3359, n3048 );
dff WX3423_reg ( clk, reset, WX3423, n3208 );
dff CRC_OUT_7_31_reg ( clk, reset, CRC_OUT_7_31, n3492 );
dff CRC_OUT_7_0_reg ( clk, reset, CRC_OUT_7_0, n3368 );
dff CRC_OUT_7_1_reg ( clk, reset, CRC_OUT_7_1, n3372 );
dff CRC_OUT_7_2_reg ( clk, reset, CRC_OUT_7_2, n3376 );
dff CRC_OUT_7_3_reg ( clk, reset, CRC_OUT_7_3, n3380 );
dff CRC_OUT_7_4_reg ( clk, reset, CRC_OUT_7_4, n3384 );
dff CRC_OUT_7_5_reg ( clk, reset, CRC_OUT_7_5, n3388 );
dff CRC_OUT_7_6_reg ( clk, reset, CRC_OUT_7_6, n3392 );
dff CRC_OUT_7_7_reg ( clk, reset, CRC_OUT_7_7, n3396 );
dff CRC_OUT_7_8_reg ( clk, reset, CRC_OUT_7_8, n3400 );
dff CRC_OUT_7_9_reg ( clk, reset, CRC_OUT_7_9, n3404 );
dff CRC_OUT_7_10_reg ( clk, reset, CRC_OUT_7_10, n3408 );
dff CRC_OUT_7_11_reg ( clk, reset, CRC_OUT_7_11, n3412 );
dff CRC_OUT_7_12_reg ( clk, reset, CRC_OUT_7_12, n3416 );
dff CRC_OUT_7_13_reg ( clk, reset, CRC_OUT_7_13, n3420 );
dff CRC_OUT_7_14_reg ( clk, reset, CRC_OUT_7_14, n3424 );
dff CRC_OUT_7_15_reg ( clk, reset, CRC_OUT_7_15, n3428 );
dff CRC_OUT_7_16_reg ( clk, reset, CRC_OUT_7_16, n3432 );
dff CRC_OUT_7_17_reg ( clk, reset, CRC_OUT_7_17, n3436 );
dff CRC_OUT_7_18_reg ( clk, reset, CRC_OUT_7_18, n3440 );
dff CRC_OUT_7_19_reg ( clk, reset, CRC_OUT_7_19, n3444 );
dff CRC_OUT_7_20_reg ( clk, reset, CRC_OUT_7_20, n3448 );
dff CRC_OUT_7_21_reg ( clk, reset, CRC_OUT_7_21, n3452 );
dff CRC_OUT_7_22_reg ( clk, reset, CRC_OUT_7_22, n3456 );
dff CRC_OUT_7_23_reg ( clk, reset, CRC_OUT_7_23, n3460 );
dff CRC_OUT_7_24_reg ( clk, reset, CRC_OUT_7_24, n3464 );
dff CRC_OUT_7_25_reg ( clk, reset, CRC_OUT_7_25, n3468 );
dff CRC_OUT_7_26_reg ( clk, reset, CRC_OUT_7_26, n3472 );
dff CRC_OUT_7_27_reg ( clk, reset, CRC_OUT_7_27, n3476 );
dff CRC_OUT_7_28_reg ( clk, reset, CRC_OUT_7_28, n3480 );
dff CRC_OUT_7_29_reg ( clk, reset, CRC_OUT_7_29, n3484 );
dff CRC_OUT_7_30_reg ( clk, reset, CRC_OUT_7_30, n3488 );
dff WX3233_reg ( clk, reset, WX3233, n2733 );
dff WX3297_reg ( clk, reset, WX3297, n2893 );
dff WX3361_reg ( clk, reset, WX3361, n3053 );
dff WX3425_reg ( clk, reset, WX3425, n3213 );
dff WX3235_reg ( clk, reset, WX3235, n2738 );
dff WX3299_reg ( clk, reset, WX3299, n2898 );
dff WX3363_reg ( clk, reset, WX3363, n3058 );
dff WX3427_reg ( clk, reset, WX3427, n3218 );
dff WX3237_reg ( clk, reset, WX3237, n2743 );
dff WX3301_reg ( clk, reset, WX3301, n2903 );
dff WX3365_reg ( clk, reset, WX3365, n3063 );
dff WX3429_reg ( clk, reset, WX3429, n3223 );
dff WX3239_reg ( clk, reset, WX3239, n2748 );
dff WX3303_reg ( clk, reset, WX3303, n2908 );
dff WX3367_reg ( clk, reset, WX3367, n3068 );
dff WX3431_reg ( clk, reset, WX3431, n3228 );
dff WX3241_reg ( clk, reset, WX3241, n2753 );
dff WX3305_reg ( clk, reset, WX3305, n2913 );
dff WX3369_reg ( clk, reset, WX3369, n3073 );
dff WX3433_reg ( clk, reset, WX3433, n3233 );
dff WX3243_reg ( clk, reset, WX3243, n2758 );
dff WX3307_reg ( clk, reset, WX3307, n2918 );
dff WX3371_reg ( clk, reset, WX3371, n3078 );
dff WX3435_reg ( clk, reset, WX3435, n3238 );
dff WX3245_reg ( clk, reset, WX3245, n2763 );
dff WX3309_reg ( clk, reset, WX3309, n2923 );
dff WX3373_reg ( clk, reset, WX3373, n3083 );
dff WX3437_reg ( clk, reset, WX3437, n3243 );
dff WX3247_reg ( clk, reset, WX3247, n2768 );
dff WX3311_reg ( clk, reset, WX3311, n2928 );
dff WX3375_reg ( clk, reset, WX3375, n3088 );
dff WX3439_reg ( clk, reset, WX3439, n3248 );
dff WX3249_reg ( clk, reset, WX3249, n2773 );
dff WX3313_reg ( clk, reset, WX3313, n2933 );
dff WX3377_reg ( clk, reset, WX3377, n3093 );
dff WX3441_reg ( clk, reset, WX3441, n3253 );
dff WX3251_reg ( clk, reset, WX3251, n2778 );
dff WX3315_reg ( clk, reset, WX3315, n2938 );
dff WX3379_reg ( clk, reset, WX3379, n3098 );
dff WX3443_reg ( clk, reset, WX3443, n3258 );
dff WX3253_reg ( clk, reset, WX3253, n2783 );
dff WX3317_reg ( clk, reset, WX3317, n2943 );
dff WX3381_reg ( clk, reset, WX3381, n3103 );
dff WX3445_reg ( clk, reset, WX3445, n3263 );
dff WX3255_reg ( clk, reset, WX3255, n2788 );
dff WX3319_reg ( clk, reset, WX3319, n2948 );
dff WX3383_reg ( clk, reset, WX3383, n3108 );
dff WX3447_reg ( clk, reset, WX3447, n3268 );
dff WX3257_reg ( clk, reset, WX3257, n2793 );
dff WX3321_reg ( clk, reset, WX3321, n2953 );
dff WX3385_reg ( clk, reset, WX3385, n3113 );
dff WX3449_reg ( clk, reset, WX3449, n3273 );
dff WX3259_reg ( clk, reset, WX3259, n2798 );
dff WX3323_reg ( clk, reset, WX3323, n2958 );
dff WX3387_reg ( clk, reset, WX3387, n3118 );
dff WX3451_reg ( clk, reset, WX3451, n3278 );
dff WX3261_reg ( clk, reset, WX3261, n2803 );
dff WX3325_reg ( clk, reset, WX3325, n2963 );
dff WX3389_reg ( clk, reset, WX3389, n3123 );
dff WX3453_reg ( clk, reset, WX3453, n3283 );
dff WX3263_reg ( clk, reset, WX3263, n2808 );
dff WX3327_reg ( clk, reset, WX3327, n2968 );
dff WX3391_reg ( clk, reset, WX3391, n3128 );
dff WX3455_reg ( clk, reset, WX3455, n3288 );
dff WX3265_reg ( clk, reset, WX3265, n2813 );
dff WX3329_reg ( clk, reset, WX3329, n2973 );
dff WX3393_reg ( clk, reset, WX3393, n3133 );
dff WX3457_reg ( clk, reset, WX3457, n3293 );
dff WX3267_reg ( clk, reset, WX3267, n2818 );
dff WX3331_reg ( clk, reset, WX3331, n2978 );
dff WX3395_reg ( clk, reset, WX3395, n3138 );
dff WX3459_reg ( clk, reset, WX3459, n3298 );
dff WX3269_reg ( clk, reset, WX3269, n2823 );
dff WX3333_reg ( clk, reset, WX3333, n2983 );
dff WX3397_reg ( clk, reset, WX3397, n3143 );
dff WX3461_reg ( clk, reset, WX3461, n3303 );
dff WX3271_reg ( clk, reset, WX3271, n2828 );
dff WX3335_reg ( clk, reset, WX3335, n2988 );
dff WX3399_reg ( clk, reset, WX3399, n3148 );
dff WX3463_reg ( clk, reset, WX3463, n3308 );
dff WX3273_reg ( clk, reset, WX3273, n2833 );
dff WX3337_reg ( clk, reset, WX3337, n2993 );
dff WX3401_reg ( clk, reset, WX3401, n3153 );
dff WX3465_reg ( clk, reset, WX3465, n3313 );
dff WX3275_reg ( clk, reset, WX3275, n2838 );
dff WX3339_reg ( clk, reset, WX3339, n2998 );
dff WX3403_reg ( clk, reset, WX3403, n3158 );
dff WX3467_reg ( clk, reset, WX3467, n3318 );
dff WX3277_reg ( clk, reset, WX3277, n2843 );
dff WX3341_reg ( clk, reset, WX3341, n3003 );
dff WX3405_reg ( clk, reset, WX3405, n3163 );
dff WX3469_reg ( clk, reset, WX3469, n3323 );
dff WX3279_reg ( clk, reset, WX3279, n2848 );
dff WX3343_reg ( clk, reset, WX3343, n3008 );
dff WX3407_reg ( clk, reset, WX3407, n3168 );
dff WX3471_reg ( clk, reset, WX3471, n3328 );
dff WX3281_reg ( clk, reset, WX3281, n2853 );
dff WX3345_reg ( clk, reset, WX3345, n3013 );
dff WX3409_reg ( clk, reset, WX3409, n3173 );
dff WX3473_reg ( clk, reset, WX3473, n3333 );
dff WX3283_reg ( clk, reset, WX3283, n2858 );
dff WX3347_reg ( clk, reset, WX3347, n3018 );
dff WX3411_reg ( clk, reset, WX3411, n3178 );
dff WX3475_reg ( clk, reset, WX3475, n3338 );
dff WX3285_reg ( clk, reset, WX3285, n2863 );
dff WX3349_reg ( clk, reset, WX3349, n3023 );
dff WX3413_reg ( clk, reset, WX3413, n3183 );
dff WX3477_reg ( clk, reset, WX3477, n3343 );
dff WX3287_reg ( clk, reset, WX3287, n2868 );
dff WX3351_reg ( clk, reset, WX3351, n3028 );
dff WX3415_reg ( clk, reset, WX3415, n3188 );
dff WX3479_reg ( clk, reset, WX3479, n3348 );
dff WX3289_reg ( clk, reset, WX3289, n2873 );
dff WX3353_reg ( clk, reset, WX3353, n3033 );
dff WX3417_reg ( clk, reset, WX3417, n3193 );
dff WX3481_reg ( clk, reset, WX3481, n3353 );
dff WX3291_reg ( clk, reset, WX3291, n2878 );
dff WX3355_reg ( clk, reset, WX3355, n3038 );
dff WX3419_reg ( clk, reset, WX3419, n3198 );
dff WX3483_reg ( clk, reset, WX3483, n3358 );
dff WX3293_reg ( clk, reset, WX3293, n2883 );
dff WX3357_reg ( clk, reset, WX3357, n3043 );
dff WX3421_reg ( clk, reset, WX3421, n3203 );
dff WX3485_reg ( clk, reset, WX3485, n3363 );
dff WX1938_reg ( clk, reset, WX1938, n1800 );
dff WX2002_reg ( clk, reset, WX2002, n1960 );
dff WX2066_reg ( clk, reset, WX2066, n2120 );
dff WX2130_reg ( clk, reset, WX2130, n2280 );
dff CRC_OUT_8_31_reg ( clk, reset, CRC_OUT_8_31, n2564 );
dff CRC_OUT_8_0_reg ( clk, reset, CRC_OUT_8_0, n2440 );
dff CRC_OUT_8_1_reg ( clk, reset, CRC_OUT_8_1, n2444 );
dff CRC_OUT_8_2_reg ( clk, reset, CRC_OUT_8_2, n2448 );
dff CRC_OUT_8_3_reg ( clk, reset, CRC_OUT_8_3, n2452 );
dff CRC_OUT_8_4_reg ( clk, reset, CRC_OUT_8_4, n2456 );
dff CRC_OUT_8_5_reg ( clk, reset, CRC_OUT_8_5, n2460 );
dff CRC_OUT_8_6_reg ( clk, reset, CRC_OUT_8_6, n2464 );
dff CRC_OUT_8_7_reg ( clk, reset, CRC_OUT_8_7, n2468 );
dff CRC_OUT_8_8_reg ( clk, reset, CRC_OUT_8_8, n2472 );
dff CRC_OUT_8_9_reg ( clk, reset, CRC_OUT_8_9, n2476 );
dff CRC_OUT_8_10_reg ( clk, reset, CRC_OUT_8_10, n2480 );
dff CRC_OUT_8_11_reg ( clk, reset, CRC_OUT_8_11, n2484 );
dff CRC_OUT_8_12_reg ( clk, reset, CRC_OUT_8_12, n2488 );
dff CRC_OUT_8_13_reg ( clk, reset, CRC_OUT_8_13, n2492 );
dff CRC_OUT_8_14_reg ( clk, reset, CRC_OUT_8_14, n2496 );
dff CRC_OUT_8_15_reg ( clk, reset, CRC_OUT_8_15, n2500 );
dff CRC_OUT_8_16_reg ( clk, reset, CRC_OUT_8_16, n2504 );
dff CRC_OUT_8_17_reg ( clk, reset, CRC_OUT_8_17, n2508 );
dff CRC_OUT_8_18_reg ( clk, reset, CRC_OUT_8_18, n2512 );
dff CRC_OUT_8_19_reg ( clk, reset, CRC_OUT_8_19, n2516 );
dff CRC_OUT_8_20_reg ( clk, reset, CRC_OUT_8_20, n2520 );
dff CRC_OUT_8_21_reg ( clk, reset, CRC_OUT_8_21, n2524 );
dff CRC_OUT_8_22_reg ( clk, reset, CRC_OUT_8_22, n2528 );
dff CRC_OUT_8_23_reg ( clk, reset, CRC_OUT_8_23, n2532 );
dff CRC_OUT_8_24_reg ( clk, reset, CRC_OUT_8_24, n2536 );
dff CRC_OUT_8_25_reg ( clk, reset, CRC_OUT_8_25, n2540 );
dff CRC_OUT_8_26_reg ( clk, reset, CRC_OUT_8_26, n2544 );
dff CRC_OUT_8_27_reg ( clk, reset, CRC_OUT_8_27, n2548 );
dff CRC_OUT_8_28_reg ( clk, reset, CRC_OUT_8_28, n2552 );
dff CRC_OUT_8_29_reg ( clk, reset, CRC_OUT_8_29, n2556 );
dff CRC_OUT_8_30_reg ( clk, reset, CRC_OUT_8_30, n2560 );
dff WX1940_reg ( clk, reset, WX1940, n1805 );
dff WX2004_reg ( clk, reset, WX2004, n1965 );
dff WX2068_reg ( clk, reset, WX2068, n2125 );
dff WX2132_reg ( clk, reset, WX2132, n2285 );
dff WX1942_reg ( clk, reset, WX1942, n1810 );
dff WX2006_reg ( clk, reset, WX2006, n1970 );
dff WX2070_reg ( clk, reset, WX2070, n2130 );
dff WX2134_reg ( clk, reset, WX2134, n2290 );
dff WX1944_reg ( clk, reset, WX1944, n1815 );
dff WX2008_reg ( clk, reset, WX2008, n1975 );
dff WX2072_reg ( clk, reset, WX2072, n2135 );
dff WX2136_reg ( clk, reset, WX2136, n2295 );
dff WX1946_reg ( clk, reset, WX1946, n1820 );
dff WX2010_reg ( clk, reset, WX2010, n1980 );
dff WX2074_reg ( clk, reset, WX2074, n2140 );
dff WX2138_reg ( clk, reset, WX2138, n2300 );
dff WX1948_reg ( clk, reset, WX1948, n1825 );
dff WX2012_reg ( clk, reset, WX2012, n1985 );
dff WX2076_reg ( clk, reset, WX2076, n2145 );
dff WX2140_reg ( clk, reset, WX2140, n2305 );
dff WX1950_reg ( clk, reset, WX1950, n1830 );
dff WX2014_reg ( clk, reset, WX2014, n1990 );
dff WX2078_reg ( clk, reset, WX2078, n2150 );
dff WX2142_reg ( clk, reset, WX2142, n2310 );
dff WX1952_reg ( clk, reset, WX1952, n1835 );
dff WX2016_reg ( clk, reset, WX2016, n1995 );
dff WX2080_reg ( clk, reset, WX2080, n2155 );
dff WX2144_reg ( clk, reset, WX2144, n2315 );
dff WX1954_reg ( clk, reset, WX1954, n1840 );
dff WX2018_reg ( clk, reset, WX2018, n2000 );
dff WX2082_reg ( clk, reset, WX2082, n2160 );
dff WX2146_reg ( clk, reset, WX2146, n2320 );
dff WX1956_reg ( clk, reset, WX1956, n1845 );
dff WX2020_reg ( clk, reset, WX2020, n2005 );
dff WX2084_reg ( clk, reset, WX2084, n2165 );
dff WX2148_reg ( clk, reset, WX2148, n2325 );
dff WX1958_reg ( clk, reset, WX1958, n1850 );
dff WX2022_reg ( clk, reset, WX2022, n2010 );
dff WX2086_reg ( clk, reset, WX2086, n2170 );
dff WX2150_reg ( clk, reset, WX2150, n2330 );
dff WX1960_reg ( clk, reset, WX1960, n1855 );
dff WX2024_reg ( clk, reset, WX2024, n2015 );
dff WX2088_reg ( clk, reset, WX2088, n2175 );
dff WX2152_reg ( clk, reset, WX2152, n2335 );
dff WX1962_reg ( clk, reset, WX1962, n1860 );
dff WX2026_reg ( clk, reset, WX2026, n2020 );
dff WX2090_reg ( clk, reset, WX2090, n2180 );
dff WX2154_reg ( clk, reset, WX2154, n2340 );
dff WX1964_reg ( clk, reset, WX1964, n1865 );
dff WX2028_reg ( clk, reset, WX2028, n2025 );
dff WX2092_reg ( clk, reset, WX2092, n2185 );
dff WX2156_reg ( clk, reset, WX2156, n2345 );
dff WX1966_reg ( clk, reset, WX1966, n1870 );
dff WX2030_reg ( clk, reset, WX2030, n2030 );
dff WX2094_reg ( clk, reset, WX2094, n2190 );
dff WX2158_reg ( clk, reset, WX2158, n2350 );
dff WX1968_reg ( clk, reset, WX1968, n1875 );
dff WX2032_reg ( clk, reset, WX2032, n2035 );
dff WX2096_reg ( clk, reset, WX2096, n2195 );
dff WX2160_reg ( clk, reset, WX2160, n2355 );
dff WX1970_reg ( clk, reset, WX1970, n1880 );
dff WX2034_reg ( clk, reset, WX2034, n2040 );
dff WX2098_reg ( clk, reset, WX2098, n2200 );
dff WX2162_reg ( clk, reset, WX2162, n2360 );
dff WX1972_reg ( clk, reset, WX1972, n1885 );
dff WX2036_reg ( clk, reset, WX2036, n2045 );
dff WX2100_reg ( clk, reset, WX2100, n2205 );
dff WX2164_reg ( clk, reset, WX2164, n2365 );
dff WX1974_reg ( clk, reset, WX1974, n1890 );
dff WX2038_reg ( clk, reset, WX2038, n2050 );
dff WX2102_reg ( clk, reset, WX2102, n2210 );
dff WX2166_reg ( clk, reset, WX2166, n2370 );
dff WX1976_reg ( clk, reset, WX1976, n1895 );
dff WX2040_reg ( clk, reset, WX2040, n2055 );
dff WX2104_reg ( clk, reset, WX2104, n2215 );
dff WX2168_reg ( clk, reset, WX2168, n2375 );
dff WX1978_reg ( clk, reset, WX1978, n1900 );
dff WX2042_reg ( clk, reset, WX2042, n2060 );
dff WX2106_reg ( clk, reset, WX2106, n2220 );
dff WX2170_reg ( clk, reset, WX2170, n2380 );
dff WX1980_reg ( clk, reset, WX1980, n1905 );
dff WX2044_reg ( clk, reset, WX2044, n2065 );
dff WX2108_reg ( clk, reset, WX2108, n2225 );
dff WX2172_reg ( clk, reset, WX2172, n2385 );
dff WX1982_reg ( clk, reset, WX1982, n1910 );
dff WX2046_reg ( clk, reset, WX2046, n2070 );
dff WX2110_reg ( clk, reset, WX2110, n2230 );
dff WX2174_reg ( clk, reset, WX2174, n2390 );
dff WX1984_reg ( clk, reset, WX1984, n1915 );
dff WX2048_reg ( clk, reset, WX2048, n2075 );
dff WX2112_reg ( clk, reset, WX2112, n2235 );
dff WX2176_reg ( clk, reset, WX2176, n2395 );
dff WX1986_reg ( clk, reset, WX1986, n1920 );
dff WX2050_reg ( clk, reset, WX2050, n2080 );
dff WX2114_reg ( clk, reset, WX2114, n2240 );
dff WX2178_reg ( clk, reset, WX2178, n2400 );
dff WX1988_reg ( clk, reset, WX1988, n1925 );
dff WX2052_reg ( clk, reset, WX2052, n2085 );
dff WX2116_reg ( clk, reset, WX2116, n2245 );
dff WX2180_reg ( clk, reset, WX2180, n2405 );
dff WX1990_reg ( clk, reset, WX1990, n1930 );
dff WX2054_reg ( clk, reset, WX2054, n2090 );
dff WX2118_reg ( clk, reset, WX2118, n2250 );
dff WX2182_reg ( clk, reset, WX2182, n2410 );
dff WX1992_reg ( clk, reset, WX1992, n1935 );
dff WX2056_reg ( clk, reset, WX2056, n2095 );
dff WX2120_reg ( clk, reset, WX2120, n2255 );
dff WX2184_reg ( clk, reset, WX2184, n2415 );
dff WX1994_reg ( clk, reset, WX1994, n1940 );
dff WX2058_reg ( clk, reset, WX2058, n2100 );
dff WX2122_reg ( clk, reset, WX2122, n2260 );
dff WX2186_reg ( clk, reset, WX2186, n2420 );
dff WX1996_reg ( clk, reset, WX1996, n1945 );
dff WX2060_reg ( clk, reset, WX2060, n2105 );
dff WX2124_reg ( clk, reset, WX2124, n2265 );
dff WX2188_reg ( clk, reset, WX2188, n2425 );
dff WX1998_reg ( clk, reset, WX1998, n1950 );
dff WX2062_reg ( clk, reset, WX2062, n2110 );
dff WX2126_reg ( clk, reset, WX2126, n2270 );
dff WX2190_reg ( clk, reset, WX2190, n2430 );
dff WX2000_reg ( clk, reset, WX2000, n1955 );
dff WX2064_reg ( clk, reset, WX2064, n2115 );
dff WX2128_reg ( clk, reset, WX2128, n2275 );
dff WX2192_reg ( clk, reset, WX2192, n2435 );
dff WX645_reg ( clk, reset, WX645, n872 );
dff WX709_reg ( clk, reset, WX709, n1032 );
dff WX773_reg ( clk, reset, WX773, n1192 );
dff WX837_reg ( clk, reset, WX837, n1352 );
dff CRC_OUT_9_31_reg ( clk, reset, CRC_OUT_9_31, n1636 );
dff CRC_OUT_9_0_reg ( clk, reset, CRC_OUT_9_0, n1512 );
dff CRC_OUT_9_1_reg ( clk, reset, CRC_OUT_9_1, n1516 );
dff CRC_OUT_9_2_reg ( clk, reset, CRC_OUT_9_2, n1520 );
dff CRC_OUT_9_3_reg ( clk, reset, CRC_OUT_9_3, n1524 );
dff CRC_OUT_9_4_reg ( clk, reset, CRC_OUT_9_4, n1528 );
dff CRC_OUT_9_5_reg ( clk, reset, CRC_OUT_9_5, n1532 );
dff CRC_OUT_9_6_reg ( clk, reset, CRC_OUT_9_6, n1536 );
dff WX695_reg ( clk, reset, WX695, n997 );
dff WX759_reg ( clk, reset, WX759, n1157 );
dff WX823_reg ( clk, reset, WX823, n1317 );
dff WX887_reg ( clk, reset, WX887, n1477 );
dff CRC_OUT_9_7_reg ( clk, reset, CRC_OUT_9_7, n1540 );
dff WX693_reg ( clk, reset, WX693, n992 );
dff WX757_reg ( clk, reset, WX757, n1152 );
dff WX821_reg ( clk, reset, WX821, n1312 );
dff WX885_reg ( clk, reset, WX885, n1472 );
dff CRC_OUT_9_8_reg ( clk, reset, CRC_OUT_9_8, n1544 );
dff WX691_reg ( clk, reset, WX691, n987 );
dff WX755_reg ( clk, reset, WX755, n1147 );
dff WX819_reg ( clk, reset, WX819, n1307 );
dff WX883_reg ( clk, reset, WX883, n1467 );
dff CRC_OUT_9_9_reg ( clk, reset, CRC_OUT_9_9, n1548 );
dff WX689_reg ( clk, reset, WX689, n982 );
dff WX753_reg ( clk, reset, WX753, n1142 );
dff WX817_reg ( clk, reset, WX817, n1302 );
dff WX881_reg ( clk, reset, WX881, n1462 );
dff CRC_OUT_9_10_reg ( clk, reset, CRC_OUT_9_10, n1552 );
dff WX687_reg ( clk, reset, WX687, n977 );
dff WX751_reg ( clk, reset, WX751, n1137 );
dff WX815_reg ( clk, reset, WX815, n1297 );
dff WX879_reg ( clk, reset, WX879, n1457 );
dff CRC_OUT_9_11_reg ( clk, reset, CRC_OUT_9_11, n1556 );
dff WX685_reg ( clk, reset, WX685, n972 );
dff WX749_reg ( clk, reset, WX749, n1132 );
dff WX813_reg ( clk, reset, WX813, n1292 );
dff WX877_reg ( clk, reset, WX877, n1452 );
dff CRC_OUT_9_12_reg ( clk, reset, CRC_OUT_9_12, n1560 );
dff WX683_reg ( clk, reset, WX683, n967 );
dff WX747_reg ( clk, reset, WX747, n1127 );
dff WX811_reg ( clk, reset, WX811, n1287 );
dff WX875_reg ( clk, reset, WX875, n1447 );
dff CRC_OUT_9_13_reg ( clk, reset, CRC_OUT_9_13, n1564 );
dff WX681_reg ( clk, reset, WX681, n962 );
dff WX745_reg ( clk, reset, WX745, n1122 );
dff WX809_reg ( clk, reset, WX809, n1282 );
dff WX873_reg ( clk, reset, WX873, n1442 );
dff CRC_OUT_9_14_reg ( clk, reset, CRC_OUT_9_14, n1568 );
dff WX679_reg ( clk, reset, WX679, n957 );
dff WX743_reg ( clk, reset, WX743, n1117 );
dff WX807_reg ( clk, reset, WX807, n1277 );
dff WX871_reg ( clk, reset, WX871, n1437 );
dff CRC_OUT_9_15_reg ( clk, reset, CRC_OUT_9_15, n1572 );
dff WX677_reg ( clk, reset, WX677, n952 );
dff WX741_reg ( clk, reset, WX741, n1112 );
dff WX805_reg ( clk, reset, WX805, n1272 );
dff WX869_reg ( clk, reset, WX869, n1432 );
dff CRC_OUT_9_16_reg ( clk, reset, CRC_OUT_9_16, n1576 );
dff WX675_reg ( clk, reset, WX675, n947 );
dff WX739_reg ( clk, reset, WX739, n1107 );
dff WX803_reg ( clk, reset, WX803, n1267 );
dff WX867_reg ( clk, reset, WX867, n1427 );
dff CRC_OUT_9_17_reg ( clk, reset, CRC_OUT_9_17, n1580 );
dff WX673_reg ( clk, reset, WX673, n942 );
dff WX737_reg ( clk, reset, WX737, n1102 );
dff WX801_reg ( clk, reset, WX801, n1262 );
dff WX865_reg ( clk, reset, WX865, n1422 );
dff CRC_OUT_9_18_reg ( clk, reset, CRC_OUT_9_18, n1584 );
dff WX671_reg ( clk, reset, WX671, n937 );
dff WX735_reg ( clk, reset, WX735, n1097 );
dff WX799_reg ( clk, reset, WX799, n1257 );
dff WX863_reg ( clk, reset, WX863, n1417 );
dff CRC_OUT_9_19_reg ( clk, reset, CRC_OUT_9_19, n1588 );
dff WX669_reg ( clk, reset, WX669, n932 );
dff WX733_reg ( clk, reset, WX733, n1092 );
dff WX797_reg ( clk, reset, WX797, n1252 );
dff WX861_reg ( clk, reset, WX861, n1412 );
dff CRC_OUT_9_20_reg ( clk, reset, CRC_OUT_9_20, n1592 );
dff WX667_reg ( clk, reset, WX667, n927 );
dff WX731_reg ( clk, reset, WX731, n1087 );
dff WX795_reg ( clk, reset, WX795, n1247 );
dff WX859_reg ( clk, reset, WX859, n1407 );
dff CRC_OUT_9_21_reg ( clk, reset, CRC_OUT_9_21, n1596 );
dff WX665_reg ( clk, reset, WX665, n922 );
dff WX729_reg ( clk, reset, WX729, n1082 );
dff WX793_reg ( clk, reset, WX793, n1242 );
dff WX857_reg ( clk, reset, WX857, n1402 );
dff CRC_OUT_9_22_reg ( clk, reset, CRC_OUT_9_22, n1600 );
dff WX663_reg ( clk, reset, WX663, n917 );
dff WX727_reg ( clk, reset, WX727, n1077 );
dff WX791_reg ( clk, reset, WX791, n1237 );
dff WX855_reg ( clk, reset, WX855, n1397 );
dff CRC_OUT_9_23_reg ( clk, reset, CRC_OUT_9_23, n1604 );
dff WX661_reg ( clk, reset, WX661, n912 );
dff WX725_reg ( clk, reset, WX725, n1072 );
dff WX789_reg ( clk, reset, WX789, n1232 );
dff WX853_reg ( clk, reset, WX853, n1392 );
dff CRC_OUT_9_24_reg ( clk, reset, CRC_OUT_9_24, n1608 );
dff WX659_reg ( clk, reset, WX659, n907 );
dff WX723_reg ( clk, reset, WX723, n1067 );
dff WX787_reg ( clk, reset, WX787, n1227 );
dff WX851_reg ( clk, reset, WX851, n1387 );
dff CRC_OUT_9_25_reg ( clk, reset, CRC_OUT_9_25, n1612 );
dff WX657_reg ( clk, reset, WX657, n902 );
dff WX721_reg ( clk, reset, WX721, n1062 );
dff WX785_reg ( clk, reset, WX785, n1222 );
dff WX849_reg ( clk, reset, WX849, n1382 );
dff CRC_OUT_9_26_reg ( clk, reset, CRC_OUT_9_26, n1616 );
dff WX655_reg ( clk, reset, WX655, n897 );
dff WX719_reg ( clk, reset, WX719, n1057 );
dff WX783_reg ( clk, reset, WX783, n1217 );
dff WX847_reg ( clk, reset, WX847, n1377 );
dff CRC_OUT_9_27_reg ( clk, reset, CRC_OUT_9_27, n1620 );
dff WX653_reg ( clk, reset, WX653, n892 );
dff WX717_reg ( clk, reset, WX717, n1052 );
dff WX781_reg ( clk, reset, WX781, n1212 );
dff WX845_reg ( clk, reset, WX845, n1372 );
dff CRC_OUT_9_28_reg ( clk, reset, CRC_OUT_9_28, n1624 );
dff WX651_reg ( clk, reset, WX651, n887 );
dff WX715_reg ( clk, reset, WX715, n1047 );
dff WX779_reg ( clk, reset, WX779, n1207 );
dff WX843_reg ( clk, reset, WX843, n1367 );
dff CRC_OUT_9_29_reg ( clk, reset, CRC_OUT_9_29, n1628 );
dff WX649_reg ( clk, reset, WX649, n882 );
dff WX713_reg ( clk, reset, WX713, n1042 );
dff WX777_reg ( clk, reset, WX777, n1202 );
dff WX841_reg ( clk, reset, WX841, n1362 );
dff CRC_OUT_9_30_reg ( clk, reset, CRC_OUT_9_30, n1632 );
dff WX647_reg ( clk, reset, WX647, n877 );
dff WX711_reg ( clk, reset, WX711, n1037 );
dff WX775_reg ( clk, reset, WX775, n1197 );
dff WX839_reg ( clk, reset, WX839, n1357 );
dff WX697_reg ( clk, reset, WX697, n1002 );
dff WX761_reg ( clk, reset, WX761, n1162 );
dff WX825_reg ( clk, reset, WX825, n1322 );
dff WX889_reg ( clk, reset, WX889, n1482 );
dff WX699_reg ( clk, reset, WX699, n1007 );
dff WX763_reg ( clk, reset, WX763, n1167 );
dff WX827_reg ( clk, reset, WX827, n1327 );
dff WX891_reg ( clk, reset, WX891, n1487 );
dff WX701_reg ( clk, reset, WX701, n1012 );
dff WX765_reg ( clk, reset, WX765, n1172 );
dff WX829_reg ( clk, reset, WX829, n1332 );
dff WX893_reg ( clk, reset, WX893, n1492 );
dff WX703_reg ( clk, reset, WX703, n1017 );
dff WX767_reg ( clk, reset, WX767, n1177 );
dff WX831_reg ( clk, reset, WX831, n1337 );
dff WX895_reg ( clk, reset, WX895, n1497 );
dff WX705_reg ( clk, reset, WX705, n1022 );
dff WX769_reg ( clk, reset, WX769, n1182 );
dff WX833_reg ( clk, reset, WX833, n1342 );
dff WX897_reg ( clk, reset, WX897, n1502 );
dff WX707_reg ( clk, reset, WX707, n1027 );
dff WX771_reg ( clk, reset, WX771, n1187 );
dff WX835_reg ( clk, reset, WX835, n1347 );
dff WX899_reg ( clk, reset, WX899, n1507 );
buf U5152 ( n4387, n4389 );
buf U5153 ( n4339, n4342 );
buf U5154 ( n4335, n4343 );
buf U5155 ( n4337, n4343 );
buf U5156 ( n4338, n4343 );
buf U5157 ( n4425, n4435 );
buf U5158 ( n4428, n4434 );
buf U5159 ( n4427, n4434 );
buf U5160 ( n4432, n4433 );
buf U5161 ( n4431, n4433 );
buf U5162 ( n4429, n4434 );
buf U5163 ( n4430, n4433 );
buf U5164 ( n4426, n4435 );
buf U5165 ( n4386, n4389 );
buf U5166 ( n4385, n4389 );
buf U5167 ( n4383, n4390 );
buf U5168 ( n4382, n4390 );
buf U5169 ( n4381, n4390 );
buf U5170 ( n4378, n4391 );
buf U5171 ( n4379, n4391 );
buf U5172 ( n4389, n4345 );
buf U5173 ( n4342, n4319 );
buf U5174 ( n4343, n4319 );
buf U5175 ( n4466, n4468 );
buf U5176 ( n4463, n4469 );
buf U5177 ( n4464, n4469 );
buf U5178 ( n4434, n4393 );
buf U5179 ( n4433, n4393 );
buf U5180 ( n4462, n4469 );
buf U5181 ( n4465, n4468 );
buf U5182 ( n4461, n4470 );
buf U5183 ( n4460, n4470 );
buf U5184 ( n4390, n4345 );
buf U5185 ( n4345, n360 );
buf U5186 ( n4393, n356 );
buf U5187 ( n4468, n4436 );
buf U5188 ( n4469, n4436 );
buf U5189 ( n4477, n4494 );
buf U5190 ( n4475, n4495 );
buf U5191 ( n4436, n352 );
buf U5192 ( n4480, n4494 );
buf U5193 ( n4479, n4494 );
buf U5194 ( n4474, n4495 );
buf U5195 ( n4491, n4492 );
buf U5196 ( n4478, n4494 );
buf U5197 ( n4476, n4495 );
buf U5198 ( n4486, n4493 );
buf U5199 ( n4487, n4492 );
buf U5200 ( n4488, n4492 );
buf U5201 ( n4489, n4492 );
buf U5202 ( n4490, n4492 );
buf U5203 ( n4482, n4493 );
buf U5204 ( n4481, n4494 );
buf U5205 ( n4483, n4493 );
buf U5206 ( n4484, n4493 );
buf U5207 ( n4485, n4493 );
buf U5208 ( n4494, RESET );
buf U5209 ( n4472, TM1 );
buf U5210 ( n4492, RESET );
buf U5211 ( n4493, RESET );
buf U5212 ( n4346, n4387 );
buf U5213 ( n4349, n4387 );
buf U5214 ( n4347, n4387 );
buf U5215 ( n4351, n4386 );
buf U5216 ( n4350, n4386 );
buf U5217 ( n4355, n4385 );
buf U5218 ( n4354, n4385 );
buf U5219 ( n4353, n4386 );
buf U5220 ( n4358, n4383 );
buf U5221 ( n4357, n4385 );
buf U5222 ( n4362, n4382 );
buf U5223 ( n4361, n4383 );
buf U5224 ( n4359, n4383 );
buf U5225 ( n4366, n4381 );
buf U5226 ( n4365, n4382 );
buf U5227 ( n4363, n4382 );
buf U5228 ( n4369, n4381 );
buf U5229 ( n4367, n4381 );
buf U5230 ( n4375, n4378 );
buf U5231 ( n4374, n4378 );
buf U5232 ( n4373, n4379 );
buf U5233 ( n4371, n4379 );
buf U5234 ( n4370, n4379 );
buf U5235 ( n4377, n4378 );
not U5236 ( n4321, n4339 );
not U5237 ( n4322, n4339 );
not U5238 ( n4333, n4335 );
not U5239 ( n4330, n4337 );
not U5240 ( n4326, n4338 );
not U5241 ( n4325, n4338 );
not U5242 ( n4334, n4335 );
not U5243 ( n4331, n4335 );
not U5244 ( n4329, n4337 );
not U5245 ( n4327, n4337 );
not U5246 ( n4323, n4338 );
buf U5247 ( n4407, n4429 );
buf U5248 ( n4409, n4429 );
buf U5249 ( n4413, n4428 );
buf U5250 ( n4411, n4428 );
buf U5251 ( n4410, n4428 );
buf U5252 ( n4415, n4427 );
buf U5253 ( n4414, n4427 );
buf U5254 ( n4417, n4427 );
buf U5255 ( n4394, n4432 );
buf U5256 ( n4398, n4431 );
buf U5257 ( n4397, n4432 );
buf U5258 ( n4395, n4432 );
buf U5259 ( n4402, n4430 );
buf U5260 ( n4401, n4431 );
buf U5261 ( n4399, n4431 );
buf U5262 ( n4406, n4429 );
buf U5263 ( n4405, n4430 );
buf U5264 ( n4403, n4430 );
buf U5265 ( n4419, n4426 );
buf U5266 ( n4418, n4426 );
buf U5267 ( n4423, n4425 );
buf U5268 ( n4422, n4425 );
buf U5269 ( n4421, n4426 );
buf U5270 ( n4424, n4425 );
buf U5271 ( n4447, n4464 );
buf U5272 ( n4450, n4463 );
buf U5273 ( n4449, n4463 );
buf U5274 ( n4448, n4463 );
buf U5275 ( n4452, n4462 );
buf U5276 ( n4451, n4462 );
buf U5277 ( n4453, n4462 );
buf U5278 ( n4442, n4465 );
buf U5279 ( n4441, n4466 );
buf U5280 ( n4440, n4466 );
buf U5281 ( n4446, n4464 );
buf U5282 ( n4445, n4464 );
buf U5283 ( n4444, n4465 );
buf U5284 ( n4443, n4465 );
buf U5285 ( n4439, n4466 );
buf U5286 ( n4455, n4461 );
buf U5287 ( n4454, n4461 );
buf U5288 ( n4457, n4460 );
buf U5289 ( n4456, n4461 );
buf U5290 ( n4458, n4460 );
buf U5291 ( n4459, n4460 );
buf U5292 ( n4438, n4467 );
buf U5293 ( n4437, n4467 );
buf U5294 ( n4341, n4342 );
nor U5295 ( n666, n4346, n4675 );
buf U5296 ( n4391, n4345 );
not U5297 ( n4588, n4608 );
buf U5298 ( n4467, n4468 );
buf U5299 ( n4435, n4393 );
not U5300 ( n4523, n4601 );
not U5301 ( n4587, n4627 );
not U5302 ( n4585, n4626 );
not U5303 ( n4586, n4626 );
not U5304 ( n4522, n4600 );
not U5305 ( n4521, n4600 );
not U5306 ( n4520, n4600 );
not U5307 ( n4508, n4595 );
not U5308 ( n4512, n4596 );
not U5309 ( n4517, n4598 );
not U5310 ( n4516, n4597 );
not U5311 ( n4513, n4596 );
not U5312 ( n4514, n4597 );
not U5313 ( n4515, n4597 );
not U5314 ( n4507, n4593 );
not U5315 ( n4506, n4593 );
not U5316 ( n4505, n4593 );
not U5317 ( n4504, n4592 );
not U5318 ( n4518, n4598 );
not U5319 ( n4519, n4598 );
not U5320 ( n4511, n4596 );
not U5321 ( n4510, n4595 );
not U5322 ( n4509, n4595 );
not U5323 ( n4524, n4601 );
not U5324 ( n4565, n4618 );
not U5325 ( n4560, n4616 );
not U5326 ( n4562, n4617 );
not U5327 ( n4564, n4618 );
not U5328 ( n4561, n4617 );
not U5329 ( n4563, n4617 );
not U5330 ( n4556, n4615 );
not U5331 ( n4551, n4612 );
not U5332 ( n4553, n4613 );
not U5333 ( n4555, n4615 );
not U5334 ( n4554, n4613 );
not U5335 ( n4552, n4613 );
not U5336 ( n4566, n4618 );
not U5337 ( n4559, n4616 );
not U5338 ( n4578, n4623 );
not U5339 ( n4558, n4616 );
not U5340 ( n4581, n4625 );
not U5341 ( n4580, n4625 );
not U5342 ( n4577, n4623 );
not U5343 ( n4557, n4615 );
not U5344 ( n4567, n4620 );
not U5345 ( n4582, n4625 );
not U5346 ( n4572, n4621 );
not U5347 ( n4569, n4620 );
not U5348 ( n4571, n4621 );
not U5349 ( n4570, n4621 );
not U5350 ( n4568, n4620 );
not U5351 ( n4583, n4626 );
not U5352 ( n4574, n4622 );
not U5353 ( n4576, n4623 );
not U5354 ( n4575, n4622 );
not U5355 ( n4573, n4622 );
not U5356 ( n4547, n4611 );
not U5357 ( n4548, n4611 );
not U5358 ( n4543, n4610 );
not U5359 ( n4541, n4608 );
not U5360 ( n4546, n4611 );
not U5361 ( n4545, n4610 );
not U5362 ( n4550, n4612 );
not U5363 ( n4544, n4610 );
not U5364 ( n4549, n4612 );
not U5365 ( n4542, n4608 );
not U5366 ( n4500, n4591 );
not U5367 ( n4497, n4590 );
not U5368 ( n4502, n4592 );
not U5369 ( n4496, n4590 );
not U5370 ( n4499, n4591 );
not U5371 ( n4498, n4590 );
not U5372 ( n4501, n4591 );
not U5373 ( n4503, n4592 );
not U5374 ( n4534, n4605 );
not U5375 ( n4535, n4606 );
not U5376 ( n4539, n4607 );
not U5377 ( n4537, n4606 );
not U5378 ( n4540, n4607 );
not U5379 ( n4538, n4607 );
not U5380 ( n4536, n4606 );
not U5381 ( n4529, n4603 );
not U5382 ( n4526, n4602 );
not U5383 ( n4533, n4605 );
not U5384 ( n4532, n4605 );
not U5385 ( n4528, n4602 );
not U5386 ( n4527, n4602 );
not U5387 ( n4531, n4603 );
not U5388 ( n4525, n4601 );
not U5389 ( n4530, n4603 );
nand U5390 ( n360, n4472, TM0 );
nand U5391 ( n4267, n4588, n4473 );
not U5392 ( n4608, n4477 );
buf U5393 ( n4319, n680 );
nor U5394 ( n680, n4267, TM0 );
buf U5395 ( n4470, n4436 );
nand U5396 ( n356, n4273, n4523 );
nor U5397 ( n4273, TM0, n4473 );
not U5398 ( n4601, n4475 );
not U5399 ( n4627, n4480 );
not U5400 ( n4626, n4479 );
not U5401 ( n4600, n4475 );
not U5402 ( n4597, n4475 );
not U5403 ( n4593, n4474 );
not U5404 ( n4592, n4474 );
not U5405 ( n4598, n4475 );
not U5406 ( n4596, n4475 );
not U5407 ( n4595, n4474 );
not U5408 ( n4675, n4491 );
not U5409 ( n4617, n4478 );
not U5410 ( n4613, n4477 );
not U5411 ( n4618, n4478 );
not U5412 ( n4616, n4478 );
not U5413 ( n4615, n4478 );
not U5414 ( n4625, n4479 );
not U5415 ( n4621, n4479 );
not U5416 ( n4620, n4478 );
not U5417 ( n4623, n4479 );
not U5418 ( n4622, n4479 );
not U5419 ( n4611, n4477 );
not U5420 ( n4610, n4477 );
not U5421 ( n4612, n4477 );
not U5422 ( n4590, n4474 );
not U5423 ( n4591, n4474 );
not U5424 ( n4607, n4476 );
not U5425 ( n4606, n4476 );
not U5426 ( n4605, n4476 );
not U5427 ( n4602, n4476 );
not U5428 ( n4603, n4476 );
not U5429 ( n4673, n4491 );
not U5430 ( n4653, n4486 );
not U5431 ( n4652, n4486 );
not U5432 ( n4651, n4486 );
not U5433 ( n4650, n4486 );
not U5434 ( n4648, n4486 );
not U5435 ( n4661, n4488 );
not U5436 ( n4660, n4488 );
not U5437 ( n4658, n4487 );
not U5438 ( n4657, n4487 );
not U5439 ( n4656, n4487 );
not U5440 ( n4655, n4487 );
not U5441 ( n4666, n4489 );
not U5442 ( n4665, n4489 );
not U5443 ( n4663, n4489 );
not U5444 ( n4662, n4488 );
not U5445 ( n4670, n4490 );
not U5446 ( n4668, n4490 );
not U5447 ( n4667, n4490 );
not U5448 ( n4637, n4482 );
not U5449 ( n4638, n4482 );
not U5450 ( n4640, n4482 );
not U5451 ( n4672, n4491 );
not U5452 ( n4671, n4491 );
not U5453 ( n4633, n4481 );
not U5454 ( n4635, n4481 );
not U5455 ( n4636, n4481 );
not U5456 ( n4632, n4481 );
not U5457 ( n4641, n4483 );
not U5458 ( n4628, n4480 );
not U5459 ( n4630, n4480 );
not U5460 ( n4631, n4480 );
not U5461 ( n4642, n4483 );
not U5462 ( n4645, n4484 );
not U5463 ( n4643, n4484 );
not U5464 ( n4647, n4485 );
not U5465 ( n4646, n4485 );
not U5466 ( n4473, TM1 );
nand U5467 ( n872, n661, n662 );
nor U5468 ( n661, n667, n668 );
nor U5469 ( n662, n663, n664 );
nor U5470 ( n668, n347, n4406 );
nand U5471 ( n1800, n4134, n4135 );
nor U5472 ( n4134, n4143, n4144 );
nor U5473 ( n4135, n4137, n4138 );
nor U5474 ( n4144, n665, n4410 );
nand U5475 ( n2728, n3627, n3628 );
nor U5476 ( n3627, n3634, n3635 );
nor U5477 ( n3628, n3629, n3630 );
nor U5478 ( n3635, n3636, n4414 );
nand U5479 ( n3656, n3190, n3191 );
nor U5480 ( n3190, n3199, n3200 );
nor U5481 ( n3191, n3192, n3194 );
nor U5482 ( n3200, n3201, n4417 );
nand U5483 ( n4584, n2727, n2729 );
nor U5484 ( n2727, n2736, n2737 );
nor U5485 ( n2729, n2730, n2731 );
nor U5486 ( n2737, n2739, n4421 );
nand U5487 ( n5512, n2296, n2297 );
nor U5488 ( n2296, n2304, n2306 );
nor U5489 ( n2297, n2298, n2299 );
nor U5490 ( n2306, n2307, n4424 );
nand U5491 ( n6440, n1833, n1834 );
nor U5492 ( n1833, n1842, n1843 );
nor U5493 ( n1834, n1836, n1837 );
nor U5494 ( n1843, n1844, n4395 );
nand U5495 ( n7368, n1401, n1403 );
nor U5496 ( n1401, n1410, n1411 );
nor U5497 ( n1403, n1404, n1405 );
nor U5498 ( n1411, n1413, n4399 );
or U5499 ( n8296, n943, n944 );
nand U5500 ( n944, n945, n946 );
nand U5501 ( n943, n949, n950 );
or U5502 ( n945, n4424, n948 );
nor U5503 ( n4200, n4346, n672 );
nor U5504 ( n4214, n4346, n673 );
nor U5505 ( n4228, n4346, n674 );
nor U5506 ( n4242, n4346, n675 );
nor U5507 ( n4255, n4346, n733 );
nor U5508 ( n4270, n4346, n814 );
nor U5509 ( n3685, n4350, n3689 );
nor U5510 ( n3698, n4350, n3702 );
nor U5511 ( n3710, n4349, n3714 );
nor U5512 ( n3723, n4349, n3727 );
nor U5513 ( n3735, n4349, n3739 );
nor U5514 ( n3748, n4349, n3752 );
nor U5515 ( n3760, n4349, n3765 );
nor U5516 ( n3774, n4349, n3779 );
nor U5517 ( n3788, n4349, n3793 );
nor U5518 ( n3802, n4349, n3807 );
nor U5519 ( n3815, n4349, n3820 );
nor U5520 ( n3829, n4349, n3834 );
nor U5521 ( n3843, n4349, n3848 );
nor U5522 ( n3857, n4349, n3862 );
nor U5523 ( n3870, n4347, n3875 );
nor U5524 ( n3884, n4347, n3889 );
nor U5525 ( n3899, n4347, n3905 );
nor U5526 ( n3915, n4347, n3922 );
nor U5527 ( n3932, n4347, n3938 );
nor U5528 ( n3948, n4347, n3954 );
nor U5529 ( n3964, n4347, n3970 );
nor U5530 ( n3980, n4347, n3987 );
nor U5531 ( n3997, n4347, n4003 );
nor U5532 ( n4013, n4347, n4019 );
nor U5533 ( n4029, n4347, n4035 );
nor U5534 ( n4045, n4347, n4052 );
nor U5535 ( n4062, n4346, n4068 );
nor U5536 ( n4078, n4346, n4084 );
nor U5537 ( n4094, n4346, n4100 );
nor U5538 ( n4110, n4346, n4117 );
nor U5539 ( n4127, n4346, n4133 );
nor U5540 ( n3254, n4353, n3257 );
nor U5541 ( n3266, n4353, n3270 );
nor U5542 ( n3279, n4353, n3282 );
nor U5543 ( n3291, n4353, n3295 );
nor U5544 ( n3304, n4353, n3307 );
nor U5545 ( n3316, n4353, n3320 );
nor U5546 ( n3329, n4353, n3332 );
nor U5547 ( n3341, n4353, n3345 );
nor U5548 ( n3354, n4353, n3357 );
nor U5549 ( n3366, n4351, n3370 );
nor U5550 ( n3379, n4351, n3383 );
nor U5551 ( n3393, n4351, n3397 );
nor U5552 ( n3406, n4351, n3410 );
nor U5553 ( n3419, n4351, n3423 );
nor U5554 ( n3433, n4351, n3437 );
nor U5555 ( n3446, n4351, n3450 );
nor U5556 ( n3461, n4351, n3465 );
nor U5557 ( n3475, n4351, n3479 );
nor U5558 ( n3490, n4351, n3494 );
nor U5559 ( n3502, n4351, n3505 );
nor U5560 ( n3513, n4351, n3516 );
nor U5561 ( n3524, n4350, n3527 );
nor U5562 ( n3535, n4350, n3538 );
nor U5563 ( n3546, n4350, n3549 );
nor U5564 ( n3557, n4350, n3560 );
nor U5565 ( n3568, n4350, n3571 );
nor U5566 ( n3579, n4350, n3582 );
nor U5567 ( n3590, n4350, n3593 );
nor U5568 ( n3601, n4350, n3604 );
nor U5569 ( n3612, n4350, n3615 );
nor U5570 ( n3623, n4350, n3626 );
nor U5571 ( n2791, n4357, n2795 );
nor U5572 ( n2804, n4357, n2807 );
nor U5573 ( n2816, n4357, n2820 );
nor U5574 ( n2829, n4357, n2832 );
nor U5575 ( n2841, n4355, n2845 );
nor U5576 ( n2854, n4355, n2857 );
nor U5577 ( n2866, n4355, n2870 );
nor U5578 ( n2879, n4355, n2882 );
nor U5579 ( n2891, n4355, n2895 );
nor U5580 ( n2904, n4355, n2907 );
nor U5581 ( n2916, n4355, n2920 );
nor U5582 ( n2929, n4355, n2932 );
nor U5583 ( n2941, n4355, n2945 );
nor U5584 ( n2954, n4355, n2957 );
nor U5585 ( n2966, n4355, n2970 );
nor U5586 ( n2979, n4355, n2982 );
nor U5587 ( n2992, n4354, n2996 );
nor U5588 ( n3006, n4354, n3010 );
nor U5589 ( n3020, n4354, n3024 );
nor U5590 ( n3034, n4354, n3037 );
nor U5591 ( n3047, n4354, n3051 );
nor U5592 ( n3061, n4354, n3065 );
nor U5593 ( n3075, n4354, n3079 );
nor U5594 ( n3089, n4354, n3092 );
nor U5595 ( n3102, n4354, n3106 );
nor U5596 ( n3116, n4354, n3120 );
nor U5597 ( n3130, n4354, n3134 );
nor U5598 ( n3144, n4354, n3147 );
nor U5599 ( n3157, n4353, n3161 );
nor U5600 ( n3171, n4353, n3175 );
nor U5601 ( n3185, n4353, n3189 );
nor U5602 ( n2359, n4359, n2363 );
nor U5603 ( n2372, n4359, n2376 );
nor U5604 ( n2384, n4359, n2388 );
nor U5605 ( n2397, n4359, n2401 );
nor U5606 ( n2409, n4359, n2413 );
nor U5607 ( n2422, n4359, n2426 );
nor U5608 ( n2434, n4359, n2438 );
nor U5609 ( n2447, n4359, n2451 );
nor U5610 ( n2461, n4359, n2465 );
nor U5611 ( n2474, n4359, n2478 );
nor U5612 ( n2487, n4359, n2491 );
nor U5613 ( n2501, n4358, n2505 );
nor U5614 ( n2514, n4358, n2518 );
nor U5615 ( n2527, n4358, n2531 );
nor U5616 ( n2541, n4358, n2545 );
nor U5617 ( n2554, n4358, n2558 );
nor U5618 ( n2568, n4358, n2571 );
nor U5619 ( n2579, n4358, n2582 );
nor U5620 ( n2590, n4358, n2593 );
nor U5621 ( n2601, n4358, n2604 );
nor U5622 ( n2612, n4358, n2615 );
nor U5623 ( n2623, n4358, n2626 );
nor U5624 ( n2634, n4358, n2637 );
nor U5625 ( n2645, n4357, n2648 );
nor U5626 ( n2656, n4357, n2659 );
nor U5627 ( n2667, n4357, n2670 );
nor U5628 ( n2678, n4357, n2681 );
nor U5629 ( n2689, n4357, n2692 );
nor U5630 ( n2700, n4357, n2703 );
nor U5631 ( n2711, n4357, n2714 );
nor U5632 ( n2722, n4357, n2726 );
nor U5633 ( n1897, n4363, n1901 );
nor U5634 ( n1909, n4363, n1913 );
nor U5635 ( n1922, n4363, n1926 );
nor U5636 ( n1934, n4363, n1938 );
nor U5637 ( n1947, n4363, n1951 );
nor U5638 ( n1959, n4363, n1963 );
nor U5639 ( n1972, n4362, n1976 );
nor U5640 ( n1984, n4362, n1988 );
nor U5641 ( n1997, n4362, n2001 );
nor U5642 ( n2009, n4362, n2013 );
nor U5643 ( n2022, n4362, n2026 );
nor U5644 ( n2034, n4362, n2038 );
nor U5645 ( n2047, n4362, n2051 );
nor U5646 ( n2059, n4362, n2063 );
nor U5647 ( n2072, n4362, n2076 );
nor U5648 ( n2084, n4362, n2088 );
nor U5649 ( n2098, n4362, n2102 );
nor U5650 ( n2112, n4362, n2116 );
nor U5651 ( n2126, n4361, n2129 );
nor U5652 ( n2139, n4361, n2143 );
nor U5653 ( n2153, n4361, n2157 );
nor U5654 ( n2167, n4361, n2171 );
nor U5655 ( n2181, n4361, n2184 );
nor U5656 ( n2194, n4361, n2198 );
nor U5657 ( n2208, n4361, n2212 );
nor U5658 ( n2222, n4361, n2226 );
nor U5659 ( n2236, n4361, n2239 );
nor U5660 ( n2249, n4361, n2253 );
nor U5661 ( n2263, n4361, n2267 );
nor U5662 ( n2277, n4361, n2281 );
nor U5663 ( n2291, n4359, n2294 );
nor U5664 ( n1465, n4367, n1469 );
nor U5665 ( n1478, n4366, n1481 );
nor U5666 ( n1490, n4366, n1494 );
nor U5667 ( n1503, n4366, n1506 );
nor U5668 ( n1515, n4366, n1519 );
nor U5669 ( n1529, n4366, n1533 );
nor U5670 ( n1542, n4366, n1546 );
nor U5671 ( n1555, n4366, n1559 );
nor U5672 ( n1569, n4366, n1573 );
nor U5673 ( n1582, n4366, n1586 );
nor U5674 ( n1595, n4366, n1599 );
nor U5675 ( n1609, n4366, n1613 );
nor U5676 ( n1622, n4366, n1626 );
nor U5677 ( n1635, n4365, n1639 );
nor U5678 ( n1646, n4365, n1649 );
nor U5679 ( n1656, n4365, n1659 );
nor U5680 ( n1667, n4365, n1670 );
nor U5681 ( n1678, n4365, n1681 );
nor U5682 ( n1689, n4365, n1692 );
nor U5683 ( n1700, n4365, n1703 );
nor U5684 ( n1711, n4365, n1714 );
nor U5685 ( n1722, n4365, n1725 );
nor U5686 ( n1733, n4365, n1736 );
nor U5687 ( n1744, n4365, n1747 );
nor U5688 ( n1755, n4365, n1758 );
nor U5689 ( n1766, n4363, n1769 );
nor U5690 ( n1777, n4363, n1780 );
nor U5691 ( n1788, n4363, n1791 );
nor U5692 ( n1801, n4363, n1804 );
nor U5693 ( n1814, n4363, n1818 );
nor U5694 ( n1828, n4363, n1832 );
nor U5695 ( n1103, n4369, n1106 );
nor U5696 ( n1115, n4369, n1119 );
nor U5697 ( n1128, n4369, n1131 );
nor U5698 ( n1140, n4369, n1144 );
nor U5699 ( n1153, n4369, n1156 );
nor U5700 ( n1165, n4369, n1169 );
nor U5701 ( n1178, n4369, n1181 );
nor U5702 ( n1190, n4369, n1194 );
nor U5703 ( n1204, n4369, n1208 );
nor U5704 ( n1218, n4369, n1221 );
nor U5705 ( n1231, n4369, n1235 );
nor U5706 ( n1245, n4369, n1249 );
nor U5707 ( n1259, n4367, n1263 );
nor U5708 ( n1273, n4367, n1276 );
nor U5709 ( n1286, n4367, n1290 );
nor U5710 ( n1300, n4367, n1304 );
nor U5711 ( n1314, n4367, n1318 );
nor U5712 ( n1328, n4367, n1331 );
nor U5713 ( n1341, n4367, n1345 );
nor U5714 ( n1355, n4367, n1359 );
nor U5715 ( n1369, n4367, n1373 );
nor U5716 ( n1383, n4367, n1386 );
nor U5717 ( n1396, n4367, n1400 );
nand U5718 ( n1845, n3988, n3989 );
nor U5719 ( n3989, n3990, n3992 );
nor U5720 ( n3988, n3997, n3998 );
nor U5721 ( n3990, n3537, n4334 );
nand U5722 ( n1840, n4004, n4005 );
nor U5723 ( n4005, n4007, n4008 );
nor U5724 ( n4004, n4013, n4014 );
nor U5725 ( n4007, n3548, n4331 );
nand U5726 ( n1835, n4020, n4022 );
nor U5727 ( n4022, n4023, n4024 );
nor U5728 ( n4020, n4029, n4030 );
nor U5729 ( n4023, n3559, n4333 );
nand U5730 ( n1830, n4037, n4038 );
nor U5731 ( n4038, n4039, n4040 );
nor U5732 ( n4037, n4045, n4047 );
nor U5733 ( n4039, n3570, n4323 );
nor U5734 ( n655, n4374, n660 );
nor U5735 ( n644, n4374, n649 );
nor U5736 ( n633, n4374, n638 );
nor U5737 ( n622, n4374, n627 );
nor U5738 ( n601, n4374, n606 );
nor U5739 ( n576, n4374, n581 );
nor U5740 ( n554, n4374, n559 );
nor U5741 ( n543, n4374, n548 );
nor U5742 ( n532, n4374, n537 );
nor U5743 ( n521, n4375, n526 );
nor U5744 ( n510, n4375, n515 );
nor U5745 ( n499, n4375, n504 );
nor U5746 ( n488, n4375, n493 );
nor U5747 ( n477, n4375, n482 );
nor U5748 ( n466, n4375, n471 );
nor U5749 ( n455, n4375, n460 );
nor U5750 ( n444, n4375, n449 );
nor U5751 ( n433, n4375, n438 );
nor U5752 ( n422, n4375, n427 );
nor U5753 ( n411, n4375, n416 );
nor U5754 ( n400, n4375, n405 );
nor U5755 ( n1003, n4370, n1006 );
nor U5756 ( n1015, n4370, n1019 );
nor U5757 ( n1028, n4370, n1031 );
nor U5758 ( n1040, n4370, n1044 );
nor U5759 ( n1053, n4370, n1056 );
nor U5760 ( n1065, n4370, n1069 );
nor U5761 ( n1078, n4370, n1081 );
nor U5762 ( n1090, n4370, n1094 );
nor U5763 ( n681, n4374, n684 );
nor U5764 ( n689, n4374, n692 );
nor U5765 ( n697, n4374, n700 );
nor U5766 ( n705, n4373, n708 );
nor U5767 ( n713, n4373, n716 );
nor U5768 ( n721, n4373, n724 );
nor U5769 ( n729, n4373, n732 );
nor U5770 ( n738, n4373, n741 );
nor U5771 ( n746, n4373, n749 );
nor U5772 ( n754, n4373, n757 );
nor U5773 ( n762, n4373, n765 );
nor U5774 ( n770, n4373, n773 );
nor U5775 ( n778, n4373, n781 );
nor U5776 ( n786, n4373, n789 );
nor U5777 ( n794, n4373, n797 );
nor U5778 ( n802, n4371, n805 );
nor U5779 ( n810, n4371, n813 );
nor U5780 ( n819, n4371, n822 );
nor U5781 ( n827, n4371, n830 );
nor U5782 ( n835, n4371, n838 );
nor U5783 ( n843, n4371, n846 );
nor U5784 ( n851, n4371, n854 );
nor U5785 ( n859, n4371, n862 );
nor U5786 ( n868, n4371, n871 );
nor U5787 ( n878, n4371, n881 );
nor U5788 ( n888, n4371, n891 );
nor U5789 ( n898, n4371, n901 );
nor U5790 ( n908, n4370, n911 );
nor U5791 ( n918, n4370, n921 );
nor U5792 ( n928, n4370, n931 );
nor U5793 ( n938, n4370, n941 );
nor U5794 ( n389, n4377, n394 );
nor U5795 ( n378, n4377, n383 );
nor U5796 ( n367, n4377, n372 );
nor U5797 ( n354, n4377, n361 );
nor U5798 ( n518, n520, n4321 );
nor U5799 ( n507, n509, n4321 );
nor U5800 ( n496, n498, n4321 );
nor U5801 ( n485, n487, n4321 );
nor U5802 ( n474, n476, n4321 );
nor U5803 ( n463, n465, n4321 );
nor U5804 ( n452, n454, n4321 );
nor U5805 ( n441, n443, n4321 );
nor U5806 ( n430, n432, n4321 );
nor U5807 ( n419, n421, n4321 );
nor U5808 ( n408, n410, n4321 );
nor U5809 ( n397, n399, n4321 );
nor U5810 ( n386, n388, n4322 );
nor U5811 ( n375, n377, n4322 );
nor U5812 ( n364, n366, n4322 );
nor U5813 ( n350, n353, n4322 );
nor U5814 ( n1023, n699, n4322 );
nor U5815 ( n1035, n707, n4322 );
nor U5816 ( n1048, n715, n4322 );
nor U5817 ( n1060, n723, n4322 );
nor U5818 ( n1073, n731, n4322 );
nor U5819 ( n1085, n740, n4322 );
nor U5820 ( n1098, n748, n4322 );
nor U5821 ( n1110, n756, n4322 );
nor U5822 ( n664, n665, n4325 );
nor U5823 ( n4138, n3636, n4333 );
nor U5824 ( n3630, n3201, n4333 );
nor U5825 ( n3194, n2739, n4330 );
nor U5826 ( n2731, n2307, n4326 );
nor U5827 ( n2299, n1844, n4326 );
nor U5828 ( n1837, n1413, n4325 );
nor U5829 ( n1405, n948, n4323 );
nor U5830 ( n4195, n3688, n4333 );
nor U5831 ( n4209, n3700, n4333 );
nor U5832 ( n4223, n3713, n4334 );
nor U5833 ( n4237, n3725, n4334 );
nor U5834 ( n4250, n3738, n4334 );
nor U5835 ( n4264, n3750, n4334 );
nor U5836 ( n652, n654, n4327 );
nor U5837 ( n641, n643, n4326 );
nor U5838 ( n630, n632, n4325 );
nor U5839 ( n619, n621, n4323 );
nor U5840 ( n598, n600, n4329 );
nor U5841 ( n573, n575, n4327 );
nor U5842 ( n551, n553, n4327 );
nor U5843 ( n540, n542, n4330 );
nor U5844 ( n529, n531, n4325 );
nor U5845 ( n3680, n3256, n4333 );
nor U5846 ( n3693, n3269, n4333 );
nor U5847 ( n3705, n3281, n4331 );
nor U5848 ( n3718, n3294, n4331 );
nor U5849 ( n3730, n3306, n4331 );
nor U5850 ( n3743, n3319, n4331 );
nor U5851 ( n3755, n3331, n4331 );
nor U5852 ( n3769, n3344, n4331 );
nor U5853 ( n3783, n3356, n4331 );
nor U5854 ( n3797, n3369, n4331 );
nor U5855 ( n3810, n3382, n4326 );
nor U5856 ( n3824, n3395, n4323 );
nor U5857 ( n3838, n3409, n4329 );
nor U5858 ( n3852, n3422, n4327 );
nor U5859 ( n3865, n3435, n4334 );
nor U5860 ( n3879, n3449, n4334 );
nor U5861 ( n3893, n3463, n4334 );
nor U5862 ( n3909, n3478, n4334 );
nor U5863 ( n3925, n3493, n4334 );
nor U5864 ( n3942, n3504, n4334 );
nor U5865 ( n3958, n3515, n4334 );
nor U5866 ( n3974, n3526, n4334 );
nor U5867 ( n4055, n3581, n4333 );
nor U5868 ( n4072, n3592, n4333 );
nor U5869 ( n4088, n3603, n4333 );
nor U5870 ( n4104, n3614, n4333 );
nor U5871 ( n4120, n3625, n4333 );
nor U5872 ( n3249, n2794, n4330 );
nor U5873 ( n3261, n2806, n4330 );
nor U5874 ( n3274, n2819, n4330 );
nor U5875 ( n3286, n2831, n4330 );
nor U5876 ( n3299, n2844, n4330 );
nor U5877 ( n3311, n2856, n4330 );
nor U5878 ( n3324, n2869, n4331 );
nor U5879 ( n3336, n2881, n4331 );
nor U5880 ( n3349, n2894, n4331 );
nor U5881 ( n3361, n2906, n4331 );
nor U5882 ( n3374, n2919, n4329 );
nor U5883 ( n3387, n2931, n4329 );
nor U5884 ( n3401, n2944, n4329 );
nor U5885 ( n3414, n2956, n4329 );
nor U5886 ( n3427, n2969, n4329 );
nor U5887 ( n3441, n2981, n4329 );
nor U5888 ( n3454, n2995, n4329 );
nor U5889 ( n3469, n3009, n4329 );
nor U5890 ( n3483, n3022, n4330 );
nor U5891 ( n3497, n3036, n4330 );
nor U5892 ( n3508, n3050, n4330 );
nor U5893 ( n3519, n3064, n4330 );
nor U5894 ( n3530, n3077, n4331 );
nor U5895 ( n3541, n3091, n4327 );
nor U5896 ( n3552, n3105, n4326 );
nor U5897 ( n3563, n3119, n4325 );
nor U5898 ( n3574, n3132, n4333 );
nor U5899 ( n3585, n3146, n4333 );
nor U5900 ( n3596, n3160, n4330 );
nor U5901 ( n3607, n3174, n4334 );
nor U5902 ( n3618, n3187, n4333 );
nor U5903 ( n2786, n2362, n4326 );
nor U5904 ( n2799, n2374, n4326 );
nor U5905 ( n2811, n2387, n4330 );
nor U5906 ( n2824, n2399, n4326 );
nor U5907 ( n2836, n2412, n4325 );
nor U5908 ( n2849, n2424, n4329 );
nor U5909 ( n2861, n2437, n4327 );
nor U5910 ( n2874, n2450, n4327 );
nor U5911 ( n2886, n2463, n4327 );
nor U5912 ( n2899, n2477, n4327 );
nor U5913 ( n2911, n2490, n4327 );
nor U5914 ( n2924, n2503, n4327 );
nor U5915 ( n2936, n2517, n4327 );
nor U5916 ( n2949, n2530, n4327 );
nor U5917 ( n2961, n2543, n4329 );
nor U5918 ( n2974, n2557, n4329 );
nor U5919 ( n2986, n2570, n4329 );
nor U5920 ( n3000, n2581, n4329 );
nor U5921 ( n3014, n2592, n4334 );
nor U5922 ( n3027, n2603, n4329 );
nor U5923 ( n3041, n2614, n4327 );
nor U5924 ( n3055, n2625, n4330 );
nor U5925 ( n3069, n2636, n4334 );
nor U5926 ( n3082, n2647, n4331 );
nor U5927 ( n3096, n2658, n4323 );
nor U5928 ( n3110, n2669, n4330 );
nor U5929 ( n3124, n2680, n4327 );
nor U5930 ( n3137, n2691, n4327 );
nor U5931 ( n3151, n2702, n4327 );
nor U5932 ( n3165, n2713, n4327 );
nor U5933 ( n3179, n2725, n4330 );
nor U5934 ( n2354, n1899, n4326 );
nor U5935 ( n2367, n1912, n4326 );
nor U5936 ( n2379, n1924, n4327 );
nor U5937 ( n2392, n1937, n4334 );
nor U5938 ( n2404, n1949, n4329 );
nor U5939 ( n2417, n1962, n4327 );
nor U5940 ( n2429, n1974, n4326 );
nor U5941 ( n2442, n1987, n4325 );
nor U5942 ( n2455, n1999, n4330 );
nor U5943 ( n2469, n2012, n4334 );
nor U5944 ( n2482, n2024, n4325 );
nor U5945 ( n2495, n2037, n4323 );
nor U5946 ( n2509, n2049, n4333 );
nor U5947 ( n2522, n2062, n4329 );
nor U5948 ( n2535, n2074, n4334 );
nor U5949 ( n2549, n2087, n4331 );
nor U5950 ( n2562, n2101, n4329 );
nor U5951 ( n2574, n2114, n4327 );
nor U5952 ( n2585, n2128, n4323 );
nor U5953 ( n2596, n2142, n4333 );
nor U5954 ( n2607, n2156, n4330 );
nor U5955 ( n2618, n2169, n4326 );
nor U5956 ( n2629, n2183, n4333 );
nor U5957 ( n2640, n2197, n4326 );
nor U5958 ( n2651, n2211, n4325 );
nor U5959 ( n2662, n2224, n4331 );
nor U5960 ( n2673, n2238, n4326 );
nor U5961 ( n2684, n2252, n4326 );
nor U5962 ( n2695, n2266, n4326 );
nor U5963 ( n2706, n2279, n4326 );
nor U5964 ( n2717, n2293, n4326 );
nor U5965 ( n1892, n1468, n4325 );
nor U5966 ( n1904, n1480, n4325 );
nor U5967 ( n1917, n1493, n4325 );
nor U5968 ( n1929, n1505, n4325 );
nor U5969 ( n1942, n1518, n4325 );
nor U5970 ( n1954, n1531, n4325 );
nor U5971 ( n1967, n1545, n4331 );
nor U5972 ( n1979, n1558, n4323 );
nor U5973 ( n1992, n1571, n4333 );
nor U5974 ( n2004, n1585, n4329 );
nor U5975 ( n2017, n1598, n4326 );
nor U5976 ( n2029, n1611, n4326 );
nor U5977 ( n2042, n1625, n4325 );
nor U5978 ( n2054, n1638, n4323 );
nor U5979 ( n2067, n1648, n4326 );
nor U5980 ( n2079, n1658, n4334 );
nor U5981 ( n2092, n1669, n4334 );
nor U5982 ( n2106, n1680, n4331 );
nor U5983 ( n2119, n1691, n4325 );
nor U5984 ( n2133, n1702, n4325 );
nor U5985 ( n2147, n1713, n4325 );
nor U5986 ( n2161, n1724, n4325 );
nor U5987 ( n2174, n1735, n4327 );
nor U5988 ( n2188, n1746, n4329 );
nor U5989 ( n2202, n1757, n4327 );
nor U5990 ( n2216, n1768, n4326 );
nor U5991 ( n2229, n1779, n4325 );
nor U5992 ( n2243, n1790, n4330 );
nor U5993 ( n2257, n1803, n4334 );
nor U5994 ( n2271, n1817, n4331 );
nor U5995 ( n2284, n1831, n4326 );
nor U5996 ( n1460, n1005, n4333 );
nor U5997 ( n1473, n1018, n4330 );
nor U5998 ( n1485, n1030, n4331 );
nor U5999 ( n1498, n1043, n4330 );
nor U6000 ( n1510, n1055, n4326 );
nor U6001 ( n1523, n1068, n4325 );
nor U6002 ( n1537, n1080, n4323 );
nor U6003 ( n1550, n1093, n4323 );
nor U6004 ( n1563, n1105, n4323 );
nor U6005 ( n1577, n1118, n4323 );
nor U6006 ( n1590, n1130, n4323 );
nor U6007 ( n1603, n1143, n4323 );
nor U6008 ( n1617, n1155, n4323 );
nor U6009 ( n1630, n1168, n4323 );
nor U6010 ( n1642, n1180, n4334 );
nor U6011 ( n1652, n1193, n4333 );
nor U6012 ( n1662, n1206, n4325 );
nor U6013 ( n1673, n1220, n4330 );
nor U6014 ( n1684, n1234, n4333 );
nor U6015 ( n1695, n1248, n4323 );
nor U6016 ( n1706, n1261, n4333 );
nor U6017 ( n1717, n1275, n4329 );
nor U6018 ( n1728, n1289, n4329 );
nor U6019 ( n1739, n1303, n4327 );
nor U6020 ( n1750, n1316, n4333 );
nor U6021 ( n1761, n1330, n4325 );
nor U6022 ( n1772, n1344, n4323 );
nor U6023 ( n1783, n1358, n4323 );
nor U6024 ( n1794, n1371, n4323 );
nor U6025 ( n1808, n1385, n4323 );
nor U6026 ( n1822, n1399, n4325 );
nor U6027 ( n998, n683, n4321 );
nor U6028 ( n1010, n691, n4322 );
nor U6029 ( n1123, n764, n4334 );
nor U6030 ( n1135, n772, n4331 );
nor U6031 ( n1148, n780, n4330 );
nor U6032 ( n1160, n788, n4331 );
nor U6033 ( n1173, n796, n4334 );
nor U6034 ( n1185, n804, n4331 );
nor U6035 ( n1198, n812, n4331 );
nor U6036 ( n1211, n821, n4323 );
nor U6037 ( n1225, n829, n4326 );
nor U6038 ( n1239, n837, n4333 );
nor U6039 ( n1253, n845, n4329 );
nor U6040 ( n1266, n853, n4327 );
nor U6041 ( n1280, n861, n4329 );
nor U6042 ( n1294, n870, n4330 );
nor U6043 ( n1308, n880, n4323 );
nor U6044 ( n1321, n890, n4323 );
nor U6045 ( n1335, n900, n4321 );
nor U6046 ( n1349, n910, n4322 );
nor U6047 ( n1363, n920, n4321 );
nor U6048 ( n1376, n930, n4322 );
nor U6049 ( n1390, n940, n4321 );
nor U6050 ( n352, n4267, n4471 );
nor U6051 ( n3687, n3688, n4413 );
nor U6052 ( n3699, n3700, n4413 );
nor U6053 ( n3712, n3713, n4413 );
nor U6054 ( n3724, n3725, n4413 );
nor U6055 ( n3737, n3738, n4413 );
nor U6056 ( n3749, n3750, n4413 );
nor U6057 ( n3762, n353, n4413 );
nor U6058 ( n3775, n366, n4413 );
nor U6059 ( n3789, n377, n4413 );
nor U6060 ( n3803, n388, n4413 );
nor U6061 ( n3817, n399, n4413 );
nor U6062 ( n3830, n410, n4413 );
nor U6063 ( n3844, n421, n4411 );
nor U6064 ( n3858, n432, n4411 );
nor U6065 ( n3872, n443, n4411 );
nor U6066 ( n3885, n454, n4411 );
nor U6067 ( n3900, n465, n4411 );
nor U6068 ( n3917, n476, n4411 );
nor U6069 ( n3933, n487, n4411 );
nor U6070 ( n3949, n498, n4411 );
nor U6071 ( n3965, n509, n4411 );
nor U6072 ( n3982, n520, n4411 );
nor U6073 ( n3998, n531, n4411 );
nor U6074 ( n4014, n542, n4411 );
nor U6075 ( n4030, n553, n4410 );
nor U6076 ( n4047, n575, n4410 );
nor U6077 ( n4063, n600, n4410 );
nor U6078 ( n4079, n621, n4410 );
nor U6079 ( n4095, n632, n4410 );
nor U6080 ( n4112, n643, n4410 );
nor U6081 ( n4128, n654, n4410 );
nor U6082 ( n3255, n3256, n4417 );
nor U6083 ( n3267, n3269, n4417 );
nor U6084 ( n3280, n3281, n4417 );
nor U6085 ( n3292, n3294, n4417 );
nor U6086 ( n3305, n3306, n4417 );
nor U6087 ( n3317, n3319, n4417 );
nor U6088 ( n3330, n3331, n4417 );
nor U6089 ( n3342, n3344, n4417 );
nor U6090 ( n3355, n3356, n4415 );
nor U6091 ( n3367, n3369, n4415 );
nor U6092 ( n3381, n3382, n4415 );
nor U6093 ( n3394, n3395, n4415 );
nor U6094 ( n3407, n3409, n4415 );
nor U6095 ( n3421, n3422, n4415 );
nor U6096 ( n3434, n3435, n4415 );
nor U6097 ( n3447, n3449, n4415 );
nor U6098 ( n3462, n3463, n4415 );
nor U6099 ( n3477, n3478, n4415 );
nor U6100 ( n3491, n3493, n4415 );
nor U6101 ( n3503, n3504, n4415 );
nor U6102 ( n3514, n3515, n4414 );
nor U6103 ( n3525, n3526, n4414 );
nor U6104 ( n3536, n3537, n4414 );
nor U6105 ( n3547, n3548, n4414 );
nor U6106 ( n3558, n3559, n4414 );
nor U6107 ( n3569, n3570, n4414 );
nor U6108 ( n3580, n3581, n4414 );
nor U6109 ( n3591, n3592, n4414 );
nor U6110 ( n3602, n3603, n4414 );
nor U6111 ( n3613, n3614, n4414 );
nor U6112 ( n3624, n3625, n4414 );
nor U6113 ( n3172, n3174, n4417 );
nor U6114 ( n3186, n3187, n4417 );
nor U6115 ( n1898, n1899, n4395 );
nor U6116 ( n1911, n1912, n4395 );
nor U6117 ( n1923, n1924, n4395 );
nor U6118 ( n1936, n1937, n4395 );
nor U6119 ( n1948, n1949, n4395 );
nor U6120 ( n1961, n1962, n4395 );
nor U6121 ( n1973, n1974, n4395 );
nor U6122 ( n1986, n1987, n4395 );
nor U6123 ( n1998, n1999, n4395 );
nor U6124 ( n2011, n2012, n4395 );
nor U6125 ( n2023, n2024, n4394 );
nor U6126 ( n2036, n2037, n4394 );
nor U6127 ( n2048, n2049, n4394 );
nor U6128 ( n2061, n2062, n4394 );
nor U6129 ( n2073, n2074, n4394 );
nor U6130 ( n2086, n2087, n4394 );
nor U6131 ( n2099, n2101, n4394 );
nor U6132 ( n2113, n2114, n4394 );
nor U6133 ( n2127, n2128, n4394 );
nor U6134 ( n2141, n2142, n4394 );
nor U6135 ( n2154, n2156, n4394 );
nor U6136 ( n2168, n2169, n4401 );
nor U6137 ( n1466, n1468, n4399 );
nor U6138 ( n1479, n1480, n4399 );
nor U6139 ( n1491, n1493, n4399 );
nor U6140 ( n1504, n1505, n4399 );
nor U6141 ( n1517, n1518, n4399 );
nor U6142 ( n1530, n1531, n4399 );
nor U6143 ( n1543, n1545, n4398 );
nor U6144 ( n1557, n1558, n4398 );
nor U6145 ( n1570, n1571, n4398 );
nor U6146 ( n1583, n1585, n4398 );
nor U6147 ( n1597, n1598, n4398 );
nor U6148 ( n1610, n1611, n4398 );
nor U6149 ( n1623, n1625, n4398 );
nor U6150 ( n1637, n1638, n4398 );
nor U6151 ( n1647, n1648, n4398 );
nor U6152 ( n1657, n1658, n4398 );
nor U6153 ( n1668, n1669, n4398 );
nor U6154 ( n1679, n1680, n4398 );
nor U6155 ( n1690, n1691, n4397 );
nor U6156 ( n1701, n1702, n4397 );
nor U6157 ( n1712, n1713, n4397 );
nor U6158 ( n1723, n1724, n4397 );
nor U6159 ( n1734, n1735, n4397 );
nor U6160 ( n1745, n1746, n4397 );
nor U6161 ( n1756, n1757, n4397 );
nor U6162 ( n1767, n1768, n4397 );
nor U6163 ( n1778, n1779, n4397 );
nor U6164 ( n1789, n1790, n4397 );
nor U6165 ( n1802, n1803, n4397 );
nor U6166 ( n1816, n1817, n4397 );
nor U6167 ( n1829, n1831, n4395 );
nor U6168 ( n1004, n1005, n4403 );
nor U6169 ( n1016, n1018, n4403 );
nor U6170 ( n1029, n1030, n4403 );
nor U6171 ( n1041, n1043, n4402 );
nor U6172 ( n1054, n1055, n4402 );
nor U6173 ( n1066, n1068, n4402 );
nor U6174 ( n1079, n1080, n4402 );
nor U6175 ( n1091, n1093, n4402 );
nor U6176 ( n1104, n1105, n4402 );
nor U6177 ( n1116, n1118, n4402 );
nor U6178 ( n1129, n1130, n4402 );
nor U6179 ( n1141, n1143, n4402 );
nor U6180 ( n1154, n1155, n4402 );
nor U6181 ( n1166, n1168, n4402 );
nor U6182 ( n1179, n1180, n4402 );
nor U6183 ( n1191, n1193, n4401 );
nor U6184 ( n1205, n1206, n4401 );
nor U6185 ( n1219, n1220, n4401 );
nor U6186 ( n1233, n1234, n4401 );
nor U6187 ( n1246, n1248, n4401 );
nor U6188 ( n1260, n1261, n4401 );
nor U6189 ( n1274, n1275, n4401 );
nor U6190 ( n1288, n1289, n4401 );
nor U6191 ( n1301, n1303, n4401 );
nor U6192 ( n1315, n1316, n4401 );
nor U6193 ( n1329, n1330, n4401 );
nor U6194 ( n1343, n1344, n4399 );
nor U6195 ( n1356, n1358, n4399 );
nor U6196 ( n1370, n1371, n4399 );
nor U6197 ( n1384, n1385, n4399 );
nor U6198 ( n1398, n1399, n4399 );
nor U6199 ( n682, n683, n4406 );
nor U6200 ( n690, n691, n4406 );
nor U6201 ( n698, n699, n4406 );
nor U6202 ( n706, n707, n4406 );
nor U6203 ( n714, n715, n4406 );
nor U6204 ( n722, n723, n4406 );
nor U6205 ( n730, n731, n4406 );
nor U6206 ( n739, n740, n4406 );
nor U6207 ( n747, n748, n4406 );
nor U6208 ( n755, n756, n4406 );
nor U6209 ( n763, n764, n4405 );
nor U6210 ( n771, n772, n4405 );
nor U6211 ( n779, n780, n4405 );
nor U6212 ( n787, n788, n4405 );
nor U6213 ( n795, n796, n4405 );
nor U6214 ( n803, n804, n4405 );
nor U6215 ( n811, n812, n4405 );
nor U6216 ( n820, n821, n4405 );
nor U6217 ( n828, n829, n4405 );
nor U6218 ( n836, n837, n4405 );
nor U6219 ( n844, n845, n4405 );
nor U6220 ( n852, n853, n4405 );
nor U6221 ( n860, n861, n4403 );
nor U6222 ( n869, n870, n4403 );
nor U6223 ( n879, n880, n4403 );
nor U6224 ( n889, n890, n4403 );
nor U6225 ( n899, n900, n4403 );
nor U6226 ( n909, n910, n4403 );
nor U6227 ( n919, n920, n4403 );
nor U6228 ( n929, n930, n4403 );
nor U6229 ( n939, n940, n4403 );
nor U6230 ( n4202, n285, n4410 );
nor U6231 ( n4215, n287, n4410 );
nor U6232 ( n4229, n289, n4410 );
nor U6233 ( n4243, n291, n4410 );
nor U6234 ( n4257, n293, n4417 );
nor U6235 ( n4272, n295, n4394 );
nor U6236 ( n656, n345, n4406 );
nor U6237 ( n645, n343, n4407 );
nor U6238 ( n634, n341, n4407 );
nor U6239 ( n623, n339, n4407 );
nor U6240 ( n602, n337, n4407 );
nor U6241 ( n577, n335, n4407 );
nor U6242 ( n555, n333, n4407 );
nor U6243 ( n544, n331, n4407 );
nor U6244 ( n533, n329, n4407 );
nor U6245 ( n522, n327, n4407 );
nor U6246 ( n511, n325, n4407 );
nor U6247 ( n500, n323, n4407 );
nor U6248 ( n489, n321, n4407 );
nor U6249 ( n478, n319, n4409 );
nor U6250 ( n467, n317, n4409 );
nor U6251 ( n456, n315, n4409 );
nor U6252 ( n445, n313, n4409 );
nor U6253 ( n434, n311, n4409 );
nor U6254 ( n423, n309, n4409 );
nor U6255 ( n412, n307, n4409 );
nor U6256 ( n401, n305, n4409 );
nor U6257 ( n390, n303, n4409 );
nor U6258 ( n379, n301, n4409 );
nor U6259 ( n368, n299, n4409 );
nor U6260 ( n355, n297, n4409 );
nor U6261 ( n2792, n2794, n4421 );
nor U6262 ( n2805, n2806, n4421 );
nor U6263 ( n2817, n2819, n4421 );
nor U6264 ( n2830, n2831, n4421 );
nor U6265 ( n2842, n2844, n4421 );
nor U6266 ( n2855, n2856, n4419 );
nor U6267 ( n2867, n2869, n4419 );
nor U6268 ( n2880, n2881, n4419 );
nor U6269 ( n2892, n2894, n4419 );
nor U6270 ( n2905, n2906, n4419 );
nor U6271 ( n2917, n2919, n4419 );
nor U6272 ( n2930, n2931, n4419 );
nor U6273 ( n2942, n2944, n4419 );
nor U6274 ( n2955, n2956, n4419 );
nor U6275 ( n2967, n2969, n4419 );
nor U6276 ( n2980, n2981, n4419 );
nor U6277 ( n2994, n2995, n4419 );
nor U6278 ( n3007, n3009, n4418 );
nor U6279 ( n3021, n3022, n4418 );
nor U6280 ( n3035, n3036, n4418 );
nor U6281 ( n3049, n3050, n4418 );
nor U6282 ( n3062, n3064, n4418 );
nor U6283 ( n3076, n3077, n4418 );
nor U6284 ( n3090, n3091, n4418 );
nor U6285 ( n3104, n3105, n4418 );
nor U6286 ( n3117, n3119, n4418 );
nor U6287 ( n3131, n3132, n4418 );
nor U6288 ( n3145, n3146, n4418 );
nor U6289 ( n3159, n3160, n4418 );
nor U6290 ( n2373, n2374, n4423 );
nor U6291 ( n2386, n2387, n4423 );
nor U6292 ( n2398, n2399, n4423 );
nor U6293 ( n2411, n2412, n4423 );
nor U6294 ( n2423, n2424, n4423 );
nor U6295 ( n2436, n2437, n4423 );
nor U6296 ( n2449, n2450, n4423 );
nor U6297 ( n2462, n2463, n4423 );
nor U6298 ( n2475, n2477, n4423 );
nor U6299 ( n2489, n2490, n4423 );
nor U6300 ( n2502, n2503, n4423 );
nor U6301 ( n2515, n2517, n4423 );
nor U6302 ( n2529, n2530, n4422 );
nor U6303 ( n2542, n2543, n4422 );
nor U6304 ( n2555, n2557, n4422 );
nor U6305 ( n2569, n2570, n4422 );
nor U6306 ( n2580, n2581, n4422 );
nor U6307 ( n2591, n2592, n4422 );
nor U6308 ( n2602, n2603, n4422 );
nor U6309 ( n2613, n2614, n4422 );
nor U6310 ( n2624, n2625, n4422 );
nor U6311 ( n2635, n2636, n4422 );
nor U6312 ( n2646, n2647, n4422 );
nor U6313 ( n2657, n2658, n4422 );
nor U6314 ( n2668, n2669, n4421 );
nor U6315 ( n2679, n2680, n4421 );
nor U6316 ( n2690, n2691, n4421 );
nor U6317 ( n2701, n2702, n4421 );
nor U6318 ( n2712, n2713, n4421 );
nor U6319 ( n2724, n2725, n4421 );
nor U6320 ( n2361, n2362, n4424 );
nor U6321 ( n2182, n2183, n4424 );
nor U6322 ( n2196, n2197, n4424 );
nor U6323 ( n2209, n2211, n4424 );
nor U6324 ( n2223, n2224, n4424 );
nor U6325 ( n2237, n2238, n4424 );
nor U6326 ( n2251, n2252, n4424 );
nor U6327 ( n2264, n2266, n4424 );
nor U6328 ( n2278, n2279, n4424 );
nor U6329 ( n2292, n2293, n4424 );
not U6330 ( n5, n606 );
not U6331 ( n7, n559 );
not U6332 ( n8, n548 );
not U6333 ( n9, n537 );
not U6334 ( n10, n526 );
not U6335 ( n11, n515 );
not U6336 ( n17, n449 );
not U6337 ( n19, n427 );
not U6338 ( n21, n405 );
not U6339 ( n22, n394 );
not U6340 ( n29, n674 );
not U6341 ( n30, n673 );
not U6342 ( n31, n672 );
not U6343 ( n2, n649 );
not U6344 ( n14, n482 );
not U6345 ( n1, n660 );
not U6346 ( n3, n638 );
not U6347 ( n4, n627 );
not U6348 ( n6, n581 );
not U6349 ( n12, n504 );
not U6350 ( n13, n493 );
not U6351 ( n15, n471 );
not U6352 ( n16, n460 );
not U6353 ( n18, n438 );
not U6354 ( n23, n383 );
not U6355 ( n24, n372 );
not U6356 ( n25, n361 );
not U6357 ( n26, n814 );
not U6358 ( n249, n941 );
not U6359 ( n250, n931 );
not U6360 ( n251, n921 );
not U6361 ( n252, n911 );
not U6362 ( n253, n901 );
not U6363 ( n254, n891 );
not U6364 ( n255, n881 );
not U6365 ( n256, n871 );
not U6366 ( n257, n862 );
not U6367 ( n258, n854 );
not U6368 ( n259, n846 );
not U6369 ( n260, n838 );
not U6370 ( n261, n830 );
not U6371 ( n262, n822 );
not U6372 ( n263, n813 );
not U6373 ( n264, n805 );
not U6374 ( n265, n797 );
not U6375 ( n266, n789 );
not U6376 ( n267, n781 );
not U6377 ( n268, n773 );
not U6378 ( n269, n765 );
not U6379 ( n270, n757 );
not U6380 ( n271, n749 );
not U6381 ( n272, n741 );
not U6382 ( n273, n732 );
not U6383 ( n274, n724 );
not U6384 ( n275, n716 );
not U6385 ( n276, n708 );
not U6386 ( n277, n700 );
not U6387 ( n278, n692 );
not U6388 ( n279, n684 );
not U6389 ( n218, n1400 );
not U6390 ( n219, n1386 );
not U6391 ( n220, n1373 );
not U6392 ( n221, n1359 );
not U6393 ( n222, n1345 );
not U6394 ( n223, n1331 );
not U6395 ( n224, n1318 );
not U6396 ( n225, n1304 );
not U6397 ( n226, n1290 );
not U6398 ( n227, n1276 );
not U6399 ( n228, n1263 );
not U6400 ( n229, n1249 );
not U6401 ( n230, n1235 );
not U6402 ( n231, n1221 );
not U6403 ( n232, n1208 );
not U6404 ( n233, n1194 );
not U6405 ( n234, n1181 );
not U6406 ( n235, n1169 );
not U6407 ( n236, n1156 );
not U6408 ( n237, n1144 );
not U6409 ( n238, n1131 );
not U6410 ( n239, n1119 );
not U6411 ( n240, n1106 );
not U6412 ( n241, n1094 );
not U6413 ( n242, n1081 );
not U6414 ( n243, n1069 );
not U6415 ( n244, n1056 );
not U6416 ( n245, n1044 );
not U6417 ( n246, n1031 );
not U6418 ( n247, n1019 );
not U6419 ( n248, n1006 );
not U6420 ( n187, n1832 );
not U6421 ( n188, n1818 );
not U6422 ( n189, n1804 );
not U6423 ( n190, n1791 );
not U6424 ( n191, n1780 );
not U6425 ( n192, n1769 );
not U6426 ( n193, n1758 );
not U6427 ( n194, n1747 );
not U6428 ( n195, n1736 );
not U6429 ( n196, n1725 );
not U6430 ( n197, n1714 );
not U6431 ( n198, n1703 );
not U6432 ( n199, n1692 );
not U6433 ( n200, n1681 );
not U6434 ( n201, n1670 );
not U6435 ( n202, n1659 );
not U6436 ( n203, n1649 );
not U6437 ( n204, n1639 );
not U6438 ( n205, n1626 );
not U6439 ( n206, n1613 );
not U6440 ( n207, n1599 );
not U6441 ( n208, n1586 );
not U6442 ( n209, n1573 );
not U6443 ( n210, n1559 );
not U6444 ( n211, n1546 );
not U6445 ( n212, n1533 );
not U6446 ( n213, n1519 );
not U6447 ( n214, n1506 );
not U6448 ( n215, n1494 );
not U6449 ( n216, n1481 );
not U6450 ( n217, n1469 );
not U6451 ( n156, n2294 );
not U6452 ( n157, n2281 );
not U6453 ( n158, n2267 );
not U6454 ( n159, n2253 );
not U6455 ( n160, n2239 );
not U6456 ( n161, n2226 );
not U6457 ( n162, n2212 );
not U6458 ( n163, n2198 );
not U6459 ( n164, n2184 );
not U6460 ( n165, n2171 );
not U6461 ( n166, n2157 );
not U6462 ( n167, n2143 );
not U6463 ( n168, n2129 );
not U6464 ( n169, n2116 );
not U6465 ( n170, n2102 );
not U6466 ( n171, n2088 );
not U6467 ( n172, n2076 );
not U6468 ( n173, n2063 );
not U6469 ( n174, n2051 );
not U6470 ( n175, n2038 );
not U6471 ( n176, n2026 );
not U6472 ( n177, n2013 );
not U6473 ( n178, n2001 );
not U6474 ( n179, n1988 );
not U6475 ( n180, n1976 );
not U6476 ( n181, n1963 );
not U6477 ( n182, n1951 );
not U6478 ( n183, n1938 );
not U6479 ( n184, n1926 );
not U6480 ( n185, n1913 );
not U6481 ( n186, n1901 );
not U6482 ( n125, n2726 );
not U6483 ( n126, n2714 );
not U6484 ( n127, n2703 );
not U6485 ( n128, n2692 );
not U6486 ( n129, n2681 );
not U6487 ( n130, n2670 );
not U6488 ( n131, n2659 );
not U6489 ( n132, n2648 );
not U6490 ( n133, n2637 );
not U6491 ( n134, n2626 );
not U6492 ( n135, n2615 );
not U6493 ( n136, n2604 );
not U6494 ( n137, n2593 );
not U6495 ( n138, n2582 );
not U6496 ( n139, n2571 );
not U6497 ( n140, n2558 );
not U6498 ( n141, n2545 );
not U6499 ( n142, n2531 );
not U6500 ( n143, n2518 );
not U6501 ( n144, n2505 );
not U6502 ( n145, n2491 );
not U6503 ( n146, n2478 );
not U6504 ( n147, n2465 );
not U6505 ( n148, n2451 );
not U6506 ( n149, n2438 );
not U6507 ( n150, n2426 );
not U6508 ( n151, n2413 );
not U6509 ( n152, n2401 );
not U6510 ( n153, n2388 );
not U6511 ( n154, n2376 );
not U6512 ( n155, n2363 );
not U6513 ( n94, n3189 );
not U6514 ( n95, n3175 );
not U6515 ( n96, n3161 );
not U6516 ( n97, n3147 );
not U6517 ( n98, n3134 );
not U6518 ( n99, n3120 );
not U6519 ( n100, n3106 );
not U6520 ( n101, n3092 );
not U6521 ( n102, n3079 );
not U6522 ( n103, n3065 );
not U6523 ( n104, n3051 );
not U6524 ( n105, n3037 );
not U6525 ( n106, n3024 );
not U6526 ( n107, n3010 );
not U6527 ( n108, n2996 );
not U6528 ( n109, n2982 );
not U6529 ( n110, n2970 );
not U6530 ( n111, n2957 );
not U6531 ( n112, n2945 );
not U6532 ( n113, n2932 );
not U6533 ( n114, n2920 );
not U6534 ( n115, n2907 );
not U6535 ( n116, n2895 );
not U6536 ( n117, n2882 );
not U6537 ( n118, n2870 );
not U6538 ( n119, n2857 );
not U6539 ( n120, n2845 );
not U6540 ( n121, n2832 );
not U6541 ( n122, n2820 );
not U6542 ( n123, n2807 );
not U6543 ( n124, n2795 );
not U6544 ( n63, n3626 );
not U6545 ( n64, n3615 );
not U6546 ( n65, n3604 );
not U6547 ( n66, n3593 );
not U6548 ( n67, n3582 );
not U6549 ( n68, n3571 );
not U6550 ( n69, n3560 );
not U6551 ( n70, n3549 );
not U6552 ( n71, n3538 );
not U6553 ( n72, n3527 );
not U6554 ( n73, n3516 );
not U6555 ( n74, n3505 );
not U6556 ( n75, n3494 );
not U6557 ( n76, n3479 );
not U6558 ( n77, n3465 );
not U6559 ( n78, n3450 );
not U6560 ( n79, n3437 );
not U6561 ( n80, n3423 );
not U6562 ( n81, n3410 );
not U6563 ( n82, n3397 );
not U6564 ( n83, n3383 );
not U6565 ( n84, n3370 );
not U6566 ( n85, n3357 );
not U6567 ( n86, n3345 );
not U6568 ( n87, n3332 );
not U6569 ( n88, n3320 );
not U6570 ( n89, n3307 );
not U6571 ( n90, n3295 );
not U6572 ( n91, n3282 );
not U6573 ( n92, n3270 );
not U6574 ( n93, n3257 );
not U6575 ( n32, n4133 );
not U6576 ( n33, n4117 );
not U6577 ( n34, n4100 );
not U6578 ( n35, n4084 );
not U6579 ( n36, n4068 );
not U6580 ( n37, n4052 );
not U6581 ( n38, n4035 );
not U6582 ( n39, n4019 );
not U6583 ( n40, n4003 );
not U6584 ( n41, n3987 );
not U6585 ( n42, n3970 );
not U6586 ( n43, n3954 );
not U6587 ( n44, n3938 );
not U6588 ( n45, n3922 );
not U6589 ( n46, n3905 );
not U6590 ( n47, n3889 );
not U6591 ( n48, n3875 );
not U6592 ( n49, n3862 );
not U6593 ( n50, n3848 );
not U6594 ( n51, n3834 );
not U6595 ( n52, n3820 );
not U6596 ( n53, n3807 );
not U6597 ( n54, n3793 );
not U6598 ( n55, n3779 );
not U6599 ( n56, n3765 );
not U6600 ( n57, n3752 );
not U6601 ( n58, n3739 );
not U6602 ( n59, n3727 );
not U6603 ( n60, n3714 );
not U6604 ( n61, n3702 );
not U6605 ( n62, n3689 );
not U6606 ( n20, n416 );
not U6607 ( n27, n733 );
not U6608 ( n28, n675 );
xor U6609 ( n345, n657, n658 );
xnor U6610 ( n657, WX711, n659 );
xor U6611 ( n658, WX647, TM1 );
xor U6612 ( n659, WX839, WX775 );
xor U6613 ( n343, n646, n647 );
xnor U6614 ( n646, WX713, n648 );
xor U6615 ( n647, WX649, TM1 );
xor U6616 ( n648, WX841, WX777 );
xor U6617 ( n341, n635, n636 );
xnor U6618 ( n635, WX715, n637 );
xor U6619 ( n636, WX651, TM1 );
xor U6620 ( n637, WX843, WX779 );
xor U6621 ( n347, n669, n670 );
xnor U6622 ( n669, WX709, n671 );
xor U6623 ( n670, WX645, TM1 );
xor U6624 ( n671, WX837, WX773 );
xor U6625 ( DATA_9_28, n4278, n341 );
nand U6626 ( n4278, TM0, WX491 );
xor U6627 ( DATA_9_29, n4279, n343 );
nand U6628 ( n4279, TM0, WX489 );
xor U6629 ( DATA_9_30, n4280, n345 );
nand U6630 ( n4280, TM0, WX487 );
xor U6631 ( DATA_9_31, n4282, n347 );
nand U6632 ( n4282, TM0, WX485 );
xor U6633 ( n339, n624, n625 );
xnor U6634 ( n624, WX717, n626 );
xor U6635 ( n625, WX653, TM1 );
xor U6636 ( n626, WX845, WX781 );
xor U6637 ( n337, n603, n604 );
xnor U6638 ( n603, WX719, n605 );
xor U6639 ( n604, WX655, TM1 );
xor U6640 ( n605, WX847, WX783 );
xor U6641 ( n335, n578, n579 );
xnor U6642 ( n578, WX721, n580 );
xor U6643 ( n579, WX657, TM1 );
xor U6644 ( n580, WX849, WX785 );
xor U6645 ( n333, n556, n557 );
xnor U6646 ( n556, WX723, n558 );
xor U6647 ( n557, WX659, TM1 );
xor U6648 ( n558, WX851, WX787 );
xor U6649 ( n331, n545, n546 );
xnor U6650 ( n545, WX725, n547 );
xor U6651 ( n546, WX661, TM1 );
xor U6652 ( n547, WX853, WX789 );
xor U6653 ( n329, n534, n535 );
xnor U6654 ( n534, WX727, n536 );
xor U6655 ( n535, WX663, TM1 );
xor U6656 ( n536, WX855, WX791 );
xor U6657 ( n327, n523, n524 );
xnor U6658 ( n523, WX729, n525 );
xor U6659 ( n524, WX665, TM1 );
xor U6660 ( n525, WX857, WX793 );
xor U6661 ( n325, n512, n513 );
xnor U6662 ( n512, WX731, n514 );
xor U6663 ( n513, WX667, TM1 );
xor U6664 ( n514, WX859, WX795 );
xor U6665 ( n323, n501, n502 );
xnor U6666 ( n501, WX733, n503 );
xor U6667 ( n502, WX669, TM1 );
xor U6668 ( n503, WX861, WX797 );
xor U6669 ( n321, n490, n491 );
xnor U6670 ( n490, WX735, n492 );
xor U6671 ( n491, WX671, TM1 );
xor U6672 ( n492, WX863, WX799 );
xor U6673 ( n319, n479, n480 );
xnor U6674 ( n479, WX737, n481 );
xor U6675 ( n480, WX673, TM1 );
xor U6676 ( n481, WX865, WX801 );
xor U6677 ( n317, n468, n469 );
xnor U6678 ( n468, WX739, n470 );
xor U6679 ( n469, WX675, TM1 );
xor U6680 ( n470, WX867, WX803 );
xor U6681 ( DATA_9_16, n4283, n317 );
nand U6682 ( n4283, TM0, WX515 );
xor U6683 ( DATA_9_17, n4284, n319 );
nand U6684 ( n4284, TM0, WX513 );
xor U6685 ( DATA_9_18, n4285, n321 );
nand U6686 ( n4285, TM0, WX511 );
xor U6687 ( DATA_9_19, n4287, n323 );
nand U6688 ( n4287, TM0, WX509 );
xor U6689 ( DATA_9_20, n4288, n325 );
nand U6690 ( n4288, TM0, WX507 );
xor U6691 ( DATA_9_21, n4289, n327 );
nand U6692 ( n4289, TM0, WX505 );
xor U6693 ( DATA_9_22, n4290, n329 );
nand U6694 ( n4290, TM0, WX503 );
xor U6695 ( DATA_9_23, n4292, n331 );
nand U6696 ( n4292, TM0, WX501 );
xor U6697 ( DATA_9_24, n4293, n333 );
nand U6698 ( n4293, TM0, WX499 );
xor U6699 ( DATA_9_25, n4294, n335 );
nand U6700 ( n4294, TM0, WX497 );
xor U6701 ( DATA_9_26, n4295, n337 );
nand U6702 ( n4295, TM0, WX495 );
xor U6703 ( DATA_9_27, n4297, n339 );
nand U6704 ( n4297, TM0, WX493 );
and U6705 ( n663, WX485, n666 );
and U6706 ( n4137, n666, WX1778 );
and U6707 ( n3629, n666, WX3071 );
and U6708 ( n3192, n666, WX4364 );
and U6709 ( n2730, n666, WX5657 );
and U6710 ( n2298, n666, WX6950 );
and U6711 ( n1836, n666, WX8243 );
and U6712 ( n1404, n666, WX9536 );
nand U6713 ( n950, WX10829, n666 );
nand U6714 ( n1027, n4193, n4194 );
nor U6715 ( n4194, n4195, n4197 );
nor U6716 ( n4193, n4200, n4202 );
and U6717 ( n4197, n4448, CRC_OUT_9_0 );
nand U6718 ( n1022, n4207, n4208 );
nor U6719 ( n4208, n4209, n4210 );
nor U6720 ( n4207, n4214, n4215 );
and U6721 ( n4210, n4448, CRC_OUT_9_1 );
nand U6722 ( n1017, n4220, n4222 );
nor U6723 ( n4222, n4223, n4224 );
nor U6724 ( n4220, n4228, n4229 );
and U6725 ( n4224, n4448, CRC_OUT_9_2 );
nand U6726 ( n1012, n4234, n4235 );
nor U6727 ( n4235, n4237, n4238 );
nor U6728 ( n4234, n4242, n4243 );
and U6729 ( n4238, n4448, CRC_OUT_9_3 );
nand U6730 ( n1007, n4248, n4249 );
nor U6731 ( n4249, n4250, n4252 );
nor U6732 ( n4248, n4255, n4257 );
and U6733 ( n4252, n4453, CRC_OUT_9_4 );
nand U6734 ( n1002, n4262, n4263 );
nor U6735 ( n4263, n4264, n4265 );
nor U6736 ( n4262, n4270, n4272 );
and U6737 ( n4265, n4440, CRC_OUT_9_5 );
nand U6738 ( n1955, n3678, n3679 );
nor U6739 ( n3679, n3680, n3682 );
nor U6740 ( n3678, n3685, n3687 );
and U6741 ( n3682, n4451, CRC_OUT_8_0 );
nand U6742 ( n1950, n3690, n3692 );
nor U6743 ( n3692, n3693, n3694 );
nor U6744 ( n3690, n3698, n3699 );
and U6745 ( n3694, n4451, CRC_OUT_8_1 );
nand U6746 ( n1945, n3703, n3704 );
nor U6747 ( n3704, n3705, n3707 );
nor U6748 ( n3703, n3710, n3712 );
and U6749 ( n3707, n4450, CRC_OUT_8_2 );
nand U6750 ( n1940, n3715, n3717 );
nor U6751 ( n3717, n3718, n3719 );
nor U6752 ( n3715, n3723, n3724 );
and U6753 ( n3719, n4450, CRC_OUT_8_3 );
nand U6754 ( n1935, n3728, n3729 );
nor U6755 ( n3729, n3730, n3732 );
nor U6756 ( n3728, n3735, n3737 );
and U6757 ( n3732, n4450, CRC_OUT_8_4 );
nand U6758 ( n1930, n3740, n3742 );
nor U6759 ( n3742, n3743, n3744 );
nor U6760 ( n3740, n3748, n3749 );
and U6761 ( n3744, n4450, CRC_OUT_8_5 );
nand U6762 ( n1925, n3753, n3754 );
nor U6763 ( n3754, n3755, n3757 );
nor U6764 ( n3753, n3760, n3762 );
and U6765 ( n3757, n4450, CRC_OUT_8_6 );
nand U6766 ( n1920, n3767, n3768 );
nor U6767 ( n3768, n3769, n3770 );
nor U6768 ( n3767, n3774, n3775 );
and U6769 ( n3770, n4450, CRC_OUT_8_7 );
nand U6770 ( n1915, n3780, n3782 );
nor U6771 ( n3782, n3783, n3784 );
nor U6772 ( n3780, n3788, n3789 );
and U6773 ( n3784, n4450, CRC_OUT_8_8 );
nand U6774 ( n1910, n3794, n3795 );
nor U6775 ( n3795, n3797, n3798 );
nor U6776 ( n3794, n3802, n3803 );
and U6777 ( n3798, n4450, CRC_OUT_8_9 );
nand U6778 ( n1905, n3808, n3809 );
nor U6779 ( n3809, n3810, n3812 );
nor U6780 ( n3808, n3815, n3817 );
and U6781 ( n3812, n4450, CRC_OUT_8_10 );
nand U6782 ( n1900, n3822, n3823 );
nor U6783 ( n3823, n3824, n3825 );
nor U6784 ( n3822, n3829, n3830 );
and U6785 ( n3825, n4450, CRC_OUT_8_11 );
nand U6786 ( n1895, n3835, n3837 );
nor U6787 ( n3837, n3838, n3839 );
nor U6788 ( n3835, n3843, n3844 );
and U6789 ( n3839, n4450, CRC_OUT_8_12 );
nand U6790 ( n1890, n3849, n3850 );
nor U6791 ( n3850, n3852, n3853 );
nor U6792 ( n3849, n3857, n3858 );
and U6793 ( n3853, n4450, CRC_OUT_8_13 );
nand U6794 ( n1885, n3863, n3864 );
nor U6795 ( n3864, n3865, n3867 );
nor U6796 ( n3863, n3870, n3872 );
and U6797 ( n3867, n4450, CRC_OUT_8_14 );
nand U6798 ( n1880, n3877, n3878 );
nor U6799 ( n3878, n3879, n3880 );
nor U6800 ( n3877, n3884, n3885 );
and U6801 ( n3880, n4449, CRC_OUT_8_15 );
nand U6802 ( n1875, n3890, n3892 );
nor U6803 ( n3892, n3893, n3894 );
nor U6804 ( n3890, n3899, n3900 );
and U6805 ( n3894, n4449, CRC_OUT_8_16 );
nand U6806 ( n1870, n3907, n3908 );
nor U6807 ( n3908, n3909, n3910 );
nor U6808 ( n3907, n3915, n3917 );
and U6809 ( n3910, n4449, CRC_OUT_8_17 );
nand U6810 ( n1865, n3923, n3924 );
nor U6811 ( n3924, n3925, n3927 );
nor U6812 ( n3923, n3932, n3933 );
and U6813 ( n3927, n4449, CRC_OUT_8_18 );
nand U6814 ( n1860, n3939, n3940 );
nor U6815 ( n3940, n3942, n3943 );
nor U6816 ( n3939, n3948, n3949 );
and U6817 ( n3943, n4449, CRC_OUT_8_19 );
nand U6818 ( n1855, n3955, n3957 );
nor U6819 ( n3957, n3958, n3959 );
nor U6820 ( n3955, n3964, n3965 );
and U6821 ( n3959, n4449, CRC_OUT_8_20 );
nand U6822 ( n1850, n3972, n3973 );
nor U6823 ( n3973, n3974, n3975 );
nor U6824 ( n3972, n3980, n3982 );
and U6825 ( n3975, n4449, CRC_OUT_8_21 );
nand U6826 ( n1825, n4053, n4054 );
nor U6827 ( n4054, n4055, n4057 );
nor U6828 ( n4053, n4062, n4063 );
and U6829 ( n4057, n4449, CRC_OUT_8_26 );
nand U6830 ( n1820, n4069, n4070 );
nor U6831 ( n4070, n4072, n4073 );
nor U6832 ( n4069, n4078, n4079 );
and U6833 ( n4073, n4449, CRC_OUT_8_27 );
nand U6834 ( n1815, n4085, n4087 );
nor U6835 ( n4087, n4088, n4089 );
nor U6836 ( n4085, n4094, n4095 );
and U6837 ( n4089, n4448, CRC_OUT_8_28 );
nand U6838 ( n1810, n4102, n4103 );
nor U6839 ( n4103, n4104, n4105 );
nor U6840 ( n4102, n4110, n4112 );
and U6841 ( n4105, n4448, CRC_OUT_8_29 );
nand U6842 ( n1805, n4118, n4119 );
nor U6843 ( n4119, n4120, n4122 );
nor U6844 ( n4118, n4127, n4128 );
and U6845 ( n4122, n4448, CRC_OUT_8_30 );
nand U6846 ( n2883, n3246, n3247 );
nor U6847 ( n3247, n3249, n3250 );
nor U6848 ( n3246, n3254, n3255 );
and U6849 ( n3250, n4453, CRC_OUT_7_0 );
nand U6850 ( n2878, n3259, n3260 );
nor U6851 ( n3260, n3261, n3262 );
nor U6852 ( n3259, n3266, n3267 );
and U6853 ( n3262, n4453, CRC_OUT_7_1 );
nand U6854 ( n2873, n3271, n3272 );
nor U6855 ( n3272, n3274, n3275 );
nor U6856 ( n3271, n3279, n3280 );
and U6857 ( n3275, n4453, CRC_OUT_7_2 );
nand U6858 ( n2868, n3284, n3285 );
nor U6859 ( n3285, n3286, n3287 );
nor U6860 ( n3284, n3291, n3292 );
and U6861 ( n3287, n4453, CRC_OUT_7_3 );
nand U6862 ( n2863, n3296, n3297 );
nor U6863 ( n3297, n3299, n3300 );
nor U6864 ( n3296, n3304, n3305 );
and U6865 ( n3300, n4453, CRC_OUT_7_4 );
nand U6866 ( n2858, n3309, n3310 );
nor U6867 ( n3310, n3311, n3312 );
nor U6868 ( n3309, n3316, n3317 );
and U6869 ( n3312, n4453, CRC_OUT_7_5 );
nand U6870 ( n2853, n3321, n3322 );
nor U6871 ( n3322, n3324, n3325 );
nor U6872 ( n3321, n3329, n3330 );
and U6873 ( n3325, n4453, CRC_OUT_7_6 );
nand U6874 ( n2848, n3334, n3335 );
nor U6875 ( n3335, n3336, n3337 );
nor U6876 ( n3334, n3341, n3342 );
and U6877 ( n3337, n4453, CRC_OUT_7_7 );
nand U6878 ( n2843, n3346, n3347 );
nor U6879 ( n3347, n3349, n3350 );
nor U6880 ( n3346, n3354, n3355 );
and U6881 ( n3350, n4452, CRC_OUT_7_8 );
nand U6882 ( n2838, n3359, n3360 );
nor U6883 ( n3360, n3361, n3362 );
nor U6884 ( n3359, n3366, n3367 );
and U6885 ( n3362, n4452, CRC_OUT_7_9 );
nand U6886 ( n2833, n3371, n3373 );
nor U6887 ( n3373, n3374, n3375 );
nor U6888 ( n3371, n3379, n3381 );
and U6889 ( n3375, n4452, CRC_OUT_7_10 );
nand U6890 ( n2828, n3385, n3386 );
nor U6891 ( n3386, n3387, n3389 );
nor U6892 ( n3385, n3393, n3394 );
and U6893 ( n3389, n4452, CRC_OUT_7_11 );
nand U6894 ( n2823, n3398, n3399 );
nor U6895 ( n3399, n3401, n3402 );
nor U6896 ( n3398, n3406, n3407 );
and U6897 ( n3402, n4452, CRC_OUT_7_12 );
nand U6898 ( n2818, n3411, n3413 );
nor U6899 ( n3413, n3414, n3415 );
nor U6900 ( n3411, n3419, n3421 );
and U6901 ( n3415, n4452, CRC_OUT_7_13 );
nand U6902 ( n2813, n3425, n3426 );
nor U6903 ( n3426, n3427, n3429 );
nor U6904 ( n3425, n3433, n3434 );
and U6905 ( n3429, n4452, CRC_OUT_7_14 );
nand U6906 ( n2808, n3438, n3439 );
nor U6907 ( n3439, n3441, n3442 );
nor U6908 ( n3438, n3446, n3447 );
and U6909 ( n3442, n4452, CRC_OUT_7_15 );
nand U6910 ( n2803, n3451, n3453 );
nor U6911 ( n3453, n3454, n3455 );
nor U6912 ( n3451, n3461, n3462 );
and U6913 ( n3455, n4452, CRC_OUT_7_16 );
nand U6914 ( n2798, n3466, n3467 );
nor U6915 ( n3467, n3469, n3470 );
nor U6916 ( n3466, n3475, n3477 );
and U6917 ( n3470, n4452, CRC_OUT_7_17 );
nand U6918 ( n2793, n3481, n3482 );
nor U6919 ( n3482, n3483, n3485 );
nor U6920 ( n3481, n3490, n3491 );
and U6921 ( n3485, n4452, CRC_OUT_7_18 );
nand U6922 ( n2788, n3495, n3496 );
nor U6923 ( n3496, n3497, n3498 );
nor U6924 ( n3495, n3502, n3503 );
and U6925 ( n3498, n4452, CRC_OUT_7_19 );
nand U6926 ( n2783, n3506, n3507 );
nor U6927 ( n3507, n3508, n3509 );
nor U6928 ( n3506, n3513, n3514 );
and U6929 ( n3509, n4452, CRC_OUT_7_20 );
nand U6930 ( n2778, n3517, n3518 );
nor U6931 ( n3518, n3519, n3520 );
nor U6932 ( n3517, n3524, n3525 );
and U6933 ( n3520, n4451, CRC_OUT_7_21 );
nand U6934 ( n2773, n3528, n3529 );
nor U6935 ( n3529, n3530, n3531 );
nor U6936 ( n3528, n3535, n3536 );
and U6937 ( n3531, n4451, CRC_OUT_7_22 );
nand U6938 ( n2768, n3539, n3540 );
nor U6939 ( n3540, n3541, n3542 );
nor U6940 ( n3539, n3546, n3547 );
and U6941 ( n3542, n4451, CRC_OUT_7_23 );
nand U6942 ( n2763, n3550, n3551 );
nor U6943 ( n3551, n3552, n3553 );
nor U6944 ( n3550, n3557, n3558 );
and U6945 ( n3553, n4451, CRC_OUT_7_24 );
nand U6946 ( n2758, n3561, n3562 );
nor U6947 ( n3562, n3563, n3564 );
nor U6948 ( n3561, n3568, n3569 );
and U6949 ( n3564, n4451, CRC_OUT_7_25 );
nand U6950 ( n2753, n3572, n3573 );
nor U6951 ( n3573, n3574, n3575 );
nor U6952 ( n3572, n3579, n3580 );
and U6953 ( n3575, n4451, CRC_OUT_7_26 );
nand U6954 ( n2748, n3583, n3584 );
nor U6955 ( n3584, n3585, n3586 );
nor U6956 ( n3583, n3590, n3591 );
and U6957 ( n3586, n4451, CRC_OUT_7_27 );
nand U6958 ( n2743, n3594, n3595 );
nor U6959 ( n3595, n3596, n3597 );
nor U6960 ( n3594, n3601, n3602 );
and U6961 ( n3597, n4451, CRC_OUT_7_28 );
nand U6962 ( n2738, n3605, n3606 );
nor U6963 ( n3606, n3607, n3608 );
nor U6964 ( n3605, n3612, n3613 );
and U6965 ( n3608, n4451, CRC_OUT_7_29 );
nand U6966 ( n2733, n3616, n3617 );
nor U6967 ( n3617, n3618, n3619 );
nor U6968 ( n3616, n3623, n3624 );
and U6969 ( n3619, n4451, CRC_OUT_7_30 );
nand U6970 ( n3811, n2784, n2785 );
nor U6971 ( n2785, n2786, n2787 );
nor U6972 ( n2784, n2791, n2792 );
and U6973 ( n2787, n4456, CRC_OUT_6_0 );
nand U6974 ( n3806, n2796, n2797 );
nor U6975 ( n2797, n2799, n2800 );
nor U6976 ( n2796, n2804, n2805 );
and U6977 ( n2800, n4456, CRC_OUT_6_1 );
nand U6978 ( n3801, n2809, n2810 );
nor U6979 ( n2810, n2811, n2812 );
nor U6980 ( n2809, n2816, n2817 );
and U6981 ( n2812, n4455, CRC_OUT_6_2 );
nand U6982 ( n3796, n2821, n2822 );
nor U6983 ( n2822, n2824, n2825 );
nor U6984 ( n2821, n2829, n2830 );
and U6985 ( n2825, n4455, CRC_OUT_6_3 );
nand U6986 ( n3791, n2834, n2835 );
nor U6987 ( n2835, n2836, n2837 );
nor U6988 ( n2834, n2841, n2842 );
and U6989 ( n2837, n4455, CRC_OUT_6_4 );
nand U6990 ( n3786, n2846, n2847 );
nor U6991 ( n2847, n2849, n2850 );
nor U6992 ( n2846, n2854, n2855 );
and U6993 ( n2850, n4455, CRC_OUT_6_5 );
nand U6994 ( n3781, n2859, n2860 );
nor U6995 ( n2860, n2861, n2862 );
nor U6996 ( n2859, n2866, n2867 );
and U6997 ( n2862, n4455, CRC_OUT_6_6 );
nand U6998 ( n3776, n2871, n2872 );
nor U6999 ( n2872, n2874, n2875 );
nor U7000 ( n2871, n2879, n2880 );
and U7001 ( n2875, n4455, CRC_OUT_6_7 );
nand U7002 ( n3771, n2884, n2885 );
nor U7003 ( n2885, n2886, n2887 );
nor U7004 ( n2884, n2891, n2892 );
and U7005 ( n2887, n4455, CRC_OUT_6_8 );
nand U7006 ( n3766, n2896, n2897 );
nor U7007 ( n2897, n2899, n2900 );
nor U7008 ( n2896, n2904, n2905 );
and U7009 ( n2900, n4455, CRC_OUT_6_9 );
nand U7010 ( n3761, n2909, n2910 );
nor U7011 ( n2910, n2911, n2912 );
nor U7012 ( n2909, n2916, n2917 );
and U7013 ( n2912, n4455, CRC_OUT_6_10 );
nand U7014 ( n3756, n2921, n2922 );
nor U7015 ( n2922, n2924, n2925 );
nor U7016 ( n2921, n2929, n2930 );
and U7017 ( n2925, n4455, CRC_OUT_6_11 );
nand U7018 ( n3751, n2934, n2935 );
nor U7019 ( n2935, n2936, n2937 );
nor U7020 ( n2934, n2941, n2942 );
and U7021 ( n2937, n4455, CRC_OUT_6_12 );
nand U7022 ( n3746, n2946, n2947 );
nor U7023 ( n2947, n2949, n2950 );
nor U7024 ( n2946, n2954, n2955 );
and U7025 ( n2950, n4455, CRC_OUT_6_13 );
nand U7026 ( n3741, n2959, n2960 );
nor U7027 ( n2960, n2961, n2962 );
nor U7028 ( n2959, n2966, n2967 );
and U7029 ( n2962, n4455, CRC_OUT_6_14 );
nand U7030 ( n3736, n2971, n2972 );
nor U7031 ( n2972, n2974, n2975 );
nor U7032 ( n2971, n2979, n2980 );
and U7033 ( n2975, n4454, CRC_OUT_6_15 );
nand U7034 ( n3731, n2984, n2985 );
nor U7035 ( n2985, n2986, n2987 );
nor U7036 ( n2984, n2992, n2994 );
and U7037 ( n2987, n4454, CRC_OUT_6_16 );
nand U7038 ( n3726, n2997, n2999 );
nor U7039 ( n2999, n3000, n3001 );
nor U7040 ( n2997, n3006, n3007 );
and U7041 ( n3001, n4454, CRC_OUT_6_17 );
nand U7042 ( n3721, n3011, n3012 );
nor U7043 ( n3012, n3014, n3015 );
nor U7044 ( n3011, n3020, n3021 );
and U7045 ( n3015, n4454, CRC_OUT_6_18 );
nand U7046 ( n3716, n3025, n3026 );
nor U7047 ( n3026, n3027, n3029 );
nor U7048 ( n3025, n3034, n3035 );
and U7049 ( n3029, n4454, CRC_OUT_6_19 );
nand U7050 ( n3711, n3039, n3040 );
nor U7051 ( n3040, n3041, n3042 );
nor U7052 ( n3039, n3047, n3049 );
and U7053 ( n3042, n4454, CRC_OUT_6_20 );
nand U7054 ( n3706, n3052, n3054 );
nor U7055 ( n3054, n3055, n3056 );
nor U7056 ( n3052, n3061, n3062 );
and U7057 ( n3056, n4454, CRC_OUT_6_21 );
nand U7058 ( n3701, n3066, n3067 );
nor U7059 ( n3067, n3069, n3070 );
nor U7060 ( n3066, n3075, n3076 );
and U7061 ( n3070, n4454, CRC_OUT_6_22 );
nand U7062 ( n3696, n3080, n3081 );
nor U7063 ( n3081, n3082, n3084 );
nor U7064 ( n3080, n3089, n3090 );
and U7065 ( n3084, n4454, CRC_OUT_6_23 );
nand U7066 ( n3691, n3094, n3095 );
nor U7067 ( n3095, n3096, n3097 );
nor U7068 ( n3094, n3102, n3104 );
and U7069 ( n3097, n4454, CRC_OUT_6_24 );
nand U7070 ( n3686, n3107, n3109 );
nor U7071 ( n3109, n3110, n3111 );
nor U7072 ( n3107, n3116, n3117 );
and U7073 ( n3111, n4454, CRC_OUT_6_25 );
nand U7074 ( n3681, n3121, n3122 );
nor U7075 ( n3122, n3124, n3125 );
nor U7076 ( n3121, n3130, n3131 );
and U7077 ( n3125, n4454, CRC_OUT_6_26 );
nand U7078 ( n3676, n3135, n3136 );
nor U7079 ( n3136, n3137, n3139 );
nor U7080 ( n3135, n3144, n3145 );
and U7081 ( n3139, n4454, CRC_OUT_6_27 );
nand U7082 ( n3671, n3149, n3150 );
nor U7083 ( n3150, n3151, n3152 );
nor U7084 ( n3149, n3157, n3159 );
and U7085 ( n3152, n4453, CRC_OUT_6_28 );
nand U7086 ( n3666, n3162, n3164 );
nor U7087 ( n3164, n3165, n3166 );
nor U7088 ( n3162, n3171, n3172 );
and U7089 ( n3166, n4453, CRC_OUT_6_29 );
nand U7090 ( n3661, n3176, n3177 );
nor U7091 ( n3177, n3179, n3180 );
nor U7092 ( n3176, n3185, n3186 );
and U7093 ( n3180, n4453, CRC_OUT_6_30 );
nand U7094 ( n4739, n2352, n2353 );
nor U7095 ( n2353, n2354, n2356 );
nor U7096 ( n2352, n2359, n2361 );
and U7097 ( n2356, n4458, CRC_OUT_5_0 );
nand U7098 ( n4734, n2364, n2366 );
nor U7099 ( n2366, n2367, n2368 );
nor U7100 ( n2364, n2372, n2373 );
and U7101 ( n2368, n4458, CRC_OUT_5_1 );
nand U7102 ( n4729, n2377, n2378 );
nor U7103 ( n2378, n2379, n2381 );
nor U7104 ( n2377, n2384, n2386 );
and U7105 ( n2381, n4458, CRC_OUT_5_2 );
nand U7106 ( n4724, n2389, n2391 );
nor U7107 ( n2391, n2392, n2393 );
nor U7108 ( n2389, n2397, n2398 );
and U7109 ( n2393, n4458, CRC_OUT_5_3 );
nand U7110 ( n4719, n2402, n2403 );
nor U7111 ( n2403, n2404, n2406 );
nor U7112 ( n2402, n2409, n2411 );
and U7113 ( n2406, n4458, CRC_OUT_5_4 );
nand U7114 ( n4714, n2414, n2416 );
nor U7115 ( n2416, n2417, n2418 );
nor U7116 ( n2414, n2422, n2423 );
and U7117 ( n2418, n4458, CRC_OUT_5_5 );
nand U7118 ( n4709, n2427, n2428 );
nor U7119 ( n2428, n2429, n2431 );
nor U7120 ( n2427, n2434, n2436 );
and U7121 ( n2431, n4458, CRC_OUT_5_6 );
nand U7122 ( n4704, n2439, n2441 );
nor U7123 ( n2441, n2442, n2443 );
nor U7124 ( n2439, n2447, n2449 );
and U7125 ( n2443, n4458, CRC_OUT_5_7 );
nand U7126 ( n4699, n2453, n2454 );
nor U7127 ( n2454, n2455, n2457 );
nor U7128 ( n2453, n2461, n2462 );
and U7129 ( n2457, n4457, CRC_OUT_5_8 );
nand U7130 ( n4694, n2466, n2467 );
nor U7131 ( n2467, n2469, n2470 );
nor U7132 ( n2466, n2474, n2475 );
and U7133 ( n2470, n4457, CRC_OUT_5_9 );
nand U7134 ( n4689, n2479, n2481 );
nor U7135 ( n2481, n2482, n2483 );
nor U7136 ( n2479, n2487, n2489 );
and U7137 ( n2483, n4457, CRC_OUT_5_10 );
nand U7138 ( n4684, n2493, n2494 );
nor U7139 ( n2494, n2495, n2497 );
nor U7140 ( n2493, n2501, n2502 );
and U7141 ( n2497, n4457, CRC_OUT_5_11 );
nand U7142 ( n4679, n2506, n2507 );
nor U7143 ( n2507, n2509, n2510 );
nor U7144 ( n2506, n2514, n2515 );
and U7145 ( n2510, n4457, CRC_OUT_5_12 );
nand U7146 ( n4674, n2519, n2521 );
nor U7147 ( n2521, n2522, n2523 );
nor U7148 ( n2519, n2527, n2529 );
and U7149 ( n2523, n4457, CRC_OUT_5_13 );
nand U7150 ( n4669, n2533, n2534 );
nor U7151 ( n2534, n2535, n2537 );
nor U7152 ( n2533, n2541, n2542 );
and U7153 ( n2537, n4457, CRC_OUT_5_14 );
nand U7154 ( n4664, n2546, n2547 );
nor U7155 ( n2547, n2549, n2550 );
nor U7156 ( n2546, n2554, n2555 );
and U7157 ( n2550, n4457, CRC_OUT_5_15 );
nand U7158 ( n4659, n2559, n2561 );
nor U7159 ( n2561, n2562, n2563 );
nor U7160 ( n2559, n2568, n2569 );
and U7161 ( n2563, n4457, CRC_OUT_5_16 );
nand U7162 ( n4654, n2572, n2573 );
nor U7163 ( n2573, n2574, n2575 );
nor U7164 ( n2572, n2579, n2580 );
and U7165 ( n2575, n4457, CRC_OUT_5_17 );
nand U7166 ( n4649, n2583, n2584 );
nor U7167 ( n2584, n2585, n2586 );
nor U7168 ( n2583, n2590, n2591 );
and U7169 ( n2586, n4457, CRC_OUT_5_18 );
nand U7170 ( n4644, n2594, n2595 );
nor U7171 ( n2595, n2596, n2597 );
nor U7172 ( n2594, n2601, n2602 );
and U7173 ( n2597, n4457, CRC_OUT_5_19 );
nand U7174 ( n4639, n2605, n2606 );
nor U7175 ( n2606, n2607, n2608 );
nor U7176 ( n2605, n2612, n2613 );
and U7177 ( n2608, n4457, CRC_OUT_5_20 );
nand U7178 ( n4634, n2616, n2617 );
nor U7179 ( n2617, n2618, n2619 );
nor U7180 ( n2616, n2623, n2624 );
and U7181 ( n2619, n4456, CRC_OUT_5_21 );
nand U7182 ( n4629, n2627, n2628 );
nor U7183 ( n2628, n2629, n2630 );
nor U7184 ( n2627, n2634, n2635 );
and U7185 ( n2630, n4456, CRC_OUT_5_22 );
nand U7186 ( n4624, n2638, n2639 );
nor U7187 ( n2639, n2640, n2641 );
nor U7188 ( n2638, n2645, n2646 );
and U7189 ( n2641, n4456, CRC_OUT_5_23 );
nand U7190 ( n4619, n2649, n2650 );
nor U7191 ( n2650, n2651, n2652 );
nor U7192 ( n2649, n2656, n2657 );
and U7193 ( n2652, n4456, CRC_OUT_5_24 );
nand U7194 ( n4614, n2660, n2661 );
nor U7195 ( n2661, n2662, n2663 );
nor U7196 ( n2660, n2667, n2668 );
and U7197 ( n2663, n4456, CRC_OUT_5_25 );
nand U7198 ( n4609, n2671, n2672 );
nor U7199 ( n2672, n2673, n2674 );
nor U7200 ( n2671, n2678, n2679 );
and U7201 ( n2674, n4456, CRC_OUT_5_26 );
nand U7202 ( n4604, n2682, n2683 );
nor U7203 ( n2683, n2684, n2685 );
nor U7204 ( n2682, n2689, n2690 );
and U7205 ( n2685, n4456, CRC_OUT_5_27 );
nand U7206 ( n4599, n2693, n2694 );
nor U7207 ( n2694, n2695, n2696 );
nor U7208 ( n2693, n2700, n2701 );
and U7209 ( n2696, n4456, CRC_OUT_5_28 );
nand U7210 ( n4594, n2704, n2705 );
nor U7211 ( n2705, n2706, n2707 );
nor U7212 ( n2704, n2711, n2712 );
and U7213 ( n2707, n4456, CRC_OUT_5_29 );
nand U7214 ( n4589, n2715, n2716 );
nor U7215 ( n2716, n2717, n2718 );
nor U7216 ( n2715, n2722, n2724 );
and U7217 ( n2718, n4456, CRC_OUT_5_30 );
nand U7218 ( n5667, n1889, n1891 );
nor U7219 ( n1891, n1892, n1893 );
nor U7220 ( n1889, n1897, n1898 );
and U7221 ( n1893, n4441, CRC_OUT_4_0 );
nand U7222 ( n5662, n1902, n1903 );
nor U7223 ( n1903, n1904, n1906 );
nor U7224 ( n1902, n1909, n1911 );
and U7225 ( n1906, n4440, CRC_OUT_4_1 );
nand U7226 ( n5657, n1914, n1916 );
nor U7227 ( n1916, n1917, n1918 );
nor U7228 ( n1914, n1922, n1923 );
and U7229 ( n1918, n4441, CRC_OUT_4_2 );
nand U7230 ( n5652, n1927, n1928 );
nor U7231 ( n1928, n1929, n1931 );
nor U7232 ( n1927, n1934, n1936 );
and U7233 ( n1931, n4441, CRC_OUT_4_3 );
nand U7234 ( n5647, n1939, n1941 );
nor U7235 ( n1941, n1942, n1943 );
nor U7236 ( n1939, n1947, n1948 );
and U7237 ( n1943, n4441, CRC_OUT_4_4 );
nand U7238 ( n5642, n1952, n1953 );
nor U7239 ( n1953, n1954, n1956 );
nor U7240 ( n1952, n1959, n1961 );
and U7241 ( n1956, n4440, CRC_OUT_4_5 );
nand U7242 ( n5637, n1964, n1966 );
nor U7243 ( n1966, n1967, n1968 );
nor U7244 ( n1964, n1972, n1973 );
and U7245 ( n1968, n4441, CRC_OUT_4_6 );
nand U7246 ( n5632, n1977, n1978 );
nor U7247 ( n1978, n1979, n1981 );
nor U7248 ( n1977, n1984, n1986 );
and U7249 ( n1981, n4440, CRC_OUT_4_7 );
nand U7250 ( n5627, n1989, n1991 );
nor U7251 ( n1991, n1992, n1993 );
nor U7252 ( n1989, n1997, n1998 );
and U7253 ( n1993, n4440, CRC_OUT_4_8 );
nand U7254 ( n5622, n2002, n2003 );
nor U7255 ( n2003, n2004, n2006 );
nor U7256 ( n2002, n2009, n2011 );
and U7257 ( n2006, n4441, CRC_OUT_4_9 );
nand U7258 ( n5617, n2014, n2016 );
nor U7259 ( n2016, n2017, n2018 );
nor U7260 ( n2014, n2022, n2023 );
and U7261 ( n2018, n4440, CRC_OUT_4_10 );
nand U7262 ( n5612, n2027, n2028 );
nor U7263 ( n2028, n2029, n2031 );
nor U7264 ( n2027, n2034, n2036 );
and U7265 ( n2031, n4440, CRC_OUT_4_11 );
nand U7266 ( n5607, n2039, n2041 );
nor U7267 ( n2041, n2042, n2043 );
nor U7268 ( n2039, n2047, n2048 );
and U7269 ( n2043, n4441, CRC_OUT_4_12 );
nand U7270 ( n5602, n2052, n2053 );
nor U7271 ( n2053, n2054, n2056 );
nor U7272 ( n2052, n2059, n2061 );
and U7273 ( n2056, n4440, CRC_OUT_4_13 );
nand U7274 ( n5597, n2064, n2066 );
nor U7275 ( n2066, n2067, n2068 );
nor U7276 ( n2064, n2072, n2073 );
and U7277 ( n2068, n4439, CRC_OUT_4_14 );
nand U7278 ( n5592, n2077, n2078 );
nor U7279 ( n2078, n2079, n2081 );
nor U7280 ( n2077, n2084, n2086 );
and U7281 ( n2081, n4440, CRC_OUT_4_15 );
nand U7282 ( n5587, n2089, n2091 );
nor U7283 ( n2091, n2092, n2093 );
nor U7284 ( n2089, n2098, n2099 );
and U7285 ( n2093, n4439, CRC_OUT_4_16 );
nand U7286 ( n5582, n2103, n2104 );
nor U7287 ( n2104, n2106, n2107 );
nor U7288 ( n2103, n2112, n2113 );
and U7289 ( n2107, n4439, CRC_OUT_4_17 );
nand U7290 ( n5577, n2117, n2118 );
nor U7291 ( n2118, n2119, n2121 );
nor U7292 ( n2117, n2126, n2127 );
and U7293 ( n2121, n4440, CRC_OUT_4_18 );
nand U7294 ( n5572, n2131, n2132 );
nor U7295 ( n2132, n2133, n2134 );
nor U7296 ( n2131, n2139, n2141 );
and U7297 ( n2134, n4441, CRC_OUT_4_19 );
nand U7298 ( n5567, n2144, n2146 );
nor U7299 ( n2146, n2147, n2148 );
nor U7300 ( n2144, n2153, n2154 );
and U7301 ( n2148, n4439, CRC_OUT_4_20 );
nand U7302 ( n5562, n2158, n2159 );
nor U7303 ( n2159, n2161, n2162 );
nor U7304 ( n2158, n2167, n2168 );
and U7305 ( n2162, n4444, CRC_OUT_4_21 );
nand U7306 ( n5557, n2172, n2173 );
nor U7307 ( n2173, n2174, n2176 );
nor U7308 ( n2172, n2181, n2182 );
and U7309 ( n2176, n4459, CRC_OUT_4_22 );
nand U7310 ( n5552, n2186, n2187 );
nor U7311 ( n2187, n2188, n2189 );
nor U7312 ( n2186, n2194, n2196 );
and U7313 ( n2189, n4459, CRC_OUT_4_23 );
nand U7314 ( n5547, n2199, n2201 );
nor U7315 ( n2201, n2202, n2203 );
nor U7316 ( n2199, n2208, n2209 );
and U7317 ( n2203, n4459, CRC_OUT_4_24 );
nand U7318 ( n5542, n2213, n2214 );
nor U7319 ( n2214, n2216, n2217 );
nor U7320 ( n2213, n2222, n2223 );
and U7321 ( n2217, n4459, CRC_OUT_4_25 );
nand U7322 ( n5537, n2227, n2228 );
nor U7323 ( n2228, n2229, n2231 );
nor U7324 ( n2227, n2236, n2237 );
and U7325 ( n2231, n4459, CRC_OUT_4_26 );
nand U7326 ( n5532, n2241, n2242 );
nor U7327 ( n2242, n2243, n2244 );
nor U7328 ( n2241, n2249, n2251 );
and U7329 ( n2244, n4458, CRC_OUT_4_27 );
nand U7330 ( n5527, n2254, n2256 );
nor U7331 ( n2256, n2257, n2258 );
nor U7332 ( n2254, n2263, n2264 );
and U7333 ( n2258, n4458, CRC_OUT_4_28 );
nand U7334 ( n5522, n2268, n2269 );
nor U7335 ( n2269, n2271, n2272 );
nor U7336 ( n2268, n2277, n2278 );
and U7337 ( n2272, n4458, CRC_OUT_4_29 );
nand U7338 ( n5517, n2282, n2283 );
nor U7339 ( n2283, n2284, n2286 );
nor U7340 ( n2282, n2291, n2292 );
and U7341 ( n2286, n4458, CRC_OUT_4_30 );
nand U7342 ( n6595, n1458, n1459 );
nor U7343 ( n1459, n1460, n1461 );
nor U7344 ( n1458, n1465, n1466 );
and U7345 ( n1461, n4443, CRC_OUT_3_0 );
nand U7346 ( n6590, n1470, n1471 );
nor U7347 ( n1471, n1473, n1474 );
nor U7348 ( n1470, n1478, n1479 );
and U7349 ( n1474, n4443, CRC_OUT_3_1 );
nand U7350 ( n6585, n1483, n1484 );
nor U7351 ( n1484, n1485, n1486 );
nor U7352 ( n1483, n1490, n1491 );
and U7353 ( n1486, n4443, CRC_OUT_3_2 );
nand U7354 ( n6580, n1495, n1496 );
nor U7355 ( n1496, n1498, n1499 );
nor U7356 ( n1495, n1503, n1504 );
and U7357 ( n1499, n4443, CRC_OUT_3_3 );
nand U7358 ( n6575, n1508, n1509 );
nor U7359 ( n1509, n1510, n1511 );
nor U7360 ( n1508, n1515, n1517 );
and U7361 ( n1511, n4443, CRC_OUT_3_4 );
nand U7362 ( n6570, n1521, n1522 );
nor U7363 ( n1522, n1523, n1525 );
nor U7364 ( n1521, n1529, n1530 );
and U7365 ( n1525, n4443, CRC_OUT_3_5 );
nand U7366 ( n6565, n1534, n1535 );
nor U7367 ( n1535, n1537, n1538 );
nor U7368 ( n1534, n1542, n1543 );
and U7369 ( n1538, n4443, CRC_OUT_3_6 );
nand U7370 ( n6560, n1547, n1549 );
nor U7371 ( n1549, n1550, n1551 );
nor U7372 ( n1547, n1555, n1557 );
and U7373 ( n1551, n4443, CRC_OUT_3_7 );
nand U7374 ( n6555, n1561, n1562 );
nor U7375 ( n1562, n1563, n1565 );
nor U7376 ( n1561, n1569, n1570 );
and U7377 ( n1565, n4443, CRC_OUT_3_8 );
nand U7378 ( n6550, n1574, n1575 );
nor U7379 ( n1575, n1577, n1578 );
nor U7380 ( n1574, n1582, n1583 );
and U7381 ( n1578, n4443, CRC_OUT_3_9 );
nand U7382 ( n6545, n1587, n1589 );
nor U7383 ( n1589, n1590, n1591 );
nor U7384 ( n1587, n1595, n1597 );
and U7385 ( n1591, n4443, CRC_OUT_3_10 );
nand U7386 ( n6540, n1601, n1602 );
nor U7387 ( n1602, n1603, n1605 );
nor U7388 ( n1601, n1609, n1610 );
and U7389 ( n1605, n4442, CRC_OUT_3_11 );
nand U7390 ( n6535, n1614, n1615 );
nor U7391 ( n1615, n1617, n1618 );
nor U7392 ( n1614, n1622, n1623 );
and U7393 ( n1618, n4442, CRC_OUT_3_12 );
nand U7394 ( n6530, n1627, n1629 );
nor U7395 ( n1629, n1630, n1631 );
nor U7396 ( n1627, n1635, n1637 );
and U7397 ( n1631, n4442, CRC_OUT_3_13 );
nand U7398 ( n6525, n1640, n1641 );
nor U7399 ( n1641, n1642, n1643 );
nor U7400 ( n1640, n1646, n1647 );
and U7401 ( n1643, n4442, CRC_OUT_3_14 );
nand U7402 ( n6520, n1650, n1651 );
nor U7403 ( n1651, n1652, n1653 );
nor U7404 ( n1650, n1656, n1657 );
and U7405 ( n1653, n4442, CRC_OUT_3_15 );
nand U7406 ( n6515, n1660, n1661 );
nor U7407 ( n1661, n1662, n1663 );
nor U7408 ( n1660, n1667, n1668 );
and U7409 ( n1663, n4442, CRC_OUT_3_16 );
nand U7410 ( n6510, n1671, n1672 );
nor U7411 ( n1672, n1673, n1674 );
nor U7412 ( n1671, n1678, n1679 );
and U7413 ( n1674, n4442, CRC_OUT_3_17 );
nand U7414 ( n6505, n1682, n1683 );
nor U7415 ( n1683, n1684, n1685 );
nor U7416 ( n1682, n1689, n1690 );
and U7417 ( n1685, n4442, CRC_OUT_3_18 );
nand U7418 ( n6500, n1693, n1694 );
nor U7419 ( n1694, n1695, n1696 );
nor U7420 ( n1693, n1700, n1701 );
and U7421 ( n1696, n4442, CRC_OUT_3_19 );
nand U7422 ( n6495, n1704, n1705 );
nor U7423 ( n1705, n1706, n1707 );
nor U7424 ( n1704, n1711, n1712 );
and U7425 ( n1707, n4442, CRC_OUT_3_20 );
nand U7426 ( n6490, n1715, n1716 );
nor U7427 ( n1716, n1717, n1718 );
nor U7428 ( n1715, n1722, n1723 );
and U7429 ( n1718, n4442, CRC_OUT_3_21 );
nand U7430 ( n6485, n1726, n1727 );
nor U7431 ( n1727, n1728, n1729 );
nor U7432 ( n1726, n1733, n1734 );
and U7433 ( n1729, n4442, CRC_OUT_3_22 );
nand U7434 ( n6480, n1737, n1738 );
nor U7435 ( n1738, n1739, n1740 );
nor U7436 ( n1737, n1744, n1745 );
and U7437 ( n1740, n4442, CRC_OUT_3_23 );
nand U7438 ( n6475, n1748, n1749 );
nor U7439 ( n1749, n1750, n1751 );
nor U7440 ( n1748, n1755, n1756 );
and U7441 ( n1751, n4441, CRC_OUT_3_24 );
nand U7442 ( n6470, n1759, n1760 );
nor U7443 ( n1760, n1761, n1762 );
nor U7444 ( n1759, n1766, n1767 );
and U7445 ( n1762, n4441, CRC_OUT_3_25 );
nand U7446 ( n6465, n1770, n1771 );
nor U7447 ( n1771, n1772, n1773 );
nor U7448 ( n1770, n1777, n1778 );
and U7449 ( n1773, n4441, CRC_OUT_3_26 );
nand U7450 ( n6460, n1781, n1782 );
nor U7451 ( n1782, n1783, n1784 );
nor U7452 ( n1781, n1788, n1789 );
and U7453 ( n1784, n4441, CRC_OUT_3_27 );
nand U7454 ( n6455, n1792, n1793 );
nor U7455 ( n1793, n1794, n1796 );
nor U7456 ( n1792, n1801, n1802 );
and U7457 ( n1796, n4440, CRC_OUT_3_28 );
nand U7458 ( n6450, n1806, n1807 );
nor U7459 ( n1807, n1808, n1809 );
nor U7460 ( n1806, n1814, n1816 );
and U7461 ( n1809, n4441, CRC_OUT_3_29 );
nand U7462 ( n6445, n1819, n1821 );
nor U7463 ( n1821, n1822, n1823 );
nor U7464 ( n1819, n1828, n1829 );
and U7465 ( n1823, n4440, CRC_OUT_3_30 );
nand U7466 ( n7483, n1095, n1096 );
nor U7467 ( n1096, n1098, n1099 );
nor U7468 ( n1095, n1103, n1104 );
and U7469 ( n1099, n4445, CRC_OUT_2_8 );
nand U7470 ( n7478, n1108, n1109 );
nor U7471 ( n1109, n1110, n1111 );
nor U7472 ( n1108, n1115, n1116 );
and U7473 ( n1111, n4445, CRC_OUT_2_9 );
nand U7474 ( n7473, n1120, n1121 );
nor U7475 ( n1121, n1123, n1124 );
nor U7476 ( n1120, n1128, n1129 );
and U7477 ( n1124, n4445, CRC_OUT_2_10 );
nand U7478 ( n7468, n1133, n1134 );
nor U7479 ( n1134, n1135, n1136 );
nor U7480 ( n1133, n1140, n1141 );
and U7481 ( n1136, n4445, CRC_OUT_2_11 );
nand U7482 ( n7463, n1145, n1146 );
nor U7483 ( n1146, n1148, n1149 );
nor U7484 ( n1145, n1153, n1154 );
and U7485 ( n1149, n4445, CRC_OUT_2_12 );
nand U7486 ( n7458, n1158, n1159 );
nor U7487 ( n1159, n1160, n1161 );
nor U7488 ( n1158, n1165, n1166 );
and U7489 ( n1161, n4445, CRC_OUT_2_13 );
nand U7490 ( n7453, n1170, n1171 );
nor U7491 ( n1171, n1173, n1174 );
nor U7492 ( n1170, n1178, n1179 );
and U7493 ( n1174, n4445, CRC_OUT_2_14 );
nand U7494 ( n7448, n1183, n1184 );
nor U7495 ( n1184, n1185, n1186 );
nor U7496 ( n1183, n1190, n1191 );
and U7497 ( n1186, n4445, CRC_OUT_2_15 );
nand U7498 ( n7443, n1195, n1196 );
nor U7499 ( n1196, n1198, n1199 );
nor U7500 ( n1195, n1204, n1205 );
and U7501 ( n1199, n4445, CRC_OUT_2_16 );
nand U7502 ( n7438, n1209, n1210 );
nor U7503 ( n1210, n1211, n1213 );
nor U7504 ( n1209, n1218, n1219 );
and U7505 ( n1213, n4445, CRC_OUT_2_17 );
nand U7506 ( n7433, n1223, n1224 );
nor U7507 ( n1224, n1225, n1226 );
nor U7508 ( n1223, n1231, n1233 );
and U7509 ( n1226, n4444, CRC_OUT_2_18 );
nand U7510 ( n7428, n1236, n1238 );
nor U7511 ( n1238, n1239, n1240 );
nor U7512 ( n1236, n1245, n1246 );
and U7513 ( n1240, n4444, CRC_OUT_2_19 );
nand U7514 ( n7423, n1250, n1251 );
nor U7515 ( n1251, n1253, n1254 );
nor U7516 ( n1250, n1259, n1260 );
and U7517 ( n1254, n4444, CRC_OUT_2_20 );
nand U7518 ( n7418, n1264, n1265 );
nor U7519 ( n1265, n1266, n1268 );
nor U7520 ( n1264, n1273, n1274 );
and U7521 ( n1268, n4444, CRC_OUT_2_21 );
nand U7522 ( n7413, n1278, n1279 );
nor U7523 ( n1279, n1280, n1281 );
nor U7524 ( n1278, n1286, n1288 );
and U7525 ( n1281, n4444, CRC_OUT_2_22 );
nand U7526 ( n7408, n1291, n1293 );
nor U7527 ( n1293, n1294, n1295 );
nor U7528 ( n1291, n1300, n1301 );
and U7529 ( n1295, n4444, CRC_OUT_2_23 );
nand U7530 ( n7403, n1305, n1306 );
nor U7531 ( n1306, n1308, n1309 );
nor U7532 ( n1305, n1314, n1315 );
and U7533 ( n1309, n4444, CRC_OUT_2_24 );
nand U7534 ( n7398, n1319, n1320 );
nor U7535 ( n1320, n1321, n1323 );
nor U7536 ( n1319, n1328, n1329 );
and U7537 ( n1323, n4444, CRC_OUT_2_25 );
nand U7538 ( n7393, n1333, n1334 );
nor U7539 ( n1334, n1335, n1336 );
nor U7540 ( n1333, n1341, n1343 );
and U7541 ( n1336, n4444, CRC_OUT_2_26 );
nand U7542 ( n7388, n1346, n1348 );
nor U7543 ( n1348, n1349, n1350 );
nor U7544 ( n1346, n1355, n1356 );
and U7545 ( n1350, n4444, CRC_OUT_2_27 );
nand U7546 ( n7383, n1360, n1361 );
nor U7547 ( n1361, n1363, n1364 );
nor U7548 ( n1360, n1369, n1370 );
and U7549 ( n1364, n4444, CRC_OUT_2_28 );
nand U7550 ( n7378, n1374, n1375 );
nor U7551 ( n1375, n1376, n1378 );
nor U7552 ( n1374, n1383, n1384 );
and U7553 ( n1378, n4444, CRC_OUT_2_29 );
nand U7554 ( n7373, n1388, n1389 );
nor U7555 ( n1389, n1390, n1391 );
nor U7556 ( n1388, n1396, n1398 );
and U7557 ( n1391, n4443, CRC_OUT_2_30 );
nand U7558 ( n877, n650, n651 );
nor U7559 ( n651, n652, n653 );
nor U7560 ( n650, n655, n656 );
and U7561 ( n653, n4446, CRC_OUT_9_30 );
nand U7562 ( n882, n639, n640 );
nor U7563 ( n640, n641, n642 );
nor U7564 ( n639, n644, n645 );
and U7565 ( n642, n4446, CRC_OUT_9_29 );
nand U7566 ( n887, n628, n629 );
nor U7567 ( n629, n630, n631 );
nor U7568 ( n628, n633, n634 );
and U7569 ( n631, n4446, CRC_OUT_9_28 );
nand U7570 ( n892, n617, n618 );
nor U7571 ( n618, n619, n620 );
nor U7572 ( n617, n622, n623 );
and U7573 ( n620, n4446, CRC_OUT_9_27 );
nand U7574 ( n897, n596, n597 );
nor U7575 ( n597, n598, n599 );
nor U7576 ( n596, n601, n602 );
and U7577 ( n599, n4446, CRC_OUT_9_26 );
nand U7578 ( n902, n571, n572 );
nor U7579 ( n572, n573, n574 );
nor U7580 ( n571, n576, n577 );
and U7581 ( n574, n4446, CRC_OUT_9_25 );
nand U7582 ( n907, n549, n550 );
nor U7583 ( n550, n551, n552 );
nor U7584 ( n549, n554, n555 );
and U7585 ( n552, n4446, CRC_OUT_9_24 );
nand U7586 ( n912, n538, n539 );
nor U7587 ( n539, n540, n541 );
nor U7588 ( n538, n543, n544 );
and U7589 ( n541, n4447, CRC_OUT_9_23 );
nand U7590 ( n917, n527, n528 );
nor U7591 ( n528, n529, n530 );
nor U7592 ( n527, n532, n533 );
and U7593 ( n530, n4447, CRC_OUT_9_22 );
nand U7594 ( n922, n516, n517 );
nor U7595 ( n517, n518, n519 );
nor U7596 ( n516, n521, n522 );
and U7597 ( n519, n4447, CRC_OUT_9_21 );
nand U7598 ( n927, n505, n506 );
nor U7599 ( n506, n507, n508 );
nor U7600 ( n505, n510, n511 );
and U7601 ( n508, n4447, CRC_OUT_9_20 );
nand U7602 ( n932, n494, n495 );
nor U7603 ( n495, n496, n497 );
nor U7604 ( n494, n499, n500 );
and U7605 ( n497, n4447, CRC_OUT_9_19 );
nand U7606 ( n937, n483, n484 );
nor U7607 ( n484, n485, n486 );
nor U7608 ( n483, n488, n489 );
and U7609 ( n486, n4447, CRC_OUT_9_18 );
nand U7610 ( n942, n472, n473 );
nor U7611 ( n473, n474, n475 );
nor U7612 ( n472, n477, n478 );
and U7613 ( n475, n4447, CRC_OUT_9_17 );
nand U7614 ( n947, n461, n462 );
nor U7615 ( n462, n463, n464 );
nor U7616 ( n461, n466, n467 );
and U7617 ( n464, n4447, CRC_OUT_9_16 );
nand U7618 ( n952, n450, n451 );
nor U7619 ( n451, n452, n453 );
nor U7620 ( n450, n455, n456 );
and U7621 ( n453, n4447, CRC_OUT_9_15 );
nand U7622 ( n957, n439, n440 );
nor U7623 ( n440, n441, n442 );
nor U7624 ( n439, n444, n445 );
and U7625 ( n442, n4447, CRC_OUT_9_14 );
nand U7626 ( n962, n428, n429 );
nor U7627 ( n429, n430, n431 );
nor U7628 ( n428, n433, n434 );
and U7629 ( n431, n4447, CRC_OUT_9_13 );
nand U7630 ( n967, n417, n418 );
nor U7631 ( n418, n419, n420 );
nor U7632 ( n417, n422, n423 );
and U7633 ( n420, n4447, CRC_OUT_9_12 );
nand U7634 ( n972, n406, n407 );
nor U7635 ( n407, n408, n409 );
nor U7636 ( n406, n411, n412 );
and U7637 ( n409, n4447, CRC_OUT_9_11 );
nand U7638 ( n977, n395, n396 );
nor U7639 ( n396, n397, n398 );
nor U7640 ( n395, n400, n401 );
and U7641 ( n398, n4448, CRC_OUT_9_10 );
nand U7642 ( n7523, n995, n996 );
nor U7643 ( n996, n998, n999 );
nor U7644 ( n995, n1003, n1004 );
and U7645 ( n999, n4446, CRC_OUT_2_0 );
nand U7646 ( n7518, n1008, n1009 );
nor U7647 ( n1009, n1010, n1011 );
nor U7648 ( n1008, n1015, n1016 );
and U7649 ( n1011, n4446, CRC_OUT_2_1 );
nand U7650 ( n7513, n1020, n1021 );
nor U7651 ( n1021, n1023, n1024 );
nor U7652 ( n1020, n1028, n1029 );
and U7653 ( n1024, n4446, CRC_OUT_2_2 );
nand U7654 ( n7508, n1033, n1034 );
nor U7655 ( n1034, n1035, n1036 );
nor U7656 ( n1033, n1040, n1041 );
and U7657 ( n1036, n4446, CRC_OUT_2_3 );
nand U7658 ( n7503, n1045, n1046 );
nor U7659 ( n1046, n1048, n1049 );
nor U7660 ( n1045, n1053, n1054 );
and U7661 ( n1049, n4446, CRC_OUT_2_4 );
nand U7662 ( n7498, n1058, n1059 );
nor U7663 ( n1059, n1060, n1061 );
nor U7664 ( n1058, n1065, n1066 );
and U7665 ( n1061, n4445, CRC_OUT_2_5 );
nand U7666 ( n7493, n1070, n1071 );
nor U7667 ( n1071, n1073, n1074 );
nor U7668 ( n1070, n1078, n1079 );
and U7669 ( n1074, n4445, CRC_OUT_2_6 );
nand U7670 ( n7488, n1083, n1084 );
nor U7671 ( n1084, n1085, n1086 );
nor U7672 ( n1083, n1090, n1091 );
and U7673 ( n1086, n4445, CRC_OUT_2_7 );
nand U7674 ( n8451, n676, n677 );
and U7675 ( n677, n678, n679 );
nor U7676 ( n676, n681, n682 );
nand U7677 ( n679, DATA_0_0, n4341 );
nand U7678 ( n8446, n685, n686 );
and U7679 ( n686, n687, n688 );
nor U7680 ( n685, n689, n690 );
nand U7681 ( n688, DATA_0_1, n4341 );
nand U7682 ( n8441, n693, n694 );
and U7683 ( n694, n695, n696 );
nor U7684 ( n693, n697, n698 );
nand U7685 ( n696, DATA_0_2, n4341 );
nand U7686 ( n8436, n701, n702 );
and U7687 ( n702, n703, n704 );
nor U7688 ( n701, n705, n706 );
nand U7689 ( n704, DATA_0_3, n4341 );
nand U7690 ( n8431, n709, n710 );
and U7691 ( n710, n711, n712 );
nor U7692 ( n709, n713, n714 );
nand U7693 ( n712, DATA_0_4, n4341 );
nand U7694 ( n8426, n717, n718 );
and U7695 ( n718, n719, n720 );
nor U7696 ( n717, n721, n722 );
nand U7697 ( n720, DATA_0_5, n4341 );
nand U7698 ( n8421, n725, n726 );
and U7699 ( n726, n727, n728 );
nor U7700 ( n725, n729, n730 );
nand U7701 ( n728, DATA_0_6, n4341 );
nand U7702 ( n8416, n734, n735 );
and U7703 ( n735, n736, n737 );
nor U7704 ( n734, n738, n739 );
nand U7705 ( n737, DATA_0_7, n4341 );
nand U7706 ( n8411, n742, n743 );
and U7707 ( n743, n744, n745 );
nor U7708 ( n742, n746, n747 );
nand U7709 ( n745, DATA_0_8, n4341 );
nand U7710 ( n8406, n750, n751 );
and U7711 ( n751, n752, n753 );
nor U7712 ( n750, n754, n755 );
nand U7713 ( n753, DATA_0_9, n4341 );
nand U7714 ( n8401, n758, n759 );
and U7715 ( n759, n760, n761 );
nor U7716 ( n758, n762, n763 );
nand U7717 ( n761, DATA_0_10, n4341 );
nand U7718 ( n8396, n766, n767 );
and U7719 ( n767, n768, n769 );
nor U7720 ( n766, n770, n771 );
nand U7721 ( n769, DATA_0_11, n4341 );
nand U7722 ( n8391, n774, n775 );
and U7723 ( n775, n776, n777 );
nor U7724 ( n774, n778, n779 );
nand U7725 ( n777, DATA_0_12, n4341 );
nand U7726 ( n8386, n782, n783 );
and U7727 ( n783, n784, n785 );
nor U7728 ( n782, n786, n787 );
nand U7729 ( n785, DATA_0_13, n4339 );
nand U7730 ( n8381, n790, n791 );
and U7731 ( n791, n792, n793 );
nor U7732 ( n790, n794, n795 );
nand U7733 ( n793, DATA_0_14, n4339 );
nand U7734 ( n8376, n798, n799 );
and U7735 ( n799, n800, n801 );
nor U7736 ( n798, n802, n803 );
nand U7737 ( n801, DATA_0_15, n4339 );
nand U7738 ( n8371, n806, n807 );
and U7739 ( n807, n808, n809 );
nor U7740 ( n806, n810, n811 );
nand U7741 ( n809, DATA_0_16, n4339 );
nand U7742 ( n8366, n815, n816 );
and U7743 ( n816, n817, n818 );
nor U7744 ( n815, n819, n820 );
nand U7745 ( n818, DATA_0_17, n4339 );
nand U7746 ( n8361, n823, n824 );
and U7747 ( n824, n825, n826 );
nor U7748 ( n823, n827, n828 );
nand U7749 ( n826, DATA_0_18, n4339 );
nand U7750 ( n8356, n831, n832 );
and U7751 ( n832, n833, n834 );
nor U7752 ( n831, n835, n836 );
nand U7753 ( n834, DATA_0_19, n4339 );
nand U7754 ( n8351, n839, n840 );
and U7755 ( n840, n841, n842 );
nor U7756 ( n839, n843, n844 );
nand U7757 ( n842, DATA_0_20, n4339 );
nand U7758 ( n8346, n847, n848 );
and U7759 ( n848, n849, n850 );
nor U7760 ( n847, n851, n852 );
nand U7761 ( n850, DATA_0_21, n4339 );
nand U7762 ( n8341, n855, n856 );
and U7763 ( n856, n857, n858 );
nor U7764 ( n855, n859, n860 );
nand U7765 ( n858, DATA_0_22, n4339 );
nand U7766 ( n8336, n863, n864 );
and U7767 ( n864, n865, n866 );
nor U7768 ( n863, n868, n869 );
nand U7769 ( n866, DATA_0_23, n4339 );
nand U7770 ( n8331, n873, n874 );
and U7771 ( n874, n875, n876 );
nor U7772 ( n873, n878, n879 );
nand U7773 ( n876, DATA_0_24, n4339 );
nand U7774 ( n8326, n883, n884 );
and U7775 ( n884, n885, n886 );
nor U7776 ( n883, n888, n889 );
nand U7777 ( n886, DATA_0_25, n4339 );
nand U7778 ( n8321, n893, n894 );
and U7779 ( n894, n895, n896 );
nor U7780 ( n893, n898, n899 );
nand U7781 ( n896, DATA_0_26, n4339 );
nand U7782 ( n8316, n903, n904 );
and U7783 ( n904, n905, n906 );
nor U7784 ( n903, n908, n909 );
nand U7785 ( n906, DATA_0_27, n4339 );
nand U7786 ( n8311, n913, n914 );
and U7787 ( n914, n915, n916 );
nor U7788 ( n913, n918, n919 );
nand U7789 ( n916, DATA_0_28, n4339 );
nand U7790 ( n8306, n923, n924 );
and U7791 ( n924, n925, n926 );
nor U7792 ( n923, n928, n929 );
nand U7793 ( n926, DATA_0_29, n4339 );
nand U7794 ( n8301, n933, n934 );
and U7795 ( n934, n935, n936 );
nor U7796 ( n933, n938, n939 );
nand U7797 ( n936, DATA_0_30, n4339 );
nand U7798 ( n982, n384, n385 );
nor U7799 ( n385, n386, n387 );
nor U7800 ( n384, n389, n390 );
and U7801 ( n387, n4448, CRC_OUT_9_9 );
nand U7802 ( n987, n373, n374 );
nor U7803 ( n374, n375, n376 );
nor U7804 ( n373, n378, n379 );
and U7805 ( n376, n4448, CRC_OUT_9_8 );
nand U7806 ( n992, n362, n363 );
nor U7807 ( n363, n364, n365 );
nor U7808 ( n362, n367, n368 );
and U7809 ( n365, n4448, CRC_OUT_9_7 );
nand U7810 ( n997, n348, n349 );
nor U7811 ( n349, n350, n351 );
nor U7812 ( n348, n354, n355 );
and U7813 ( n351, n4448, CRC_OUT_9_6 );
not U7814 ( n4471, TM0 );
xor U7815 ( n299, n369, n370 );
xnor U7816 ( n369, WX757, n371 );
xor U7817 ( n370, WX693, TM0 );
xor U7818 ( n371, WX885, WX821 );
xor U7819 ( n297, n357, n358 );
xnor U7820 ( n357, WX759, n359 );
xor U7821 ( n358, WX695, TM0 );
xor U7822 ( n359, WX887, WX823 );
xor U7823 ( DATA_9_6, n4298, n297 );
nand U7824 ( n4298, TM0, WX535 );
xor U7825 ( DATA_9_7, n4299, n299 );
nand U7826 ( n4299, TM0, WX533 );
and U7827 ( n3992, n4449, CRC_OUT_8_22 );
and U7828 ( n4008, n4449, CRC_OUT_8_23 );
and U7829 ( n4024, n4449, CRC_OUT_8_24 );
and U7830 ( n4040, n4449, CRC_OUT_8_25 );
and U7831 ( n667, n4446, CRC_OUT_9_31 );
and U7832 ( n4143, n4448, CRC_OUT_8_31 );
and U7833 ( n3634, n4451, CRC_OUT_7_31 );
and U7834 ( n3199, n4453, CRC_OUT_6_31 );
and U7835 ( n1842, n4440, CRC_OUT_3_31 );
and U7836 ( n1410, n4443, CRC_OUT_2_31 );
xor U7837 ( n285, n4203, n4204 );
xnor U7838 ( n4203, WX771, n4205 );
xor U7839 ( n4204, WX707, TM0 );
xor U7840 ( n4205, WX899, WX835 );
xor U7841 ( n287, n4217, n4218 );
xnor U7842 ( n4217, WX769, n4219 );
xor U7843 ( n4218, WX705, TM0 );
xor U7844 ( n4219, WX897, WX833 );
xor U7845 ( n289, n4230, n4232 );
xnor U7846 ( n4230, WX767, n4233 );
xor U7847 ( n4232, WX703, TM0 );
xor U7848 ( n4233, WX895, WX831 );
xor U7849 ( n291, n4244, n4245 );
xnor U7850 ( n4244, WX765, n4247 );
xor U7851 ( n4245, WX701, TM0 );
xor U7852 ( n4247, WX893, WX829 );
xor U7853 ( n293, n4258, n4259 );
xnor U7854 ( n4258, WX763, n4260 );
xor U7855 ( n4259, WX699, TM0 );
xor U7856 ( n4260, WX891, WX827 );
xor U7857 ( n295, n4274, n4275 );
xnor U7858 ( n4274, WX761, n4277 );
xor U7859 ( n4275, WX697, TM0 );
xor U7860 ( n4277, WX889, WX825 );
xor U7861 ( n315, n457, n458 );
xnor U7862 ( n457, WX741, n459 );
xor U7863 ( n458, WX677, TM0 );
xor U7864 ( n459, WX869, WX805 );
xor U7865 ( n313, n446, n447 );
xnor U7866 ( n446, WX743, n448 );
xor U7867 ( n447, WX679, TM0 );
xor U7868 ( n448, WX871, WX807 );
xor U7869 ( n311, n435, n436 );
xnor U7870 ( n435, WX745, n437 );
xor U7871 ( n436, WX681, TM0 );
xor U7872 ( n437, WX873, WX809 );
xor U7873 ( n309, n424, n425 );
xnor U7874 ( n424, WX747, n426 );
xor U7875 ( n425, WX683, TM0 );
xor U7876 ( n426, WX875, WX811 );
xor U7877 ( n307, n413, n414 );
xnor U7878 ( n413, WX749, n415 );
xor U7879 ( n414, WX685, TM0 );
xor U7880 ( n415, WX877, WX813 );
xor U7881 ( n305, n402, n403 );
xnor U7882 ( n402, WX751, n404 );
xor U7883 ( n403, WX687, TM0 );
xor U7884 ( n404, WX879, WX815 );
xor U7885 ( n303, n391, n392 );
xnor U7886 ( n391, WX753, n393 );
xor U7887 ( n392, WX689, TM0 );
xor U7888 ( n393, WX881, WX817 );
xor U7889 ( n301, n380, n381 );
xnor U7890 ( n380, WX755, n382 );
xor U7891 ( n381, WX691, TM0 );
xor U7892 ( n382, WX883, WX819 );
xor U7893 ( DATA_9_0, n4301, n285 );
nand U7894 ( n4301, TM0, WX547 );
xor U7895 ( DATA_9_1, n4302, n287 );
nand U7896 ( n4302, TM0, WX545 );
xor U7897 ( DATA_9_2, n4303, n289 );
nand U7898 ( n4303, TM0, WX543 );
xor U7899 ( DATA_9_3, n4305, n291 );
nand U7900 ( n4305, TM0, WX541 );
xor U7901 ( DATA_9_4, n4306, n293 );
nand U7902 ( n4306, TM0, WX539 );
xor U7903 ( DATA_9_5, n4307, n295 );
nand U7904 ( n4307, TM0, WX537 );
xor U7905 ( DATA_9_8, n4309, n301 );
nand U7906 ( n4309, TM0, WX531 );
xor U7907 ( DATA_9_9, n4310, n303 );
nand U7908 ( n4310, TM0, WX529 );
xor U7909 ( DATA_9_10, n4311, n305 );
nand U7910 ( n4311, TM0, WX527 );
xor U7911 ( DATA_9_11, n4313, n307 );
nand U7912 ( n4313, TM0, WX525 );
xor U7913 ( DATA_9_12, n4314, n309 );
nand U7914 ( n4314, TM0, WX523 );
xor U7915 ( DATA_9_13, n4315, n311 );
nand U7916 ( n4315, TM0, WX521 );
xor U7917 ( DATA_9_14, n4317, n313 );
nand U7918 ( n4317, TM0, WX519 );
xor U7919 ( DATA_9_15, n4318, n315 );
nand U7920 ( n4318, TM0, WX517 );
nand U7921 ( n817, CRC_OUT_1_17, n4439 );
nand U7922 ( n825, CRC_OUT_1_18, n4439 );
nand U7923 ( n841, CRC_OUT_1_20, n4439 );
nand U7924 ( n849, CRC_OUT_1_21, n4439 );
nand U7925 ( n865, CRC_OUT_1_23, n4439 );
nand U7926 ( n875, CRC_OUT_1_24, n4439 );
nand U7927 ( n925, CRC_OUT_1_29, n4439 );
nand U7928 ( n935, CRC_OUT_1_30, n4439 );
and U7929 ( n2736, n4456, CRC_OUT_5_31 );
and U7930 ( n2304, n4458, CRC_OUT_4_31 );
nand U7931 ( n946, CRC_OUT_1_31, n4438 );
nand U7932 ( n678, CRC_OUT_1_0, n4438 );
nand U7933 ( n687, CRC_OUT_1_1, n4437 );
nand U7934 ( n695, CRC_OUT_1_2, n4438 );
nand U7935 ( n711, CRC_OUT_1_4, n4437 );
nand U7936 ( n719, CRC_OUT_1_5, n4437 );
nand U7937 ( n727, CRC_OUT_1_6, n4438 );
nand U7938 ( n736, CRC_OUT_1_7, n4437 );
nand U7939 ( n744, CRC_OUT_1_8, n4438 );
nand U7940 ( n752, CRC_OUT_1_9, n4438 );
nand U7941 ( n768, CRC_OUT_1_11, n4438 );
nand U7942 ( n776, CRC_OUT_1_12, n4437 );
nand U7943 ( n784, CRC_OUT_1_13, n4437 );
nand U7944 ( n792, CRC_OUT_1_14, n4438 );
nand U7945 ( n808, CRC_OUT_1_16, n4437 );
nand U7946 ( n833, CRC_OUT_1_19, n4437 );
nand U7947 ( n857, CRC_OUT_1_22, n4437 );
nand U7948 ( n885, CRC_OUT_1_25, n4438 );
nand U7949 ( n895, CRC_OUT_1_26, n4437 );
nand U7950 ( n905, CRC_OUT_1_27, n4437 );
nand U7951 ( n915, CRC_OUT_1_28, n4438 );
nand U7952 ( n703, CRC_OUT_1_3, n4438 );
nand U7953 ( n760, CRC_OUT_1_10, n4437 );
nand U7954 ( n800, CRC_OUT_1_15, n4438 );
buf U7955 ( n4495, RESET );
nand U7956 ( n949, DATA_0_31, n4339 );
xor U7957 ( n665, n4145, n4147 );
xnor U7958 ( n4145, WX2002, n4148 );
xor U7959 ( n4147, WX1938, TM1 );
xor U7960 ( n4148, WX2130, WX2066 );
xor U7961 ( n3636, n4139, n4140 );
xnor U7962 ( n4139, WX3295, n4142 );
xor U7963 ( n4140, WX3231, TM1 );
xor U7964 ( n4142, WX3423, WX3359 );
xor U7965 ( n3201, n3631, n3632 );
xnor U7966 ( n3631, WX4588, n3633 );
xor U7967 ( n3632, WX4524, TM1 );
xor U7968 ( n3633, WX4716, WX4652 );
xor U7969 ( n2739, n3195, n3196 );
xnor U7970 ( n3195, WX5881, n3197 );
xor U7971 ( n3196, WX5817, TM1 );
xor U7972 ( n3197, WX6009, WX5945 );
xor U7973 ( n2307, n2732, n2734 );
xnor U7974 ( n2732, WX7174, n2735 );
xor U7975 ( n2734, WX7110, TM1 );
xor U7976 ( n2735, WX7302, WX7238 );
xor U7977 ( n1844, n2301, n2302 );
xnor U7978 ( n2301, WX8467, n2303 );
xor U7979 ( n2302, WX8403, TM1 );
xor U7980 ( n2303, WX8595, WX8531 );
xor U7981 ( n465, n3902, n3903 );
xnor U7982 ( n3902, WX2032, n3904 );
xor U7983 ( n3903, WX1968, TM1 );
xor U7984 ( n3904, WX2160, WX2096 );
xor U7985 ( n476, n3918, n3919 );
xnor U7986 ( n3918, WX2030, n3920 );
xor U7987 ( n3919, WX1966, TM1 );
xor U7988 ( n3920, WX2158, WX2094 );
xor U7989 ( n487, n3934, n3935 );
xnor U7990 ( n3934, WX2028, n3937 );
xor U7991 ( n3935, WX1964, TM1 );
xor U7992 ( n3937, WX2156, WX2092 );
xor U7993 ( n498, n3950, n3952 );
xnor U7994 ( n3950, WX2026, n3953 );
xor U7995 ( n3952, WX1962, TM1 );
xor U7996 ( n3953, WX2154, WX2090 );
xor U7997 ( n509, n3967, n3968 );
xnor U7998 ( n3967, WX2024, n3969 );
xor U7999 ( n3968, WX1960, TM1 );
xor U8000 ( n3969, WX2152, WX2088 );
xor U8001 ( n520, n3983, n3984 );
xnor U8002 ( n3983, WX2022, n3985 );
xor U8003 ( n3984, WX1958, TM1 );
xor U8004 ( n3985, WX2150, WX2086 );
xor U8005 ( n531, n3999, n4000 );
xnor U8006 ( n3999, WX2020, n4002 );
xor U8007 ( n4000, WX1956, TM1 );
xor U8008 ( n4002, WX2148, WX2084 );
xor U8009 ( n542, n4015, n4017 );
xnor U8010 ( n4015, WX2018, n4018 );
xor U8011 ( n4017, WX1954, TM1 );
xor U8012 ( n4018, WX2146, WX2082 );
xor U8013 ( n553, n4032, n4033 );
xnor U8014 ( n4032, WX2016, n4034 );
xor U8015 ( n4033, WX1952, TM1 );
xor U8016 ( n4034, WX2144, WX2080 );
xor U8017 ( n575, n4048, n4049 );
xnor U8018 ( n4048, WX2014, n4050 );
xor U8019 ( n4049, WX1950, TM1 );
xor U8020 ( n4050, WX2142, WX2078 );
xor U8021 ( n600, n4064, n4065 );
xnor U8022 ( n4064, WX2012, n4067 );
xor U8023 ( n4065, WX1948, TM1 );
xor U8024 ( n4067, WX2140, WX2076 );
xor U8025 ( n621, n4080, n4082 );
xnor U8026 ( n4080, WX2010, n4083 );
xor U8027 ( n4082, WX1946, TM1 );
xor U8028 ( n4083, WX2138, WX2074 );
xor U8029 ( n632, n4097, n4098 );
xnor U8030 ( n4097, WX2008, n4099 );
xor U8031 ( n4098, WX1944, TM1 );
xor U8032 ( n4099, WX2136, WX2072 );
xor U8033 ( n643, n4113, n4114 );
xnor U8034 ( n4113, WX2006, n4115 );
xor U8035 ( n4114, WX1942, TM1 );
xor U8036 ( n4115, WX2134, WX2070 );
xor U8037 ( n654, n4129, n4130 );
xnor U8038 ( n4129, WX2004, n4132 );
xor U8039 ( n4130, WX1940, TM1 );
xor U8040 ( n4132, WX2132, WX2068 );
xor U8041 ( n3463, n3895, n3897 );
xnor U8042 ( n3895, WX3325, n3898 );
xor U8043 ( n3897, WX3261, TM1 );
xor U8044 ( n3898, WX3453, WX3389 );
xor U8045 ( n3478, n3912, n3913 );
xnor U8046 ( n3912, WX3323, n3914 );
xor U8047 ( n3913, WX3259, TM1 );
xor U8048 ( n3914, WX3451, WX3387 );
xor U8049 ( n3493, n3928, n3929 );
xnor U8050 ( n3928, WX3321, n3930 );
xor U8051 ( n3929, WX3257, TM1 );
xor U8052 ( n3930, WX3449, WX3385 );
xor U8053 ( n3504, n3944, n3945 );
xnor U8054 ( n3944, WX3319, n3947 );
xor U8055 ( n3945, WX3255, TM1 );
xor U8056 ( n3947, WX3447, WX3383 );
xor U8057 ( n3515, n3960, n3962 );
xnor U8058 ( n3960, WX3317, n3963 );
xor U8059 ( n3962, WX3253, TM1 );
xor U8060 ( n3963, WX3445, WX3381 );
xor U8061 ( n3526, n3977, n3978 );
xnor U8062 ( n3977, WX3315, n3979 );
xor U8063 ( n3978, WX3251, TM1 );
xor U8064 ( n3979, WX3443, WX3379 );
xor U8065 ( n3537, n3993, n3994 );
xnor U8066 ( n3993, WX3313, n3995 );
xor U8067 ( n3994, WX3249, TM1 );
xor U8068 ( n3995, WX3441, WX3377 );
xor U8069 ( n3548, n4009, n4010 );
xnor U8070 ( n4009, WX3311, n4012 );
xor U8071 ( n4010, WX3247, TM1 );
xor U8072 ( n4012, WX3439, WX3375 );
xor U8073 ( n3559, n4025, n4027 );
xnor U8074 ( n4025, WX3309, n4028 );
xor U8075 ( n4027, WX3245, TM1 );
xor U8076 ( n4028, WX3437, WX3373 );
xor U8077 ( n3570, n4042, n4043 );
xnor U8078 ( n4042, WX3307, n4044 );
xor U8079 ( n4043, WX3243, TM1 );
xor U8080 ( n4044, WX3435, WX3371 );
xor U8081 ( n3581, n4058, n4059 );
xnor U8082 ( n4058, WX3305, n4060 );
xor U8083 ( n4059, WX3241, TM1 );
xor U8084 ( n4060, WX3433, WX3369 );
xor U8085 ( n3592, n4074, n4075 );
xnor U8086 ( n4074, WX3303, n4077 );
xor U8087 ( n4075, WX3239, TM1 );
xor U8088 ( n4077, WX3431, WX3367 );
xor U8089 ( n3603, n4090, n4092 );
xnor U8090 ( n4090, WX3301, n4093 );
xor U8091 ( n4092, WX3237, TM1 );
xor U8092 ( n4093, WX3429, WX3365 );
xor U8093 ( n3614, n4107, n4108 );
xnor U8094 ( n4107, WX3299, n4109 );
xor U8095 ( n4108, WX3235, TM1 );
xor U8096 ( n4109, WX3427, WX3363 );
xor U8097 ( n3625, n4123, n4124 );
xnor U8098 ( n4123, WX3297, n4125 );
xor U8099 ( n4124, WX3233, TM1 );
xor U8100 ( n4125, WX3425, WX3361 );
xor U8101 ( n2995, n3457, n3458 );
xnor U8102 ( n3457, WX4618, n3459 );
xor U8103 ( n3458, WX4554, TM1 );
xor U8104 ( n3459, WX4746, WX4682 );
xor U8105 ( n3009, n3471, n3473 );
xnor U8106 ( n3471, WX4616, n3474 );
xor U8107 ( n3473, WX4552, TM1 );
xor U8108 ( n3474, WX4744, WX4680 );
xor U8109 ( n3022, n3486, n3487 );
xnor U8110 ( n3486, WX4614, n3489 );
xor U8111 ( n3487, WX4550, TM1 );
xor U8112 ( n3489, WX4742, WX4678 );
xor U8113 ( n3036, n3499, n3500 );
xnor U8114 ( n3499, WX4612, n3501 );
xor U8115 ( n3500, WX4548, TM1 );
xor U8116 ( n3501, WX4740, WX4676 );
xor U8117 ( n3050, n3510, n3511 );
xnor U8118 ( n3510, WX4610, n3512 );
xor U8119 ( n3511, WX4546, TM1 );
xor U8120 ( n3512, WX4738, WX4674 );
xor U8121 ( n3064, n3521, n3522 );
xnor U8122 ( n3521, WX4608, n3523 );
xor U8123 ( n3522, WX4544, n4472 );
xor U8124 ( n3523, WX4736, WX4672 );
xor U8125 ( n3077, n3532, n3533 );
xnor U8126 ( n3532, WX4606, n3534 );
xor U8127 ( n3533, WX4542, n4472 );
xor U8128 ( n3534, WX4734, WX4670 );
xor U8129 ( n3091, n3543, n3544 );
xnor U8130 ( n3543, WX4604, n3545 );
xor U8131 ( n3544, WX4540, n4472 );
xor U8132 ( n3545, WX4732, WX4668 );
xor U8133 ( n3105, n3554, n3555 );
xnor U8134 ( n3554, WX4602, n3556 );
xor U8135 ( n3555, WX4538, n4472 );
xor U8136 ( n3556, WX4730, WX4666 );
xor U8137 ( n3119, n3565, n3566 );
xnor U8138 ( n3565, WX4600, n3567 );
xor U8139 ( n3566, WX4536, n4472 );
xor U8140 ( n3567, WX4728, WX4664 );
xor U8141 ( n3132, n3576, n3577 );
xnor U8142 ( n3576, WX4598, n3578 );
xor U8143 ( n3577, WX4534, n4472 );
xor U8144 ( n3578, WX4726, WX4662 );
xor U8145 ( n3146, n3587, n3588 );
xnor U8146 ( n3587, WX4596, n3589 );
xor U8147 ( n3588, WX4532, n4472 );
xor U8148 ( n3589, WX4724, WX4660 );
xor U8149 ( n3160, n3598, n3599 );
xnor U8150 ( n3598, WX4594, n3600 );
xor U8151 ( n3599, WX4530, TM1 );
xor U8152 ( n3600, WX4722, WX4658 );
xor U8153 ( n3174, n3609, n3610 );
xnor U8154 ( n3609, WX4592, n3611 );
xor U8155 ( n3610, WX4528, TM1 );
xor U8156 ( n3611, WX4720, WX4656 );
xor U8157 ( n3187, n3620, n3621 );
xnor U8158 ( n3620, WX4590, n3622 );
xor U8159 ( n3621, WX4526, TM1 );
xor U8160 ( n3622, WX4718, WX4654 );
xor U8161 ( n2570, n2989, n2990 );
xnor U8162 ( n2989, WX5911, n2991 );
xor U8163 ( n2990, WX5847, TM1 );
xor U8164 ( n2991, WX6039, WX5975 );
xor U8165 ( n2581, n3002, n3004 );
xnor U8166 ( n3002, WX5909, n3005 );
xor U8167 ( n3004, WX5845, TM1 );
xor U8168 ( n3005, WX6037, WX5973 );
xor U8169 ( n2592, n3016, n3017 );
xnor U8170 ( n3016, WX5907, n3019 );
xor U8171 ( n3017, WX5843, TM1 );
xor U8172 ( n3019, WX6035, WX5971 );
xor U8173 ( n2603, n3030, n3031 );
xnor U8174 ( n3030, WX5905, n3032 );
xor U8175 ( n3031, WX5841, TM1 );
xor U8176 ( n3032, WX6033, WX5969 );
xor U8177 ( n2614, n3044, n3045 );
xnor U8178 ( n3044, WX5903, n3046 );
xor U8179 ( n3045, WX5839, TM1 );
xor U8180 ( n3046, WX6031, WX5967 );
xor U8181 ( n2625, n3057, n3059 );
xnor U8182 ( n3057, WX5901, n3060 );
xor U8183 ( n3059, WX5837, TM1 );
xor U8184 ( n3060, WX6029, WX5965 );
xor U8185 ( n2636, n3071, n3072 );
xnor U8186 ( n3071, WX5899, n3074 );
xor U8187 ( n3072, WX5835, TM1 );
xor U8188 ( n3074, WX6027, WX5963 );
xor U8189 ( n2647, n3085, n3086 );
xnor U8190 ( n3085, WX5897, n3087 );
xor U8191 ( n3086, WX5833, TM1 );
xor U8192 ( n3087, WX6025, WX5961 );
xor U8193 ( n2658, n3099, n3100 );
xnor U8194 ( n3099, WX5895, n3101 );
xor U8195 ( n3100, WX5831, TM1 );
xor U8196 ( n3101, WX6023, WX5959 );
xor U8197 ( n2669, n3112, n3114 );
xnor U8198 ( n3112, WX5893, n3115 );
xor U8199 ( n3114, WX5829, TM1 );
xor U8200 ( n3115, WX6021, WX5957 );
xor U8201 ( n2680, n3126, n3127 );
xnor U8202 ( n3126, WX5891, n3129 );
xor U8203 ( n3127, WX5827, TM1 );
xor U8204 ( n3129, WX6019, WX5955 );
xor U8205 ( n2691, n3140, n3141 );
xnor U8206 ( n3140, WX5889, n3142 );
xor U8207 ( n3141, WX5825, TM1 );
xor U8208 ( n3142, WX6017, WX5953 );
xor U8209 ( n2702, n3154, n3155 );
xnor U8210 ( n3154, WX5887, n3156 );
xor U8211 ( n3155, WX5823, TM1 );
xor U8212 ( n3156, WX6015, WX5951 );
xor U8213 ( n2713, n3167, n3169 );
xnor U8214 ( n3167, WX5885, n3170 );
xor U8215 ( n3169, WX5821, TM1 );
xor U8216 ( n3170, WX6013, WX5949 );
xor U8217 ( n2725, n3181, n3182 );
xnor U8218 ( n3181, WX5883, n3184 );
xor U8219 ( n3182, WX5819, TM1 );
xor U8220 ( n3184, WX6011, WX5947 );
xor U8221 ( n2101, n2565, n2566 );
xnor U8222 ( n2565, WX7204, n2567 );
xor U8223 ( n2566, WX7140, TM1 );
xor U8224 ( n2567, WX7332, WX7268 );
xor U8225 ( n2114, n2576, n2577 );
xnor U8226 ( n2576, WX7202, n2578 );
xor U8227 ( n2577, WX7138, TM1 );
xor U8228 ( n2578, WX7330, WX7266 );
xor U8229 ( n2128, n2587, n2588 );
xnor U8230 ( n2587, WX7200, n2589 );
xor U8231 ( n2588, WX7136, n4472 );
xor U8232 ( n2589, WX7328, WX7264 );
xor U8233 ( n2142, n2598, n2599 );
xnor U8234 ( n2598, WX7198, n2600 );
xor U8235 ( n2599, WX7134, TM1 );
xor U8236 ( n2600, WX7326, WX7262 );
xor U8237 ( n2156, n2609, n2610 );
xnor U8238 ( n2609, WX7196, n2611 );
xor U8239 ( n2610, WX7132, TM1 );
xor U8240 ( n2611, WX7324, WX7260 );
xor U8241 ( n2169, n2620, n2621 );
xnor U8242 ( n2620, WX7194, n2622 );
xor U8243 ( n2621, WX7130, TM1 );
xor U8244 ( n2622, WX7322, WX7258 );
xor U8245 ( n2183, n2631, n2632 );
xnor U8246 ( n2631, WX7192, n2633 );
xor U8247 ( n2632, WX7128, TM1 );
xor U8248 ( n2633, WX7320, WX7256 );
xor U8249 ( n2197, n2642, n2643 );
xnor U8250 ( n2642, WX7190, n2644 );
xor U8251 ( n2643, WX7126, TM1 );
xor U8252 ( n2644, WX7318, WX7254 );
xor U8253 ( n2211, n2653, n2654 );
xnor U8254 ( n2653, WX7188, n2655 );
xor U8255 ( n2654, WX7124, TM1 );
xor U8256 ( n2655, WX7316, WX7252 );
xor U8257 ( n2224, n2664, n2665 );
xnor U8258 ( n2664, WX7186, n2666 );
xor U8259 ( n2665, WX7122, TM1 );
xor U8260 ( n2666, WX7314, WX7250 );
xor U8261 ( n2238, n2675, n2676 );
xnor U8262 ( n2675, WX7184, n2677 );
xor U8263 ( n2676, WX7120, TM1 );
xor U8264 ( n2677, WX7312, WX7248 );
xor U8265 ( n2252, n2686, n2687 );
xnor U8266 ( n2686, WX7182, n2688 );
xor U8267 ( n2687, WX7118, TM1 );
xor U8268 ( n2688, WX7310, WX7246 );
xor U8269 ( n2266, n2697, n2698 );
xnor U8270 ( n2697, WX7180, n2699 );
xor U8271 ( n2698, WX7116, TM1 );
xor U8272 ( n2699, WX7308, WX7244 );
xor U8273 ( n2279, n2708, n2709 );
xnor U8274 ( n2708, WX7178, n2710 );
xor U8275 ( n2709, WX7114, TM1 );
xor U8276 ( n2710, WX7306, WX7242 );
xor U8277 ( n2293, n2719, n2720 );
xnor U8278 ( n2719, WX7176, n2721 );
xor U8279 ( n2720, WX7112, TM1 );
xor U8280 ( n2721, WX7304, WX7240 );
xor U8281 ( n1669, n2094, n2096 );
xnor U8282 ( n2094, WX8497, n2097 );
xor U8283 ( n2096, WX8433, n4472 );
xor U8284 ( n2097, WX8625, WX8561 );
xor U8285 ( n1680, n2108, n2109 );
xnor U8286 ( n2108, WX8495, n2111 );
xor U8287 ( n2109, WX8431, n4472 );
xor U8288 ( n2111, WX8623, WX8559 );
xor U8289 ( n1691, n2122, n2123 );
xnor U8290 ( n2122, WX8493, n2124 );
xor U8291 ( n2123, WX8429, n4472 );
xor U8292 ( n2124, WX8621, WX8557 );
xor U8293 ( n1702, n2136, n2137 );
xnor U8294 ( n2136, WX8491, n2138 );
xor U8295 ( n2137, WX8427, n4472 );
xor U8296 ( n2138, WX8619, WX8555 );
xor U8297 ( n1713, n2149, n2151 );
xnor U8298 ( n2149, WX8489, n2152 );
xor U8299 ( n2151, WX8425, n4472 );
xor U8300 ( n2152, WX8617, WX8553 );
xor U8301 ( n1724, n2163, n2164 );
xnor U8302 ( n2163, WX8487, n2166 );
xor U8303 ( n2164, WX8423, TM1 );
xor U8304 ( n2166, WX8615, WX8551 );
xor U8305 ( n1735, n2177, n2178 );
xnor U8306 ( n2177, WX8485, n2179 );
xor U8307 ( n2178, WX8421, TM1 );
xor U8308 ( n2179, WX8613, WX8549 );
xor U8309 ( n1746, n2191, n2192 );
xnor U8310 ( n2191, WX8483, n2193 );
xor U8311 ( n2192, WX8419, TM1 );
xor U8312 ( n2193, WX8611, WX8547 );
xor U8313 ( n1757, n2204, n2206 );
xnor U8314 ( n2204, WX8481, n2207 );
xor U8315 ( n2206, WX8417, TM1 );
xor U8316 ( n2207, WX8609, WX8545 );
xor U8317 ( n1768, n2218, n2219 );
xnor U8318 ( n2218, WX8479, n2221 );
xor U8319 ( n2219, WX8415, TM1 );
xor U8320 ( n2221, WX8607, WX8543 );
xor U8321 ( n1779, n2232, n2233 );
xnor U8322 ( n2232, WX8477, n2234 );
xor U8323 ( n2233, WX8413, TM1 );
xor U8324 ( n2234, WX8605, WX8541 );
xor U8325 ( n1790, n2246, n2247 );
xnor U8326 ( n2246, WX8475, n2248 );
xor U8327 ( n2247, WX8411, TM1 );
xor U8328 ( n2248, WX8603, WX8539 );
xor U8329 ( n1803, n2259, n2261 );
xnor U8330 ( n2259, WX8473, n2262 );
xor U8331 ( n2261, WX8409, TM1 );
xor U8332 ( n2262, WX8601, WX8537 );
xor U8333 ( n1817, n2273, n2274 );
xnor U8334 ( n2273, WX8471, n2276 );
xor U8335 ( n2274, WX8407, TM1 );
xor U8336 ( n2276, WX8599, WX8535 );
xor U8337 ( n1831, n2287, n2288 );
xnor U8338 ( n2287, WX8469, n2289 );
xor U8339 ( n2288, WX8405, TM1 );
xor U8340 ( n2289, WX8597, WX8533 );
xor U8341 ( n1413, n1838, n1839 );
xnor U8342 ( n1838, WX9760, n1841 );
xor U8343 ( n1839, WX9696, TM1 );
xor U8344 ( n1841, WX9888, WX9824 );
xor U8345 ( n1206, n1664, n1665 );
xnor U8346 ( n1664, WX9790, n1666 );
xor U8347 ( n1665, WX9726, TM1 );
xor U8348 ( n1666, WX9918, WX9854 );
xor U8349 ( n1220, n1675, n1676 );
xnor U8350 ( n1675, WX9788, n1677 );
xor U8351 ( n1676, WX9724, TM1 );
xor U8352 ( n1677, WX9916, WX9852 );
xor U8353 ( n1234, n1686, n1687 );
xnor U8354 ( n1686, WX9786, n1688 );
xor U8355 ( n1687, WX9722, TM1 );
xor U8356 ( n1688, WX9914, WX9850 );
xor U8357 ( n1248, n1697, n1698 );
xnor U8358 ( n1697, WX9784, n1699 );
xor U8359 ( n1698, WX9720, n4472 );
xor U8360 ( n1699, WX9912, WX9848 );
xor U8361 ( n1261, n1708, n1709 );
xnor U8362 ( n1708, WX9782, n1710 );
xor U8363 ( n1709, WX9718, TM1 );
xor U8364 ( n1710, WX9910, WX9846 );
xor U8365 ( n1275, n1719, n1720 );
xnor U8366 ( n1719, WX9780, n1721 );
xor U8367 ( n1720, WX9716, TM1 );
xor U8368 ( n1721, WX9908, WX9844 );
xor U8369 ( n1289, n1730, n1731 );
xnor U8370 ( n1730, WX9778, n1732 );
xor U8371 ( n1731, WX9714, n4472 );
xor U8372 ( n1732, WX9906, WX9842 );
xor U8373 ( n1303, n1741, n1742 );
xnor U8374 ( n1741, WX9776, n1743 );
xor U8375 ( n1742, WX9712, TM1 );
xor U8376 ( n1743, WX9904, WX9840 );
xor U8377 ( n1316, n1752, n1753 );
xnor U8378 ( n1752, WX9774, n1754 );
xor U8379 ( n1753, WX9710, TM1 );
xor U8380 ( n1754, WX9902, WX9838 );
xor U8381 ( n1330, n1763, n1764 );
xnor U8382 ( n1763, WX9772, n1765 );
xor U8383 ( n1764, WX9708, TM1 );
xor U8384 ( n1765, WX9900, WX9836 );
xor U8385 ( n1344, n1774, n1775 );
xnor U8386 ( n1774, WX9770, n1776 );
xor U8387 ( n1775, WX9706, TM1 );
xor U8388 ( n1776, WX9898, WX9834 );
xor U8389 ( n1358, n1785, n1786 );
xnor U8390 ( n1785, WX9768, n1787 );
xor U8391 ( n1786, WX9704, TM1 );
xor U8392 ( n1787, WX9896, WX9832 );
xor U8393 ( n1371, n1797, n1798 );
xnor U8394 ( n1797, WX9766, n1799 );
xor U8395 ( n1798, WX9702, TM1 );
xor U8396 ( n1799, WX9894, WX9830 );
xor U8397 ( n1385, n1811, n1812 );
xnor U8398 ( n1811, WX9764, n1813 );
xor U8399 ( n1812, WX9700, TM1 );
xor U8400 ( n1813, WX9892, WX9828 );
xor U8401 ( n1399, n1824, n1826 );
xnor U8402 ( n1824, WX9762, n1827 );
xor U8403 ( n1826, WX9698, n4472 );
xor U8404 ( n1827, WX9890, WX9826 );
xor U8405 ( n812, n1200, n1201 );
xnor U8406 ( n1200, WX11083, n1203 );
xor U8407 ( n1201, WX11019, TM1 );
xor U8408 ( n1203, WX11211, WX11147 );
xor U8409 ( n821, n1214, n1215 );
xnor U8410 ( n1214, WX11081, n1216 );
xor U8411 ( n1215, WX11017, TM1 );
xor U8412 ( n1216, WX11209, WX11145 );
xor U8413 ( n829, n1228, n1229 );
xnor U8414 ( n1228, WX11079, n1230 );
xor U8415 ( n1229, WX11015, TM1 );
xor U8416 ( n1230, WX11207, WX11143 );
xor U8417 ( n837, n1241, n1243 );
xnor U8418 ( n1241, WX11077, n1244 );
xor U8419 ( n1243, WX11013, TM1 );
xor U8420 ( n1244, WX11205, WX11141 );
xor U8421 ( n845, n1255, n1256 );
xnor U8422 ( n1255, WX11075, n1258 );
xor U8423 ( n1256, WX11011, TM1 );
xor U8424 ( n1258, WX11203, WX11139 );
xor U8425 ( n853, n1269, n1270 );
xnor U8426 ( n1269, WX11073, n1271 );
xor U8427 ( n1270, WX11009, TM1 );
xor U8428 ( n1271, WX11201, WX11137 );
xor U8429 ( n861, n1283, n1284 );
xnor U8430 ( n1283, WX11071, n1285 );
xor U8431 ( n1284, WX11007, TM1 );
xor U8432 ( n1285, WX11199, WX11135 );
xor U8433 ( n870, n1296, n1298 );
xnor U8434 ( n1296, WX11069, n1299 );
xor U8435 ( n1298, WX11005, TM1 );
xor U8436 ( n1299, WX11197, WX11133 );
xor U8437 ( n880, n1310, n1311 );
xnor U8438 ( n1310, WX11067, n1313 );
xor U8439 ( n1311, WX11003, n4472 );
xor U8440 ( n1313, WX11195, WX11131 );
xor U8441 ( n890, n1324, n1325 );
xnor U8442 ( n1324, WX11065, n1326 );
xor U8443 ( n1325, WX11001, TM1 );
xor U8444 ( n1326, WX11193, WX11129 );
xor U8445 ( n900, n1338, n1339 );
xnor U8446 ( n1338, WX11063, n1340 );
xor U8447 ( n1339, WX10999, TM1 );
xor U8448 ( n1340, WX11191, WX11127 );
xor U8449 ( n910, n1351, n1353 );
xnor U8450 ( n1351, WX11061, n1354 );
xor U8451 ( n1353, WX10997, TM1 );
xor U8452 ( n1354, WX11189, WX11125 );
xor U8453 ( n920, n1365, n1366 );
xnor U8454 ( n1365, WX11059, n1368 );
xor U8455 ( n1366, WX10995, TM1 );
xor U8456 ( n1368, WX11187, WX11123 );
xor U8457 ( n930, n1379, n1380 );
xnor U8458 ( n1379, WX11057, n1381 );
xor U8459 ( n1380, WX10993, n4472 );
xor U8460 ( n1381, WX11185, WX11121 );
xor U8461 ( n940, n1393, n1394 );
xnor U8462 ( n1393, WX11055, n1395 );
xor U8463 ( n1394, WX10991, TM1 );
xor U8464 ( n1395, WX11183, WX11119 );
xor U8465 ( n948, n1406, n1408 );
xnor U8466 ( n1406, WX11053, n1409 );
xor U8467 ( n1408, WX10989, n4472 );
xor U8468 ( n1409, WX11181, WX11117 );
nand U8469 ( n672, n4587, WX547 );
nand U8470 ( n673, n4587, WX545 );
nand U8471 ( n674, n4587, WX543 );
nand U8472 ( n606, n4587, WX495 );
nand U8473 ( n559, n4587, WX499 );
nand U8474 ( n548, n4587, WX501 );
nand U8475 ( n537, n4587, WX503 );
nand U8476 ( n526, n4587, WX505 );
nand U8477 ( n515, n4587, WX507 );
nand U8478 ( n449, n4587, WX519 );
nand U8479 ( n427, n4587, WX523 );
nand U8480 ( n405, n4587, WX527 );
nand U8481 ( n394, n4587, WX529 );
nand U8482 ( n649, n4585, WX489 );
nand U8483 ( n482, n4585, WX513 );
nand U8484 ( n814, n4586, WX537 );
nand U8485 ( n660, n4586, WX487 );
nand U8486 ( n638, n4586, WX491 );
nand U8487 ( n627, n4586, WX493 );
nand U8488 ( n581, n4586, WX497 );
nand U8489 ( n504, n4586, WX509 );
nand U8490 ( n493, n4586, WX511 );
nand U8491 ( n471, n4586, WX515 );
nand U8492 ( n460, n4586, WX517 );
nand U8493 ( n438, n4586, WX521 );
nand U8494 ( n383, n4586, WX531 );
nand U8495 ( n372, n4586, WX533 );
nand U8496 ( n361, n4586, WX535 );
nand U8497 ( n3689, WX1840, n4518 );
nand U8498 ( n3702, WX1838, n4518 );
nand U8499 ( n3714, WX1836, n4518 );
nand U8500 ( n3727, WX1834, n4518 );
nand U8501 ( n3739, WX1832, n4518 );
nand U8502 ( n3752, WX1830, n4518 );
nand U8503 ( n3765, WX1828, n4518 );
nand U8504 ( n3779, WX1826, n4521 );
nand U8505 ( n3793, WX1824, n4521 );
nand U8506 ( n3807, WX1822, n4521 );
nand U8507 ( n3820, WX1820, n4521 );
nand U8508 ( n3834, WX1818, n4521 );
nand U8509 ( n3848, WX1816, n4521 );
nand U8510 ( n3862, WX1814, n4521 );
nand U8511 ( n3875, WX1812, n4521 );
nand U8512 ( n3889, WX1810, n4521 );
nand U8513 ( n3905, WX1808, n4522 );
nand U8514 ( n3922, WX1806, n4522 );
nand U8515 ( n3938, WX1804, n4522 );
nand U8516 ( n3954, WX1802, n4522 );
nand U8517 ( n3970, WX1800, n4523 );
nand U8518 ( n3987, WX1798, n4522 );
nand U8519 ( n4003, WX1796, n4522 );
nand U8520 ( n4019, WX1794, n4522 );
nand U8521 ( n4035, WX1792, n4522 );
nand U8522 ( n4052, WX1790, n4522 );
nand U8523 ( n4068, WX1788, n4522 );
nand U8524 ( n4084, WX1786, n4522 );
nand U8525 ( n4100, WX1784, n4522 );
nand U8526 ( n4117, WX1782, n4523 );
nand U8527 ( n4133, WX1780, n4523 );
nand U8528 ( n3257, WX3133, n4524 );
nand U8529 ( n3270, WX3131, n4523 );
nand U8530 ( n3282, WX3129, n4523 );
nand U8531 ( n3295, WX3127, n4524 );
nand U8532 ( n3307, WX3125, n4524 );
nand U8533 ( n3320, WX3123, n4523 );
nand U8534 ( n3332, WX3121, n4523 );
nand U8535 ( n3345, WX3119, n4524 );
nand U8536 ( n3357, WX3117, n4523 );
nand U8537 ( n3370, WX3115, n4524 );
nand U8538 ( n3383, WX3113, n4524 );
nand U8539 ( n3397, WX3111, n4521 );
nand U8540 ( n3410, WX3109, n4521 );
nand U8541 ( n3423, WX3107, n4521 );
nand U8542 ( n3437, WX3105, n4520 );
nand U8543 ( n3450, WX3103, n4520 );
nand U8544 ( n3465, WX3101, n4520 );
nand U8545 ( n3479, WX3099, n4520 );
nand U8546 ( n3494, WX3097, n4520 );
nand U8547 ( n3505, WX3095, n4520 );
nand U8548 ( n3516, WX3093, n4520 );
nand U8549 ( n3527, WX3091, n4520 );
nand U8550 ( n3538, WX3089, n4520 );
nand U8551 ( n3549, WX3087, n4520 );
nand U8552 ( n3560, WX3085, n4520 );
nand U8553 ( n3571, WX3083, n4520 );
nand U8554 ( n3582, WX3081, n4519 );
nand U8555 ( n3593, WX3079, n4519 );
nand U8556 ( n3604, WX3077, n4519 );
nand U8557 ( n3615, WX3075, n4519 );
nand U8558 ( n3626, WX3073, n4519 );
nand U8559 ( n2795, WX4426, n4507 );
nand U8560 ( n2807, WX4424, n4507 );
nand U8561 ( n2820, WX4422, n4507 );
nand U8562 ( n2832, WX4420, n4507 );
nand U8563 ( n2845, WX4418, n4507 );
nand U8564 ( n2857, WX4416, n4507 );
nand U8565 ( n2870, WX4414, n4507 );
nand U8566 ( n2882, WX4412, n4507 );
nand U8567 ( n2895, WX4410, n4507 );
nand U8568 ( n2907, WX4408, n4507 );
nand U8569 ( n2920, WX4406, n4508 );
nand U8570 ( n2932, WX4404, n4508 );
nand U8571 ( n2945, WX4402, n4508 );
nand U8572 ( n2957, WX4400, n4508 );
nand U8573 ( n2970, WX4398, n4508 );
nand U8574 ( n2982, WX4396, n4508 );
nand U8575 ( n2996, WX4394, n4508 );
nand U8576 ( n3010, WX4392, n4508 );
nand U8577 ( n3024, WX4390, n4508 );
nand U8578 ( n3037, WX4388, n4508 );
nand U8579 ( n3051, WX4386, n4508 );
nand U8580 ( n3065, WX4384, n4508 );
nand U8581 ( n3079, WX4382, n4509 );
nand U8582 ( n3092, WX4380, n4509 );
nand U8583 ( n3106, WX4378, n4509 );
nand U8584 ( n3120, WX4376, n4509 );
nand U8585 ( n3134, WX4374, n4509 );
nand U8586 ( n3147, WX4372, n4509 );
nand U8587 ( n3161, WX4370, n4509 );
nand U8588 ( n3175, WX4368, n4509 );
nand U8589 ( n3189, WX4366, n4509 );
nand U8590 ( n2363, WX5719, n4513 );
nand U8591 ( n2376, WX5717, n4513 );
nand U8592 ( n2388, WX5715, n4512 );
nand U8593 ( n2401, WX5713, n4512 );
nand U8594 ( n2413, WX5711, n4512 );
nand U8595 ( n2426, WX5709, n4512 );
nand U8596 ( n2438, WX5707, n4512 );
nand U8597 ( n2451, WX5705, n4512 );
nand U8598 ( n2465, WX5703, n4512 );
nand U8599 ( n2478, WX5701, n4512 );
nand U8600 ( n2491, WX5699, n4512 );
nand U8601 ( n2505, WX5697, n4512 );
nand U8602 ( n2518, WX5695, n4512 );
nand U8603 ( n2531, WX5693, n4512 );
nand U8604 ( n2545, WX5691, n4511 );
nand U8605 ( n2558, WX5689, n4511 );
nand U8606 ( n2571, WX5687, n4511 );
nand U8607 ( n2582, WX5685, n4511 );
nand U8608 ( n2593, WX5683, n4511 );
nand U8609 ( n2604, WX5681, n4511 );
nand U8610 ( n2615, WX5679, n4511 );
nand U8611 ( n2626, WX5677, n4511 );
nand U8612 ( n2637, WX5675, n4511 );
nand U8613 ( n2648, WX5673, n4511 );
nand U8614 ( n2659, WX5671, n4504 );
nand U8615 ( n2670, WX5669, n4504 );
nand U8616 ( n2681, WX5667, n4504 );
nand U8617 ( n2692, WX5665, n4504 );
nand U8618 ( n2703, WX5663, n4504 );
nand U8619 ( n2714, WX5661, n4504 );
nand U8620 ( n2726, WX5659, n4504 );
nand U8621 ( n1901, WX7012, n4507 );
nand U8622 ( n1913, WX7010, n4518 );
nand U8623 ( n1926, WX7008, n4518 );
nand U8624 ( n1938, WX7006, n4518 );
nand U8625 ( n1951, WX7004, n4517 );
nand U8626 ( n1963, WX7002, n4517 );
nand U8627 ( n1976, WX7000, n4517 );
nand U8628 ( n1988, WX6998, n4517 );
nand U8629 ( n2001, WX6996, n4517 );
nand U8630 ( n2013, WX6994, n4517 );
nand U8631 ( n2026, WX6992, n4517 );
nand U8632 ( n2038, WX6990, n4517 );
nand U8633 ( n2051, WX6988, n4517 );
nand U8634 ( n2063, WX6986, n4517 );
nand U8635 ( n2076, WX6984, n4517 );
nand U8636 ( n2088, WX6982, n4517 );
nand U8637 ( n2102, WX6980, n4516 );
nand U8638 ( n2116, WX6978, n4516 );
nand U8639 ( n2129, WX6976, n4516 );
nand U8640 ( n2143, WX6974, n4516 );
nand U8641 ( n2157, WX6972, n4516 );
nand U8642 ( n2171, WX6970, n4516 );
nand U8643 ( n2184, WX6968, n4516 );
nand U8644 ( n2198, WX6966, n4516 );
nand U8645 ( n2212, WX6964, n4516 );
nand U8646 ( n2226, WX6962, n4516 );
nand U8647 ( n2239, WX6960, n4516 );
nand U8648 ( n2253, WX6958, n4516 );
nand U8649 ( n2267, WX6956, n4515 );
nand U8650 ( n2281, WX6954, n4515 );
nand U8651 ( n2294, WX6952, n4515 );
nand U8652 ( n1469, WX8305, n4513 );
nand U8653 ( n1481, WX8303, n4513 );
nand U8654 ( n1494, WX8301, n4513 );
nand U8655 ( n1506, WX8299, n4513 );
nand U8656 ( n1519, WX8297, n4513 );
nand U8657 ( n1533, WX8295, n4513 );
nand U8658 ( n1546, WX8293, n4513 );
nand U8659 ( n1559, WX8291, n4513 );
nand U8660 ( n1573, WX8289, n4513 );
nand U8661 ( n1586, WX8287, n4513 );
nand U8662 ( n1599, WX8285, n4514 );
nand U8663 ( n1613, WX8283, n4514 );
nand U8664 ( n1626, WX8281, n4514 );
nand U8665 ( n1639, WX8279, n4514 );
nand U8666 ( n1649, WX8277, n4514 );
nand U8667 ( n1659, WX8275, n4514 );
nand U8668 ( n1670, WX8273, n4514 );
nand U8669 ( n1681, WX8271, n4514 );
nand U8670 ( n1692, WX8269, n4514 );
nand U8671 ( n1703, WX8267, n4514 );
nand U8672 ( n1714, WX8265, n4514 );
nand U8673 ( n1725, WX8263, n4514 );
nand U8674 ( n1736, WX8261, n4515 );
nand U8675 ( n1747, WX8259, n4515 );
nand U8676 ( n1758, WX8257, n4515 );
nand U8677 ( n1769, WX8255, n4515 );
nand U8678 ( n1780, WX8253, n4515 );
nand U8679 ( n1791, WX8251, n4515 );
nand U8680 ( n1804, WX8249, n4515 );
nand U8681 ( n1818, WX8247, n4515 );
nand U8682 ( n1832, WX8245, n4515 );
nand U8683 ( n1006, WX9598, n4507 );
nand U8684 ( n1019, WX9596, n4506 );
nand U8685 ( n1031, WX9594, n4506 );
nand U8686 ( n1044, WX9592, n4506 );
nand U8687 ( n1056, WX9590, n4506 );
nand U8688 ( n1069, WX9588, n4506 );
nand U8689 ( n1081, WX9586, n4506 );
nand U8690 ( n1094, WX9584, n4506 );
nand U8691 ( n1106, WX9582, n4506 );
nand U8692 ( n1119, WX9580, n4506 );
nand U8693 ( n1131, WX9578, n4506 );
nand U8694 ( n1144, WX9576, n4506 );
nand U8695 ( n1156, WX9574, n4506 );
nand U8696 ( n1169, WX9572, n4505 );
nand U8697 ( n1181, WX9570, n4505 );
nand U8698 ( n1194, WX9568, n4518 );
nand U8699 ( n1208, WX9566, n4505 );
nand U8700 ( n1221, WX9564, n4505 );
nand U8701 ( n1235, WX9562, n4505 );
nand U8702 ( n1249, WX9560, n4505 );
nand U8703 ( n1263, WX9558, n4505 );
nand U8704 ( n1276, WX9556, n4505 );
nand U8705 ( n1290, WX9554, n4505 );
nand U8706 ( n1304, WX9552, n4505 );
nand U8707 ( n1318, WX9550, n4505 );
nand U8708 ( n1331, WX9548, n4505 );
nand U8709 ( n1345, WX9546, n4504 );
nand U8710 ( n1359, WX9544, n4504 );
nand U8711 ( n1373, WX9542, n4504 );
nand U8712 ( n1386, WX9540, n4504 );
nand U8713 ( n1400, WX9538, n4504 );
nand U8714 ( n684, WX10891, n4518 );
nand U8715 ( n692, WX10889, n4519 );
nand U8716 ( n700, WX10887, n4519 );
nand U8717 ( n708, WX10885, n4519 );
nand U8718 ( n716, WX10883, n4519 );
nand U8719 ( n724, WX10881, n4519 );
nand U8720 ( n732, WX10879, n4519 );
nand U8721 ( n741, WX10877, n4519 );
nand U8722 ( n749, WX10875, n4524 );
nand U8723 ( n757, WX10873, n4523 );
nand U8724 ( n765, WX10871, n4524 );
nand U8725 ( n773, WX10869, n4523 );
nand U8726 ( n781, WX10867, n4524 );
nand U8727 ( n789, WX10865, n4523 );
nand U8728 ( n797, WX10863, n4511 );
nand U8729 ( n805, WX10861, n4510 );
nand U8730 ( n813, WX10859, n4510 );
nand U8731 ( n822, WX10857, n4510 );
nand U8732 ( n830, WX10855, n4510 );
nand U8733 ( n838, WX10853, n4510 );
nand U8734 ( n846, WX10851, n4510 );
nand U8735 ( n854, WX10849, n4511 );
nand U8736 ( n862, WX10847, n4510 );
nand U8737 ( n871, WX10845, n4510 );
nand U8738 ( n881, WX10843, n4510 );
nand U8739 ( n891, WX10841, n4510 );
nand U8740 ( n901, WX10839, n4510 );
nand U8741 ( n911, WX10837, n4510 );
nand U8742 ( n921, WX10835, n4509 );
nand U8743 ( n931, WX10833, n4509 );
nand U8744 ( n941, WX10831, n4509 );
nand U8745 ( n675, n4588, WX541 );
nand U8746 ( n733, n4588, WX539 );
nand U8747 ( n416, n4588, WX525 );
and U8748 ( n2275, n4564, WX2064 );
and U8749 ( n2270, n4564, WX2062 );
and U8750 ( n2265, n4564, WX2060 );
and U8751 ( n2260, n4563, WX2058 );
and U8752 ( n2255, n4563, WX2056 );
and U8753 ( n2250, n4563, WX2054 );
and U8754 ( n2245, n4563, WX2052 );
and U8755 ( n2240, n4563, WX2050 );
and U8756 ( n2235, n4563, WX2048 );
and U8757 ( n2230, n4563, WX2046 );
and U8758 ( n2225, n4563, WX2044 );
and U8759 ( n2220, n4563, WX2042 );
and U8760 ( n2215, n4563, WX2040 );
and U8761 ( n2210, n4563, WX2038 );
and U8762 ( n2205, n4563, WX2036 );
and U8763 ( n2200, n4562, WX2034 );
and U8764 ( n3203, n4554, WX3357 );
and U8765 ( n3198, n4554, WX3355 );
and U8766 ( n3193, n4554, WX3353 );
and U8767 ( n3188, n4554, WX3351 );
and U8768 ( n3183, n4554, WX3349 );
and U8769 ( n3178, n4554, WX3347 );
and U8770 ( n3173, n4554, WX3345 );
and U8771 ( n3168, n4554, WX3343 );
and U8772 ( n3163, n4554, WX3341 );
and U8773 ( n3158, n4554, WX3339 );
and U8774 ( n3153, n4554, WX3337 );
and U8775 ( n3148, n4554, WX3335 );
and U8776 ( n3143, n4553, WX3333 );
and U8777 ( n3138, n4553, WX3331 );
and U8778 ( n3133, n4553, WX3329 );
and U8779 ( n3128, n4553, WX3327 );
and U8780 ( n4131, n4580, WX4650 );
and U8781 ( n4126, n4580, WX4648 );
and U8782 ( n4121, n4580, WX4646 );
and U8783 ( n4116, n4580, WX4644 );
and U8784 ( n4111, n4580, WX4642 );
and U8785 ( n4106, n4580, WX4640 );
and U8786 ( n4101, n4580, WX4638 );
and U8787 ( n4096, n4578, WX4636 );
and U8788 ( n4091, n4578, WX4634 );
and U8789 ( n4086, n4578, WX4632 );
and U8790 ( n4081, n4578, WX4630 );
and U8791 ( n4076, n4578, WX4628 );
and U8792 ( n4071, n4578, WX4626 );
and U8793 ( n4066, n4578, WX4624 );
and U8794 ( n4061, n4578, WX4622 );
and U8795 ( n4056, n4578, WX4620 );
and U8796 ( n5059, n4570, WX5943 );
and U8797 ( n5054, n4570, WX5941 );
and U8798 ( n5049, n4570, WX5939 );
and U8799 ( n5044, n4570, WX5937 );
and U8800 ( n5039, n4570, WX5935 );
and U8801 ( n5034, n4570, WX5933 );
and U8802 ( n5029, n4570, WX5931 );
and U8803 ( n5024, n4570, WX5929 );
and U8804 ( n5019, n4570, WX5927 );
and U8805 ( n5014, n4569, WX5925 );
and U8806 ( n5009, n4569, WX5923 );
and U8807 ( n5004, n4569, WX5921 );
and U8808 ( n4999, n4569, WX5919 );
and U8809 ( n4994, n4569, WX5917 );
and U8810 ( n4989, n4569, WX5915 );
and U8811 ( n4984, n4569, WX5913 );
and U8812 ( n6915, n4549, WX8529 );
and U8813 ( n6910, n4549, WX8527 );
and U8814 ( n6905, n4549, WX8525 );
and U8815 ( n6900, n4549, WX8523 );
and U8816 ( n6895, n4549, WX8521 );
and U8817 ( n6890, n4549, WX8519 );
and U8818 ( n6885, n4549, WX8517 );
and U8819 ( n6880, n4549, WX8515 );
and U8820 ( n6875, n4549, WX8513 );
and U8821 ( n6870, n4549, WX8511 );
and U8822 ( n2435, n4566, WX2128 );
and U8823 ( n2430, n4566, WX2126 );
and U8824 ( n2425, n4566, WX2124 );
and U8825 ( n2420, n4566, WX2122 );
and U8826 ( n2415, n4566, WX2120 );
and U8827 ( n2410, n4566, WX2118 );
and U8828 ( n2405, n4566, WX2116 );
and U8829 ( n2400, n4566, WX2114 );
and U8830 ( n2395, n4566, WX2112 );
and U8831 ( n2390, n4565, WX2110 );
and U8832 ( n2385, n4565, WX2108 );
and U8833 ( n2380, n4565, WX2106 );
and U8834 ( n2375, n4565, WX2104 );
and U8835 ( n2370, n4565, WX2102 );
and U8836 ( n2365, n4565, WX2100 );
and U8837 ( n2360, n4565, WX2098 );
and U8838 ( n2355, n4565, WX2096 );
and U8839 ( n2035, n4560, WX1968 );
and U8840 ( n2350, n4565, WX2094 );
and U8841 ( n2030, n4560, WX1966 );
and U8842 ( n2345, n4565, WX2092 );
and U8843 ( n2025, n4560, WX1964 );
and U8844 ( n2340, n4565, WX2090 );
and U8845 ( n2020, n4560, WX1962 );
and U8846 ( n2335, n4565, WX2088 );
and U8847 ( n2015, n4560, WX1960 );
and U8848 ( n2330, n4565, WX2086 );
and U8849 ( n2010, n4560, WX1958 );
and U8850 ( n2325, n4564, WX2084 );
and U8851 ( n2005, n4559, WX1956 );
and U8852 ( n2320, n4564, WX2082 );
and U8853 ( n2000, n4559, WX1954 );
and U8854 ( n2315, n4564, WX2080 );
and U8855 ( n1995, n4559, WX1952 );
and U8856 ( n2310, n4564, WX2078 );
and U8857 ( n1990, n4559, WX1950 );
and U8858 ( n2305, n4564, WX2076 );
and U8859 ( n1985, n4559, WX1948 );
and U8860 ( n2300, n4564, WX2074 );
and U8861 ( n1980, n4559, WX1946 );
and U8862 ( n2295, n4564, WX2072 );
and U8863 ( n1975, n4559, WX1944 );
and U8864 ( n2290, n4564, WX2070 );
and U8865 ( n1970, n4559, WX1942 );
and U8866 ( n2285, n4564, WX2068 );
and U8867 ( n1965, n4559, WX1940 );
and U8868 ( n2280, n4564, WX2066 );
and U8869 ( n1960, n4563, WX1938 );
and U8870 ( n3363, n4557, WX3421 );
and U8871 ( n3358, n4557, WX3419 );
and U8872 ( n3353, n4557, WX3417 );
and U8873 ( n3348, n4557, WX3415 );
and U8874 ( n3343, n4557, WX3413 );
and U8875 ( n3338, n4557, WX3411 );
and U8876 ( n3333, n4556, WX3409 );
and U8877 ( n3328, n4556, WX3407 );
and U8878 ( n3323, n4556, WX3405 );
and U8879 ( n3318, n4556, WX3403 );
and U8880 ( n3313, n4556, WX3401 );
and U8881 ( n3308, n4556, WX3399 );
and U8882 ( n3303, n4556, WX3397 );
and U8883 ( n3298, n4556, WX3395 );
and U8884 ( n3293, n4556, WX3393 );
and U8885 ( n3288, n4556, WX3391 );
and U8886 ( n3283, n4556, WX3389 );
and U8887 ( n2963, n4551, WX3261 );
and U8888 ( n3278, n4556, WX3387 );
and U8889 ( n2958, n4551, WX3259 );
and U8890 ( n3273, n4556, WX3385 );
and U8891 ( n2953, n4551, WX3257 );
and U8892 ( n3268, n4555, WX3383 );
and U8893 ( n2948, n4555, WX3255 );
and U8894 ( n3263, n4555, WX3381 );
and U8895 ( n2943, n4567, WX3253 );
and U8896 ( n3258, n4555, WX3379 );
and U8897 ( n2938, n4567, WX3251 );
and U8898 ( n3253, n4555, WX3377 );
and U8899 ( n2933, n4567, WX3249 );
and U8900 ( n3248, n4555, WX3375 );
and U8901 ( n2928, n4567, WX3247 );
and U8902 ( n3243, n4555, WX3373 );
and U8903 ( n2923, n4567, WX3245 );
and U8904 ( n3238, n4555, WX3371 );
and U8905 ( n2918, n4567, WX3243 );
and U8906 ( n3233, n4555, WX3369 );
and U8907 ( n2913, n4567, WX3241 );
and U8908 ( n3228, n4555, WX3367 );
and U8909 ( n2908, n4567, WX3239 );
and U8910 ( n3223, n4555, WX3365 );
and U8911 ( n2903, n4566, WX3237 );
and U8912 ( n3218, n4555, WX3363 );
and U8913 ( n2898, n4566, WX3235 );
and U8914 ( n3213, n4555, WX3361 );
and U8915 ( n2893, n4566, WX3233 );
and U8916 ( n3208, n4554, WX3359 );
and U8917 ( n2888, n4566, WX3231 );
and U8918 ( n4291, n4583, WX4714 );
and U8919 ( n4286, n4583, WX4712 );
and U8920 ( n4281, n4582, WX4710 );
and U8921 ( n4276, n4582, WX4708 );
and U8922 ( n4271, n4582, WX4706 );
and U8923 ( n4266, n4582, WX4704 );
and U8924 ( n4261, n4582, WX4702 );
and U8925 ( n4256, n4582, WX4700 );
and U8926 ( n4251, n4582, WX4698 );
and U8927 ( n4246, n4582, WX4696 );
and U8928 ( n4241, n4582, WX4694 );
and U8929 ( n4236, n4582, WX4692 );
and U8930 ( n4231, n4581, WX4690 );
and U8931 ( n4226, n4582, WX4688 );
and U8932 ( n4221, n4582, WX4686 );
and U8933 ( n4216, n4581, WX4684 );
and U8934 ( n4211, n4581, WX4682 );
and U8935 ( n3891, n4558, WX4554 );
and U8936 ( n4206, n4581, WX4680 );
and U8937 ( n3886, n4558, WX4552 );
and U8938 ( n4201, n4581, WX4678 );
and U8939 ( n3881, n4558, WX4550 );
and U8940 ( n4196, n4581, WX4676 );
and U8941 ( n3876, n4558, WX4548 );
and U8942 ( n4191, n4581, WX4674 );
and U8943 ( n3871, n4558, WX4546 );
and U8944 ( n4186, n4581, WX4672 );
and U8945 ( n3866, n4558, WX4544 );
and U8946 ( n4181, n4581, WX4670 );
and U8947 ( n3861, n4558, WX4542 );
and U8948 ( n4176, n4581, WX4668 );
and U8949 ( n3856, n4558, WX4540 );
and U8950 ( n4171, n4581, WX4666 );
and U8951 ( n3851, n4558, WX4538 );
and U8952 ( n4166, n4581, WX4664 );
and U8953 ( n3846, n4557, WX4536 );
and U8954 ( n4161, n4580, WX4662 );
and U8955 ( n3841, n4557, WX4534 );
and U8956 ( n4156, n4580, WX4660 );
and U8957 ( n3836, n4557, WX4532 );
and U8958 ( n4151, n4580, WX4658 );
and U8959 ( n3831, n4557, WX4530 );
and U8960 ( n4146, n4580, WX4656 );
and U8961 ( n3826, n4557, WX4528 );
and U8962 ( n4141, n4580, WX4654 );
and U8963 ( n3821, n4557, WX4526 );
and U8964 ( n4136, n4580, WX4652 );
and U8965 ( n3816, n4557, WX4524 );
and U8966 ( n5219, n4573, WX6007 );
and U8967 ( n5214, n4573, WX6005 );
and U8968 ( n5209, n4573, WX6003 );
and U8969 ( n5204, n4572, WX6001 );
and U8970 ( n5199, n4572, WX5999 );
and U8971 ( n5194, n4572, WX5997 );
and U8972 ( n5189, n4572, WX5995 );
and U8973 ( n5184, n4572, WX5993 );
and U8974 ( n5179, n4572, WX5991 );
and U8975 ( n5174, n4572, WX5989 );
and U8976 ( n5169, n4572, WX5987 );
and U8977 ( n5164, n4572, WX5985 );
and U8978 ( n5159, n4572, WX5983 );
and U8979 ( n5154, n4572, WX5981 );
and U8980 ( n5149, n4572, WX5979 );
and U8981 ( n5144, n4571, WX5977 );
and U8982 ( n5139, n4571, WX5975 );
and U8983 ( n4819, n4585, WX5847 );
and U8984 ( n5134, n4571, WX5973 );
and U8985 ( n4814, n4583, WX5845 );
and U8986 ( n5129, n4571, WX5971 );
and U8987 ( n4809, n4583, WX5843 );
and U8988 ( n5124, n4571, WX5969 );
and U8989 ( n4804, n4585, WX5841 );
and U8990 ( n5119, n4571, WX5967 );
and U8991 ( n4799, n4585, WX5839 );
and U8992 ( n5114, n4571, WX5965 );
and U8993 ( n4794, n4585, WX5837 );
and U8994 ( n5109, n4571, WX5963 );
and U8995 ( n4789, n4583, WX5835 );
and U8996 ( n5104, n4571, WX5961 );
and U8997 ( n4784, n4585, WX5833 );
and U8998 ( n5099, n4571, WX5959 );
and U8999 ( n4779, n4583, WX5831 );
and U9000 ( n5094, n4571, WX5957 );
and U9001 ( n4774, n4583, WX5829 );
and U9002 ( n5089, n4571, WX5955 );
and U9003 ( n4769, n4583, WX5827 );
and U9004 ( n5084, n4571, WX5953 );
and U9005 ( n4764, n4583, WX5825 );
and U9006 ( n5079, n4570, WX5951 );
and U9007 ( n4759, n4583, WX5823 );
and U9008 ( n5074, n4570, WX5949 );
and U9009 ( n4754, n4583, WX5821 );
and U9010 ( n5069, n4570, WX5947 );
and U9011 ( n4749, n4583, WX5819 );
and U9012 ( n5064, n4570, WX5945 );
and U9013 ( n4744, n4583, WX5817 );
and U9014 ( n5747, n4574, WX7140 );
and U9015 ( n5742, n4574, WX7138 );
and U9016 ( n5737, n4574, WX7136 );
and U9017 ( n5732, n4574, WX7134 );
and U9018 ( n5727, n4574, WX7132 );
and U9019 ( n5722, n4574, WX7130 );
and U9020 ( n5717, n4573, WX7128 );
and U9021 ( n5712, n4573, WX7126 );
and U9022 ( n5707, n4573, WX7124 );
and U9023 ( n5702, n4573, WX7122 );
and U9024 ( n5697, n4573, WX7120 );
and U9025 ( n5692, n4573, WX7118 );
and U9026 ( n5687, n4573, WX7116 );
and U9027 ( n5682, n4573, WX7114 );
and U9028 ( n5677, n4573, WX7112 );
and U9029 ( n5672, n4573, WX7110 );
and U9030 ( n7075, n4546, WX8593 );
and U9031 ( n7070, n4546, WX8591 );
and U9032 ( n7065, n4546, WX8589 );
and U9033 ( n7060, n4546, WX8587 );
and U9034 ( n7055, n4546, WX8585 );
and U9035 ( n7050, n4547, WX8583 );
and U9036 ( n7045, n4547, WX8581 );
and U9037 ( n7040, n4547, WX8579 );
and U9038 ( n7035, n4547, WX8577 );
and U9039 ( n7030, n4547, WX8575 );
and U9040 ( n7025, n4547, WX8573 );
and U9041 ( n7020, n4547, WX8571 );
and U9042 ( n7015, n4547, WX8569 );
and U9043 ( n7010, n4547, WX8567 );
and U9044 ( n7005, n4547, WX8565 );
and U9045 ( n7000, n4547, WX8563 );
and U9046 ( n6995, n4547, WX8561 );
and U9047 ( n6990, n4547, WX8559 );
and U9048 ( n6985, n4548, WX8557 );
and U9049 ( n6980, n4548, WX8555 );
and U9050 ( n6975, n4548, WX8553 );
and U9051 ( n6970, n4548, WX8551 );
and U9052 ( n6965, n4548, WX8549 );
and U9053 ( n6960, n4548, WX8547 );
and U9054 ( n6955, n4548, WX8545 );
and U9055 ( n6950, n4548, WX8543 );
and U9056 ( n6945, n4548, WX8541 );
and U9057 ( n6940, n4548, WX8539 );
and U9058 ( n6935, n4548, WX8537 );
and U9059 ( n6930, n4548, WX8535 );
and U9060 ( n6925, n4548, WX8533 );
and U9061 ( n6920, n4549, WX8531 );
and U9062 ( n7998, n4543, WX9884 );
and U9063 ( n7603, n4542, WX9726 );
and U9064 ( n7598, n4543, WX9724 );
and U9065 ( n7593, n4543, WX9722 );
and U9066 ( n7588, n4543, WX9720 );
and U9067 ( n7583, n4543, WX9718 );
and U9068 ( n7578, n4543, WX9716 );
and U9069 ( n7573, n4543, WX9714 );
and U9070 ( n7568, n4543, WX9712 );
and U9071 ( n7563, n4543, WX9710 );
and U9072 ( n7558, n4543, WX9708 );
and U9073 ( n7553, n4543, WX9706 );
and U9074 ( n7548, n4543, WX9704 );
and U9075 ( n7543, n4543, WX9702 );
and U9076 ( n7538, n4544, WX9700 );
and U9077 ( n7533, n4544, WX9698 );
and U9078 ( n7528, n4544, WX9696 );
and U9079 ( n8456, n4542, WX10989 );
and U9080 ( n8931, n4550, WX11179 );
and U9081 ( n8531, n4545, WX11019 );
and U9082 ( n8526, n4545, WX11017 );
and U9083 ( n8521, n4545, WX11015 );
and U9084 ( n8516, n4544, WX11013 );
and U9085 ( n8511, n4544, WX11011 );
and U9086 ( n8506, n4544, WX11009 );
and U9087 ( n8501, n4544, WX11007 );
and U9088 ( n8496, n4544, WX11005 );
and U9089 ( n8491, n4544, WX11003 );
and U9090 ( n8486, n4544, WX11001 );
and U9091 ( n8481, n4544, WX10999 );
and U9092 ( n8476, n4544, WX10997 );
and U9093 ( n8471, n4544, WX10995 );
and U9094 ( n8466, n4542, WX10993 );
and U9095 ( n8461, n4542, WX10991 );
and U9096 ( n2115, n4561, WX2000 );
and U9097 ( n2110, n4561, WX1998 );
and U9098 ( n2105, n4561, WX1996 );
and U9099 ( n2100, n4561, WX1994 );
and U9100 ( n2095, n4561, WX1992 );
and U9101 ( n2090, n4561, WX1990 );
and U9102 ( n2085, n4561, WX1988 );
and U9103 ( n2080, n4561, WX1986 );
and U9104 ( n2075, n4561, WX1984 );
and U9105 ( n2070, n4560, WX1982 );
and U9106 ( n2065, n4560, WX1980 );
and U9107 ( n2060, n4560, WX1978 );
and U9108 ( n2055, n4560, WX1976 );
and U9109 ( n2050, n4560, WX1974 );
and U9110 ( n2045, n4560, WX1972 );
and U9111 ( n2040, n4560, WX1970 );
and U9112 ( n2195, n4562, WX2032 );
and U9113 ( n2190, n4562, WX2030 );
and U9114 ( n2185, n4562, WX2028 );
and U9115 ( n2180, n4562, WX2026 );
and U9116 ( n2175, n4562, WX2024 );
and U9117 ( n2170, n4562, WX2022 );
and U9118 ( n2165, n4562, WX2020 );
and U9119 ( n2160, n4562, WX2018 );
and U9120 ( n2155, n4562, WX2016 );
and U9121 ( n2150, n4562, WX2014 );
and U9122 ( n2145, n4562, WX2012 );
and U9123 ( n2140, n4562, WX2010 );
and U9124 ( n2135, n4561, WX2008 );
and U9125 ( n2130, n4561, WX2006 );
and U9126 ( n2125, n4561, WX2004 );
and U9127 ( n2120, n4561, WX2002 );
and U9128 ( n3043, n4552, WX3293 );
and U9129 ( n3038, n4552, WX3291 );
and U9130 ( n3033, n4552, WX3289 );
and U9131 ( n3028, n4552, WX3287 );
and U9132 ( n3023, n4552, WX3285 );
and U9133 ( n3018, n4552, WX3283 );
and U9134 ( n3013, n4551, WX3281 );
and U9135 ( n3008, n4551, WX3279 );
and U9136 ( n3003, n4551, WX3277 );
and U9137 ( n2998, n4551, WX3275 );
and U9138 ( n2993, n4551, WX3273 );
and U9139 ( n2988, n4551, WX3271 );
and U9140 ( n2983, n4551, WX3269 );
and U9141 ( n2978, n4551, WX3267 );
and U9142 ( n2973, n4551, WX3265 );
and U9143 ( n2968, n4551, WX3263 );
and U9144 ( n3123, n4553, WX3325 );
and U9145 ( n3118, n4553, WX3323 );
and U9146 ( n3113, n4553, WX3321 );
and U9147 ( n3108, n4553, WX3319 );
and U9148 ( n3103, n4553, WX3317 );
and U9149 ( n3098, n4553, WX3315 );
and U9150 ( n3093, n4553, WX3313 );
and U9151 ( n3088, n4553, WX3311 );
and U9152 ( n3083, n4553, WX3309 );
and U9153 ( n3078, n4552, WX3307 );
and U9154 ( n3073, n4552, WX3305 );
and U9155 ( n3068, n4552, WX3303 );
and U9156 ( n3063, n4552, WX3301 );
and U9157 ( n3058, n4552, WX3299 );
and U9158 ( n3053, n4552, WX3297 );
and U9159 ( n3048, n4552, WX3295 );
and U9160 ( n3971, n4577, WX4586 );
and U9161 ( n3966, n4577, WX4584 );
and U9162 ( n3961, n4576, WX4582 );
and U9163 ( n3956, n4576, WX4580 );
and U9164 ( n3951, n4576, WX4578 );
and U9165 ( n3946, n4576, WX4576 );
and U9166 ( n3941, n4576, WX4574 );
and U9167 ( n3936, n4576, WX4572 );
and U9168 ( n3931, n4559, WX4570 );
and U9169 ( n3926, n4559, WX4568 );
and U9170 ( n3921, n4559, WX4566 );
and U9171 ( n3916, n4559, WX4564 );
and U9172 ( n3911, n4558, WX4562 );
and U9173 ( n3906, n4558, WX4560 );
and U9174 ( n3901, n4558, WX4558 );
and U9175 ( n3896, n4558, WX4556 );
and U9176 ( n4051, n4578, WX4618 );
and U9177 ( n4046, n4578, WX4616 );
and U9178 ( n4041, n4578, WX4614 );
and U9179 ( n4036, n4578, WX4612 );
and U9180 ( n4031, n4577, WX4610 );
and U9181 ( n4026, n4581, WX4608 );
and U9182 ( n4021, n4577, WX4606 );
and U9183 ( n4016, n4577, WX4604 );
and U9184 ( n4011, n4577, WX4602 );
and U9185 ( n4006, n4577, WX4600 );
and U9186 ( n4001, n4577, WX4598 );
and U9187 ( n3996, n4577, WX4596 );
and U9188 ( n3991, n4577, WX4594 );
and U9189 ( n3986, n4577, WX4592 );
and U9190 ( n3981, n4577, WX4590 );
and U9191 ( n3976, n4577, WX4588 );
and U9192 ( n4899, n4568, WX5879 );
and U9193 ( n4894, n4568, WX5877 );
and U9194 ( n4889, n4568, WX5875 );
and U9195 ( n4884, n4567, WX5873 );
and U9196 ( n4879, n4567, WX5871 );
and U9197 ( n4874, n4567, WX5869 );
and U9198 ( n4869, n4567, WX5867 );
and U9199 ( n4864, n4567, WX5865 );
and U9200 ( n4859, n4572, WX5863 );
and U9201 ( n4854, n4582, WX5861 );
and U9202 ( n4849, n4585, WX5859 );
and U9203 ( n4844, n4585, WX5857 );
and U9204 ( n4839, n4585, WX5855 );
and U9205 ( n4834, n4585, WX5853 );
and U9206 ( n4829, n4585, WX5851 );
and U9207 ( n4824, n4585, WX5849 );
and U9208 ( n4979, n4569, WX5911 );
and U9209 ( n4974, n4569, WX5909 );
and U9210 ( n4969, n4569, WX5907 );
and U9211 ( n4964, n4569, WX5905 );
and U9212 ( n4959, n4569, WX5903 );
and U9213 ( n4954, n4569, WX5901 );
and U9214 ( n4949, n4568, WX5899 );
and U9215 ( n4944, n4568, WX5897 );
and U9216 ( n4939, n4568, WX5895 );
and U9217 ( n4934, n4568, WX5893 );
and U9218 ( n4929, n4568, WX5891 );
and U9219 ( n4924, n4568, WX5889 );
and U9220 ( n4919, n4568, WX5887 );
and U9221 ( n4914, n4568, WX5885 );
and U9222 ( n4909, n4568, WX5883 );
and U9223 ( n4904, n4568, WX5881 );
and U9224 ( n5827, n4575, WX7172 );
and U9225 ( n5822, n4575, WX7170 );
and U9226 ( n5817, n4575, WX7168 );
and U9227 ( n5812, n4575, WX7166 );
and U9228 ( n5807, n4575, WX7164 );
and U9229 ( n5802, n4575, WX7162 );
and U9230 ( n5797, n4575, WX7160 );
and U9231 ( n5792, n4575, WX7158 );
and U9232 ( n5787, n4575, WX7156 );
and U9233 ( n5782, n4574, WX7154 );
and U9234 ( n5777, n4574, WX7152 );
and U9235 ( n5772, n4574, WX7150 );
and U9236 ( n5767, n4574, WX7148 );
and U9237 ( n5762, n4574, WX7146 );
and U9238 ( n5757, n4574, WX7144 );
and U9239 ( n5752, n4574, WX7142 );
and U9240 ( n5887, n4545, WX7196 );
and U9241 ( n5882, n4576, WX7194 );
and U9242 ( n5877, n4576, WX7192 );
and U9243 ( n5872, n4576, WX7190 );
and U9244 ( n5867, n4576, WX7188 );
and U9245 ( n5862, n4576, WX7186 );
and U9246 ( n5857, n4576, WX7184 );
and U9247 ( n5852, n4576, WX7182 );
and U9248 ( n5847, n4575, WX7180 );
and U9249 ( n5842, n4575, WX7178 );
and U9250 ( n5837, n4575, WX7176 );
and U9251 ( n5832, n4575, WX7174 );
and U9252 ( n7683, n4541, WX9758 );
and U9253 ( n7678, n4541, WX9756 );
and U9254 ( n7673, n4541, WX9754 );
and U9255 ( n7668, n4541, WX9752 );
and U9256 ( n7663, n4541, WX9750 );
and U9257 ( n7658, n4541, WX9748 );
and U9258 ( n7653, n4541, WX9746 );
and U9259 ( n7648, n4542, WX9744 );
and U9260 ( n7643, n4542, WX9742 );
and U9261 ( n7638, n4542, WX9740 );
and U9262 ( n7633, n4542, WX9738 );
and U9263 ( n7628, n4542, WX9736 );
and U9264 ( n7623, n4542, WX9734 );
and U9265 ( n7618, n4542, WX9732 );
and U9266 ( n7613, n4542, WX9730 );
and U9267 ( n7608, n4542, WX9728 );
and U9268 ( n7713, n4541, WX9770 );
and U9269 ( n7708, n4541, WX9768 );
and U9270 ( n7703, n4541, WX9766 );
and U9271 ( n7698, n4541, WX9764 );
and U9272 ( n7693, n4541, WX9762 );
and U9273 ( n7688, n4541, WX9760 );
and U9274 ( n8616, n4546, WX11053 );
and U9275 ( n8611, n4546, WX11051 );
and U9276 ( n8606, n4546, WX11049 );
and U9277 ( n8601, n4546, WX11047 );
and U9278 ( n8596, n4546, WX11045 );
and U9279 ( n8591, n4546, WX11043 );
and U9280 ( n8586, n4546, WX11041 );
and U9281 ( n8581, n4546, WX11039 );
and U9282 ( n8576, n4545, WX11037 );
and U9283 ( n8571, n4545, WX11035 );
and U9284 ( n8566, n4545, WX11033 );
and U9285 ( n8561, n4545, WX11031 );
and U9286 ( n8556, n4545, WX11029 );
and U9287 ( n8551, n4545, WX11027 );
and U9288 ( n8546, n4545, WX11025 );
and U9289 ( n8541, n4545, WX11023 );
and U9290 ( n8536, n4545, WX11021 );
and U9291 ( n8686, n4550, WX11081 );
and U9292 ( n8681, n4550, WX11079 );
and U9293 ( n8676, n4550, WX11077 );
and U9294 ( n8671, n4550, WX11075 );
and U9295 ( n8666, n4550, WX11073 );
and U9296 ( n8661, n4550, WX11071 );
and U9297 ( n8656, n4550, WX11069 );
and U9298 ( n8651, n4550, WX11067 );
and U9299 ( n8646, n4550, WX11065 );
and U9300 ( n8641, n4550, WX11063 );
and U9301 ( n8636, n4550, WX11061 );
and U9302 ( n8631, n4550, WX11059 );
and U9303 ( n8626, n4549, WX11057 );
and U9304 ( n8621, n4549, WX11055 );
and U9305 ( n1507, WX835, n4496 );
and U9306 ( n1502, WX833, n4496 );
and U9307 ( n1497, WX831, n4496 );
and U9308 ( n1492, WX829, n4496 );
and U9309 ( n1487, WX827, n4496 );
and U9310 ( n1482, WX825, n4496 );
and U9311 ( n1357, WX775, n4498 );
and U9312 ( n1362, WX777, n4498 );
and U9313 ( n1367, WX779, n4498 );
and U9314 ( n1372, WX781, n4498 );
and U9315 ( n1377, WX783, n4498 );
and U9316 ( n1382, WX785, n4498 );
and U9317 ( n1387, WX787, n4498 );
and U9318 ( n1392, WX789, n4497 );
and U9319 ( n1397, WX791, n4497 );
and U9320 ( n1402, WX793, n4497 );
and U9321 ( n1407, WX795, n4497 );
and U9322 ( n1412, WX797, n4497 );
and U9323 ( n1417, WX799, n4497 );
and U9324 ( n1422, WX801, n4497 );
and U9325 ( n1427, WX803, n4497 );
and U9326 ( n1432, WX805, n4497 );
and U9327 ( n1437, WX807, n4497 );
and U9328 ( n1442, WX809, n4497 );
and U9329 ( n1447, WX811, n4497 );
and U9330 ( n1452, WX813, n4496 );
and U9331 ( n1457, WX815, n4496 );
and U9332 ( n1462, WX817, n4496 );
and U9333 ( n1467, WX819, n4496 );
and U9334 ( n1472, WX821, n4496 );
and U9335 ( n1477, WX823, n4496 );
and U9336 ( n1352, WX773, n4498 );
and U9337 ( n1187, WX707, n4501 );
and U9338 ( n1182, WX705, n4501 );
and U9339 ( n1177, WX703, n4501 );
and U9340 ( n1172, WX701, n4501 );
and U9341 ( n1167, WX699, n4501 );
and U9342 ( n1162, WX697, n4501 );
and U9343 ( n1037, WX647, n4503 );
and U9344 ( n1042, WX649, n4503 );
and U9345 ( n1047, WX651, n4503 );
and U9346 ( n1052, WX653, n4503 );
and U9347 ( n1057, WX655, n4503 );
and U9348 ( n1062, WX657, n4503 );
and U9349 ( n1067, WX659, n4503 );
and U9350 ( n1072, WX661, n4502 );
and U9351 ( n1077, WX663, n4503 );
and U9352 ( n1082, WX665, n4503 );
and U9353 ( n1087, WX667, n4503 );
and U9354 ( n1092, WX669, n4503 );
and U9355 ( n1097, WX671, n4502 );
and U9356 ( n1102, WX673, n4502 );
and U9357 ( n1107, WX675, n4502 );
and U9358 ( n1112, WX677, n4502 );
and U9359 ( n1117, WX679, n4502 );
and U9360 ( n1122, WX681, n4502 );
and U9361 ( n1127, WX683, n4502 );
and U9362 ( n1132, WX685, n4502 );
and U9363 ( n1137, WX687, n4502 );
and U9364 ( n1142, WX689, n4501 );
and U9365 ( n1147, WX691, n4502 );
and U9366 ( n1152, WX693, n4502 );
and U9367 ( n1157, WX695, n4501 );
and U9368 ( n1032, WX645, n4503 );
and U9369 ( n1347, WX771, n4498 );
and U9370 ( n1342, WX769, n4498 );
and U9371 ( n1337, WX767, n4498 );
and U9372 ( n1332, WX765, n4498 );
and U9373 ( n1327, WX763, n4499 );
and U9374 ( n1322, WX761, n4499 );
and U9375 ( n1197, WX711, n4501 );
and U9376 ( n1202, WX713, n4501 );
and U9377 ( n1207, WX715, n4501 );
and U9378 ( n1212, WX717, n4500 );
and U9379 ( n1217, WX719, n4500 );
and U9380 ( n1222, WX721, n4500 );
and U9381 ( n1227, WX723, n4500 );
and U9382 ( n1232, WX725, n4500 );
and U9383 ( n1237, WX727, n4500 );
and U9384 ( n1242, WX729, n4500 );
and U9385 ( n1247, WX731, n4500 );
and U9386 ( n1252, WX733, n4500 );
and U9387 ( n1257, WX735, n4500 );
and U9388 ( n1262, WX737, n4500 );
and U9389 ( n1267, WX739, n4500 );
and U9390 ( n1272, WX741, n4499 );
and U9391 ( n1277, WX743, n4499 );
and U9392 ( n1282, WX745, n4499 );
and U9393 ( n1287, WX747, n4499 );
and U9394 ( n1292, WX749, n4499 );
and U9395 ( n1297, WX751, n4499 );
and U9396 ( n1302, WX753, n4499 );
and U9397 ( n1307, WX755, n4499 );
and U9398 ( n1312, WX757, n4499 );
and U9399 ( n1317, WX759, n4499 );
and U9400 ( n1192, WX709, n4501 );
and U9401 ( n5987, n4535, WX7236 );
and U9402 ( n5982, n4535, WX7234 );
and U9403 ( n5977, n4535, WX7232 );
and U9404 ( n5972, n4535, WX7230 );
and U9405 ( n5967, n4535, WX7228 );
and U9406 ( n5962, n4535, WX7226 );
and U9407 ( n5957, n4535, WX7224 );
and U9408 ( n5952, n4535, WX7222 );
and U9409 ( n5947, n4535, WX7220 );
and U9410 ( n5942, n4535, WX7218 );
and U9411 ( n5937, n4535, WX7216 );
and U9412 ( n5932, n4535, WX7214 );
and U9413 ( n5927, n4536, WX7212 );
and U9414 ( n5922, n4536, WX7210 );
and U9415 ( n5917, n4536, WX7208 );
and U9416 ( n5912, n4536, WX7206 );
and U9417 ( n6865, n4526, WX8509 );
and U9418 ( n6860, n4527, WX8507 );
and U9419 ( n6855, n4528, WX8505 );
and U9420 ( n6850, n4526, WX8503 );
and U9421 ( n6845, n4527, WX8501 );
and U9422 ( n6840, n4526, WX8499 );
and U9423 ( n7843, n4539, WX9822 );
and U9424 ( n7838, n4539, WX9820 );
and U9425 ( n7833, n4539, WX9818 );
and U9426 ( n7828, n4539, WX9816 );
and U9427 ( n7823, n4539, WX9814 );
and U9428 ( n7818, n4539, WX9812 );
and U9429 ( n7813, n4539, WX9810 );
and U9430 ( n7808, n4539, WX9808 );
and U9431 ( n7803, n4539, WX9806 );
and U9432 ( n7798, n4539, WX9804 );
and U9433 ( n7793, n4539, WX9802 );
and U9434 ( n7788, n4539, WX9800 );
and U9435 ( n7783, n4539, WX9798 );
and U9436 ( n7778, n4540, WX9796 );
and U9437 ( n7773, n4540, WX9794 );
and U9438 ( n7768, n4540, WX9792 );
and U9439 ( n8771, n4526, WX11115 );
and U9440 ( n8766, n4527, WX11113 );
and U9441 ( n8761, n4526, WX11111 );
and U9442 ( n8756, n4526, WX11109 );
and U9443 ( n8751, n4529, WX11107 );
and U9444 ( n8746, n4527, WX11105 );
and U9445 ( n8741, n4526, WX11103 );
and U9446 ( n8736, n4527, WX11101 );
and U9447 ( n8731, n4527, WX11099 );
and U9448 ( n8726, n4527, WX11097 );
and U9449 ( n8721, n4528, WX11095 );
and U9450 ( n8716, n4527, WX11093 );
and U9451 ( n8711, n4527, WX11091 );
and U9452 ( n8706, n4528, WX11089 );
and U9453 ( n8701, n4527, WX11087 );
and U9454 ( n8696, n4527, WX11085 );
and U9455 ( n6147, n4532, WX7300 );
and U9456 ( n6142, n4532, WX7298 );
and U9457 ( n6137, n4532, WX7296 );
and U9458 ( n6132, n4532, WX7294 );
and U9459 ( n6127, n4532, WX7292 );
and U9460 ( n6122, n4532, WX7290 );
and U9461 ( n6117, n4532, WX7288 );
and U9462 ( n6112, n4532, WX7286 );
and U9463 ( n6107, n4532, WX7284 );
and U9464 ( n6102, n4532, WX7282 );
and U9465 ( n6097, n4532, WX7280 );
and U9466 ( n6092, n4533, WX7278 );
and U9467 ( n6087, n4533, WX7276 );
and U9468 ( n6082, n4533, WX7274 );
and U9469 ( n6077, n4533, WX7272 );
and U9470 ( n6072, n4533, WX7270 );
and U9471 ( n6067, n4533, WX7268 );
and U9472 ( n6062, n4533, WX7266 );
and U9473 ( n6057, n4534, WX7264 );
and U9474 ( n6052, n4534, WX7262 );
and U9475 ( n6047, n4534, WX7260 );
and U9476 ( n6042, n4534, WX7258 );
and U9477 ( n6037, n4534, WX7256 );
and U9478 ( n6032, n4534, WX7254 );
and U9479 ( n6027, n4534, WX7252 );
and U9480 ( n6022, n4534, WX7250 );
and U9481 ( n6017, n4534, WX7248 );
and U9482 ( n6012, n4534, WX7246 );
and U9483 ( n6007, n4534, WX7244 );
and U9484 ( n6002, n4534, WX7242 );
and U9485 ( n5997, n4534, WX7240 );
and U9486 ( n5992, n4535, WX7238 );
and U9487 ( n6675, n4528, WX8433 );
and U9488 ( n6670, n4529, WX8431 );
and U9489 ( n6665, n4528, WX8429 );
and U9490 ( n6660, n4528, WX8427 );
and U9491 ( n6655, n4529, WX8425 );
and U9492 ( n6650, n4529, WX8423 );
and U9493 ( n6645, n4529, WX8421 );
and U9494 ( n6640, n4529, WX8419 );
and U9495 ( n6635, n4529, WX8417 );
and U9496 ( n6630, n4529, WX8415 );
and U9497 ( n6625, n4529, WX8413 );
and U9498 ( n6620, n4529, WX8411 );
and U9499 ( n6615, n4529, WX8409 );
and U9500 ( n6610, n4530, WX8407 );
and U9501 ( n6605, n4530, WX8405 );
and U9502 ( n6600, n4530, WX8403 );
and U9503 ( n8003, n4528, WX9886 );
and U9504 ( n7993, n4536, WX9882 );
and U9505 ( n7988, n4536, WX9880 );
and U9506 ( n7983, n4536, WX9878 );
and U9507 ( n7978, n4536, WX9876 );
and U9508 ( n7973, n4537, WX9874 );
and U9509 ( n7968, n4537, WX9872 );
and U9510 ( n7963, n4537, WX9870 );
and U9511 ( n7958, n4537, WX9868 );
and U9512 ( n7953, n4537, WX9866 );
and U9513 ( n7948, n4537, WX9864 );
and U9514 ( n7943, n4537, WX9862 );
and U9515 ( n7938, n4537, WX9860 );
and U9516 ( n7933, n4537, WX9858 );
and U9517 ( n7928, n4537, WX9856 );
and U9518 ( n7923, n4537, WX9854 );
and U9519 ( n7918, n4537, WX9852 );
and U9520 ( n7913, n4537, WX9850 );
and U9521 ( n7908, n4538, WX9848 );
and U9522 ( n7903, n4538, WX9846 );
and U9523 ( n7898, n4538, WX9844 );
and U9524 ( n7893, n4538, WX9842 );
and U9525 ( n7888, n4538, WX9840 );
and U9526 ( n7883, n4538, WX9838 );
and U9527 ( n7878, n4538, WX9836 );
and U9528 ( n7873, n4538, WX9834 );
and U9529 ( n7868, n4538, WX9832 );
and U9530 ( n7863, n4538, WX9830 );
and U9531 ( n7858, n4538, WX9828 );
and U9532 ( n7853, n4538, WX9826 );
and U9533 ( n7848, n4538, WX9824 );
and U9534 ( n8776, n4530, WX11117 );
and U9535 ( n8926, n4536, WX11177 );
and U9536 ( n8921, n4533, WX11175 );
and U9537 ( n8916, n4533, WX11173 );
and U9538 ( n8911, n4533, WX11171 );
and U9539 ( n8906, n4533, WX11169 );
and U9540 ( n8901, n4533, WX11167 );
and U9541 ( n8896, n4533, WX11165 );
and U9542 ( n8891, n4532, WX11163 );
and U9543 ( n8886, n4532, WX11161 );
and U9544 ( n8881, n4531, WX11159 );
and U9545 ( n8876, n4531, WX11157 );
and U9546 ( n8871, n4531, WX11155 );
and U9547 ( n8866, n4531, WX11153 );
and U9548 ( n8861, n4531, WX11151 );
and U9549 ( n8856, n4531, WX11149 );
and U9550 ( n8851, n4531, WX11147 );
and U9551 ( n8846, n4531, WX11145 );
and U9552 ( n8841, n4531, WX11143 );
and U9553 ( n8836, n4531, WX11141 );
and U9554 ( n8831, n4531, WX11139 );
and U9555 ( n8826, n4531, WX11137 );
and U9556 ( n8821, n4531, WX11135 );
and U9557 ( n8816, n4530, WX11133 );
and U9558 ( n8811, n4530, WX11131 );
and U9559 ( n8806, n4530, WX11129 );
and U9560 ( n8801, n4525, WX11127 );
and U9561 ( n8796, n4530, WX11125 );
and U9562 ( n8791, n4530, WX11123 );
and U9563 ( n8786, n4530, WX11121 );
and U9564 ( n8781, n4530, WX11119 );
and U9565 ( n5907, n4536, WX7204 );
and U9566 ( n5902, n4536, WX7202 );
and U9567 ( n5897, n4536, WX7200 );
and U9568 ( n5892, n4536, WX7198 );
and U9569 ( n6755, n4525, WX8465 );
and U9570 ( n6750, n4525, WX8463 );
and U9571 ( n6745, n4526, WX8461 );
and U9572 ( n6740, n4525, WX8459 );
and U9573 ( n6725, n4525, WX8453 );
and U9574 ( n6715, n4527, WX8449 );
and U9575 ( n6710, n4528, WX8447 );
and U9576 ( n6705, n4528, WX8445 );
and U9577 ( n6700, n4528, WX8443 );
and U9578 ( n6695, n4529, WX8441 );
and U9579 ( n6690, n4528, WX8439 );
and U9580 ( n6685, n4529, WX8437 );
and U9581 ( n6680, n4528, WX8435 );
and U9582 ( n6835, n4525, WX8497 );
and U9583 ( n6830, n4527, WX8495 );
and U9584 ( n6825, n4525, WX8493 );
and U9585 ( n6820, n4525, WX8491 );
and U9586 ( n6815, n4526, WX8489 );
and U9587 ( n6810, n4525, WX8487 );
and U9588 ( n6805, n4525, WX8485 );
and U9589 ( n6800, n4526, WX8483 );
and U9590 ( n6795, n4528, WX8481 );
and U9591 ( n6790, n4526, WX8479 );
and U9592 ( n6785, n4525, WX8477 );
and U9593 ( n6780, n4526, WX8475 );
and U9594 ( n6775, n4526, WX8473 );
and U9595 ( n6770, n4525, WX8471 );
and U9596 ( n6765, n4525, WX8469 );
and U9597 ( n6760, n4530, WX8467 );
and U9598 ( n7763, n4540, WX9790 );
and U9599 ( n7758, n4540, WX9788 );
and U9600 ( n7753, n4540, WX9786 );
and U9601 ( n7748, n4540, WX9784 );
and U9602 ( n7743, n4540, WX9782 );
and U9603 ( n7738, n4540, WX9780 );
and U9604 ( n7733, n4540, WX9778 );
and U9605 ( n7728, n4540, WX9776 );
and U9606 ( n7723, n4540, WX9774 );
and U9607 ( n7718, n4540, WX9772 );
and U9608 ( n8691, n4530, WX11083 );
and U9609 ( n6735, n4524, WX8457 );
and U9610 ( n6730, n4524, WX8455 );
and U9611 ( n6720, n4524, WX8451 );
nor U9612 ( n867, WX485, n4675 );
nor U9613 ( n7363, WX9536, n4675 );
nor U9614 ( n6435, WX8243, n4673 );
nor U9615 ( n5507, WX6950, n4675 );
nor U9616 ( n4579, WX5657, n4675 );
nor U9617 ( n3651, WX4364, n4673 );
nor U9618 ( n2723, WX3071, n4673 );
nor U9619 ( n1795, WX1778, n4673 );
nor U9620 ( n8291, WX10829, n4673 );
nor U9621 ( n2440, n4655, n3677 );
xor U9622 ( n3677, WX2192, CRC_OUT_8_31 );
nor U9623 ( n3368, n4662, n3245 );
xor U9624 ( n3245, WX3485, CRC_OUT_7_31 );
nor U9625 ( n4296, n4665, n2782 );
xor U9626 ( n2782, WX4778, CRC_OUT_6_31 );
nor U9627 ( n5224, n4673, n2351 );
xor U9628 ( n2351, WX6071, CRC_OUT_5_31 );
nor U9629 ( n6152, n4637, n1888 );
xor U9630 ( n1888, WX7364, CRC_OUT_4_31 );
nor U9631 ( n7080, n4630, n1456 );
xor U9632 ( n1456, WX8657, CRC_OUT_3_31 );
nor U9633 ( n8008, n4641, n994 );
xor U9634 ( n994, WX9950, CRC_OUT_2_31 );
nor U9635 ( n8936, n4645, n616 );
xor U9636 ( n616, WX11243, CRC_OUT_1_31 );
nor U9637 ( n1632, n4655, n4150 );
xor U9638 ( n4150, WX839, CRC_OUT_9_29 );
nor U9639 ( n1628, n4655, n4152 );
xor U9640 ( n4152, WX841, CRC_OUT_9_28 );
nor U9641 ( n1624, n4655, n4153 );
xor U9642 ( n4153, WX843, CRC_OUT_9_27 );
nor U9643 ( n1620, n4653, n4154 );
xor U9644 ( n4154, WX845, CRC_OUT_9_26 );
nor U9645 ( n1616, n4653, n4155 );
xor U9646 ( n4155, WX847, CRC_OUT_9_25 );
nor U9647 ( n1612, n4653, n4157 );
xor U9648 ( n4157, WX849, CRC_OUT_9_24 );
nor U9649 ( n1608, n4653, n4158 );
xor U9650 ( n4158, WX851, CRC_OUT_9_23 );
nor U9651 ( n1604, n4653, n4159 );
xor U9652 ( n4159, WX853, CRC_OUT_9_22 );
nor U9653 ( n1600, n4652, n4160 );
xor U9654 ( n4160, WX855, CRC_OUT_9_21 );
nor U9655 ( n1596, n4652, n4162 );
xor U9656 ( n4162, WX857, CRC_OUT_9_20 );
nor U9657 ( n1592, n4652, n4163 );
xor U9658 ( n4163, WX859, CRC_OUT_9_19 );
nor U9659 ( n1588, n4652, n4164 );
xor U9660 ( n4164, WX861, CRC_OUT_9_18 );
nor U9661 ( n1584, n4652, n4165 );
xor U9662 ( n4165, WX863, CRC_OUT_9_17 );
nor U9663 ( n1580, n4651, n4167 );
xor U9664 ( n4167, WX865, CRC_OUT_9_16 );
nor U9665 ( n1576, n4651, n4168 );
xor U9666 ( n4168, CRC_OUT_9_15, n4169 );
xor U9667 ( n4169, WX867, CRC_OUT_9_31 );
nor U9668 ( n1572, n4651, n4170 );
xor U9669 ( n4170, WX869, CRC_OUT_9_14 );
nor U9670 ( n1568, n4651, n4172 );
xor U9671 ( n4172, WX871, CRC_OUT_9_13 );
nor U9672 ( n1564, n4651, n4173 );
xor U9673 ( n4173, WX873, CRC_OUT_9_12 );
nor U9674 ( n1560, n4650, n4174 );
xor U9675 ( n4174, WX875, CRC_OUT_9_11 );
nor U9676 ( n1556, n4650, n4175 );
xor U9677 ( n4175, CRC_OUT_9_10, n4177 );
xor U9678 ( n4177, WX877, CRC_OUT_9_31 );
nor U9679 ( n1552, n4650, n4178 );
xor U9680 ( n4178, WX879, CRC_OUT_9_9 );
nor U9681 ( n1548, n4650, n4179 );
xor U9682 ( n4179, WX881, CRC_OUT_9_8 );
nor U9683 ( n1544, n4650, n4180 );
xor U9684 ( n4180, WX883, CRC_OUT_9_7 );
nor U9685 ( n1540, n4648, n4182 );
xor U9686 ( n4182, WX885, CRC_OUT_9_6 );
nor U9687 ( n1536, n4648, n4183 );
xor U9688 ( n4183, WX887, CRC_OUT_9_5 );
nor U9689 ( n1532, n4648, n4184 );
xor U9690 ( n4184, WX889, CRC_OUT_9_4 );
nor U9691 ( n1528, n4648, n4185 );
xor U9692 ( n4185, CRC_OUT_9_3, n4187 );
xor U9693 ( n4187, WX891, CRC_OUT_9_31 );
nor U9694 ( n1524, n4648, n4188 );
xor U9695 ( n4188, WX893, CRC_OUT_9_2 );
nor U9696 ( n1520, n4647, n4189 );
xor U9697 ( n4189, WX895, CRC_OUT_9_1 );
nor U9698 ( n1516, n4662, n4190 );
xor U9699 ( n4190, WX897, CRC_OUT_9_0 );
nor U9700 ( n1636, n4655, n4149 );
xor U9701 ( n4149, WX837, CRC_OUT_9_30 );
nor U9702 ( n2560, n4661, n3638 );
xor U9703 ( n3638, WX2132, CRC_OUT_8_29 );
nor U9704 ( n2556, n4661, n3639 );
xor U9705 ( n3639, WX2134, CRC_OUT_8_28 );
nor U9706 ( n2552, n4661, n3640 );
xor U9707 ( n3640, WX2136, CRC_OUT_8_27 );
nor U9708 ( n2548, n4661, n3641 );
xor U9709 ( n3641, WX2138, CRC_OUT_8_26 );
nor U9710 ( n2544, n4661, n3642 );
xor U9711 ( n3642, WX2140, CRC_OUT_8_25 );
nor U9712 ( n2540, n4660, n3643 );
xor U9713 ( n3643, WX2142, CRC_OUT_8_24 );
nor U9714 ( n2536, n4660, n3644 );
xor U9715 ( n3644, WX2144, CRC_OUT_8_23 );
nor U9716 ( n2532, n4660, n3645 );
xor U9717 ( n3645, WX2146, CRC_OUT_8_22 );
nor U9718 ( n2528, n4660, n3646 );
xor U9719 ( n3646, WX2148, CRC_OUT_8_21 );
nor U9720 ( n2524, n4660, n3647 );
xor U9721 ( n3647, WX2150, CRC_OUT_8_20 );
nor U9722 ( n2520, n4658, n3648 );
xor U9723 ( n3648, WX2152, CRC_OUT_8_19 );
nor U9724 ( n2516, n4658, n3649 );
xor U9725 ( n3649, WX2154, CRC_OUT_8_18 );
nor U9726 ( n2512, n4658, n3650 );
xor U9727 ( n3650, WX2156, CRC_OUT_8_17 );
nor U9728 ( n2508, n4658, n3652 );
xor U9729 ( n3652, WX2158, CRC_OUT_8_16 );
nor U9730 ( n2504, n4658, n3653 );
xor U9731 ( n3653, CRC_OUT_8_15, n3654 );
xor U9732 ( n3654, WX2160, CRC_OUT_8_31 );
nor U9733 ( n2500, n4657, n3655 );
xor U9734 ( n3655, WX2162, CRC_OUT_8_14 );
nor U9735 ( n2496, n4657, n3657 );
xor U9736 ( n3657, WX2164, CRC_OUT_8_13 );
nor U9737 ( n2492, n4657, n3658 );
xor U9738 ( n3658, WX2166, CRC_OUT_8_12 );
nor U9739 ( n2488, n4657, n3659 );
xor U9740 ( n3659, WX2168, CRC_OUT_8_11 );
nor U9741 ( n2484, n4657, n3660 );
xor U9742 ( n3660, CRC_OUT_8_10, n3662 );
xor U9743 ( n3662, WX2170, CRC_OUT_8_31 );
nor U9744 ( n2480, n4656, n3663 );
xor U9745 ( n3663, WX2172, CRC_OUT_8_9 );
nor U9746 ( n2476, n4656, n3664 );
xor U9747 ( n3664, WX2174, CRC_OUT_8_8 );
nor U9748 ( n2472, n4656, n3665 );
xor U9749 ( n3665, WX2176, CRC_OUT_8_7 );
nor U9750 ( n2468, n4656, n3667 );
xor U9751 ( n3667, WX2178, CRC_OUT_8_6 );
nor U9752 ( n2464, n4656, n3668 );
xor U9753 ( n3668, WX2180, CRC_OUT_8_5 );
nor U9754 ( n2460, n4657, n3669 );
xor U9755 ( n3669, WX2182, CRC_OUT_8_4 );
nor U9756 ( n2456, n4656, n3670 );
xor U9757 ( n3670, CRC_OUT_8_3, n3672 );
xor U9758 ( n3672, WX2184, CRC_OUT_8_31 );
nor U9759 ( n2452, n4655, n3673 );
xor U9760 ( n3673, WX2186, CRC_OUT_8_2 );
nor U9761 ( n2448, n4648, n3674 );
xor U9762 ( n3674, WX2188, CRC_OUT_8_1 );
nor U9763 ( n2444, n4641, n3675 );
xor U9764 ( n3675, WX2190, CRC_OUT_8_0 );
nor U9765 ( n2564, n4673, n3637 );
xor U9766 ( n3637, WX2130, CRC_OUT_8_30 );
nor U9767 ( n3488, n4666, n3204 );
xor U9768 ( n3204, WX3425, CRC_OUT_7_29 );
nor U9769 ( n3484, n4666, n3205 );
xor U9770 ( n3205, WX3427, CRC_OUT_7_28 );
nor U9771 ( n3480, n4665, n3206 );
xor U9772 ( n3206, WX3429, CRC_OUT_7_27 );
nor U9773 ( n3476, n4666, n3207 );
xor U9774 ( n3207, WX3431, CRC_OUT_7_26 );
nor U9775 ( n3472, n4663, n3209 );
xor U9776 ( n3209, WX3433, CRC_OUT_7_25 );
nor U9777 ( n3468, n4665, n3210 );
xor U9778 ( n3210, WX3435, CRC_OUT_7_24 );
nor U9779 ( n3464, n4666, n3211 );
xor U9780 ( n3211, WX3437, CRC_OUT_7_23 );
nor U9781 ( n3460, n4666, n3212 );
xor U9782 ( n3212, WX3439, CRC_OUT_7_22 );
nor U9783 ( n3456, n4666, n3214 );
xor U9784 ( n3214, WX3441, CRC_OUT_7_21 );
nor U9785 ( n3452, n4665, n3215 );
xor U9786 ( n3215, WX3443, CRC_OUT_7_20 );
nor U9787 ( n3448, n4665, n3216 );
xor U9788 ( n3216, WX3445, CRC_OUT_7_19 );
nor U9789 ( n3444, n4665, n3217 );
xor U9790 ( n3217, WX3447, CRC_OUT_7_18 );
nor U9791 ( n3440, n4665, n3219 );
xor U9792 ( n3219, WX3449, CRC_OUT_7_17 );
nor U9793 ( n3436, n4663, n3220 );
xor U9794 ( n3220, WX3451, CRC_OUT_7_16 );
nor U9795 ( n3432, n4663, n3221 );
xor U9796 ( n3221, CRC_OUT_7_15, n3222 );
xor U9797 ( n3222, WX3453, CRC_OUT_7_31 );
nor U9798 ( n3428, n4663, n3224 );
xor U9799 ( n3224, WX3455, CRC_OUT_7_14 );
nor U9800 ( n3424, n4663, n3225 );
xor U9801 ( n3225, WX3457, CRC_OUT_7_13 );
nor U9802 ( n3420, n4663, n3226 );
xor U9803 ( n3226, WX3459, CRC_OUT_7_12 );
nor U9804 ( n3416, n4662, n3227 );
xor U9805 ( n3227, WX3461, CRC_OUT_7_11 );
nor U9806 ( n3412, n4662, n3229 );
xor U9807 ( n3229, CRC_OUT_7_10, n3230 );
xor U9808 ( n3230, WX3463, CRC_OUT_7_31 );
nor U9809 ( n3408, n4662, n3231 );
xor U9810 ( n3231, WX3465, CRC_OUT_7_9 );
nor U9811 ( n3404, n4662, n3232 );
xor U9812 ( n3232, WX3467, CRC_OUT_7_8 );
nor U9813 ( n3400, n4637, n3234 );
xor U9814 ( n3234, WX3469, CRC_OUT_7_7 );
nor U9815 ( n3396, n4638, n3235 );
xor U9816 ( n3235, WX3471, CRC_OUT_7_6 );
nor U9817 ( n3392, n4640, n3236 );
xor U9818 ( n3236, WX3473, CRC_OUT_7_5 );
nor U9819 ( n3388, n4641, n3237 );
xor U9820 ( n3237, WX3475, CRC_OUT_7_4 );
nor U9821 ( n3384, n4642, n3239 );
xor U9822 ( n3239, CRC_OUT_7_3, n3240 );
xor U9823 ( n3240, WX3477, CRC_OUT_7_31 );
nor U9824 ( n3380, n4661, n3241 );
xor U9825 ( n3241, WX3479, CRC_OUT_7_2 );
nor U9826 ( n3376, n4660, n3242 );
xor U9827 ( n3242, WX3481, CRC_OUT_7_1 );
nor U9828 ( n3372, n4662, n3244 );
xor U9829 ( n3244, WX3483, CRC_OUT_7_0 );
nor U9830 ( n3492, n4663, n3202 );
xor U9831 ( n3202, WX3423, CRC_OUT_7_30 );
nor U9832 ( n4416, n4668, n2741 );
xor U9833 ( n2741, WX4718, CRC_OUT_6_29 );
nor U9834 ( n4412, n4671, n2742 );
xor U9835 ( n2742, WX4720, CRC_OUT_6_28 );
nor U9836 ( n4408, n4671, n2744 );
xor U9837 ( n2744, WX4722, CRC_OUT_6_27 );
nor U9838 ( n4404, n4670, n2745 );
xor U9839 ( n2745, WX4724, CRC_OUT_6_26 );
nor U9840 ( n4400, n4671, n2746 );
xor U9841 ( n2746, WX4726, CRC_OUT_6_25 );
nor U9842 ( n4396, n4668, n2747 );
xor U9843 ( n2747, WX4728, CRC_OUT_6_24 );
nor U9844 ( n4392, n4667, n2749 );
xor U9845 ( n2749, WX4730, CRC_OUT_6_23 );
nor U9846 ( n4388, n4670, n2750 );
xor U9847 ( n2750, WX4732, CRC_OUT_6_22 );
nor U9848 ( n4384, n4652, n2751 );
xor U9849 ( n2751, WX4734, CRC_OUT_6_21 );
nor U9850 ( n4380, n4670, n2752 );
xor U9851 ( n2752, WX4736, CRC_OUT_6_20 );
nor U9852 ( n4376, n4667, n2754 );
xor U9853 ( n2754, WX4738, CRC_OUT_6_19 );
nor U9854 ( n4372, n4670, n2755 );
xor U9855 ( n2755, WX4740, CRC_OUT_6_18 );
nor U9856 ( n4368, n4670, n2756 );
xor U9857 ( n2756, WX4742, CRC_OUT_6_17 );
nor U9858 ( n4364, n4668, n2757 );
xor U9859 ( n2757, WX4744, CRC_OUT_6_16 );
nor U9860 ( n4360, n4670, n2759 );
xor U9861 ( n2759, CRC_OUT_6_15, n2760 );
xor U9862 ( n2760, WX4746, CRC_OUT_6_31 );
nor U9863 ( n4356, n4667, n2761 );
xor U9864 ( n2761, WX4748, CRC_OUT_6_14 );
nor U9865 ( n4352, n4670, n2762 );
xor U9866 ( n2762, WX4750, CRC_OUT_6_13 );
nor U9867 ( n4348, n4668, n2764 );
xor U9868 ( n2764, WX4752, CRC_OUT_6_12 );
nor U9869 ( n4344, n4668, n2765 );
xor U9870 ( n2765, WX4754, CRC_OUT_6_11 );
nor U9871 ( n4340, n4667, n2766 );
xor U9872 ( n2766, CRC_OUT_6_10, n2767 );
xor U9873 ( n2767, WX4756, CRC_OUT_6_31 );
nor U9874 ( n4336, n4668, n2769 );
xor U9875 ( n2769, WX4758, CRC_OUT_6_9 );
nor U9876 ( n4332, n4655, n2770 );
xor U9877 ( n2770, WX4760, CRC_OUT_6_8 );
nor U9878 ( n4328, n4668, n2771 );
xor U9879 ( n2771, WX4762, CRC_OUT_6_7 );
nor U9880 ( n4324, n4667, n2772 );
xor U9881 ( n2772, WX4764, CRC_OUT_6_6 );
nor U9882 ( n4320, n4667, n2774 );
xor U9883 ( n2774, WX4766, CRC_OUT_6_5 );
nor U9884 ( n4316, n4661, n2775 );
xor U9885 ( n2775, WX4768, CRC_OUT_6_4 );
nor U9886 ( n4312, n4667, n2776 );
xor U9887 ( n2776, CRC_OUT_6_3, n2777 );
xor U9888 ( n2777, WX4770, CRC_OUT_6_31 );
nor U9889 ( n4308, n4666, n2779 );
xor U9890 ( n2779, WX4772, CRC_OUT_6_2 );
nor U9891 ( n4304, n4660, n2780 );
xor U9892 ( n2780, WX4774, CRC_OUT_6_1 );
nor U9893 ( n4300, n4648, n2781 );
xor U9894 ( n2781, WX4776, CRC_OUT_6_0 );
nor U9895 ( n4420, n4653, n2740 );
xor U9896 ( n2740, WX4716, CRC_OUT_6_30 );
nor U9897 ( n5344, n4638, n2309 );
xor U9898 ( n2309, WX6011, CRC_OUT_5_29 );
nor U9899 ( n5340, n4637, n2311 );
xor U9900 ( n2311, WX6013, CRC_OUT_5_28 );
nor U9901 ( n5336, n4637, n2312 );
xor U9902 ( n2312, WX6015, CRC_OUT_5_27 );
nor U9903 ( n5332, n4637, n2313 );
xor U9904 ( n2313, WX6017, CRC_OUT_5_26 );
nor U9905 ( n5328, n4637, n2314 );
xor U9906 ( n2314, WX6019, CRC_OUT_5_25 );
nor U9907 ( n5324, n4637, n2316 );
xor U9908 ( n2316, WX6021, CRC_OUT_5_24 );
nor U9909 ( n5320, n4638, n2317 );
xor U9910 ( n2317, WX6023, CRC_OUT_5_23 );
nor U9911 ( n5316, n4638, n2318 );
xor U9912 ( n2318, WX6025, CRC_OUT_5_22 );
nor U9913 ( n5312, n4638, n2319 );
xor U9914 ( n2319, WX6027, CRC_OUT_5_21 );
nor U9915 ( n5308, n4638, n2321 );
xor U9916 ( n2321, WX6029, CRC_OUT_5_20 );
nor U9917 ( n5304, n4638, n2322 );
xor U9918 ( n2322, WX6031, CRC_OUT_5_19 );
nor U9919 ( n5300, n4640, n2323 );
xor U9920 ( n2323, WX6033, CRC_OUT_5_18 );
nor U9921 ( n5296, n4640, n2324 );
xor U9922 ( n2324, WX6035, CRC_OUT_5_17 );
nor U9923 ( n5292, n4640, n2326 );
xor U9924 ( n2326, WX6037, CRC_OUT_5_16 );
nor U9925 ( n5288, n4640, n2327 );
xor U9926 ( n2327, CRC_OUT_5_15, n2328 );
xor U9927 ( n2328, WX6039, CRC_OUT_5_31 );
nor U9928 ( n5284, n4640, n2329 );
xor U9929 ( n2329, WX6041, CRC_OUT_5_14 );
nor U9930 ( n5280, n4641, n2331 );
xor U9931 ( n2331, WX6043, CRC_OUT_5_13 );
nor U9932 ( n5276, n4651, n2332 );
xor U9933 ( n2332, WX6045, CRC_OUT_5_12 );
nor U9934 ( n5272, n4672, n2333 );
xor U9935 ( n2333, WX6047, CRC_OUT_5_11 );
nor U9936 ( n5268, n4652, n2334 );
xor U9937 ( n2334, CRC_OUT_5_10, n2336 );
xor U9938 ( n2336, WX6049, CRC_OUT_5_31 );
nor U9939 ( n5264, n4672, n2337 );
xor U9940 ( n2337, WX6051, CRC_OUT_5_9 );
nor U9941 ( n5260, n4651, n2338 );
xor U9942 ( n2338, WX6053, CRC_OUT_5_8 );
nor U9943 ( n5256, n4672, n2339 );
xor U9944 ( n2339, WX6055, CRC_OUT_5_7 );
nor U9945 ( n5252, n4650, n2341 );
xor U9946 ( n2341, WX6057, CRC_OUT_5_6 );
nor U9947 ( n5248, n4672, n2342 );
xor U9948 ( n2342, WX6059, CRC_OUT_5_5 );
nor U9949 ( n5244, n4671, n2343 );
xor U9950 ( n2343, WX6061, CRC_OUT_5_4 );
nor U9951 ( n5240, n4672, n2344 );
xor U9952 ( n2344, CRC_OUT_5_3, n2346 );
xor U9953 ( n2346, WX6063, CRC_OUT_5_31 );
nor U9954 ( n5236, n4671, n2347 );
xor U9955 ( n2347, WX6065, CRC_OUT_5_2 );
nor U9956 ( n5232, n4650, n2348 );
xor U9957 ( n2348, WX6067, CRC_OUT_5_1 );
nor U9958 ( n5228, n4653, n2349 );
xor U9959 ( n2349, WX6069, CRC_OUT_5_0 );
nor U9960 ( n5348, n4640, n2308 );
xor U9961 ( n2308, WX6009, CRC_OUT_5_30 );
nor U9962 ( n6272, n4632, n1847 );
xor U9963 ( n1847, WX7304, CRC_OUT_4_29 );
nor U9964 ( n6268, n4632, n1848 );
xor U9965 ( n1848, WX7306, CRC_OUT_4_28 );
nor U9966 ( n6264, n4632, n1849 );
xor U9967 ( n1849, WX7308, CRC_OUT_4_27 );
nor U9968 ( n6260, n4632, n1851 );
xor U9969 ( n1851, WX7310, CRC_OUT_4_26 );
nor U9970 ( n6256, n4633, n1852 );
xor U9971 ( n1852, WX7312, CRC_OUT_4_25 );
nor U9972 ( n6252, n4633, n1853 );
xor U9973 ( n1853, WX7314, CRC_OUT_4_24 );
nor U9974 ( n6248, n4633, n1854 );
xor U9975 ( n1854, WX7316, CRC_OUT_4_23 );
nor U9976 ( n6244, n4633, n1856 );
xor U9977 ( n1856, WX7318, CRC_OUT_4_22 );
nor U9978 ( n6240, n4633, n1857 );
xor U9979 ( n1857, WX7320, CRC_OUT_4_21 );
nor U9980 ( n6236, n4635, n1858 );
xor U9981 ( n1858, WX7322, CRC_OUT_4_20 );
nor U9982 ( n6232, n4636, n1859 );
xor U9983 ( n1859, WX7324, CRC_OUT_4_19 );
nor U9984 ( n6228, n4632, n1861 );
xor U9985 ( n1861, WX7326, CRC_OUT_4_18 );
nor U9986 ( n6224, n4646, n1862 );
xor U9987 ( n1862, WX7328, CRC_OUT_4_17 );
nor U9988 ( n6220, n4635, n1863 );
xor U9989 ( n1863, WX7330, CRC_OUT_4_16 );
nor U9990 ( n6216, n4635, n1864 );
xor U9991 ( n1864, CRC_OUT_4_15, n1866 );
xor U9992 ( n1866, WX7332, CRC_OUT_4_31 );
nor U9993 ( n6212, n4635, n1867 );
xor U9994 ( n1867, WX7334, CRC_OUT_4_14 );
nor U9995 ( n6208, n4635, n1868 );
xor U9996 ( n1868, WX7336, CRC_OUT_4_13 );
nor U9997 ( n6204, n4635, n1869 );
xor U9998 ( n1869, WX7338, CRC_OUT_4_12 );
nor U9999 ( n6200, n4636, n1871 );
xor U10000 ( n1871, WX7340, CRC_OUT_4_11 );
nor U10001 ( n6196, n4636, n1872 );
xor U10002 ( n1872, CRC_OUT_4_10, n1873 );
xor U10003 ( n1873, WX7342, CRC_OUT_4_31 );
nor U10004 ( n6192, n4636, n1874 );
xor U10005 ( n1874, WX7344, CRC_OUT_4_9 );
nor U10006 ( n6188, n4636, n1876 );
xor U10007 ( n1876, WX7346, CRC_OUT_4_8 );
nor U10008 ( n6184, n4636, n1877 );
xor U10009 ( n1877, WX7348, CRC_OUT_4_7 );
nor U10010 ( n6180, n4638, n1878 );
xor U10011 ( n1878, WX7350, CRC_OUT_4_6 );
nor U10012 ( n6176, n4640, n1879 );
xor U10013 ( n1879, WX7352, CRC_OUT_4_5 );
nor U10014 ( n6172, n4657, n1881 );
xor U10015 ( n1881, WX7354, CRC_OUT_4_4 );
nor U10016 ( n6168, n4656, n1882 );
xor U10017 ( n1882, CRC_OUT_4_3, n1883 );
xor U10018 ( n1883, WX7356, CRC_OUT_4_31 );
nor U10019 ( n6164, n4658, n1884 );
xor U10020 ( n1884, WX7358, CRC_OUT_4_2 );
nor U10021 ( n6160, n4637, n1886 );
xor U10022 ( n1886, WX7360, CRC_OUT_4_1 );
nor U10023 ( n6156, n4658, n1887 );
xor U10024 ( n1887, WX7362, CRC_OUT_4_0 );
nor U10025 ( n6276, n4632, n1846 );
xor U10026 ( n1846, WX7302, CRC_OUT_4_30 );
nor U10027 ( n7200, n4642, n1415 );
xor U10028 ( n1415, WX8597, CRC_OUT_3_29 );
nor U10029 ( n7196, n4642, n1416 );
xor U10030 ( n1416, WX8599, CRC_OUT_3_28 );
nor U10031 ( n7192, n4642, n1418 );
xor U10032 ( n1418, WX8601, CRC_OUT_3_27 );
nor U10033 ( n7188, n4642, n1419 );
xor U10034 ( n1419, WX8603, CRC_OUT_3_26 );
nor U10035 ( n7184, n4641, n1420 );
xor U10036 ( n1420, WX8605, CRC_OUT_3_25 );
nor U10037 ( n7180, n4641, n1421 );
xor U10038 ( n1421, WX8607, CRC_OUT_3_24 );
nor U10039 ( n7176, n4641, n1423 );
xor U10040 ( n1423, WX8609, CRC_OUT_3_23 );
nor U10041 ( n7172, n4641, n1424 );
xor U10042 ( n1424, WX8611, CRC_OUT_3_22 );
nor U10043 ( n7168, n4672, n1425 );
xor U10044 ( n1425, WX8613, CRC_OUT_3_21 );
nor U10045 ( n7156, n4628, n1429 );
xor U10046 ( n1429, WX8619, CRC_OUT_3_18 );
nor U10047 ( n7152, n4628, n1430 );
xor U10048 ( n1430, WX8621, CRC_OUT_3_17 );
nor U10049 ( n7148, n4628, n1431 );
xor U10050 ( n1431, WX8623, CRC_OUT_3_16 );
nor U10051 ( n7144, n4628, n1433 );
xor U10052 ( n1433, CRC_OUT_3_15, n1434 );
xor U10053 ( n1434, WX8625, CRC_OUT_3_31 );
nor U10054 ( n7140, n4628, n1435 );
xor U10055 ( n1435, WX8627, CRC_OUT_3_14 );
nor U10056 ( n7136, n4630, n1436 );
xor U10057 ( n1436, WX8629, CRC_OUT_3_13 );
nor U10058 ( n7132, n4630, n1438 );
xor U10059 ( n1438, WX8631, CRC_OUT_3_12 );
nor U10060 ( n7128, n4630, n1439 );
xor U10061 ( n1439, WX8633, CRC_OUT_3_11 );
nor U10062 ( n7124, n4630, n1440 );
xor U10063 ( n1440, CRC_OUT_3_10, n1441 );
xor U10064 ( n1441, WX8635, CRC_OUT_3_31 );
nor U10065 ( n7120, n4630, n1443 );
xor U10066 ( n1443, WX8637, CRC_OUT_3_9 );
nor U10067 ( n7116, n4631, n1444 );
xor U10068 ( n1444, WX8639, CRC_OUT_3_8 );
nor U10069 ( n7112, n4631, n1445 );
xor U10070 ( n1445, WX8641, CRC_OUT_3_7 );
nor U10071 ( n7108, n4631, n1446 );
xor U10072 ( n1446, WX8643, CRC_OUT_3_6 );
nor U10073 ( n7104, n4631, n1448 );
xor U10074 ( n1448, WX8645, CRC_OUT_3_5 );
nor U10075 ( n7100, n4631, n1449 );
xor U10076 ( n1449, WX8647, CRC_OUT_3_4 );
nor U10077 ( n7096, n4631, n1450 );
xor U10078 ( n1450, CRC_OUT_3_3, n1451 );
xor U10079 ( n1451, WX8649, CRC_OUT_3_31 );
nor U10080 ( n7092, n4645, n1453 );
xor U10081 ( n1453, WX8651, CRC_OUT_3_2 );
nor U10082 ( n7088, n4643, n1454 );
xor U10083 ( n1454, WX8653, CRC_OUT_3_1 );
nor U10084 ( n7084, n4647, n1455 );
xor U10085 ( n1455, WX8655, CRC_OUT_3_0 );
nor U10086 ( n7204, n4642, n1414 );
xor U10087 ( n1414, WX8595, CRC_OUT_3_30 );
nor U10088 ( n8128, n4643, n953 );
xor U10089 ( n953, WX9890, CRC_OUT_2_29 );
nor U10090 ( n8124, n4645, n954 );
xor U10091 ( n954, WX9892, CRC_OUT_2_28 );
nor U10092 ( n8120, n4645, n955 );
xor U10093 ( n955, WX9894, CRC_OUT_2_27 );
nor U10094 ( n8116, n4645, n956 );
xor U10095 ( n956, WX9896, CRC_OUT_2_26 );
nor U10096 ( n8112, n4645, n958 );
xor U10097 ( n958, WX9898, CRC_OUT_2_25 );
nor U10098 ( n8108, n4645, n959 );
xor U10099 ( n959, WX9900, CRC_OUT_2_24 );
nor U10100 ( n8104, n4643, n960 );
xor U10101 ( n960, WX9902, CRC_OUT_2_23 );
nor U10102 ( n8100, n4643, n961 );
xor U10103 ( n961, WX9904, CRC_OUT_2_22 );
nor U10104 ( n8096, n4643, n963 );
xor U10105 ( n963, WX9906, CRC_OUT_2_21 );
nor U10106 ( n8092, n4643, n964 );
xor U10107 ( n964, WX9908, CRC_OUT_2_20 );
nor U10108 ( n8088, n4643, n965 );
xor U10109 ( n965, WX9910, CRC_OUT_2_19 );
nor U10110 ( n8084, n4645, n966 );
xor U10111 ( n966, WX9912, CRC_OUT_2_18 );
nor U10112 ( n8080, n4643, n968 );
xor U10113 ( n968, WX9914, CRC_OUT_2_17 );
nor U10114 ( n8076, n4667, n969 );
xor U10115 ( n969, WX9916, CRC_OUT_2_16 );
nor U10116 ( n8072, n4641, n970 );
xor U10117 ( n970, CRC_OUT_2_15, n971 );
xor U10118 ( n971, WX9918, CRC_OUT_2_31 );
nor U10119 ( n8068, n4642, n973 );
xor U10120 ( n973, WX9920, CRC_OUT_2_14 );
nor U10121 ( n8064, n4666, n974 );
xor U10122 ( n974, WX9922, CRC_OUT_2_13 );
nor U10123 ( n8060, n4665, n975 );
xor U10124 ( n975, WX9924, CRC_OUT_2_12 );
nor U10125 ( n8056, n4663, n976 );
xor U10126 ( n976, WX9926, CRC_OUT_2_11 );
nor U10127 ( n8052, n4670, n978 );
xor U10128 ( n978, CRC_OUT_2_10, n979 );
xor U10129 ( n979, WX9928, CRC_OUT_2_31 );
nor U10130 ( n8048, n4668, n980 );
xor U10131 ( n980, WX9930, CRC_OUT_2_9 );
nor U10132 ( n8044, n4642, n981 );
xor U10133 ( n981, WX9932, CRC_OUT_2_8 );
nor U10134 ( n8040, n4641, n983 );
xor U10135 ( n983, WX9934, CRC_OUT_2_7 );
nor U10136 ( n8036, n4672, n984 );
xor U10137 ( n984, WX9936, CRC_OUT_2_6 );
nor U10138 ( n8032, n4671, n985 );
xor U10139 ( n985, WX9938, CRC_OUT_2_5 );
nor U10140 ( n8028, n4671, n986 );
xor U10141 ( n986, WX9940, CRC_OUT_2_4 );
nor U10142 ( n8024, n4642, n988 );
xor U10143 ( n988, CRC_OUT_2_3, n989 );
xor U10144 ( n989, WX9942, CRC_OUT_2_31 );
nor U10145 ( n8020, n4642, n990 );
xor U10146 ( n990, WX9944, CRC_OUT_2_2 );
nor U10147 ( n8016, n4641, n991 );
xor U10148 ( n991, WX9946, CRC_OUT_2_1 );
nor U10149 ( n8012, n4633, n993 );
xor U10150 ( n993, WX9948, CRC_OUT_2_0 );
nor U10151 ( n8132, n4643, n951 );
xor U10152 ( n951, WX9888, CRC_OUT_2_30 );
nor U10153 ( n9056, n4646, n561 );
xor U10154 ( n561, WX11183, CRC_OUT_1_29 );
nor U10155 ( n9052, n4646, n562 );
xor U10156 ( n562, WX11185, CRC_OUT_1_28 );
nor U10157 ( n9048, n4647, n563 );
xor U10158 ( n563, WX11187, CRC_OUT_1_27 );
nor U10159 ( n9044, n4647, n564 );
xor U10160 ( n564, WX11189, CRC_OUT_1_26 );
nor U10161 ( n9040, n4647, n565 );
xor U10162 ( n565, WX11191, CRC_OUT_1_25 );
nor U10163 ( n9036, n4647, n566 );
xor U10164 ( n566, WX11193, CRC_OUT_1_24 );
nor U10165 ( n9032, n4647, n567 );
xor U10166 ( n567, WX11195, CRC_OUT_1_23 );
nor U10167 ( n9028, n4647, n568 );
xor U10168 ( n568, WX11197, CRC_OUT_1_22 );
nor U10169 ( n9024, n4646, n569 );
xor U10170 ( n569, WX11199, CRC_OUT_1_21 );
nor U10171 ( n9020, n4646, n570 );
xor U10172 ( n570, WX11201, CRC_OUT_1_20 );
nor U10173 ( n9016, n4646, n582 );
xor U10174 ( n582, WX11203, CRC_OUT_1_19 );
nor U10175 ( n9012, n4646, n583 );
xor U10176 ( n583, WX11205, CRC_OUT_1_18 );
nor U10177 ( n9008, n4646, n584 );
xor U10178 ( n584, WX11207, CRC_OUT_1_17 );
nor U10179 ( n9004, n4647, n585 );
xor U10180 ( n585, WX11209, CRC_OUT_1_16 );
nor U10181 ( n9000, n4646, n586 );
xor U10182 ( n586, CRC_OUT_1_15, n587 );
xor U10183 ( n587, WX11211, CRC_OUT_1_31 );
nor U10184 ( n8996, n4661, n588 );
xor U10185 ( n588, WX11213, CRC_OUT_1_14 );
nor U10186 ( n8992, n4660, n589 );
xor U10187 ( n589, WX11215, CRC_OUT_1_13 );
nor U10188 ( n8988, n4662, n590 );
xor U10189 ( n590, WX11217, CRC_OUT_1_12 );
nor U10190 ( n8984, n4646, n591 );
xor U10191 ( n591, WX11219, CRC_OUT_1_11 );
nor U10192 ( n8980, n4647, n592 );
xor U10193 ( n592, CRC_OUT_1_10, n593 );
xor U10194 ( n593, WX11221, CRC_OUT_1_31 );
nor U10195 ( n8976, n4630, n594 );
xor U10196 ( n594, WX11223, CRC_OUT_1_9 );
nor U10197 ( n8972, n4631, n595 );
xor U10198 ( n595, WX11225, CRC_OUT_1_8 );
nor U10199 ( n8968, n4628, n607 );
xor U10200 ( n607, WX11227, CRC_OUT_1_7 );
nor U10201 ( n8964, n4643, n608 );
xor U10202 ( n608, WX11229, CRC_OUT_1_6 );
nor U10203 ( n8960, n4645, n609 );
xor U10204 ( n609, WX11231, CRC_OUT_1_5 );
nor U10205 ( n8956, n4635, n610 );
xor U10206 ( n610, WX11233, CRC_OUT_1_4 );
nor U10207 ( n8952, n4636, n611 );
xor U10208 ( n611, CRC_OUT_1_3, n612 );
xor U10209 ( n612, WX11235, CRC_OUT_1_31 );
nor U10210 ( n8948, n4632, n613 );
xor U10211 ( n613, WX11237, CRC_OUT_1_2 );
nor U10212 ( n8944, n4645, n614 );
xor U10213 ( n614, WX11239, CRC_OUT_1_1 );
nor U10214 ( n8940, n4633, n615 );
xor U10215 ( n615, WX11241, CRC_OUT_1_0 );
nor U10216 ( n9060, n4628, n560 );
xor U10217 ( n560, WX11181, CRC_OUT_1_30 );
nor U10218 ( n1512, n4627, n4192 );
xor U10219 ( n4192, WX899, CRC_OUT_9_31 );
nor U10220 ( n7164, n4627, n1426 );
xor U10221 ( n1426, WX8615, CRC_OUT_3_20 );
nor U10222 ( n7160, n4627, n1428 );
xor U10223 ( n1428, WX8617, CRC_OUT_3_19 );
xor U10224 ( n3688, n4198, n4199 );
xnor U10225 ( n4198, WX2000, WX2064 );
xor U10226 ( n4199, WX2192, WX2128 );
xor U10227 ( n3700, n4212, n4213 );
xnor U10228 ( n4212, WX1998, WX2062 );
xor U10229 ( n4213, WX2190, WX2126 );
xor U10230 ( n3713, n4225, n4227 );
xnor U10231 ( n4225, WX1996, WX2060 );
xor U10232 ( n4227, WX2188, WX2124 );
xor U10233 ( n3725, n4239, n4240 );
xnor U10234 ( n4239, WX1994, WX2058 );
xor U10235 ( n4240, WX2186, WX2122 );
xor U10236 ( n3738, n4253, n4254 );
xnor U10237 ( n4253, WX1992, WX2056 );
xor U10238 ( n4254, WX2184, WX2120 );
xor U10239 ( n3750, n4268, n4269 );
xnor U10240 ( n4268, WX1990, WX2054 );
xor U10241 ( n4269, WX2182, WX2118 );
xor U10242 ( n353, n3763, n3764 );
xnor U10243 ( n3763, WX1988, WX2052 );
xor U10244 ( n3764, WX2180, WX2116 );
xor U10245 ( n366, n3777, n3778 );
xnor U10246 ( n3777, WX1986, WX2050 );
xor U10247 ( n3778, WX2178, WX2114 );
xor U10248 ( n377, n3790, n3792 );
xnor U10249 ( n3790, WX1984, WX2048 );
xor U10250 ( n3792, WX2176, WX2112 );
xor U10251 ( n388, n3804, n3805 );
xnor U10252 ( n3804, WX1982, WX2046 );
xor U10253 ( n3805, WX2174, WX2110 );
xor U10254 ( n399, n3818, n3819 );
xnor U10255 ( n3818, WX1980, WX2044 );
xor U10256 ( n3819, WX2172, WX2108 );
xor U10257 ( n410, n3832, n3833 );
xnor U10258 ( n3832, WX1978, WX2042 );
xor U10259 ( n3833, WX2170, WX2106 );
xor U10260 ( n421, n3845, n3847 );
xnor U10261 ( n3845, WX1976, WX2040 );
xor U10262 ( n3847, WX2168, WX2104 );
xor U10263 ( n432, n3859, n3860 );
xnor U10264 ( n3859, WX1974, WX2038 );
xor U10265 ( n3860, WX2166, WX2102 );
xor U10266 ( n443, n3873, n3874 );
xnor U10267 ( n3873, WX1972, WX2036 );
xor U10268 ( n3874, WX2164, WX2100 );
xor U10269 ( n454, n3887, n3888 );
xnor U10270 ( n3887, WX1970, WX2034 );
xor U10271 ( n3888, WX2162, WX2098 );
xor U10272 ( n3256, n3683, n3684 );
xnor U10273 ( n3683, WX3293, WX3357 );
xor U10274 ( n3684, WX3485, WX3421 );
xor U10275 ( n3269, n3695, n3697 );
xnor U10276 ( n3695, WX3291, WX3355 );
xor U10277 ( n3697, WX3483, WX3419 );
xor U10278 ( n3281, n3708, n3709 );
xnor U10279 ( n3708, WX3289, WX3353 );
xor U10280 ( n3709, WX3481, WX3417 );
xor U10281 ( n3294, n3720, n3722 );
xnor U10282 ( n3720, WX3287, WX3351 );
xor U10283 ( n3722, WX3479, WX3415 );
xor U10284 ( n3306, n3733, n3734 );
xnor U10285 ( n3733, WX3285, WX3349 );
xor U10286 ( n3734, WX3477, WX3413 );
xor U10287 ( n3319, n3745, n3747 );
xnor U10288 ( n3745, WX3283, WX3347 );
xor U10289 ( n3747, WX3475, WX3411 );
xor U10290 ( n3331, n3758, n3759 );
xnor U10291 ( n3758, WX3281, WX3345 );
xor U10292 ( n3759, WX3473, WX3409 );
xor U10293 ( n3344, n3772, n3773 );
xnor U10294 ( n3772, WX3279, WX3343 );
xor U10295 ( n3773, WX3471, WX3407 );
xor U10296 ( n3356, n3785, n3787 );
xnor U10297 ( n3785, WX3277, WX3341 );
xor U10298 ( n3787, WX3469, WX3405 );
xor U10299 ( n3369, n3799, n3800 );
xnor U10300 ( n3799, WX3275, WX3339 );
xor U10301 ( n3800, WX3467, WX3403 );
xor U10302 ( n3382, n3813, n3814 );
xnor U10303 ( n3813, WX3273, WX3337 );
xor U10304 ( n3814, WX3465, WX3401 );
xor U10305 ( n3395, n3827, n3828 );
xnor U10306 ( n3827, WX3271, WX3335 );
xor U10307 ( n3828, WX3463, WX3399 );
xor U10308 ( n3409, n3840, n3842 );
xnor U10309 ( n3840, WX3269, WX3333 );
xor U10310 ( n3842, WX3461, WX3397 );
xor U10311 ( n3422, n3854, n3855 );
xnor U10312 ( n3854, WX3267, WX3331 );
xor U10313 ( n3855, WX3459, WX3395 );
xor U10314 ( n3435, n3868, n3869 );
xnor U10315 ( n3868, WX3265, WX3329 );
xor U10316 ( n3869, WX3457, WX3393 );
xor U10317 ( n3449, n3882, n3883 );
xnor U10318 ( n3882, WX3263, WX3327 );
xor U10319 ( n3883, WX3455, WX3391 );
xor U10320 ( n2794, n3251, n3252 );
xnor U10321 ( n3251, WX4586, WX4650 );
xor U10322 ( n3252, WX4778, WX4714 );
xor U10323 ( n2806, n3264, n3265 );
xnor U10324 ( n3264, WX4584, WX4648 );
xor U10325 ( n3265, WX4776, WX4712 );
xor U10326 ( n2819, n3276, n3277 );
xnor U10327 ( n3276, WX4582, WX4646 );
xor U10328 ( n3277, WX4774, WX4710 );
xor U10329 ( n2831, n3289, n3290 );
xnor U10330 ( n3289, WX4580, WX4644 );
xor U10331 ( n3290, WX4772, WX4708 );
xor U10332 ( n2844, n3301, n3302 );
xnor U10333 ( n3301, WX4578, WX4642 );
xor U10334 ( n3302, WX4770, WX4706 );
xor U10335 ( n2856, n3314, n3315 );
xnor U10336 ( n3314, WX4576, WX4640 );
xor U10337 ( n3315, WX4768, WX4704 );
xor U10338 ( n2869, n3326, n3327 );
xnor U10339 ( n3326, WX4574, WX4638 );
xor U10340 ( n3327, WX4766, WX4702 );
xor U10341 ( n2881, n3339, n3340 );
xnor U10342 ( n3339, WX4572, WX4636 );
xor U10343 ( n3340, WX4764, WX4700 );
xor U10344 ( n2894, n3351, n3352 );
xnor U10345 ( n3351, WX4570, WX4634 );
xor U10346 ( n3352, WX4762, WX4698 );
xor U10347 ( n2906, n3364, n3365 );
xnor U10348 ( n3364, WX4568, WX4632 );
xor U10349 ( n3365, WX4760, WX4696 );
xor U10350 ( n2919, n3377, n3378 );
xnor U10351 ( n3377, WX4566, WX4630 );
xor U10352 ( n3378, WX4758, WX4694 );
xor U10353 ( n2931, n3390, n3391 );
xnor U10354 ( n3390, WX4564, WX4628 );
xor U10355 ( n3391, WX4756, WX4692 );
xor U10356 ( n2944, n3403, n3405 );
xnor U10357 ( n3403, WX4562, WX4626 );
xor U10358 ( n3405, WX4754, WX4690 );
xor U10359 ( n2956, n3417, n3418 );
xnor U10360 ( n3417, WX4560, WX4624 );
xor U10361 ( n3418, WX4752, WX4688 );
xor U10362 ( n2969, n3430, n3431 );
xnor U10363 ( n3430, WX4558, WX4622 );
xor U10364 ( n3431, WX4750, WX4686 );
xor U10365 ( n2981, n3443, n3445 );
xnor U10366 ( n3443, WX4556, WX4620 );
xor U10367 ( n3445, WX4748, WX4684 );
xor U10368 ( n2362, n2789, n2790 );
xnor U10369 ( n2789, WX5879, WX5943 );
xor U10370 ( n2790, WX6071, WX6007 );
xor U10371 ( n2374, n2801, n2802 );
xnor U10372 ( n2801, WX5877, WX5941 );
xor U10373 ( n2802, WX6069, WX6005 );
xor U10374 ( n2387, n2814, n2815 );
xnor U10375 ( n2814, WX5875, WX5939 );
xor U10376 ( n2815, WX6067, WX6003 );
xor U10377 ( n2399, n2826, n2827 );
xnor U10378 ( n2826, WX5873, WX5937 );
xor U10379 ( n2827, WX6065, WX6001 );
xor U10380 ( n2412, n2839, n2840 );
xnor U10381 ( n2839, WX5871, WX5935 );
xor U10382 ( n2840, WX6063, WX5999 );
xor U10383 ( n2424, n2851, n2852 );
xnor U10384 ( n2851, WX5869, WX5933 );
xor U10385 ( n2852, WX6061, WX5997 );
xor U10386 ( n2437, n2864, n2865 );
xnor U10387 ( n2864, WX5867, WX5931 );
xor U10388 ( n2865, WX6059, WX5995 );
xor U10389 ( n2450, n2876, n2877 );
xnor U10390 ( n2876, WX5865, WX5929 );
xor U10391 ( n2877, WX6057, WX5993 );
xor U10392 ( n2463, n2889, n2890 );
xnor U10393 ( n2889, WX5863, WX5927 );
xor U10394 ( n2890, WX6055, WX5991 );
xor U10395 ( n2477, n2901, n2902 );
xnor U10396 ( n2901, WX5861, WX5925 );
xor U10397 ( n2902, WX6053, WX5989 );
xor U10398 ( n2490, n2914, n2915 );
xnor U10399 ( n2914, WX5859, WX5923 );
xor U10400 ( n2915, WX6051, WX5987 );
xor U10401 ( n2503, n2926, n2927 );
xnor U10402 ( n2926, WX5857, WX5921 );
xor U10403 ( n2927, WX6049, WX5985 );
xor U10404 ( n2517, n2939, n2940 );
xnor U10405 ( n2939, WX5855, WX5919 );
xor U10406 ( n2940, WX6047, WX5983 );
xor U10407 ( n2530, n2951, n2952 );
xnor U10408 ( n2951, WX5853, WX5917 );
xor U10409 ( n2952, WX6045, WX5981 );
xor U10410 ( n2543, n2964, n2965 );
xnor U10411 ( n2964, WX5851, WX5915 );
xor U10412 ( n2965, WX6043, WX5979 );
xor U10413 ( n2557, n2976, n2977 );
xnor U10414 ( n2976, WX5849, WX5913 );
xor U10415 ( n2977, WX6041, WX5977 );
xor U10416 ( n1899, n2357, n2358 );
xnor U10417 ( n2357, WX7172, WX7236 );
xor U10418 ( n2358, WX7364, WX7300 );
xor U10419 ( n1912, n2369, n2371 );
xnor U10420 ( n2369, WX7170, WX7234 );
xor U10421 ( n2371, WX7362, WX7298 );
xor U10422 ( n1924, n2382, n2383 );
xnor U10423 ( n2382, WX7168, WX7232 );
xor U10424 ( n2383, WX7360, WX7296 );
xor U10425 ( n1937, n2394, n2396 );
xnor U10426 ( n2394, WX7166, WX7230 );
xor U10427 ( n2396, WX7358, WX7294 );
xor U10428 ( n1949, n2407, n2408 );
xnor U10429 ( n2407, WX7164, WX7228 );
xor U10430 ( n2408, WX7356, WX7292 );
xor U10431 ( n1962, n2419, n2421 );
xnor U10432 ( n2419, WX7162, WX7226 );
xor U10433 ( n2421, WX7354, WX7290 );
xor U10434 ( n1974, n2432, n2433 );
xnor U10435 ( n2432, WX7160, WX7224 );
xor U10436 ( n2433, WX7352, WX7288 );
xor U10437 ( n1987, n2445, n2446 );
xnor U10438 ( n2445, WX7158, WX7222 );
xor U10439 ( n2446, WX7350, WX7286 );
xor U10440 ( n1999, n2458, n2459 );
xnor U10441 ( n2458, WX7156, WX7220 );
xor U10442 ( n2459, WX7348, WX7284 );
xor U10443 ( n2012, n2471, n2473 );
xnor U10444 ( n2471, WX7154, WX7218 );
xor U10445 ( n2473, WX7346, WX7282 );
xor U10446 ( n2024, n2485, n2486 );
xnor U10447 ( n2485, WX7152, WX7216 );
xor U10448 ( n2486, WX7344, WX7280 );
xor U10449 ( n2037, n2498, n2499 );
xnor U10450 ( n2498, WX7150, WX7214 );
xor U10451 ( n2499, WX7342, WX7278 );
xor U10452 ( n2049, n2511, n2513 );
xnor U10453 ( n2511, WX7148, WX7212 );
xor U10454 ( n2513, WX7340, WX7276 );
xor U10455 ( n2062, n2525, n2526 );
xnor U10456 ( n2525, WX7146, WX7210 );
xor U10457 ( n2526, WX7338, WX7274 );
xor U10458 ( n2074, n2538, n2539 );
xnor U10459 ( n2538, WX7144, WX7208 );
xor U10460 ( n2539, WX7336, WX7272 );
xor U10461 ( n2087, n2551, n2553 );
xnor U10462 ( n2551, WX7142, WX7206 );
xor U10463 ( n2553, WX7334, WX7270 );
xor U10464 ( n1468, n1894, n1896 );
xnor U10465 ( n1894, WX8465, WX8529 );
xor U10466 ( n1896, WX8657, WX8593 );
xor U10467 ( n1480, n1907, n1908 );
xnor U10468 ( n1907, WX8463, WX8527 );
xor U10469 ( n1908, WX8655, WX8591 );
xor U10470 ( n1493, n1919, n1921 );
xnor U10471 ( n1919, WX8461, WX8525 );
xor U10472 ( n1921, WX8653, WX8589 );
xor U10473 ( n1505, n1932, n1933 );
xnor U10474 ( n1932, WX8459, WX8523 );
xor U10475 ( n1933, WX8651, WX8587 );
xor U10476 ( n1518, n1944, n1946 );
xnor U10477 ( n1944, WX8457, WX8521 );
xor U10478 ( n1946, WX8649, WX8585 );
xor U10479 ( n1531, n1957, n1958 );
xnor U10480 ( n1957, WX8455, WX8519 );
xor U10481 ( n1958, WX8647, WX8583 );
xor U10482 ( n1545, n1969, n1971 );
xnor U10483 ( n1969, WX8453, WX8517 );
xor U10484 ( n1971, WX8645, WX8581 );
xor U10485 ( n1558, n1982, n1983 );
xnor U10486 ( n1982, WX8451, WX8515 );
xor U10487 ( n1983, WX8643, WX8579 );
xor U10488 ( n1571, n1994, n1996 );
xnor U10489 ( n1994, WX8449, WX8513 );
xor U10490 ( n1996, WX8641, WX8577 );
xor U10491 ( n1585, n2007, n2008 );
xnor U10492 ( n2007, WX8447, WX8511 );
xor U10493 ( n2008, WX8639, WX8575 );
xor U10494 ( n1598, n2019, n2021 );
xnor U10495 ( n2019, WX8445, WX8509 );
xor U10496 ( n2021, WX8637, WX8573 );
xor U10497 ( n1611, n2032, n2033 );
xnor U10498 ( n2032, WX8443, WX8507 );
xor U10499 ( n2033, WX8635, WX8571 );
xor U10500 ( n1625, n2044, n2046 );
xnor U10501 ( n2044, WX8441, WX8505 );
xor U10502 ( n2046, WX8633, WX8569 );
xor U10503 ( n1638, n2057, n2058 );
xnor U10504 ( n2057, WX8439, WX8503 );
xor U10505 ( n2058, WX8631, WX8567 );
xor U10506 ( n1648, n2069, n2071 );
xnor U10507 ( n2069, WX8437, WX8501 );
xor U10508 ( n2071, WX8629, WX8565 );
xor U10509 ( n1658, n2082, n2083 );
xnor U10510 ( n2082, WX8435, WX8499 );
xor U10511 ( n2083, WX8627, WX8563 );
xor U10512 ( n1005, n1463, n1464 );
xnor U10513 ( n1463, WX9758, WX9822 );
xor U10514 ( n1464, WX9950, WX9886 );
xor U10515 ( n1018, n1475, n1476 );
xnor U10516 ( n1475, WX9756, WX9820 );
xor U10517 ( n1476, WX9948, WX9884 );
xor U10518 ( n1030, n1488, n1489 );
xnor U10519 ( n1488, WX9754, WX9818 );
xor U10520 ( n1489, WX9946, WX9882 );
xor U10521 ( n1043, n1500, n1501 );
xnor U10522 ( n1500, WX9752, WX9816 );
xor U10523 ( n1501, WX9944, WX9880 );
xor U10524 ( n1055, n1513, n1514 );
xnor U10525 ( n1513, WX9750, WX9814 );
xor U10526 ( n1514, WX9942, WX9878 );
xor U10527 ( n1068, n1526, n1527 );
xnor U10528 ( n1526, WX9748, WX9812 );
xor U10529 ( n1527, WX9940, WX9876 );
xor U10530 ( n1080, n1539, n1541 );
xnor U10531 ( n1539, WX9746, WX9810 );
xor U10532 ( n1541, WX9938, WX9874 );
xor U10533 ( n1093, n1553, n1554 );
xnor U10534 ( n1553, WX9744, WX9808 );
xor U10535 ( n1554, WX9936, WX9872 );
xor U10536 ( n1105, n1566, n1567 );
xnor U10537 ( n1566, WX9742, WX9806 );
xor U10538 ( n1567, WX9934, WX9870 );
xor U10539 ( n1118, n1579, n1581 );
xnor U10540 ( n1579, WX9740, WX9804 );
xor U10541 ( n1581, WX9932, WX9868 );
xor U10542 ( n1130, n1593, n1594 );
xnor U10543 ( n1593, WX9738, WX9802 );
xor U10544 ( n1594, WX9930, WX9866 );
xor U10545 ( n1143, n1606, n1607 );
xnor U10546 ( n1606, WX9736, WX9800 );
xor U10547 ( n1607, WX9928, WX9864 );
xor U10548 ( n1155, n1619, n1621 );
xnor U10549 ( n1619, WX9734, WX9798 );
xor U10550 ( n1621, WX9926, WX9862 );
xor U10551 ( n1168, n1633, n1634 );
xnor U10552 ( n1633, WX9732, WX9796 );
xor U10553 ( n1634, WX9924, WX9860 );
xor U10554 ( n1180, n1644, n1645 );
xnor U10555 ( n1644, WX9730, WX9794 );
xor U10556 ( n1645, WX9922, WX9858 );
xor U10557 ( n1193, n1654, n1655 );
xnor U10558 ( n1654, WX9728, WX9792 );
xor U10559 ( n1655, WX9920, WX9856 );
xor U10560 ( n683, n1000, n1001 );
xnor U10561 ( n1000, WX11051, WX11115 );
xor U10562 ( n1001, WX11243, WX11179 );
xor U10563 ( n691, n1013, n1014 );
xnor U10564 ( n1013, WX11049, WX11113 );
xor U10565 ( n1014, WX11241, WX11177 );
xor U10566 ( n699, n1025, n1026 );
xnor U10567 ( n1025, WX11047, WX11111 );
xor U10568 ( n1026, WX11239, WX11175 );
xor U10569 ( n707, n1038, n1039 );
xnor U10570 ( n1038, WX11045, WX11109 );
xor U10571 ( n1039, WX11237, WX11173 );
xor U10572 ( n715, n1050, n1051 );
xnor U10573 ( n1050, WX11043, WX11107 );
xor U10574 ( n1051, WX11235, WX11171 );
xor U10575 ( n723, n1063, n1064 );
xnor U10576 ( n1063, WX11041, WX11105 );
xor U10577 ( n1064, WX11233, WX11169 );
xor U10578 ( n731, n1075, n1076 );
xnor U10579 ( n1075, WX11039, WX11103 );
xor U10580 ( n1076, WX11231, WX11167 );
xor U10581 ( n740, n1088, n1089 );
xnor U10582 ( n1088, WX11037, WX11101 );
xor U10583 ( n1089, WX11229, WX11165 );
xor U10584 ( n748, n1100, n1101 );
xnor U10585 ( n1100, WX11035, WX11099 );
xor U10586 ( n1101, WX11227, WX11163 );
xor U10587 ( n756, n1113, n1114 );
xnor U10588 ( n1113, WX11033, WX11097 );
xor U10589 ( n1114, WX11225, WX11161 );
xor U10590 ( n764, n1125, n1126 );
xnor U10591 ( n1125, WX11031, WX11095 );
xor U10592 ( n1126, WX11223, WX11159 );
xor U10593 ( n772, n1138, n1139 );
xnor U10594 ( n1138, WX11029, WX11093 );
xor U10595 ( n1139, WX11221, WX11157 );
xor U10596 ( n780, n1150, n1151 );
xnor U10597 ( n1150, WX11027, WX11091 );
xor U10598 ( n1151, WX11219, WX11155 );
xor U10599 ( n788, n1163, n1164 );
xnor U10600 ( n1163, WX11025, WX11089 );
xor U10601 ( n1164, WX11217, WX11153 );
xor U10602 ( n796, n1175, n1176 );
xnor U10603 ( n1175, WX11023, WX11087 );
xor U10604 ( n1176, WX11215, WX11151 );
xor U10605 ( n804, n1188, n1189 );
xnor U10606 ( n1188, WX11021, WX11085 );
xor U10607 ( n1189, WX11213, WX11149 );
endmodule

