
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

always @(posedge clk) begin
if (reset == 1'b1) begin
Q <= 1'b0;
end
else begin
Q <= D;
end
end

endmodule


module b18_ori ( clk, reset, HOLD, NA, BS, SEL, DIN_31_, DIN_30_, DIN_29_, DIN_28_,
DIN_27_, DIN_26_, DIN_25_, DIN_24_, DIN_23_, DIN_22_, DIN_21_, DIN_20_,
DIN_19_, DIN_18_, DIN_17_, DIN_16_, DIN_15_, DIN_14_, DIN_13_, DIN_12_,
DIN_11_, DIN_10_, DIN_9_, DIN_8_, DIN_7_, DIN_6_, DIN_5_, DIN_4_,
DIN_3_, DIN_2_, DIN_1_, DIN_0_, LOGIC0, MUL_1411_U378, MUL_1411_U438,
MUL_1411_U10, MUL_1411_U439, MUL_1411_U9, MUL_1411_U440, MUL_1411_U8,
MUL_1411_U441, MUL_1411_U7, MUL_1411_U385, MUL_1411_U14, MUL_1411_U386,
MUL_1411_U13, MUL_1411_U387, MUL_1411_U12, MUL_1411_U388, MUL_1411_U11,
MUL_1411_U15, MUL_1411_U5, MUL_1421_A1_U5, U154, U39 );
input clk, reset, HOLD, NA, BS, SEL, DIN_31_, DIN_30_, DIN_29_, DIN_28_, DIN_27_,
DIN_26_, DIN_25_, DIN_24_, DIN_23_, DIN_22_, DIN_21_, DIN_20_,
DIN_19_, DIN_18_, DIN_17_, DIN_16_, DIN_15_, DIN_14_, DIN_13_,
DIN_12_, DIN_11_, DIN_10_, DIN_9_, DIN_8_, DIN_7_, DIN_6_, DIN_5_,
DIN_4_, DIN_3_, DIN_2_, DIN_1_, DIN_0_, LOGIC0;
output MUL_1411_U378, MUL_1411_U438, MUL_1411_U10, MUL_1411_U439,
MUL_1411_U9, MUL_1411_U440, MUL_1411_U8, MUL_1411_U441, MUL_1411_U7,
MUL_1411_U385, MUL_1411_U14, MUL_1411_U386, MUL_1411_U13,
MUL_1411_U387, MUL_1411_U12, MUL_1411_U388, MUL_1411_U11,
MUL_1411_U15, MUL_1411_U5, MUL_1421_A1_U5, U154, U39;
wire P3_WR_REG, P4_WR_REG, P1_P3_M_IO_N_REG, P1_P3_D_C_N_REG, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, ex_wire30, ex_wire31, ex_wire32, ex_wire33, ex_wire34, ex_wire35, ex_wire36, ex_wire37, ex_wire38, ex_wire39, ex_wire40, ex_wire41, ex_wire42, ex_wire43, ex_wire44, ex_wire45, ex_wire46, ex_wire47, ex_wire48, ex_wire49, ex_wire50, ex_wire51, ex_wire52, ex_wire53, ex_wire54, ex_wire55, ex_wire56, ex_wire57, ex_wire58, ex_wire59, ex_wire60, ex_wire61, ex_wire62, ex_wire63, ex_wire64, ex_wire65, ex_wire66, ex_wire67, ex_wire68, ex_wire69, ex_wire70, ex_wire71, ex_wire72, ex_wire73, ex_wire74, ex_wire75, ex_wire76, ex_wire77, ex_wire78, ex_wire79, ex_wire80, ex_wire81, ex_wire82, ex_wire83, ex_wire84, ex_wire85, ex_wire86, ex_wire87, ex_wire88, ex_wire89, ex_wire90, ex_wire91, ex_wire92, ex_wire93, ex_wire94, ex_wire95, ex_wire96, ex_wire97, ex_wire98, ex_wire99, ex_wire100, ex_wire101, ex_wire102, ex_wire103, ex_wire104, ex_wire105, ex_wire106, ex_wire107, ex_wire108, ex_wire109, ex_wire110, ex_wire111, ex_wire112, ex_wire113, ex_wire114, ex_wire115, ex_wire116, ex_wire117, ex_wire118, ex_wire119, ex_wire120, ex_wire121, ex_wire122, ex_wire123, ex_wire124, ex_wire125, ex_wire126, ex_wire127, ex_wire128, ex_wire129, ex_wire130, ex_wire131, ex_wire132, ex_wire133, ex_wire134, ex_wire135, ex_wire136, ex_wire137, ex_wire138, ex_wire139, ex_wire140, ex_wire141, ex_wire142, ex_wire143, ex_wire144, ex_wire145, ex_wire146, ex_wire147, ex_wire148, ex_wire149, ex_wire150, ex_wire151, ex_wire152, ex_wire153, ex_wire154, ex_wire155, ex_wire156, ex_wire157, ex_wire158, ex_wire159, ex_wire160, ex_wire161, ex_wire162, ex_wire163, ex_wire164, ex_wire165, ex_wire166, ex_wire167, ex_wire168, ex_wire169, ex_wire170, ex_wire171, ex_wire172, ex_wire173, ex_wire174, ex_wire175, ex_wire176, ex_wire177, ex_wire178, ex_wire179, ex_wire180, ex_wire181, ex_wire182, ex_wire183, ex_wire184, ex_wire185, ex_wire186, ex_wire187, ex_wire188, ex_wire189, ex_wire190, ex_wire191, ex_wire192, ex_wire193, ex_wire194, ex_wire195, ex_wire196, ex_wire197, ex_wire198, ex_wire199, ex_wire200, ex_wire201, ex_wire202, ex_wire203, ex_wire204, ex_wire205, ex_wire206, ex_wire207, ex_wire208, ex_wire209, ex_wire210, ex_wire211, ex_wire212, ex_wire213, ex_wire214, ex_wire215, ex_wire216, ex_wire217, ex_wire218, ex_wire219, ex_wire220, ex_wire221, ex_wire222, ex_wire223, ex_wire224, ex_wire225, ex_wire226, ex_wire227, ex_wire228, ex_wire229, ex_wire230, ex_wire231, ex_wire232, ex_wire233, ex_wire234, ex_wire235, ex_wire236, ex_wire237, ex_wire238, ex_wire239, ex_wire240, ex_wire241, ex_wire242, ex_wire243, ex_wire244, ex_wire245, ex_wire246, ex_wire247, ex_wire248, ex_wire249, ex_wire250, ex_wire251, ex_wire252, ex_wire253, ex_wire254, ex_wire255, ex_wire256, ex_wire257, ex_wire258, ex_wire259, ex_wire260, ex_wire261, ex_wire262, ex_wire263, ex_wire264, ex_wire265, ex_wire266, ex_wire267, ex_wire268, ex_wire269, ex_wire270, ex_wire271, ex_wire272, ex_wire273, ex_wire274, ex_wire275, ex_wire276, ex_wire277, ex_wire278, ex_wire279, ex_wire280, ex_wire281, ex_wire282, ex_wire283, ex_wire284, ex_wire285, ex_wire286, ex_wire287, ex_wire288, ex_wire289, ex_wire290, ex_wire291, ex_wire292, ex_wire293, ex_wire294, ex_wire295, ex_wire296, ex_wire297, ex_wire298, ex_wire299, ex_wire300, ex_wire301, ex_wire302, ex_wire303, ex_wire304, ex_wire305, ex_wire306, ex_wire307, ex_wire308, ex_wire309, ex_wire310, ex_wire311, ex_wire312, ex_wire313, ex_wire314, ex_wire315, ex_wire316, ex_wire317, ex_wire318, ex_wire319, ex_wire320, ex_wire321, ex_wire322, ex_wire323, ex_wire324, ex_wire325, ex_wire326, P3_RD_REG,
P1_P3_W_R_N_REG, P4_RD_REG, P2_P3_W_R_N_REG, P2_P3_M_IO_N_REG,
P2_P3_D_C_N_REG, P1_P1_ADDRESS_REG_2_, P2_P1_ADDRESS_REG_2_,
P1_P3_ADS_N_REG, P2_P3_ADS_N_REG, P1_P1_ADDRESS_REG_9_,
P1_P1_ADDRESS_REG_8_, P1_P1_ADDRESS_REG_7_, P1_P1_ADDRESS_REG_6_,
P1_P1_ADDRESS_REG_5_, P1_P1_ADDRESS_REG_4_, P4_ADDR_REG_4_,
P1_P1_ADDRESS_REG_3_, P4_ADDR_REG_2_, P1_P1_ADDRESS_REG_18_,
P1_P1_ADDRESS_REG_17_, P1_P1_ADDRESS_REG_16_, P1_P1_ADDRESS_REG_15_,
P1_P1_ADDRESS_REG_14_, P1_P1_ADDRESS_REG_13_, P1_P1_ADDRESS_REG_12_,
P1_P1_ADDRESS_REG_11_, P1_P1_ADDRESS_REG_10_, P2_P1_ADDRESS_REG_9_,
P2_P1_ADDRESS_REG_8_, P2_P1_ADDRESS_REG_7_, P2_P1_ADDRESS_REG_6_,
P2_P1_ADDRESS_REG_5_, P2_P1_ADDRESS_REG_4_, P3_ADDR_REG_4_,
P2_P1_ADDRESS_REG_3_, P3_ADDR_REG_2_, P2_P1_ADDRESS_REG_18_,
P2_P1_ADDRESS_REG_17_, P2_P1_ADDRESS_REG_16_, P2_P1_ADDRESS_REG_15_,
P2_P1_ADDRESS_REG_14_, P2_P1_ADDRESS_REG_13_, P2_P1_ADDRESS_REG_12_,
P2_P1_ADDRESS_REG_11_, P2_P1_ADDRESS_REG_10_, P1_P1_ADDRESS_REG_1_,
P4_ADDR_REG_1_, P1_P1_ADDRESS_REG_0_, P4_ADDR_REG_0_,
P2_P1_ADDRESS_REG_1_, P3_ADDR_REG_1_, P2_P1_ADDRESS_REG_0_,
P3_ADDR_REG_0_, n456, P1_P2_W_R_N_REG, P1_P2_M_IO_N_REG,
P1_READY22_REG, P1_READY11_REG, P2_P1_ADS_N_REG, P1_READY12_REG,
P1_READY21_REG, n441, n451, P1_P1_W_R_N_REG, P1_P1_M_IO_N_REG, n276,
n271, n266, n261, n256, n251, n246, n241, n236, n231, n226, n221,
n216, n211, n206, n201, n196, n191, n186, n181, n176, n171, n166,
n161, n156, n151, n146, n141, n136, n131, n126, n121, n281, n286,
n291, n296, n301, n306, n311, n316, n321, n326, n331, n336, n341,
n346, n351, n356, n361, n366, n371, n376, n381, n386, n391, n396,
n401, n406, n411, n416, n421, n426, n431, n436, P1_P1_BE_N_REG_0_,
P1_P1_ADS_N_REG, P1_P1_D_C_N_REG, P1_P1_BE_N_REG_1_,
P1_P1_BE_N_REG_3_, P1_P2_BE_N_REG_1_, P1_P2_BE_N_REG_2_,
P1_P2_BE_N_REG_0_, P1_P2_ADS_N_REG, P1_P2_D_C_N_REG,
P1_P2_BE_N_REG_3_, P1_P3_BE_N_REG_1_, P1_P3_BE_N_REG_0_,
P1_P3_BE_N_REG_3_, P1_P3_BE_N_REG_2_, P1_P1_BE_N_REG_2_,
P1_P2_DATAO_REG_0_, P1_P1_DATAO_REG_0_, P1_BUF1_REG_0_,
P1_P2_DATAO_REG_1_, P1_P1_DATAO_REG_1_, P1_BUF1_REG_1_,
P1_P2_DATAO_REG_2_, P1_P1_DATAO_REG_2_, P1_BUF1_REG_2_,
P1_P2_DATAO_REG_3_, P1_P1_DATAO_REG_3_, P1_BUF1_REG_3_,
P1_P2_DATAO_REG_4_, P1_P1_DATAO_REG_4_, P1_BUF1_REG_4_,
P1_P2_DATAO_REG_5_, P1_P1_DATAO_REG_5_, P1_BUF1_REG_5_,
P1_P2_DATAO_REG_6_, P1_P1_DATAO_REG_6_, P1_BUF1_REG_6_,
P1_P2_DATAO_REG_7_, P1_P1_DATAO_REG_7_, P1_BUF1_REG_7_,
P1_P2_DATAO_REG_8_, P1_P1_DATAO_REG_8_, P1_BUF1_REG_8_,
P1_P2_DATAO_REG_9_, P1_P1_DATAO_REG_9_, P1_BUF1_REG_9_,
P1_P2_DATAO_REG_10_, P1_P1_DATAO_REG_10_, P1_BUF1_REG_10_,
P1_P2_DATAO_REG_11_, P1_P1_DATAO_REG_11_, P1_BUF1_REG_11_,
P1_P2_DATAO_REG_12_, P1_P1_DATAO_REG_12_, P1_BUF1_REG_12_,
P1_P2_DATAO_REG_13_, P1_P1_DATAO_REG_13_, P1_BUF1_REG_13_,
P1_P2_DATAO_REG_14_, P1_P1_DATAO_REG_14_, P1_BUF1_REG_14_,
P1_P2_DATAO_REG_15_, P1_P1_DATAO_REG_15_, P1_BUF1_REG_15_,
P1_P2_DATAO_REG_16_, P1_P1_DATAO_REG_16_, P1_BUF1_REG_16_,
P1_P2_DATAO_REG_17_, P1_P1_DATAO_REG_17_, P1_BUF1_REG_17_,
P1_P2_DATAO_REG_18_, P1_P1_DATAO_REG_18_, P1_BUF1_REG_18_,
P1_P2_DATAO_REG_19_, P1_P1_DATAO_REG_19_, P1_BUF1_REG_19_,
P1_P2_DATAO_REG_20_, P1_P1_DATAO_REG_20_, P1_BUF1_REG_20_,
P1_P2_DATAO_REG_21_, P1_P1_DATAO_REG_21_, P1_BUF1_REG_21_,
P1_P2_DATAO_REG_22_, P1_P1_DATAO_REG_22_, P1_BUF1_REG_22_,
P1_P2_DATAO_REG_23_, P1_P1_DATAO_REG_23_, P1_BUF1_REG_23_,
P1_P2_DATAO_REG_24_, P1_P1_DATAO_REG_24_, P1_BUF1_REG_24_,
P1_P2_DATAO_REG_25_, P1_P1_DATAO_REG_25_, P1_BUF1_REG_25_,
P1_P2_DATAO_REG_26_, P1_P1_DATAO_REG_26_, P1_BUF1_REG_26_,
P1_P2_DATAO_REG_27_, P1_P1_DATAO_REG_27_, P1_BUF1_REG_27_,
P1_P2_DATAO_REG_28_, P1_P1_DATAO_REG_28_, P1_BUF1_REG_28_,
P1_P2_DATAO_REG_29_, P1_P1_DATAO_REG_29_, P1_BUF1_REG_29_,
P1_P2_DATAO_REG_30_, P1_P1_DATAO_REG_30_, P1_BUF1_REG_30_,
P1_P2_DATAO_REG_31_, P1_P1_DATAO_REG_31_, P1_BUF1_REG_31_,
P1_BUF2_REG_0_, P1_BUF2_REG_1_, P1_BUF2_REG_2_, P1_BUF2_REG_3_,
P1_BUF2_REG_4_, P1_BUF2_REG_5_, P1_BUF2_REG_6_, P1_BUF2_REG_7_,
P1_BUF2_REG_8_, P1_BUF2_REG_9_, P1_BUF2_REG_10_, P1_BUF2_REG_11_,
P1_BUF2_REG_12_, P1_BUF2_REG_13_, P1_BUF2_REG_14_, P1_BUF2_REG_15_,
P1_BUF2_REG_16_, P1_BUF2_REG_17_, P1_BUF2_REG_18_, P1_BUF2_REG_19_,
P1_BUF2_REG_20_, P1_BUF2_REG_21_, P1_BUF2_REG_22_, P1_BUF2_REG_23_,
P1_BUF2_REG_24_, P1_BUF2_REG_25_, P1_BUF2_REG_26_, P1_BUF2_REG_27_,
P1_BUF2_REG_28_, P1_BUF2_REG_29_, P1_BUF2_REG_30_, P1_BUF2_REG_31_,
P1_P2_ADDRESS_REG_9_, P1_P3_ADDRESS_REG_9_, P1_P2_ADDRESS_REG_8_,
P1_P3_ADDRESS_REG_8_, P1_P2_ADDRESS_REG_7_, P1_P3_ADDRESS_REG_7_,
P1_P2_ADDRESS_REG_6_, P1_P3_ADDRESS_REG_6_, P1_P2_ADDRESS_REG_5_,
P1_P3_ADDRESS_REG_5_, P1_P2_ADDRESS_REG_4_, P1_P3_ADDRESS_REG_4_,
P1_P2_ADDRESS_REG_3_, P1_P3_ADDRESS_REG_3_, P1_P2_ADDRESS_REG_2_,
P1_P3_ADDRESS_REG_2_, P1_P2_ADDRESS_REG_1_, P1_P3_ADDRESS_REG_1_,
P1_P2_ADDRESS_REG_18_, P1_P3_ADDRESS_REG_18_, P1_P2_ADDRESS_REG_17_,
P1_P3_ADDRESS_REG_17_, P1_P2_ADDRESS_REG_16_, P1_P3_ADDRESS_REG_16_,
P1_P2_ADDRESS_REG_15_, P1_P3_ADDRESS_REG_15_, P1_P2_ADDRESS_REG_14_,
P1_P3_ADDRESS_REG_14_, P1_P2_ADDRESS_REG_13_, P1_P3_ADDRESS_REG_13_,
P1_P2_ADDRESS_REG_12_, P1_P3_ADDRESS_REG_12_, P1_P2_ADDRESS_REG_11_,
P1_P3_ADDRESS_REG_11_, P1_P2_ADDRESS_REG_10_, P1_P3_ADDRESS_REG_10_,
P1_P2_ADDRESS_REG_0_, P1_P3_ADDRESS_REG_0_, n796, P2_P2_W_R_N_REG,
P2_P2_M_IO_N_REG, P2_READY22_REG, P2_READY11_REG, P2_READY12_REG,
P2_READY21_REG, n781, n791, P2_P1_W_R_N_REG, P2_P1_M_IO_N_REG, n616,
n611, n606, n601, n596, n591, n586, n581, n576, n571, n566, n561,
n556, n551, n546, n541, n536, n531, n526, n521, n516, n511, n506,
n501, n496, n491, n486, n481, n476, n471, n466, n461, n621, n626,
n631, n636, n641, n646, n651, n656, n661, n666, n671, n676, n681,
n686, n691, n696, n701, n706, n711, n716, n721, n726, n731, n736,
n741, n746, n751, n756, n761, n766, n771, n776, P2_P1_BE_N_REG_0_,
P2_P1_D_C_N_REG, P2_P1_BE_N_REG_1_, P2_P1_BE_N_REG_3_,
P2_P2_BE_N_REG_1_, P2_P2_BE_N_REG_2_, P2_P2_BE_N_REG_0_,
P2_P2_ADS_N_REG, P2_P2_D_C_N_REG, P2_P2_BE_N_REG_3_,
P2_P3_BE_N_REG_1_, P2_P3_BE_N_REG_0_, P2_P3_BE_N_REG_3_,
P2_P3_BE_N_REG_2_, P2_P1_BE_N_REG_2_, P2_P2_DATAO_REG_0_,
P2_P1_DATAO_REG_0_, P2_BUF1_REG_0_, P2_P2_DATAO_REG_1_,
P2_P1_DATAO_REG_1_, P2_BUF1_REG_1_, P2_P2_DATAO_REG_2_,
P2_P1_DATAO_REG_2_, P2_BUF1_REG_2_, P2_P2_DATAO_REG_3_,
P2_P1_DATAO_REG_3_, P2_BUF1_REG_3_, P2_P2_DATAO_REG_4_,
P2_P1_DATAO_REG_4_, P2_BUF1_REG_4_, P2_P2_DATAO_REG_5_,
P2_P1_DATAO_REG_5_, P2_BUF1_REG_5_, P2_P2_DATAO_REG_6_,
P2_P1_DATAO_REG_6_, P2_BUF1_REG_6_, P2_P2_DATAO_REG_7_,
P2_P1_DATAO_REG_7_, P2_BUF1_REG_7_, P2_P2_DATAO_REG_8_,
P2_P1_DATAO_REG_8_, P2_BUF1_REG_8_, P2_P2_DATAO_REG_9_,
P2_P1_DATAO_REG_9_, P2_BUF1_REG_9_, P2_P2_DATAO_REG_10_,
P2_P1_DATAO_REG_10_, P2_BUF1_REG_10_, P2_P2_DATAO_REG_11_,
P2_P1_DATAO_REG_11_, P2_BUF1_REG_11_, P2_P2_DATAO_REG_12_,
P2_P1_DATAO_REG_12_, P2_BUF1_REG_12_, P2_P2_DATAO_REG_13_,
P2_P1_DATAO_REG_13_, P2_BUF1_REG_13_, P2_P2_DATAO_REG_14_,
P2_P1_DATAO_REG_14_, P2_BUF1_REG_14_, P2_P2_DATAO_REG_15_,
P2_P1_DATAO_REG_15_, P2_BUF1_REG_15_, P2_P2_DATAO_REG_16_,
P2_P1_DATAO_REG_16_, P2_BUF1_REG_16_, P2_P2_DATAO_REG_17_,
P2_P1_DATAO_REG_17_, P2_BUF1_REG_17_, P2_P2_DATAO_REG_18_,
P2_P1_DATAO_REG_18_, P2_BUF1_REG_18_, P2_P2_DATAO_REG_19_,
P2_P1_DATAO_REG_19_, P2_BUF1_REG_19_, P2_P2_DATAO_REG_20_,
P2_P1_DATAO_REG_20_, P2_BUF1_REG_20_, P2_P2_DATAO_REG_21_,
P2_P1_DATAO_REG_21_, P2_BUF1_REG_21_, P2_P2_DATAO_REG_22_,
P2_P1_DATAO_REG_22_, P2_BUF1_REG_22_, P2_P2_DATAO_REG_23_,
P2_P1_DATAO_REG_23_, P2_BUF1_REG_23_, P2_P2_DATAO_REG_24_,
P2_P1_DATAO_REG_24_, P2_BUF1_REG_24_, P2_P2_DATAO_REG_25_,
P2_P1_DATAO_REG_25_, P2_BUF1_REG_25_, P2_P2_DATAO_REG_26_,
P2_P1_DATAO_REG_26_, P2_BUF1_REG_26_, P2_P2_DATAO_REG_27_,
P2_P1_DATAO_REG_27_, P2_BUF1_REG_27_, P2_P2_DATAO_REG_28_,
P2_P1_DATAO_REG_28_, P2_BUF1_REG_28_, P2_P2_DATAO_REG_29_,
P2_P1_DATAO_REG_29_, P2_BUF1_REG_29_, P2_P2_DATAO_REG_30_,
P2_P1_DATAO_REG_30_, P2_BUF1_REG_30_, P2_P2_DATAO_REG_31_,
P2_P1_DATAO_REG_31_, P2_BUF1_REG_31_, P2_BUF2_REG_0_, P2_BUF2_REG_1_,
P2_BUF2_REG_2_, P2_BUF2_REG_3_, P2_BUF2_REG_4_, P2_BUF2_REG_5_,
P2_BUF2_REG_6_, P2_BUF2_REG_7_, P2_BUF2_REG_8_, P2_BUF2_REG_9_,
P2_BUF2_REG_10_, P2_BUF2_REG_11_, P2_BUF2_REG_12_, P2_BUF2_REG_13_,
P2_BUF2_REG_14_, P2_BUF2_REG_15_, P2_BUF2_REG_16_, P2_BUF2_REG_17_,
P2_BUF2_REG_18_, P2_BUF2_REG_19_, P2_BUF2_REG_20_, P2_BUF2_REG_21_,
P2_BUF2_REG_22_, P2_BUF2_REG_23_, P2_BUF2_REG_24_, P2_BUF2_REG_25_,
P2_BUF2_REG_26_, P2_BUF2_REG_27_, P2_BUF2_REG_28_, P2_BUF2_REG_29_,
P2_BUF2_REG_30_, P2_BUF2_REG_31_, P2_P2_ADDRESS_REG_9_,
P2_P3_ADDRESS_REG_9_, P2_P2_ADDRESS_REG_8_, P2_P3_ADDRESS_REG_8_,
P2_P2_ADDRESS_REG_7_, P2_P3_ADDRESS_REG_7_, P2_P2_ADDRESS_REG_6_,
P2_P3_ADDRESS_REG_6_, P2_P2_ADDRESS_REG_5_, P2_P3_ADDRESS_REG_5_,
P2_P2_ADDRESS_REG_4_, P2_P3_ADDRESS_REG_4_, P2_P2_ADDRESS_REG_3_,
P2_P3_ADDRESS_REG_3_, P2_P2_ADDRESS_REG_2_, P2_P3_ADDRESS_REG_2_,
P2_P2_ADDRESS_REG_1_, P2_P3_ADDRESS_REG_1_, P2_P2_ADDRESS_REG_18_,
P2_P3_ADDRESS_REG_18_, P2_P2_ADDRESS_REG_17_, P2_P3_ADDRESS_REG_17_,
P2_P2_ADDRESS_REG_16_, P2_P3_ADDRESS_REG_16_, P2_P2_ADDRESS_REG_15_,
P2_P3_ADDRESS_REG_15_, P2_P2_ADDRESS_REG_14_, P2_P3_ADDRESS_REG_14_,
P2_P2_ADDRESS_REG_13_, P2_P3_ADDRESS_REG_13_, P2_P2_ADDRESS_REG_12_,
P2_P3_ADDRESS_REG_12_, P2_P2_ADDRESS_REG_11_, P2_P3_ADDRESS_REG_11_,
P2_P2_ADDRESS_REG_10_, P2_P3_ADDRESS_REG_10_, P2_P2_ADDRESS_REG_0_,
P2_P3_ADDRESS_REG_0_, P3_STATE_REG, n2016, n2006, n2001, n1996, n1991,
n1986, n1981, n1976, n1971, n1966, n1961, n1956, n1951, n1946, n1941,
n1936, n1931, n1926, n1921, n1916, n1911, n1906, n1901, n1896, n1891,
n1886, n1881, n1876, n1871, n1866, n1861, n1696, n1691, n1686, n1681,
n1676, n1671, n1666, n1661, n1656, n1651, n1646, n1641, n1636, n1631,
n1626, n1621, n1616, n1611, n1606, n1596, n1591, n1586, n1581, n1576,
n1571, n1566, n1561, n1556, n1551, n1546, n1541, n1536, n1531, n1526,
n1521, n1516, n1511, n1506, n1501, n1496, n1491, n1486, n1481, n1476,
n1471, n1466, n1461, n1456, n1451, n1446, n1441, P3_D_REG_31_, n1116,
P3_D_REG_30_, n1111, P3_D_REG_29_, n1106, P3_D_REG_28_, n1101,
P3_D_REG_27_, n1096, P3_D_REG_26_, n1091, P3_D_REG_25_, n1086,
P3_D_REG_24_, n1081, P3_D_REG_23_, n1076, n1071, P3_D_REG_21_, n1066,
P3_D_REG_20_, n1061, P3_D_REG_19_, n1056, P3_D_REG_18_, n1051,
P3_D_REG_17_, n1046, P3_D_REG_16_, n1041, P3_D_REG_15_, n1036,
P3_D_REG_14_, n1031, P3_D_REG_13_, n1026, P3_D_REG_12_, n1021,
P3_D_REG_11_, n1016, P3_D_REG_10_, n1011, P3_D_REG_9_, n1006,
P3_D_REG_8_, n1001, n996, P3_D_REG_6_, n991, P3_D_REG_5_, n986,
P3_D_REG_4_, n981, P3_D_REG_3_, n976, P3_D_REG_2_, n971, n956, n951,
n946, n941, n936, n931, n926, n921, n916, n911, n906, n901, n896,
n891, n886, n881, n876, n871, n866, n861, n856, n851, n846, n841,
n836, n831, n826, n821, n816, n811, n806, n801, P3_B_REG,
P3_REG2_REG_0_, n961, n966, n1121, n1126, n1131, n1136, n1141, n1146,
n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196,
n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246,
n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296,
n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346,
n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396,
n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1701, n1706,
n1711, n1716, n1721, n1726, n1731, n1736, n1741, n1746, n1751, n1756,
n1761, n1766, n1771, n1776, n1781, n1786, n1791, n1796, n1801, n1806,
n1811, n1816, n1821, n1826, n1831, n1836, n1841, n1846, n1851, n1856,
P3_IR_REG_31_, P1_P3_DATAO_REG_0_, P3_IR_REG_0_, P1_P3_DATAO_REG_1_,
P3_IR_REG_1_, P1_P3_DATAO_REG_2_, P3_IR_REG_2_, P1_P3_DATAO_REG_3_,
P3_IR_REG_3_, P1_P3_DATAO_REG_4_, P3_IR_REG_4_, P1_P3_DATAO_REG_5_,
P3_IR_REG_5_, P1_P3_DATAO_REG_6_, P3_IR_REG_6_, P1_P3_DATAO_REG_7_,
P3_IR_REG_7_, P1_P3_DATAO_REG_8_, P3_IR_REG_8_, P1_P3_DATAO_REG_9_,
P3_IR_REG_9_, P1_P3_DATAO_REG_10_, P3_IR_REG_10_, P1_P3_DATAO_REG_11_,
P3_IR_REG_11_, P1_P3_DATAO_REG_12_, P3_IR_REG_12_,
P1_P3_DATAO_REG_13_, P3_IR_REG_13_, P1_P3_DATAO_REG_14_,
P3_IR_REG_14_, P1_P3_DATAO_REG_15_, P3_IR_REG_15_,
P1_P3_DATAO_REG_16_, P3_IR_REG_16_, P1_P3_DATAO_REG_17_,
P3_IR_REG_17_, P1_P3_DATAO_REG_18_, P3_IR_REG_18_,
P1_P3_DATAO_REG_19_, P3_IR_REG_19_, P3_IR_REG_20_, P3_IR_REG_21_,
P3_IR_REG_22_, P3_IR_REG_23_, P3_IR_REG_24_, P3_IR_REG_25_,
P3_IR_REG_26_, P3_IR_REG_27_, P3_IR_REG_28_, P3_IR_REG_29_,
P3_IR_REG_30_, P3_REG2_REG_1_, P3_REG1_REG_1_, P3_REG0_REG_1_,
P3_REG3_REG_1_, P3_REG2_REG_2_, P3_REG1_REG_2_, P3_REG0_REG_2_,
P3_REG3_REG_2_, P3_REG0_REG_0_, P3_REG1_REG_0_, P3_REG3_REG_0_,
P3_REG2_REG_3_, P3_REG1_REG_3_, P3_REG0_REG_3_, P3_REG2_REG_4_,
P3_REG1_REG_4_, P3_REG0_REG_4_, P3_REG2_REG_5_, P3_REG1_REG_5_,
P3_REG0_REG_5_, P3_REG2_REG_6_, P3_REG1_REG_6_, P3_REG0_REG_6_,
P3_REG2_REG_7_, P3_REG1_REG_7_, P3_REG0_REG_7_, P3_REG2_REG_8_,
P3_REG1_REG_8_, P3_REG0_REG_8_, P3_REG2_REG_9_, P3_REG1_REG_9_,
P3_REG0_REG_9_, P3_REG1_REG_10_, P3_REG0_REG_10_, P3_REG2_REG_11_,
P3_REG1_REG_11_, P3_REG0_REG_11_, P3_REG2_REG_12_, P3_REG1_REG_12_,
P3_REG0_REG_12_, P3_REG2_REG_13_, P3_REG1_REG_13_, P3_REG0_REG_13_,
P3_REG2_REG_14_, P3_REG1_REG_14_, P3_REG0_REG_14_, P3_REG2_REG_15_,
P3_REG1_REG_15_, P3_REG0_REG_15_, P3_REG2_REG_16_, P3_REG1_REG_16_,
P3_REG0_REG_16_, P3_REG2_REG_17_, P3_REG1_REG_17_, P3_REG0_REG_17_,
P3_REG1_REG_18_, P3_REG0_REG_18_, P3_REG1_REG_19_, P3_REG0_REG_19_,
P3_REG1_REG_20_, P3_REG0_REG_20_, P3_REG2_REG_21_, P3_REG1_REG_21_,
P3_REG0_REG_21_, P3_REG1_REG_22_, P3_REG0_REG_22_, P3_REG2_REG_23_,
P3_REG1_REG_23_, P3_REG0_REG_23_, P3_REG2_REG_24_, P3_REG1_REG_24_,
P3_REG0_REG_24_, P3_REG1_REG_25_, P3_REG0_REG_25_, P3_REG2_REG_26_,
P3_REG1_REG_26_, P3_REG0_REG_26_, P3_REG2_REG_27_, P3_REG1_REG_27_,
P3_REG0_REG_27_, P3_REG1_REG_28_, P3_REG0_REG_28_, P3_REG1_REG_29_,
P3_REG0_REG_29_, P3_REG2_REG_30_, P3_REG1_REG_30_, P3_REG0_REG_30_,
P3_REG2_REG_31_, P3_REG1_REG_31_, P3_REG0_REG_31_, P3_REG3_REG_19_,
P3_REG3_REG_18_, P3_REG3_REG_17_, P3_REG3_REG_16_, P3_REG3_REG_15_,
P3_REG3_REG_14_, P3_REG3_REG_13_, P3_REG3_REG_12_, P3_REG3_REG_11_,
P3_REG3_REG_10_, P3_REG3_REG_9_, P3_REG3_REG_8_, P3_REG3_REG_7_,
P3_REG3_REG_6_, P3_REG3_REG_5_, P3_REG3_REG_4_, P3_REG3_REG_3_,
P3_REG3_REG_26_, P3_REG3_REG_22_, P3_REG3_REG_20_, P3_REG3_REG_24_,
P3_REG3_REG_25_, P3_REG3_REG_21_, P3_REG3_REG_28_, P3_REG3_REG_23_,
P3_REG3_REG_27_, P3_D_REG_0_, P3_D_REG_1_, P3_DATAO_REG_0_,
P3_DATAO_REG_1_, P3_DATAO_REG_2_, P3_DATAO_REG_3_, P3_DATAO_REG_4_,
P3_DATAO_REG_5_, P3_DATAO_REG_6_, P3_DATAO_REG_7_, P3_DATAO_REG_8_,
P3_DATAO_REG_9_, P3_DATAO_REG_10_, P3_DATAO_REG_11_, P3_DATAO_REG_12_,
P3_DATAO_REG_13_, P3_DATAO_REG_14_, P3_DATAO_REG_15_,
P3_DATAO_REG_16_, P3_DATAO_REG_17_, P3_DATAO_REG_18_,
P3_DATAO_REG_19_, P3_DATAO_REG_20_, P3_DATAO_REG_21_,
P3_DATAO_REG_22_, P3_DATAO_REG_23_, P3_DATAO_REG_24_,
P3_DATAO_REG_25_, P3_DATAO_REG_26_, P3_DATAO_REG_27_,
P3_DATAO_REG_28_, P3_DATAO_REG_29_, P3_DATAO_REG_30_,
P3_DATAO_REG_31_, P2_P1_INSTADDRPOINTER_REG_16_,
P2_P1_INSTADDRPOINTER_REG_25_, P2_P1_INSTADDRPOINTER_REG_7_,
P2_P1_INSTADDRPOINTER_REG_12_, P4_STATE_REG, n3241, n3231, n3226,
n3221, n3216, n3211, n3206, n3201, n3196, n3191, n3186, n3181, n3176,
n3171, n3166, n3161, n3156, n3151, n3146, n3141, n3136, n3131, n3126,
n3121, n3116, n3111, n3106, n3101, n3096, n3091, n3086, n2921, n2916,
n2911, n2906, n2901, n2896, n2891, n2886, n2881, n2876, n2871, n2866,
n2861, n2856, n2851, n2846, n2841, n2836, n2831, n2821, n2816, n2811,
n2806, n2801, n2796, n2791, n2786, n2781, n2776, n2771, n2766, n2761,
n2756, n2751, n2746, n2741, n2736, n2731, n2726, n2721, n2716, n2711,
n2706, n2701, n2696, n2691, n2686, n2681, n2676, n2671, n2666,
P4_D_REG_31_, n2341, P4_D_REG_30_, n2336, P4_D_REG_29_, n2331,
P4_D_REG_28_, n2326, P4_D_REG_27_, n2321, P4_D_REG_26_, n2316,
P4_D_REG_25_, n2311, P4_D_REG_24_, n2306, P4_D_REG_23_, n2301, n2296,
P4_D_REG_21_, n2291, P4_D_REG_20_, n2286, P4_D_REG_19_, n2281,
P4_D_REG_18_, n2276, P4_D_REG_17_, n2271, P4_D_REG_16_, n2266,
P4_D_REG_15_, n2261, P4_D_REG_14_, n2256, P4_D_REG_13_, n2251,
P4_D_REG_12_, n2246, P4_D_REG_11_, n2241, P4_D_REG_10_, n2236,
P4_D_REG_9_, n2231, P4_D_REG_8_, n2226, n2221, P4_D_REG_6_, n2216,
P4_D_REG_5_, n2211, P4_D_REG_4_, n2206, P4_D_REG_3_, n2201,
P4_D_REG_2_, n2196, n2181, n2176, n2171, n2166, n2161, n2156, n2151,
n2146, n2141, n2136, n2131, n2126, n2121, n2116, n2111, n2106, n2101,
n2096, n2091, n2086, n2081, n2076, n2071, n2066, n2061, n2056, n2051,
n2046, n2041, n2036, n2031, n2026, P4_B_REG, P4_REG2_REG_0_,
P2_P3_DATAO_REG_20_, P2_P3_DATAO_REG_21_, P2_P3_DATAO_REG_22_,
P2_P3_DATAO_REG_23_, P2_P3_DATAO_REG_24_, P2_P3_DATAO_REG_25_,
P2_P3_DATAO_REG_26_, P2_P3_DATAO_REG_27_, P2_P3_DATAO_REG_28_,
P2_P3_DATAO_REG_29_, P2_P3_DATAO_REG_30_, P2_P3_DATAO_REG_31_, n2186,
n2191, n2346, n2351, n2356, n2361, n2366, n2371, n2376, n2381, n2386,
n2391, n2396, n2401, n2406, n2411, n2416, n2421, n2426, n2431, n2436,
n2441, n2446, n2451, n2456, n2461, n2466, n2471, n2476, n2481, n2486,
n2491, n2496, n2501, n2506, n2511, n2516, n2521, n2526, n2531, n2536,
n2541, n2546, n2551, n2556, n2561, n2566, n2571, n2576, n2581, n2586,
n2591, n2596, n2601, n2606, n2611, n2616, n2621, n2626, n2631, n2636,
n2641, n2646, n2651, n2656, n2661, n2926, n2931, n2936, n2941, n2946,
n2951, n2956, n2961, n2966, n2971, n2976, n2981, n2986, n2991, n2996,
n3001, n3006, n3011, n3016, n3021, n3026, n3031, n3036, n3041, n3046,
n3051, n3056, n3061, n3066, n3071, n3076, n3081, P4_IR_REG_31_,
P2_P3_DATAO_REG_0_, P4_IR_REG_0_, P2_P3_DATAO_REG_1_, P4_IR_REG_1_,
P2_P3_DATAO_REG_2_, P4_IR_REG_2_, P2_P3_DATAO_REG_3_, P4_IR_REG_3_,
P2_P3_DATAO_REG_4_, P4_IR_REG_4_, P2_P3_DATAO_REG_5_, P4_IR_REG_5_,
P2_P3_DATAO_REG_6_, P4_IR_REG_6_, P2_P3_DATAO_REG_7_, P4_IR_REG_7_,
P2_P3_DATAO_REG_8_, P4_IR_REG_8_, P2_P3_DATAO_REG_9_, P4_IR_REG_9_,
P2_P3_DATAO_REG_10_, P4_IR_REG_10_, P2_P3_DATAO_REG_11_,
P4_IR_REG_11_, P2_P3_DATAO_REG_12_, P4_IR_REG_12_,
P2_P3_DATAO_REG_13_, P4_IR_REG_13_, P2_P3_DATAO_REG_14_,
P4_IR_REG_14_, P2_P3_DATAO_REG_15_, P4_IR_REG_15_,
P2_P3_DATAO_REG_16_, P4_IR_REG_16_, P2_P3_DATAO_REG_17_,
P4_IR_REG_17_, P2_P3_DATAO_REG_18_, P4_IR_REG_18_,
P2_P3_DATAO_REG_19_, P4_IR_REG_19_, P4_IR_REG_20_, P4_IR_REG_21_,
P4_IR_REG_22_, P4_IR_REG_23_, P4_IR_REG_24_, P4_IR_REG_25_,
P4_IR_REG_26_, P4_IR_REG_27_, P4_IR_REG_28_, P4_IR_REG_29_,
P4_IR_REG_30_, P4_REG2_REG_1_, P4_REG1_REG_1_, P4_REG0_REG_1_,
P4_REG3_REG_1_, P4_REG2_REG_2_, P4_REG1_REG_2_, P4_REG0_REG_2_,
P4_REG3_REG_2_, P4_REG0_REG_0_, P4_REG1_REG_0_, P4_REG3_REG_0_,
P4_REG2_REG_3_, P4_REG1_REG_3_, P4_REG0_REG_3_, P4_REG2_REG_4_,
P4_REG1_REG_4_, P4_REG0_REG_4_, P4_REG2_REG_5_, P4_REG1_REG_5_,
P4_REG0_REG_5_, P4_REG2_REG_6_, P4_REG1_REG_6_, P4_REG0_REG_6_,
P4_REG2_REG_7_, P4_REG1_REG_7_, P4_REG0_REG_7_, P4_REG2_REG_8_,
P4_REG1_REG_8_, P4_REG0_REG_8_, P4_REG2_REG_9_, P4_REG1_REG_9_,
P4_REG0_REG_9_, P4_REG2_REG_10_, P4_REG1_REG_10_, P4_REG0_REG_10_,
P4_REG2_REG_11_, P4_REG1_REG_11_, P4_REG0_REG_11_, P4_REG2_REG_12_,
P4_REG1_REG_12_, P4_REG0_REG_12_, P4_REG2_REG_13_, P4_REG1_REG_13_,
P4_REG0_REG_13_, P4_REG2_REG_14_, P4_REG1_REG_14_, P4_REG0_REG_14_,
P4_REG2_REG_15_, P4_REG1_REG_15_, P4_REG0_REG_15_, P4_REG2_REG_16_,
P4_REG1_REG_16_, P4_REG0_REG_16_, P4_REG2_REG_17_, P4_REG1_REG_17_,
P4_REG0_REG_17_, P4_REG1_REG_18_, P4_REG0_REG_18_, P4_REG1_REG_19_,
P4_REG0_REG_19_, P4_REG1_REG_20_, P4_REG0_REG_20_, P4_REG1_REG_21_,
P4_REG0_REG_21_, P4_REG1_REG_22_, P4_REG0_REG_22_, P4_REG1_REG_23_,
P4_REG0_REG_23_, P4_REG1_REG_24_, P4_REG0_REG_24_, P4_REG1_REG_25_,
P4_REG0_REG_25_, P4_REG1_REG_26_, P4_REG0_REG_26_, P4_REG1_REG_27_,
P4_REG0_REG_27_, P4_REG1_REG_28_, P4_REG0_REG_28_, P4_REG1_REG_29_,
P4_REG0_REG_29_, P4_REG1_REG_30_, P4_REG0_REG_30_, P4_REG1_REG_31_,
P4_REG0_REG_31_, P4_REG3_REG_19_, P4_REG3_REG_18_, P4_REG3_REG_17_,
P4_REG3_REG_16_, P4_REG3_REG_15_, P4_REG3_REG_14_, P4_REG3_REG_13_,
P4_REG3_REG_12_, P4_REG3_REG_11_, P4_REG3_REG_10_, P4_REG3_REG_9_,
P4_REG3_REG_8_, P4_REG3_REG_7_, P4_REG3_REG_6_, P4_REG3_REG_5_,
P4_REG3_REG_4_, P4_REG3_REG_3_, P4_REG3_REG_26_, P4_REG3_REG_22_,
P4_REG3_REG_20_, P4_REG3_REG_24_, P4_REG3_REG_25_, P4_REG3_REG_21_,
P4_REG3_REG_28_, P4_REG3_REG_23_, P4_REG3_REG_27_, P4_D_REG_0_,
P4_D_REG_1_, P4_DATAO_REG_0_, P4_DATAO_REG_1_, P4_DATAO_REG_2_,
P4_DATAO_REG_3_, P4_DATAO_REG_4_, P4_DATAO_REG_5_, P4_DATAO_REG_6_,
P4_DATAO_REG_7_, P4_DATAO_REG_8_, P4_DATAO_REG_9_, P4_DATAO_REG_10_,
P4_DATAO_REG_11_, P4_DATAO_REG_12_, P4_DATAO_REG_13_,
P4_DATAO_REG_14_, P4_DATAO_REG_15_, P4_DATAO_REG_16_,
P4_DATAO_REG_17_, P4_DATAO_REG_18_, P4_DATAO_REG_19_,
P4_DATAO_REG_20_, P4_DATAO_REG_21_, P4_DATAO_REG_22_,
P4_DATAO_REG_23_, P4_DATAO_REG_24_, P4_DATAO_REG_25_,
P4_DATAO_REG_26_, P4_DATAO_REG_27_, P4_DATAO_REG_28_,
P4_DATAO_REG_29_, P4_DATAO_REG_30_, P4_DATAO_REG_31_,
P2_P1_INSTADDRPOINTER_REG_21_, P2_P1_INSTADDRPOINTER_REG_28_,
P2_P1_INSTADDRPOINTER_REG_3_, P2_P1_INSTADDRPOINTER_REG_31_,
P2_P1_INSTADDRPOINTER_REG_10_, P2_P1_INSTADDRPOINTER_REG_19_,
P2_P1_INSTADDRPOINTER_REG_23_, P2_P1_INSTADDRPOINTER_REG_8_,
P2_P1_INSTADDRPOINTER_REG_5_, P2_P1_INSTADDRPOINTER_REG_14_,
P2_P1_INSTADDRPOINTER_REG_27_, P2_P1_INSTADDRPOINTER_REG_4_,
P2_P1_INSTADDRPOINTER_REG_15_, P2_P1_INSTADDRPOINTER_REG_26_,
P2_P1_INSTADDRPOINTER_REG_11_, P1_P3_STATEBS16_REG,
P1_P3_STATE2_REG_2_, P1_P3_STATE2_REG_3_, P1_P3_STATE2_REG_1_,
P1_P3_STATE2_REG_0_, P1_P3_INSTQUEUERD_ADDR_REG_3_,
P1_P3_INSTQUEUERD_ADDR_REG_2_, P1_P3_INSTQUEUERD_ADDR_REG_1_,
P1_P3_INSTQUEUERD_ADDR_REG_0_, P1_P3_INSTQUEUEWR_ADDR_REG_0_,
P1_P3_INSTQUEUEWR_ADDR_REG_2_, P1_P3_EBX_REG_31_,
P1_P3_INSTQUEUERD_ADDR_REG_4_, n5481, n5476, n5466, n5456, n5446,
n5431, n5421, n5416, n5411, n5406, n5401, n5396, n5391, n5386, n5381,
n5376, n5371, n5366, n5361, n5356, n5351, n5346, n5341, n5336, n5331,
n5326, n5321, n5316, n5311, n5306, n5301, n5296, n5291, n5286, n5281,
n5276, n5271, n5266, n5261, n5256, n5251, n5246, n5241, n5236, n5231,
n5226, n5221, n5216, n5211, n5206, n5201, n5196, n5191, n5186, n5181,
n5176, n5171, n5166, n5161, n5156, n5151, n5146, n5141, n5136, n5131,
n5126, n5121, n5116, n5111, n5106, n5101, n5091, n5086, n5081, n5076,
n5071, n5066, n5061, n5056, n5051, n5046, n5041, n5036, n5031, n5026,
n5021, n5016, n5011, n5006, n5001, n4996, n4991, n4986, n4981, n4976,
n4971, n4966, n4961, n4956, n4951, n4946, n4941, n4936, n4931, n4876,
n4871, n4866, n4861, n4856, n4851, n4846, n4841, n4836, n4831, n4826,
n4821, n4816, n4811, n4806, n4801, n4796, n4791, n4786, n4781, n4776,
n4771, n4766, n4761, n4706, n4701, n4696, n4691, n4686, n4681, n4676,
n4671, n4666, n4661, n4656, n4651, n4646, n4641, n4636, n4631, n4626,
n4621, n4616, n4611, n4606, n4601, n4596, n4591, n4586, n4581, n4576,
n4571, n4566, n4561, n4556, n4551, n4546, n4541, n4536, n4531, n4526,
n4521, n4516, n4511, n4506, n4501, n4496, n4491, n4486, n4481, n4476,
n4471, n4466, n4461, n4456, n4451, n4446, n4441, n4436, n4431, n4426,
n4421, n4416, n4411, n4406, n4401, n4396, n4391, n4386, n4381, n4376,
n4371, n4366, n4361, n4356, n4351, n4346, n4341, n4336, n4331, n4326,
n4321, n4316, n4311, n4306, n4301, n4296, n4291, n4286,
P1_P3_INSTQUEUEWR_ADDR_REG_4_, n4281, n4251, n4246, n4241, n4236,
n4231, n4226, n4221, n4216, n4211, n4206, n4201, n4196, n4191, n4186,
n4181, n4176, n4171, n4166, n4161, n4156, n4151, n4146, n4141, n4136,
n4131, n4126, n4121, n4116, n4111, n4106, n4101, n4096, n4091, n4086,
n4081, n4076, n4071, n4066, n4061, n4056, n4051, n4046, n4041, n4036,
n4031, n4026, n4021, n4016, n4011, n4006, n4001, n3996, n3991, n3986,
n3981, n3976, n3971, n3966, n3961, n3956, n3951, n3946, n3941, n3936,
n3931, n3926, n3921, n3916, n3911, n3906, n3901, n3896, n3891, n3886,
n3881, n3876, n3871, n3866, n3861, n3856, n3851, n3846, n3841, n3836,
n3831, n3826, n3821, n3816, n3811, n3806, n3801, n3796, n3791, n3786,
n3781, n3776, n3771, n3766, n3761, n3756, n3751, n3746, n3741, n3736,
n3731, n3726, n3721, n3716, n3711, n3706, n3701, n3696, n3691, n3686,
n3681, n3676, n3671, n3666, n3661, n3656, n3651, n3646, n3641, n3636,
n3631, n3626, n3621, n3616, n3611, n3606, n3601, n3591, n3586, n3581,
n3576, n3571, n3566, n3561, n3556, n3551, n3546, n3541, n3536, n3531,
n3526, n3521, n3516, n3511, n3506, n3501, n3496, n3491, n3486, n3481,
n3476, n3471, n3466, n3461, n3456, n3451, n3446, n3431, n3426, n3421,
n3416, n3411, n3406, n3401, n3396, n3391, n3386, n3381, n3376, n3371,
n3366, n3361, n3356, n3351, n3346, n3341, n3336, n3331, n3326,
P1_P3_REQUESTPENDING_REG, P1_P3_STATE_REG_1_, P1_P3_STATE_REG_2_,
P1_P3_REIP_REG_1_, P1_P3_STATE_REG_0_, P1_P3_INSTQUEUEWR_ADDR_REG_1_,
P1_P3_INSTQUEUEWR_ADDR_REG_3_, P1_P3_FLUSH_REG, P1_P3_REIP_REG_0_,
P1_P3_CODEFETCH_REG, P1_P3_READREQUEST_REG, n3251, n3256, n3261,
n3266, n3436, n3441, n3596, n4256, n4261, n4266, n4271, n4276,
P1_P3_DATAWIDTH_REG_1_, n5426, n5436, n5441, n5451, n5461, n5471,
n5486, n5491, P1_P3_DATAWIDTH_REG_0_, P1_P3_INSTADDRPOINTER_REG_31_,
P1_P3_REIP_REG_31_, P1_P3_REIP_REG_30_, P1_P3_REIP_REG_29_,
P1_P3_REIP_REG_28_, P1_P3_REIP_REG_27_, P1_P3_REIP_REG_26_,
P1_P3_REIP_REG_25_, P1_P3_REIP_REG_24_, P1_P3_REIP_REG_23_,
P1_P3_REIP_REG_22_, P1_P3_REIP_REG_21_, P1_P3_REIP_REG_20_,
P1_P3_REIP_REG_19_, P1_P3_REIP_REG_18_, P1_P3_REIP_REG_17_,
P1_P3_REIP_REG_16_, P1_P3_REIP_REG_15_, P1_P3_REIP_REG_14_,
P1_P3_REIP_REG_13_, P1_P3_REIP_REG_11_, P1_P3_REIP_REG_10_,
P1_P3_REIP_REG_8_, P1_P3_REIP_REG_7_, P1_P3_REIP_REG_5_,
P1_P3_REIP_REG_4_, P1_P3_REIP_REG_3_, P1_P3_REIP_REG_2_,
P1_P3_INSTQUEUE_REG_0__0_, P1_P3_INSTQUEUE_REG_1__0_,
P1_P3_INSTQUEUE_REG_2__0_, P1_P3_INSTQUEUE_REG_3__0_,
P1_P3_INSTQUEUE_REG_4__0_, P1_P3_INSTQUEUE_REG_5__0_,
P1_P3_INSTQUEUE_REG_6__0_, P1_P3_INSTQUEUE_REG_7__0_,
P1_P3_INSTQUEUE_REG_8__0_, P1_P3_INSTQUEUE_REG_9__0_,
P1_P3_INSTQUEUE_REG_10__0_, P1_P3_INSTQUEUE_REG_11__0_,
P1_P3_INSTQUEUE_REG_12__0_, P1_P3_INSTQUEUE_REG_13__0_,
P1_P3_INSTQUEUE_REG_14__0_, P1_P3_INSTQUEUE_REG_0__1_,
P1_P3_INSTQUEUE_REG_1__1_, P1_P3_INSTQUEUE_REG_2__1_,
P1_P3_INSTQUEUE_REG_3__1_, P1_P3_INSTQUEUE_REG_4__1_,
P1_P3_INSTQUEUE_REG_5__1_, P1_P3_INSTQUEUE_REG_6__1_,
P1_P3_INSTQUEUE_REG_7__1_, P1_P3_INSTQUEUE_REG_8__1_,
P1_P3_INSTQUEUE_REG_9__1_, P1_P3_INSTQUEUE_REG_10__1_,
P1_P3_INSTQUEUE_REG_11__1_, P1_P3_INSTQUEUE_REG_12__1_,
P1_P3_INSTQUEUE_REG_13__1_, P1_P3_INSTQUEUE_REG_14__1_,
P1_P3_INSTQUEUE_REG_0__4_, P1_P3_INSTQUEUE_REG_1__4_,
P1_P3_INSTQUEUE_REG_2__4_, P1_P3_INSTQUEUE_REG_3__4_,
P1_P3_INSTQUEUE_REG_4__4_, P1_P3_INSTQUEUE_REG_5__4_,
P1_P3_INSTQUEUE_REG_6__4_, P1_P3_INSTQUEUE_REG_7__4_,
P1_P3_INSTQUEUE_REG_8__4_, P1_P3_INSTQUEUE_REG_9__4_,
P1_P3_INSTQUEUE_REG_10__4_, P1_P3_INSTQUEUE_REG_11__4_,
P1_P3_INSTQUEUE_REG_12__4_, P1_P3_INSTQUEUE_REG_13__4_,
P1_P3_INSTQUEUE_REG_14__4_, P1_P3_INSTQUEUE_REG_0__2_,
P1_P3_INSTQUEUE_REG_1__2_, P1_P3_INSTQUEUE_REG_2__2_,
P1_P3_INSTQUEUE_REG_3__2_, P1_P3_INSTQUEUE_REG_4__2_,
P1_P3_INSTQUEUE_REG_5__2_, P1_P3_INSTQUEUE_REG_6__2_,
P1_P3_INSTQUEUE_REG_7__2_, P1_P3_INSTQUEUE_REG_8__2_,
P1_P3_INSTQUEUE_REG_9__2_, P1_P3_INSTQUEUE_REG_10__2_,
P1_P3_INSTQUEUE_REG_11__2_, P1_P3_INSTQUEUE_REG_12__2_,
P1_P3_INSTQUEUE_REG_13__2_, P1_P3_INSTQUEUE_REG_14__2_,
P1_P3_INSTQUEUE_REG_0__3_, P1_P3_INSTQUEUE_REG_1__3_,
P1_P3_INSTQUEUE_REG_2__3_, P1_P3_INSTQUEUE_REG_3__3_,
P1_P3_INSTQUEUE_REG_4__3_, P1_P3_INSTQUEUE_REG_5__3_,
P1_P3_INSTQUEUE_REG_6__3_, P1_P3_INSTQUEUE_REG_7__3_,
P1_P3_INSTQUEUE_REG_8__3_, P1_P3_INSTQUEUE_REG_9__3_,
P1_P3_INSTQUEUE_REG_10__3_, P1_P3_INSTQUEUE_REG_11__3_,
P1_P3_INSTQUEUE_REG_12__3_, P1_P3_INSTQUEUE_REG_13__3_,
P1_P3_INSTQUEUE_REG_14__3_, P1_P3_INSTQUEUE_REG_0__7_,
P1_P3_INSTQUEUE_REG_1__7_, P1_P3_INSTQUEUE_REG_2__7_,
P1_P3_INSTQUEUE_REG_3__7_, P1_P3_INSTQUEUE_REG_4__7_,
P1_P3_INSTQUEUE_REG_5__7_, P1_P3_INSTQUEUE_REG_6__7_,
P1_P3_INSTQUEUE_REG_7__7_, P1_P3_INSTQUEUE_REG_8__7_,
P1_P3_INSTQUEUE_REG_9__7_, P1_P3_INSTQUEUE_REG_10__7_,
P1_P3_INSTQUEUE_REG_11__7_, P1_P3_INSTQUEUE_REG_12__7_,
P1_P3_INSTQUEUE_REG_13__7_, P1_P3_INSTQUEUE_REG_14__7_,
P1_P3_INSTQUEUE_REG_0__5_, P1_P3_INSTQUEUE_REG_1__5_,
P1_P3_INSTQUEUE_REG_2__5_, P1_P3_INSTQUEUE_REG_3__5_,
P1_P3_INSTQUEUE_REG_4__5_, P1_P3_INSTQUEUE_REG_5__5_,
P1_P3_INSTQUEUE_REG_6__5_, P1_P3_INSTQUEUE_REG_7__5_,
P1_P3_INSTQUEUE_REG_8__5_, P1_P3_INSTQUEUE_REG_9__5_,
P1_P3_INSTQUEUE_REG_10__5_, P1_P3_INSTQUEUE_REG_11__5_,
P1_P3_INSTQUEUE_REG_12__5_, P1_P3_INSTQUEUE_REG_13__5_,
P1_P3_INSTQUEUE_REG_14__5_, P1_P3_INSTQUEUE_REG_0__6_,
P1_P3_INSTQUEUE_REG_1__6_, P1_P3_INSTQUEUE_REG_2__6_,
P1_P3_INSTQUEUE_REG_3__6_, P1_P3_INSTQUEUE_REG_4__6_,
P1_P3_INSTQUEUE_REG_5__6_, P1_P3_INSTQUEUE_REG_6__6_,
P1_P3_INSTQUEUE_REG_7__6_, P1_P3_INSTQUEUE_REG_8__6_,
P1_P3_INSTQUEUE_REG_9__6_, P1_P3_INSTQUEUE_REG_10__6_,
P1_P3_INSTQUEUE_REG_11__6_, P1_P3_INSTQUEUE_REG_12__6_,
P1_P3_INSTQUEUE_REG_13__6_, P1_P3_INSTQUEUE_REG_14__6_,
P1_P3_MORE_REG, P1_P3_INSTADDRPOINTER_REG_0_,
P1_P3_INSTADDRPOINTER_REG_1_, P1_P3_INSTADDRPOINTER_REG_2_,
P1_P3_INSTADDRPOINTER_REG_3_, P1_P3_INSTADDRPOINTER_REG_4_,
P1_P3_INSTADDRPOINTER_REG_5_, P1_P3_INSTADDRPOINTER_REG_6_,
P1_P3_INSTADDRPOINTER_REG_7_, P1_P3_INSTADDRPOINTER_REG_8_,
P1_P3_INSTADDRPOINTER_REG_9_, P1_P3_INSTADDRPOINTER_REG_10_,
P1_P3_INSTADDRPOINTER_REG_11_, P1_P3_INSTADDRPOINTER_REG_12_,
P1_P3_INSTADDRPOINTER_REG_13_, P1_P3_INSTADDRPOINTER_REG_14_,
P1_P3_INSTADDRPOINTER_REG_15_, P1_P3_INSTADDRPOINTER_REG_16_,
P1_P3_INSTADDRPOINTER_REG_17_, P1_P3_INSTADDRPOINTER_REG_18_,
P1_P3_INSTADDRPOINTER_REG_19_, P1_P3_INSTADDRPOINTER_REG_20_,
P1_P3_INSTADDRPOINTER_REG_21_, P1_P3_INSTADDRPOINTER_REG_22_,
P1_P3_INSTADDRPOINTER_REG_23_, P1_P3_INSTADDRPOINTER_REG_24_,
P1_P3_INSTADDRPOINTER_REG_25_, P1_P3_INSTADDRPOINTER_REG_26_,
P1_P3_INSTADDRPOINTER_REG_27_, P1_P3_INSTADDRPOINTER_REG_28_,
P1_P3_INSTADDRPOINTER_REG_29_, P1_P3_INSTADDRPOINTER_REG_30_,
P1_P3_PHYADDRPOINTER_REG_0_, P1_P3_PHYADDRPOINTER_REG_1_,
P1_P3_PHYADDRPOINTER_REG_2_, P1_P3_PHYADDRPOINTER_REG_3_,
P1_P3_PHYADDRPOINTER_REG_4_, P1_P3_PHYADDRPOINTER_REG_5_,
P1_P3_PHYADDRPOINTER_REG_6_, P1_P3_PHYADDRPOINTER_REG_7_,
P1_P3_PHYADDRPOINTER_REG_8_, P1_P3_PHYADDRPOINTER_REG_9_,
P1_P3_PHYADDRPOINTER_REG_10_, P1_P3_PHYADDRPOINTER_REG_11_,
P1_P3_PHYADDRPOINTER_REG_12_, P1_P3_PHYADDRPOINTER_REG_13_,
P1_P3_PHYADDRPOINTER_REG_14_, P1_P3_PHYADDRPOINTER_REG_15_,
P1_P3_PHYADDRPOINTER_REG_16_, P1_P3_PHYADDRPOINTER_REG_17_,
P1_P3_PHYADDRPOINTER_REG_18_, P1_P3_PHYADDRPOINTER_REG_19_,
P1_P3_PHYADDRPOINTER_REG_20_, P1_P3_PHYADDRPOINTER_REG_21_,
P1_P3_PHYADDRPOINTER_REG_22_, P1_P3_PHYADDRPOINTER_REG_23_,
P1_P3_PHYADDRPOINTER_REG_24_, P1_P3_PHYADDRPOINTER_REG_25_,
P1_P3_PHYADDRPOINTER_REG_26_, P1_P3_PHYADDRPOINTER_REG_27_,
P1_P3_PHYADDRPOINTER_REG_28_, P1_P3_PHYADDRPOINTER_REG_29_,
P1_P3_PHYADDRPOINTER_REG_30_, P1_P3_PHYADDRPOINTER_REG_31_,
P1_P3_EAX_REG_15_, P1_P3_LWORD_REG_15_, P1_P3_EAX_REG_14_,
P1_P3_LWORD_REG_14_, P1_P3_EAX_REG_13_, P1_P3_LWORD_REG_13_,
P1_P3_EAX_REG_12_, P1_P3_LWORD_REG_12_, P1_P3_EAX_REG_11_,
P1_P3_LWORD_REG_11_, P1_P3_LWORD_REG_10_, P1_P3_EAX_REG_9_,
P1_P3_LWORD_REG_9_, P1_P3_EAX_REG_8_, P1_P3_LWORD_REG_8_,
P1_P3_EAX_REG_7_, P1_P3_LWORD_REG_7_, P1_P3_EAX_REG_6_,
P1_P3_LWORD_REG_6_, P1_P3_EAX_REG_5_, P1_P3_LWORD_REG_5_,
P1_P3_EAX_REG_4_, P1_P3_LWORD_REG_4_, P1_P3_EAX_REG_3_,
P1_P3_LWORD_REG_3_, P1_P3_EAX_REG_2_, P1_P3_LWORD_REG_2_,
P1_P3_EAX_REG_1_, P1_P3_LWORD_REG_1_, P1_P3_EAX_REG_0_,
P1_P3_LWORD_REG_0_, P1_P3_EAX_REG_30_, P1_P3_UWORD_REG_14_,
P1_P3_EAX_REG_29_, P1_P3_EAX_REG_28_, P1_P3_EAX_REG_27_,
P1_P3_EAX_REG_26_, P1_P3_EAX_REG_25_, P1_P3_EAX_REG_24_,
P1_P3_EAX_REG_23_, P1_P3_EAX_REG_22_, P1_P3_EAX_REG_21_,
P1_P3_EAX_REG_20_, P1_P3_EAX_REG_19_, P1_P3_UWORD_REG_3_,
P1_P3_EAX_REG_18_, P1_P3_UWORD_REG_2_, P1_P3_EAX_REG_17_,
P1_P3_UWORD_REG_1_, P1_P3_EAX_REG_16_, P1_P3_UWORD_REG_0_,
P1_P3_DATAO_REG_30_, P1_P3_EBX_REG_0_, P1_P3_EBX_REG_1_,
P1_P3_EBX_REG_2_, P1_P3_EBX_REG_3_, P1_P3_EBX_REG_4_,
P1_P3_EBX_REG_5_, P1_P3_EBX_REG_6_, P1_P3_EBX_REG_7_,
P1_P3_EBX_REG_8_, P1_P3_EBX_REG_9_, P1_P3_EBX_REG_10_,
P1_P3_EBX_REG_11_, P1_P3_EBX_REG_12_, P1_P3_EBX_REG_13_,
P1_P3_EBX_REG_14_, P1_P3_EBX_REG_15_, P1_P3_EBX_REG_16_,
P1_P3_EBX_REG_17_, P1_P3_EBX_REG_18_, P1_P3_EBX_REG_19_,
P1_P3_EBX_REG_20_, P1_P3_EBX_REG_21_, P1_P3_EBX_REG_22_,
P1_P3_EBX_REG_23_, P1_P3_EBX_REG_24_, P1_P3_EBX_REG_25_,
P1_P3_EBX_REG_26_, P1_P3_EBX_REG_27_, P1_P3_EBX_REG_28_,
P1_P3_EBX_REG_29_, P1_P3_EBX_REG_30_, P1_P3_BYTEENABLE_REG_3_,
P1_P3_BYTEENABLE_REG_2_, P1_P3_BYTEENABLE_REG_1_,
P1_P3_BYTEENABLE_REG_0_, P1_P3_MEMORYFETCH_REG,
P2_P1_INSTADDRPOINTER_REG_18_, P2_P1_INSTADDRPOINTER_REG_22_,
P2_P1_INSTADDRPOINTER_REG_9_, P2_P1_INSTADDRPOINTER_REG_13_,
P2_P1_INSTADDRPOINTER_REG_20_, P2_P1_INSTADDRPOINTER_REG_1_,
P2_P1_INSTADDRPOINTER_REG_2_, P2_P1_INSTADDRPOINTER_REG_17_,
P2_P1_INSTADDRPOINTER_REG_24_, P2_P1_INSTADDRPOINTER_REG_29_,
P2_P1_INSTADDRPOINTER_REG_30_, P2_P1_INSTADDRPOINTER_REG_6_,
P1_P2_STATEBS16_REG, P1_P2_STATE2_REG_2_, P1_P2_STATE2_REG_3_,
P1_P2_STATE2_REG_1_, P1_P2_STATE2_REG_0_,
P1_P2_INSTQUEUERD_ADDR_REG_3_, P1_P2_INSTQUEUERD_ADDR_REG_2_,
P1_P2_INSTQUEUERD_ADDR_REG_1_, P1_P2_INSTQUEUERD_ADDR_REG_0_,
P1_P2_INSTQUEUEWR_ADDR_REG_0_, P1_P2_INSTQUEUEWR_ADDR_REG_2_,
P1_P2_EBX_REG_31_, P1_P2_INSTQUEUERD_ADDR_REG_4_, n7726, n7721, n7711,
n7701, n7691, n7676, n7666, n7661, n7656, n7651, n7646, n7641, n7636,
n7631, n7626, n7621, n7616, n7611, n7606, n7601, n7596, n7591, n7586,
n7581, n7576, n7571, n7566, n7561, n7556, n7551, n7546, n7541, n7536,
n7531, n7526, n7521, n7516, n7511, n7506, n7501, n7496, n7491, n7486,
n7481, n7476, n7471, n7466, n7461, n7456, n7451, n7446, n7441, n7436,
n7431, n7426, n7421, n7416, n7411, n7406, n7401, n7396, n7391, n7386,
n7381, n7376, n7371, n7366, n7361, n7356, n7351, n7346, n7336, n7331,
n7326, n7321, n7316, n7311, n7306, n7301, n7296, n7291, n7286, n7281,
n7276, n7271, n7266, n7261, n7256, n7251, n7246, n7241, n7236, n7231,
n7226, n7221, n7216, n7211, n7206, n7201, n7196, n7191, n7186, n7181,
n7176, n7171, n7166, n7161, n7156, n7151, n7146, n7141, n7136, n7131,
n7126, n7121, n7116, n7111, n7106, n7101, n7096, n7091, n7086, n7081,
n7076, n7071, n7066, n7061, n7056, n7051, n7046, n7041, n7036, n7031,
n7026, n7021, n7016, n7011, n7006, n7001, n6996, n6991, n6986, n6981,
n6976, n6971, n6966, n6961, n6956, n6951, n6946, n6941, n6936, n6931,
n6926, n6921, n6916, n6911, n6906, n6901, n6896, n6891, n6886, n6881,
n6876, n6871, n6866, n6861, n6856, n6851, n6846, n6841, n6836, n6831,
n6826, n6821, n6816, n6811, n6806, n6801, n6796, n6791, n6786, n6781,
n6776, n6771, n6766, n6761, n6756, n6751, n6746, n6741, n6736, n6731,
n6726, n6721, n6716, n6711, n6706, n6701, n6696, n6691, n6686, n6681,
n6676, n6671, n6666, n6661, n6656, n6651, n6646, n6641, n6636, n6631,
n6626, n6621, n6616, n6611, n6606, n6601, n6596, n6591, n6586, n6581,
n6576, n6571, n6566, n6561, n6556, n6551, n6546, n6541, n6536, n6531,
P1_P2_INSTQUEUEWR_ADDR_REG_4_, n6526, n6496, n6491, n6486, n6481,
n6476, n6471, n6466, n6461, n6456, n6451, n6446, n6441, n6436, n6431,
n6426, n6421, n6416, n6411, n6406, n6401, n6396, n6391, n6386, n6381,
n6376, n6371, n6366, n6361, n6356, n6351, n6346, n6341, n6336, n6331,
n6326, n6321, n6316, n6311, n6306, n6301, n6296, n6291, n6286, n6281,
n6276, n6271, n6266, n6261, n6256, n6251, n6246, n6241, n6236, n6231,
n6226, n6221, n6216, n6211, n6206, n6201, n6196, n6191, n6186, n6181,
n6176, n6171, n6166, n6161, n6156, n6151, n6146, n6141, n6136, n6131,
n6126, n6121, n6116, n6111, n6106, n6101, n6096, n6091, n6086, n6081,
n6076, n6071, n6066, n6061, n6056, n6051, n6046, n6041, n6036, n6031,
n6026, n6021, n6016, n6011, n6006, n6001, n5996, n5991, n5986, n5981,
n5976, n5971, n5966, n5961, n5956, n5951, n5946, n5941, n5936, n5931,
n5926, n5921, n5916, n5911, n5906, n5901, n5896, n5891, n5886, n5881,
n5876, n5871, n5866, n5861, n5856, n5851, n5846, n5836, n5831, n5826,
n5821, n5816, n5811, n5806, n5801, n5796, n5791, n5786, n5781, n5776,
n5771, n5766, n5761, n5756, n5751, n5746, n5741, n5736, n5731, n5726,
n5721, n5716, n5711, n5706, n5701, n5696, n5691, n5676, n5671, n5666,
n5661, n5656, n5651, n5646, n5641, n5636, n5631, n5626, n5621, n5616,
n5611, n5606, n5601, n5596, n5591, n5586, n5581, n5576, n5571, n5566,
n5561, n5556, n5551, n5546, n5541, n5536, n5531, n5526, n5521, n5516,
P1_P2_REQUESTPENDING_REG, P1_P2_STATE_REG_1_, P1_P2_STATE_REG_2_,
P1_P2_REIP_REG_1_, P1_P2_STATE_REG_0_, P1_P2_INSTQUEUEWR_ADDR_REG_1_,
P1_P2_INSTQUEUEWR_ADDR_REG_3_, P1_P2_FLUSH_REG, P1_P2_REIP_REG_0_,
P1_P2_CODEFETCH_REG, P1_P2_READREQUEST_REG, n5496, n5501, n5506,
n5511, n5681, n5686, n5841, n6501, n6506, n6511, n6516, n6521,
P1_P2_DATAWIDTH_REG_1_, n7671, n7681, n7686, n7696, n7706, n7716,
n7731, n7736, P1_P2_DATAWIDTH_REG_0_, P1_P2_INSTADDRPOINTER_REG_31_,
P1_P2_REIP_REG_31_, P1_P2_REIP_REG_30_, P1_P2_ADDRESS_REG_29_,
P1_P2_REIP_REG_29_, P1_P2_ADDRESS_REG_28_, P1_P2_REIP_REG_28_,
P1_P2_ADDRESS_REG_27_, P1_P2_REIP_REG_27_, P1_P2_ADDRESS_REG_26_,
P1_P2_REIP_REG_26_, P1_P2_ADDRESS_REG_25_, P1_P2_REIP_REG_25_,
P1_P2_ADDRESS_REG_24_, P1_P2_REIP_REG_24_, P1_P2_ADDRESS_REG_23_,
P1_P2_REIP_REG_23_, P1_P2_ADDRESS_REG_22_, P1_P2_REIP_REG_22_,
P1_P2_ADDRESS_REG_21_, P1_P2_REIP_REG_21_, P1_P2_ADDRESS_REG_20_,
P1_P2_REIP_REG_20_, P1_P2_ADDRESS_REG_19_, P1_P2_REIP_REG_19_,
P1_P2_REIP_REG_18_, P1_P2_REIP_REG_17_, P1_P2_REIP_REG_16_,
P1_P2_REIP_REG_15_, P1_P2_REIP_REG_14_, P1_P2_REIP_REG_13_,
P1_P2_REIP_REG_11_, P1_P2_REIP_REG_10_, P1_P2_REIP_REG_8_,
P1_P2_REIP_REG_7_, P1_P2_REIP_REG_5_, P1_P2_REIP_REG_4_,
P1_P2_REIP_REG_3_, P1_P2_REIP_REG_2_, P1_P2_INSTQUEUE_REG_0__0_,
P1_P2_INSTQUEUE_REG_1__0_, P1_P2_INSTQUEUE_REG_2__0_,
P1_P2_INSTQUEUE_REG_3__0_, P1_P2_INSTQUEUE_REG_4__0_,
P1_P2_INSTQUEUE_REG_5__0_, P1_P2_INSTQUEUE_REG_6__0_,
P1_P2_INSTQUEUE_REG_7__0_, P1_P2_INSTQUEUE_REG_8__0_,
P1_P2_INSTQUEUE_REG_9__0_, P1_P2_INSTQUEUE_REG_10__0_,
P1_P2_INSTQUEUE_REG_11__0_, P1_P2_INSTQUEUE_REG_12__0_,
P1_P2_INSTQUEUE_REG_13__0_, P1_P2_INSTQUEUE_REG_14__0_,
P1_P2_INSTQUEUE_REG_0__1_, P1_P2_INSTQUEUE_REG_1__1_,
P1_P2_INSTQUEUE_REG_2__1_, P1_P2_INSTQUEUE_REG_3__1_,
P1_P2_INSTQUEUE_REG_4__1_, P1_P2_INSTQUEUE_REG_5__1_,
P1_P2_INSTQUEUE_REG_6__1_, P1_P2_INSTQUEUE_REG_7__1_,
P1_P2_INSTQUEUE_REG_8__1_, P1_P2_INSTQUEUE_REG_9__1_,
P1_P2_INSTQUEUE_REG_10__1_, P1_P2_INSTQUEUE_REG_11__1_,
P1_P2_INSTQUEUE_REG_12__1_, P1_P2_INSTQUEUE_REG_13__1_,
P1_P2_INSTQUEUE_REG_14__1_, P1_P2_INSTQUEUE_REG_0__4_,
P1_P2_INSTQUEUE_REG_1__4_, P1_P2_INSTQUEUE_REG_2__4_,
P1_P2_INSTQUEUE_REG_3__4_, P1_P2_INSTQUEUE_REG_4__4_,
P1_P2_INSTQUEUE_REG_5__4_, P1_P2_INSTQUEUE_REG_6__4_,
P1_P2_INSTQUEUE_REG_7__4_, P1_P2_INSTQUEUE_REG_8__4_,
P1_P2_INSTQUEUE_REG_9__4_, P1_P2_INSTQUEUE_REG_10__4_,
P1_P2_INSTQUEUE_REG_11__4_, P1_P2_INSTQUEUE_REG_12__4_,
P1_P2_INSTQUEUE_REG_13__4_, P1_P2_INSTQUEUE_REG_14__4_,
P1_P2_INSTQUEUE_REG_0__2_, P1_P2_INSTQUEUE_REG_1__2_,
P1_P2_INSTQUEUE_REG_2__2_, P1_P2_INSTQUEUE_REG_3__2_,
P1_P2_INSTQUEUE_REG_4__2_, P1_P2_INSTQUEUE_REG_5__2_,
P1_P2_INSTQUEUE_REG_6__2_, P1_P2_INSTQUEUE_REG_7__2_,
P1_P2_INSTQUEUE_REG_8__2_, P1_P2_INSTQUEUE_REG_9__2_,
P1_P2_INSTQUEUE_REG_10__2_, P1_P2_INSTQUEUE_REG_11__2_,
P1_P2_INSTQUEUE_REG_12__2_, P1_P2_INSTQUEUE_REG_13__2_,
P1_P2_INSTQUEUE_REG_14__2_, P1_P2_INSTQUEUE_REG_0__3_,
P1_P2_INSTQUEUE_REG_1__3_, P1_P2_INSTQUEUE_REG_2__3_,
P1_P2_INSTQUEUE_REG_3__3_, P1_P2_INSTQUEUE_REG_4__3_,
P1_P2_INSTQUEUE_REG_5__3_, P1_P2_INSTQUEUE_REG_6__3_,
P1_P2_INSTQUEUE_REG_7__3_, P1_P2_INSTQUEUE_REG_8__3_,
P1_P2_INSTQUEUE_REG_9__3_, P1_P2_INSTQUEUE_REG_10__3_,
P1_P2_INSTQUEUE_REG_11__3_, P1_P2_INSTQUEUE_REG_12__3_,
P1_P2_INSTQUEUE_REG_13__3_, P1_P2_INSTQUEUE_REG_14__3_,
P1_P2_INSTQUEUE_REG_0__7_, P1_P2_INSTQUEUE_REG_1__7_,
P1_P2_INSTQUEUE_REG_2__7_, P1_P2_INSTQUEUE_REG_3__7_,
P1_P2_INSTQUEUE_REG_4__7_, P1_P2_INSTQUEUE_REG_5__7_,
P1_P2_INSTQUEUE_REG_6__7_, P1_P2_INSTQUEUE_REG_7__7_,
P1_P2_INSTQUEUE_REG_8__7_, P1_P2_INSTQUEUE_REG_9__7_,
P1_P2_INSTQUEUE_REG_10__7_, P1_P2_INSTQUEUE_REG_11__7_,
P1_P2_INSTQUEUE_REG_12__7_, P1_P2_INSTQUEUE_REG_13__7_,
P1_P2_INSTQUEUE_REG_14__7_, P1_P2_INSTQUEUE_REG_0__5_,
P1_P2_INSTQUEUE_REG_1__5_, P1_P2_INSTQUEUE_REG_2__5_,
P1_P2_INSTQUEUE_REG_3__5_, P1_P2_INSTQUEUE_REG_4__5_,
P1_P2_INSTQUEUE_REG_5__5_, P1_P2_INSTQUEUE_REG_6__5_,
P1_P2_INSTQUEUE_REG_7__5_, P1_P2_INSTQUEUE_REG_8__5_,
P1_P2_INSTQUEUE_REG_9__5_, P1_P2_INSTQUEUE_REG_10__5_,
P1_P2_INSTQUEUE_REG_11__5_, P1_P2_INSTQUEUE_REG_12__5_,
P1_P2_INSTQUEUE_REG_13__5_, P1_P2_INSTQUEUE_REG_14__5_,
P1_P2_INSTQUEUE_REG_0__6_, P1_P2_INSTQUEUE_REG_1__6_,
P1_P2_INSTQUEUE_REG_2__6_, P1_P2_INSTQUEUE_REG_3__6_,
P1_P2_INSTQUEUE_REG_4__6_, P1_P2_INSTQUEUE_REG_5__6_,
P1_P2_INSTQUEUE_REG_6__6_, P1_P2_INSTQUEUE_REG_7__6_,
P1_P2_INSTQUEUE_REG_8__6_, P1_P2_INSTQUEUE_REG_9__6_,
P1_P2_INSTQUEUE_REG_10__6_, P1_P2_INSTQUEUE_REG_11__6_,
P1_P2_INSTQUEUE_REG_12__6_, P1_P2_INSTQUEUE_REG_13__6_,
P1_P2_INSTQUEUE_REG_14__6_, P1_P2_MORE_REG,
P1_P2_INSTADDRPOINTER_REG_0_, P1_P2_INSTADDRPOINTER_REG_1_,
P1_P2_INSTADDRPOINTER_REG_2_, P1_P2_INSTADDRPOINTER_REG_3_,
P1_P2_INSTADDRPOINTER_REG_4_, P1_P2_INSTADDRPOINTER_REG_5_,
P1_P2_INSTADDRPOINTER_REG_6_, P1_P2_INSTADDRPOINTER_REG_7_,
P1_P2_INSTADDRPOINTER_REG_8_, P1_P2_INSTADDRPOINTER_REG_9_,
P1_P2_INSTADDRPOINTER_REG_10_, P1_P2_INSTADDRPOINTER_REG_11_,
P1_P2_INSTADDRPOINTER_REG_12_, P1_P2_INSTADDRPOINTER_REG_13_,
P1_P2_INSTADDRPOINTER_REG_14_, P1_P2_INSTADDRPOINTER_REG_15_,
P1_P2_INSTADDRPOINTER_REG_16_, P1_P2_INSTADDRPOINTER_REG_17_,
P1_P2_INSTADDRPOINTER_REG_18_, P1_P2_INSTADDRPOINTER_REG_19_,
P1_P2_INSTADDRPOINTER_REG_20_, P1_P2_INSTADDRPOINTER_REG_21_,
P1_P2_INSTADDRPOINTER_REG_22_, P1_P2_INSTADDRPOINTER_REG_23_,
P1_P2_INSTADDRPOINTER_REG_24_, P1_P2_INSTADDRPOINTER_REG_25_,
P1_P2_INSTADDRPOINTER_REG_26_, P1_P2_INSTADDRPOINTER_REG_27_,
P1_P2_INSTADDRPOINTER_REG_28_, P1_P2_INSTADDRPOINTER_REG_29_,
P1_P2_INSTADDRPOINTER_REG_30_, P1_P2_PHYADDRPOINTER_REG_0_,
P1_P2_PHYADDRPOINTER_REG_1_, P1_P2_PHYADDRPOINTER_REG_2_,
P1_P2_PHYADDRPOINTER_REG_3_, P1_P2_PHYADDRPOINTER_REG_4_,
P1_P2_PHYADDRPOINTER_REG_5_, P1_P2_PHYADDRPOINTER_REG_6_,
P1_P2_PHYADDRPOINTER_REG_7_, P1_P2_PHYADDRPOINTER_REG_8_,
P1_P2_PHYADDRPOINTER_REG_9_, P1_P2_PHYADDRPOINTER_REG_10_,
P1_P2_PHYADDRPOINTER_REG_11_, P1_P2_PHYADDRPOINTER_REG_12_,
P1_P2_PHYADDRPOINTER_REG_13_, P1_P2_PHYADDRPOINTER_REG_14_,
P1_P2_PHYADDRPOINTER_REG_15_, P1_P2_PHYADDRPOINTER_REG_16_,
P1_P2_PHYADDRPOINTER_REG_17_, P1_P2_PHYADDRPOINTER_REG_18_,
P1_P2_PHYADDRPOINTER_REG_19_, P1_P2_PHYADDRPOINTER_REG_20_,
P1_P2_PHYADDRPOINTER_REG_21_, P1_P2_PHYADDRPOINTER_REG_22_,
P1_P2_PHYADDRPOINTER_REG_23_, P1_P2_PHYADDRPOINTER_REG_24_,
P1_P2_PHYADDRPOINTER_REG_25_, P1_P2_PHYADDRPOINTER_REG_26_,
P1_P2_PHYADDRPOINTER_REG_27_, P1_P2_PHYADDRPOINTER_REG_28_,
P1_P2_PHYADDRPOINTER_REG_29_, P1_P2_PHYADDRPOINTER_REG_30_,
P1_P2_PHYADDRPOINTER_REG_31_, P1_P2_EAX_REG_15_, P1_P2_LWORD_REG_15_,
P1_P2_EAX_REG_14_, P1_P2_LWORD_REG_14_, P1_P2_EAX_REG_13_,
P1_P2_LWORD_REG_13_, P1_P2_EAX_REG_12_, P1_P2_LWORD_REG_12_,
P1_P2_EAX_REG_11_, P1_P2_LWORD_REG_11_, P1_P2_LWORD_REG_10_,
P1_P2_EAX_REG_9_, P1_P2_LWORD_REG_9_, P1_P2_EAX_REG_8_,
P1_P2_LWORD_REG_8_, P1_P2_EAX_REG_7_, P1_P2_LWORD_REG_7_,
P1_P2_EAX_REG_6_, P1_P2_LWORD_REG_6_, P1_P2_EAX_REG_5_,
P1_P2_LWORD_REG_5_, P1_P2_EAX_REG_4_, P1_P2_LWORD_REG_4_,
P1_P2_EAX_REG_3_, P1_P2_LWORD_REG_3_, P1_P2_EAX_REG_2_,
P1_P2_LWORD_REG_2_, P1_P2_EAX_REG_1_, P1_P2_LWORD_REG_1_,
P1_P2_EAX_REG_0_, P1_P2_LWORD_REG_0_, P1_P2_EAX_REG_30_,
P1_P2_UWORD_REG_14_, P1_P2_EAX_REG_29_, P1_P2_UWORD_REG_13_,
P1_P2_EAX_REG_28_, P1_P2_UWORD_REG_12_, P1_P2_EAX_REG_27_,
P1_P2_UWORD_REG_11_, P1_P2_EAX_REG_26_, P1_P2_UWORD_REG_10_,
P1_P2_EAX_REG_25_, P1_P2_UWORD_REG_9_, P1_P2_EAX_REG_24_,
P1_P2_UWORD_REG_8_, P1_P2_EAX_REG_23_, P1_P2_UWORD_REG_7_,
P1_P2_EAX_REG_22_, P1_P2_UWORD_REG_6_, P1_P2_EAX_REG_21_,
P1_P2_UWORD_REG_5_, P1_P2_EAX_REG_20_, P1_P2_UWORD_REG_4_,
P1_P2_EAX_REG_19_, P1_P2_UWORD_REG_3_, P1_P2_EAX_REG_18_,
P1_P2_UWORD_REG_2_, P1_P2_EAX_REG_17_, P1_P2_UWORD_REG_1_,
P1_P2_EAX_REG_16_, P1_P2_UWORD_REG_0_, P1_P2_EBX_REG_0_,
P1_P2_EBX_REG_1_, P1_P2_EBX_REG_2_, P1_P2_EBX_REG_3_,
P1_P2_EBX_REG_4_, P1_P2_EBX_REG_5_, P1_P2_EBX_REG_6_,
P1_P2_EBX_REG_7_, P1_P2_EBX_REG_8_, P1_P2_EBX_REG_9_,
P1_P2_EBX_REG_10_, P1_P2_EBX_REG_11_, P1_P2_EBX_REG_12_,
P1_P2_EBX_REG_13_, P1_P2_EBX_REG_14_, P1_P2_EBX_REG_15_,
P1_P2_EBX_REG_16_, P1_P2_EBX_REG_17_, P1_P2_EBX_REG_18_,
P1_P2_EBX_REG_19_, P1_P2_EBX_REG_20_, P1_P2_EBX_REG_21_,
P1_P2_EBX_REG_22_, P1_P2_EBX_REG_23_, P1_P2_EBX_REG_24_,
P1_P2_EBX_REG_25_, P1_P2_EBX_REG_26_, P1_P2_EBX_REG_27_,
P1_P2_EBX_REG_28_, P1_P2_EBX_REG_29_, P1_P2_EBX_REG_30_,
P1_P2_BYTEENABLE_REG_3_, P1_P2_BYTEENABLE_REG_2_,
P1_P2_BYTEENABLE_REG_1_, P1_P2_BYTEENABLE_REG_0_,
P1_P2_MEMORYFETCH_REG, P2_P1_INSTQUEUERD_ADDR_REG_3_,
P2_P1_INSTQUEUERD_ADDR_REG_1_, P2_P1_INSTQUEUERD_ADDR_REG_2_,
P2_P1_INSTQUEUERD_ADDR_REG_4_, P2_P1_INSTADDRPOINTER_REG_0_,
P1_P1_STATEBS16_REG, P1_P1_STATE2_REG_2_, P1_P1_STATE2_REG_3_,
P1_P1_STATE2_REG_1_, P1_P1_STATE2_REG_0_,
P1_P1_INSTQUEUERD_ADDR_REG_3_, P1_P1_INSTQUEUERD_ADDR_REG_2_,
P1_P1_INSTQUEUERD_ADDR_REG_1_, P1_P1_INSTQUEUERD_ADDR_REG_0_,
P1_P1_INSTQUEUEWR_ADDR_REG_0_, P1_P1_INSTQUEUEWR_ADDR_REG_2_,
P1_P1_EBX_REG_31_, P1_P1_INSTQUEUERD_ADDR_REG_4_, n9971, n9966, n9956,
n9946, n9936, n9921, n9911, n9906, n9901, n9896, n9891, n9886, n9881,
n9876, n9871, n9866, n9861, n9856, n9851, n9846, n9841, n9836, n9831,
n9826, n9821, n9816, n9811, n9806, n9801, n9796, n9791, n9786, n9781,
n9776, n9771, n9766, n9761, n9756, n9751, n9746, n9741, n9736, n9731,
n9726, n9721, n9716, n9711, n9706, n9701, n9696, n9691, n9686, n9681,
n9676, n9671, n9666, n9661, n9656, n9651, n9646, n9641, n9636, n9631,
n9626, n9621, n9616, n9611, n9606, n9601, n9596, n9591, n9581, n9576,
n9571, n9566, n9561, n9556, n9551, n9546, n9541, n9536, n9531, n9526,
n9521, n9516, n9511, n9506, n9501, n9496, n9491, n9486, n9481, n9476,
n9471, n9466, n9461, n9456, n9451, n9446, n9441, n9436, n9431, n9426,
n9421, n9416, n9411, n9406, n9401, n9396, n9391, n9386, n9381, n9376,
n9371, n9366, n9361, n9356, n9351, n9346, n9341, n9336, n9331, n9326,
n9321, n9316, n9311, n9306, n9301, n9296, n9291, n9286, n9281, n9276,
n9271, n9266, n9261, n9256, n9251, n9246, n9241, n9236, n9231, n9226,
n9221, n9216, n9211, n9206, n9201, n9196, n9191, n9186, n9181, n9176,
n9171, n9166, n9161, n9156, n9151, n9146, n9141, n9136, n9131, n9126,
n9121, n9116, n9111, n9106, n9101, n9096, n9091, n9086, n9081, n9076,
n9071, n9066, n9061, n9056, n9051, n9046, n9041, n9036, n9031, n9026,
n9021, n9016, n9011, n9006, n9001, n8996, n8991, n8986, n8981, n8976,
n8971, n8966, n8961, n8956, n8951, n8946, n8941, n8936, n8931, n8926,
n8921, n8916, n8911, n8906, n8901, n8896, n8891, n8886, n8881, n8876,
n8871, n8866, n8861, n8856, n8851, n8846, n8841, n8836, n8831, n8826,
n8821, n8816, n8811, n8806, n8801, n8796, n8791, n8786, n8781, n8776,
P1_P1_INSTQUEUEWR_ADDR_REG_4_, n8771, n8741, n8736, n8731, n8726,
n8721, n8716, n8711, n8706, n8701, n8696, n8691, n8686, n8681, n8676,
n8671, n8666, n8661, n8656, n8651, n8646, n8641, n8636, n8631, n8626,
n8621, n8616, n8611, n8606, n8601, n8596, n8591, n8586, n8581, n8576,
n8571, n8566, n8561, n8556, n8551, n8546, n8541, n8536, n8531, n8526,
n8521, n8516, n8511, n8506, n8501, n8496, n8491, n8486, n8481, n8476,
n8471, n8466, n8461, n8456, n8451, n8446, n8441, n8436, n8431, n8426,
n8421, n8416, n8411, n8406, n8401, n8396, n8391, n8386, n8381, n8376,
n8371, n8366, n8361, n8356, n8351, n8346, n8341, n8336, n8331, n8326,
n8321, n8316, n8311, n8306, n8301, n8296, n8291, n8286, n8281, n8276,
n8271, n8266, n8261, n8256, n8251, n8246, n8241, n8236, n8231, n8226,
n8221, n8216, n8211, n8206, n8201, n8196, n8191, n8186, n8181, n8176,
n8171, n8166, n8161, n8156, n8151, n8146, n8141, n8136, n8131, n8126,
n8121, n8116, n8111, n8106, n8101, n8096, n8091, n8081, n8076, n8071,
n8066, n8061, n8056, n8051, n8046, n8041, n8036, n8031, n8026, n8021,
n8016, n8011, n8006, n8001, n7996, n7991, n7986, n7981, n7976, n7971,
n7966, n7961, n7956, n7951, n7946, n7941, n7936, n7921, n7916, n7911,
n7906, n7901, n7896, n7891, n7886, n7881, n7876, n7871, n7866, n7861,
n7856, n7851, n7846, n7841, n7836, n7831, n7826, n7821, n7816, n7811,
n7806, n7801, n7796, n7791, n7786, n7781, n7776, n7771, n7766, n7761,
P1_P1_REQUESTPENDING_REG, P1_P1_STATE_REG_1_, P1_P1_STATE_REG_2_,
P1_P1_REIP_REG_1_, P1_P1_STATE_REG_0_, P1_P1_INSTQUEUEWR_ADDR_REG_1_,
P1_P1_INSTQUEUEWR_ADDR_REG_3_, P1_P1_FLUSH_REG, P1_P1_REIP_REG_0_,
P1_P1_CODEFETCH_REG, P1_P1_READREQUEST_REG, n7741, n7746, n7751,
n7756, n7926, n7931, n8086, n8746, n8751, n8756, n8761, n8766,
P1_P1_DATAWIDTH_REG_1_, n9916, n9926, n9931, n9941, n9951, n9961,
n9976, n9981, P1_P1_DATAWIDTH_REG_0_, P1_P1_INSTADDRPOINTER_REG_31_,
P1_P1_REIP_REG_31_, P1_P1_REIP_REG_30_, P1_P1_ADDRESS_REG_29_,
P1_P1_REIP_REG_29_, P1_P1_ADDRESS_REG_28_, P1_P1_REIP_REG_28_,
P1_P1_ADDRESS_REG_27_, P1_P1_REIP_REG_27_, P1_P1_ADDRESS_REG_26_,
P1_P1_REIP_REG_26_, P1_P1_ADDRESS_REG_25_, P1_P1_REIP_REG_25_,
P1_P1_ADDRESS_REG_24_, P1_P1_REIP_REG_24_, P1_P1_ADDRESS_REG_23_,
P1_P1_REIP_REG_23_, P1_P1_ADDRESS_REG_22_, P1_P1_REIP_REG_22_,
P1_P1_ADDRESS_REG_21_, P1_P1_REIP_REG_21_, P1_P1_ADDRESS_REG_20_,
P1_P1_REIP_REG_20_, P1_P1_ADDRESS_REG_19_, P1_P1_REIP_REG_19_,
P1_P1_REIP_REG_18_, P1_P1_REIP_REG_17_, P1_P1_REIP_REG_16_,
P1_P1_REIP_REG_15_, P1_P1_REIP_REG_14_, P1_P1_REIP_REG_13_,
P1_P1_REIP_REG_11_, P1_P1_REIP_REG_10_, P1_P1_REIP_REG_8_,
P1_P1_REIP_REG_7_, P1_P1_REIP_REG_5_, P1_P1_REIP_REG_4_,
P1_P1_REIP_REG_3_, P1_P1_REIP_REG_2_, P1_P1_INSTQUEUE_REG_0__0_,
P1_P1_INSTQUEUE_REG_1__0_, P1_P1_INSTQUEUE_REG_2__0_,
P1_P1_INSTQUEUE_REG_3__0_, P1_P1_INSTQUEUE_REG_4__0_,
P1_P1_INSTQUEUE_REG_5__0_, P1_P1_INSTQUEUE_REG_6__0_,
P1_P1_INSTQUEUE_REG_7__0_, P1_P1_INSTQUEUE_REG_8__0_,
P1_P1_INSTQUEUE_REG_9__0_, P1_P1_INSTQUEUE_REG_10__0_,
P1_P1_INSTQUEUE_REG_11__0_, P1_P1_INSTQUEUE_REG_12__0_,
P1_P1_INSTQUEUE_REG_13__0_, P1_P1_INSTQUEUE_REG_14__0_,
P1_P1_INSTQUEUE_REG_0__1_, P1_P1_INSTQUEUE_REG_1__1_,
P1_P1_INSTQUEUE_REG_2__1_, P1_P1_INSTQUEUE_REG_3__1_,
P1_P1_INSTQUEUE_REG_4__1_, P1_P1_INSTQUEUE_REG_5__1_,
P1_P1_INSTQUEUE_REG_6__1_, P1_P1_INSTQUEUE_REG_7__1_,
P1_P1_INSTQUEUE_REG_8__1_, P1_P1_INSTQUEUE_REG_9__1_,
P1_P1_INSTQUEUE_REG_10__1_, P1_P1_INSTQUEUE_REG_11__1_,
P1_P1_INSTQUEUE_REG_12__1_, P1_P1_INSTQUEUE_REG_13__1_,
P1_P1_INSTQUEUE_REG_14__1_, P1_P1_INSTQUEUE_REG_0__4_,
P1_P1_INSTQUEUE_REG_1__4_, P1_P1_INSTQUEUE_REG_2__4_,
P1_P1_INSTQUEUE_REG_3__4_, P1_P1_INSTQUEUE_REG_4__4_,
P1_P1_INSTQUEUE_REG_5__4_, P1_P1_INSTQUEUE_REG_6__4_,
P1_P1_INSTQUEUE_REG_7__4_, P1_P1_INSTQUEUE_REG_8__4_,
P1_P1_INSTQUEUE_REG_9__4_, P1_P1_INSTQUEUE_REG_10__4_,
P1_P1_INSTQUEUE_REG_11__4_, P1_P1_INSTQUEUE_REG_12__4_,
P1_P1_INSTQUEUE_REG_13__4_, P1_P1_INSTQUEUE_REG_14__4_,
P1_P1_INSTQUEUE_REG_0__2_, P1_P1_INSTQUEUE_REG_1__2_,
P1_P1_INSTQUEUE_REG_2__2_, P1_P1_INSTQUEUE_REG_3__2_,
P1_P1_INSTQUEUE_REG_4__2_, P1_P1_INSTQUEUE_REG_5__2_,
P1_P1_INSTQUEUE_REG_6__2_, P1_P1_INSTQUEUE_REG_7__2_,
P1_P1_INSTQUEUE_REG_8__2_, P1_P1_INSTQUEUE_REG_9__2_,
P1_P1_INSTQUEUE_REG_10__2_, P1_P1_INSTQUEUE_REG_11__2_,
P1_P1_INSTQUEUE_REG_12__2_, P1_P1_INSTQUEUE_REG_13__2_,
P1_P1_INSTQUEUE_REG_14__2_, P1_P1_INSTQUEUE_REG_0__3_,
P1_P1_INSTQUEUE_REG_1__3_, P1_P1_INSTQUEUE_REG_2__3_,
P1_P1_INSTQUEUE_REG_3__3_, P1_P1_INSTQUEUE_REG_4__3_,
P1_P1_INSTQUEUE_REG_5__3_, P1_P1_INSTQUEUE_REG_6__3_,
P1_P1_INSTQUEUE_REG_7__3_, P1_P1_INSTQUEUE_REG_8__3_,
P1_P1_INSTQUEUE_REG_9__3_, P1_P1_INSTQUEUE_REG_10__3_,
P1_P1_INSTQUEUE_REG_11__3_, P1_P1_INSTQUEUE_REG_12__3_,
P1_P1_INSTQUEUE_REG_13__3_, P1_P1_INSTQUEUE_REG_14__3_,
P1_P1_INSTQUEUE_REG_0__7_, P1_P1_INSTQUEUE_REG_1__7_,
P1_P1_INSTQUEUE_REG_2__7_, P1_P1_INSTQUEUE_REG_3__7_,
P1_P1_INSTQUEUE_REG_4__7_, P1_P1_INSTQUEUE_REG_5__7_,
P1_P1_INSTQUEUE_REG_6__7_, P1_P1_INSTQUEUE_REG_7__7_,
P1_P1_INSTQUEUE_REG_8__7_, P1_P1_INSTQUEUE_REG_9__7_,
P1_P1_INSTQUEUE_REG_10__7_, P1_P1_INSTQUEUE_REG_11__7_,
P1_P1_INSTQUEUE_REG_12__7_, P1_P1_INSTQUEUE_REG_13__7_,
P1_P1_INSTQUEUE_REG_14__7_, P1_P1_INSTQUEUE_REG_0__5_,
P1_P1_INSTQUEUE_REG_1__5_, P1_P1_INSTQUEUE_REG_2__5_,
P1_P1_INSTQUEUE_REG_3__5_, P1_P1_INSTQUEUE_REG_4__5_,
P1_P1_INSTQUEUE_REG_5__5_, P1_P1_INSTQUEUE_REG_6__5_,
P1_P1_INSTQUEUE_REG_7__5_, P1_P1_INSTQUEUE_REG_8__5_,
P1_P1_INSTQUEUE_REG_9__5_, P1_P1_INSTQUEUE_REG_10__5_,
P1_P1_INSTQUEUE_REG_11__5_, P1_P1_INSTQUEUE_REG_12__5_,
P1_P1_INSTQUEUE_REG_13__5_, P1_P1_INSTQUEUE_REG_14__5_,
P1_P1_INSTQUEUE_REG_0__6_, P1_P1_INSTQUEUE_REG_1__6_,
P1_P1_INSTQUEUE_REG_2__6_, P1_P1_INSTQUEUE_REG_3__6_,
P1_P1_INSTQUEUE_REG_4__6_, P1_P1_INSTQUEUE_REG_5__6_,
P1_P1_INSTQUEUE_REG_6__6_, P1_P1_INSTQUEUE_REG_7__6_,
P1_P1_INSTQUEUE_REG_8__6_, P1_P1_INSTQUEUE_REG_9__6_,
P1_P1_INSTQUEUE_REG_10__6_, P1_P1_INSTQUEUE_REG_11__6_,
P1_P1_INSTQUEUE_REG_12__6_, P1_P1_INSTQUEUE_REG_13__6_,
P1_P1_INSTQUEUE_REG_14__6_, P1_P1_MORE_REG,
P1_P1_INSTADDRPOINTER_REG_0_, P1_P1_INSTADDRPOINTER_REG_1_,
P1_P1_INSTADDRPOINTER_REG_2_, P1_P1_INSTADDRPOINTER_REG_3_,
P1_P1_INSTADDRPOINTER_REG_4_, P1_P1_INSTADDRPOINTER_REG_5_,
P1_P1_INSTADDRPOINTER_REG_6_, P1_P1_INSTADDRPOINTER_REG_7_,
P1_P1_INSTADDRPOINTER_REG_8_, P1_P1_INSTADDRPOINTER_REG_9_,
P1_P1_INSTADDRPOINTER_REG_10_, P1_P1_INSTADDRPOINTER_REG_11_,
P1_P1_INSTADDRPOINTER_REG_12_, P1_P1_INSTADDRPOINTER_REG_13_,
P1_P1_INSTADDRPOINTER_REG_14_, P1_P1_INSTADDRPOINTER_REG_15_,
P1_P1_INSTADDRPOINTER_REG_16_, P1_P1_INSTADDRPOINTER_REG_17_,
P1_P1_INSTADDRPOINTER_REG_18_, P1_P1_INSTADDRPOINTER_REG_19_,
P1_P1_INSTADDRPOINTER_REG_20_, P1_P1_INSTADDRPOINTER_REG_21_,
P1_P1_INSTADDRPOINTER_REG_22_, P1_P1_INSTADDRPOINTER_REG_23_,
P1_P1_INSTADDRPOINTER_REG_24_, P1_P1_INSTADDRPOINTER_REG_25_,
P1_P1_INSTADDRPOINTER_REG_26_, P1_P1_INSTADDRPOINTER_REG_27_,
P1_P1_INSTADDRPOINTER_REG_28_, P1_P1_INSTADDRPOINTER_REG_29_,
P1_P1_INSTADDRPOINTER_REG_30_, P1_P1_PHYADDRPOINTER_REG_0_,
P1_P1_PHYADDRPOINTER_REG_1_, P1_P1_PHYADDRPOINTER_REG_2_,
P1_P1_PHYADDRPOINTER_REG_3_, P1_P1_PHYADDRPOINTER_REG_4_,
P1_P1_PHYADDRPOINTER_REG_5_, P1_P1_PHYADDRPOINTER_REG_6_,
P1_P1_PHYADDRPOINTER_REG_7_, P1_P1_PHYADDRPOINTER_REG_8_,
P1_P1_PHYADDRPOINTER_REG_9_, P1_P1_PHYADDRPOINTER_REG_10_,
P1_P1_PHYADDRPOINTER_REG_11_, P1_P1_PHYADDRPOINTER_REG_12_,
P1_P1_PHYADDRPOINTER_REG_13_, P1_P1_PHYADDRPOINTER_REG_14_,
P1_P1_PHYADDRPOINTER_REG_15_, P1_P1_PHYADDRPOINTER_REG_16_,
P1_P1_PHYADDRPOINTER_REG_17_, P1_P1_PHYADDRPOINTER_REG_18_,
P1_P1_PHYADDRPOINTER_REG_19_, P1_P1_PHYADDRPOINTER_REG_20_,
P1_P1_PHYADDRPOINTER_REG_21_, P1_P1_PHYADDRPOINTER_REG_22_,
P1_P1_PHYADDRPOINTER_REG_23_, P1_P1_PHYADDRPOINTER_REG_24_,
P1_P1_PHYADDRPOINTER_REG_25_, P1_P1_PHYADDRPOINTER_REG_26_,
P1_P1_PHYADDRPOINTER_REG_27_, P1_P1_PHYADDRPOINTER_REG_28_,
P1_P1_PHYADDRPOINTER_REG_29_, P1_P1_PHYADDRPOINTER_REG_30_,
P1_P1_PHYADDRPOINTER_REG_31_, P1_P1_LWORD_REG_15_, P1_P1_EAX_REG_14_,
P1_P1_LWORD_REG_14_, P1_P1_EAX_REG_13_, P1_P1_LWORD_REG_13_,
P1_P1_LWORD_REG_12_, P1_P1_EAX_REG_11_, P1_P1_LWORD_REG_11_,
P1_P1_EAX_REG_10_, P1_P1_LWORD_REG_10_, P1_P1_LWORD_REG_9_,
P1_P1_EAX_REG_8_, P1_P1_LWORD_REG_8_, P1_P1_EAX_REG_7_,
P1_P1_LWORD_REG_7_, P1_P1_LWORD_REG_6_, P1_P1_EAX_REG_5_,
P1_P1_LWORD_REG_5_, P1_P1_EAX_REG_4_, P1_P1_LWORD_REG_4_,
P1_P1_LWORD_REG_3_, P1_P1_EAX_REG_2_, P1_P1_LWORD_REG_2_,
P1_P1_LWORD_REG_1_, P1_P1_EAX_REG_0_, P1_P1_LWORD_REG_0_,
P1_P1_EAX_REG_30_, P1_P1_UWORD_REG_14_, P1_P1_EAX_REG_29_,
P1_P1_UWORD_REG_13_, P1_P1_EAX_REG_28_, P1_P1_UWORD_REG_12_,
P1_P1_EAX_REG_27_, P1_P1_UWORD_REG_11_, P1_P1_UWORD_REG_10_,
P1_P1_EAX_REG_25_, P1_P1_UWORD_REG_9_, P1_P1_EAX_REG_24_,
P1_P1_UWORD_REG_8_, P1_P1_UWORD_REG_7_, P1_P1_EAX_REG_22_,
P1_P1_UWORD_REG_6_, P1_P1_EAX_REG_21_, P1_P1_UWORD_REG_5_,
P1_P1_UWORD_REG_4_, P1_P1_EAX_REG_19_, P1_P1_UWORD_REG_3_,
P1_P1_EAX_REG_18_, P1_P1_UWORD_REG_2_, P1_P1_UWORD_REG_1_,
P1_P1_EAX_REG_16_, P1_P1_UWORD_REG_0_, P1_P1_EBX_REG_0_,
P1_P1_EBX_REG_1_, P1_P1_EBX_REG_2_, P1_P1_EBX_REG_3_,
P1_P1_EBX_REG_4_, P1_P1_EBX_REG_5_, P1_P1_EBX_REG_6_,
P1_P1_EBX_REG_7_, P1_P1_EBX_REG_8_, P1_P1_EBX_REG_9_,
P1_P1_EBX_REG_10_, P1_P1_EBX_REG_11_, P1_P1_EBX_REG_12_,
P1_P1_EBX_REG_13_, P1_P1_EBX_REG_14_, P1_P1_EBX_REG_15_,
P1_P1_EBX_REG_16_, P1_P1_EBX_REG_17_, P1_P1_EBX_REG_18_,
P1_P1_EBX_REG_19_, P1_P1_EBX_REG_20_, P1_P1_EBX_REG_21_,
P1_P1_EBX_REG_22_, P1_P1_EBX_REG_23_, P1_P1_EBX_REG_24_,
P1_P1_EBX_REG_25_, P1_P1_EBX_REG_26_, P1_P1_EBX_REG_27_,
P1_P1_EBX_REG_28_, P1_P1_EBX_REG_29_, P1_P1_EBX_REG_30_,
P1_P1_BYTEENABLE_REG_3_, P1_P1_BYTEENABLE_REG_2_,
P1_P1_BYTEENABLE_REG_1_, P1_P1_BYTEENABLE_REG_0_,
P1_P1_MEMORYFETCH_REG, P2_P1_INSTQUEUEWR_ADDR_REG_1_,
P2_P1_INSTQUEUEWR_ADDR_REG_2_, P2_P1_INSTQUEUEWR_ADDR_REG_3_,
P2_P3_STATEBS16_REG, P2_P3_STATE2_REG_2_, P2_P3_STATE2_REG_3_,
P2_P3_STATE2_REG_1_, P2_P3_STATE2_REG_0_,
P2_P3_INSTQUEUERD_ADDR_REG_3_, P2_P3_INSTQUEUERD_ADDR_REG_2_,
P2_P3_INSTQUEUERD_ADDR_REG_1_, P2_P3_INSTQUEUERD_ADDR_REG_0_,
P2_P3_INSTQUEUEWR_ADDR_REG_0_, P2_P3_INSTQUEUEWR_ADDR_REG_2_,
P2_P3_EBX_REG_31_, P2_P3_INSTQUEUERD_ADDR_REG_4_, n12216, n12211,
n12201, n12191, n12181, n12166, n12156, n12151, n12146, n12141,
n12136, n12131, n12126, n12121, n12116, n12111, n12106, n12101,
n12096, n12091, n12086, n12081, n12076, n12071, n12066, n12061,
n12056, n12051, n12046, n12041, n12036, n12031, n12026, n12021,
n12016, n12011, n12006, n12001, n11996, n11991, n11986, n11981,
n11976, n11971, n11966, n11961, n11956, n11951, n11946, n11941,
n11936, n11931, n11926, n11921, n11916, n11911, n11906, n11901,
n11896, n11891, n11886, n11881, n11876, n11871, n11866, n11861,
n11856, n11851, n11846, n11841, n11836, n11826, n11821, n11816,
n11811, n11806, n11801, n11796, n11791, n11786, n11781, n11776,
n11771, n11766, n11761, n11756, n11751, n11746, n11741, n11736,
n11731, n11726, n11721, n11716, n11711, n11706, n11701, n11696,
n11691, n11686, n11681, n11676, n11671, n11666, n11661, n11656,
n11651, n11646, n11641, n11636, n11631, n11626, n11621, n11616,
n11611, n11606, n11601, n11596, n11591, n11586, n11581, n11576,
n11571, n11566, n11561, n11556, n11551, n11546, n11541, n11536,
n11531, n11526, n11521, n11516, n11511, n11506, n11501, n11496,
n11491, n11486, n11481, n11476, n11471, n11466, n11461, n11456,
n11451, n11446, n11441, n11436, n11431, n11426, n11421, n11416,
n11411, n11406, n11401, n11396, n11391, n11386, n11381, n11376,
n11371, n11366, n11361, n11356, n11351, n11346, n11341, n11336,
n11331, n11326, n11321, n11316, n11311, n11306, n11301, n11296,
n11291, n11286, n11281, n11276, n11271, n11266, n11261, n11256,
n11251, n11246, n11241, n11236, n11231, n11226, n11221, n11216,
n11211, n11206, n11201, n11196, n11191, n11186, n11181, n11176,
n11171, n11166, n11161, n11156, n11151, n11146, n11141, n11136,
n11131, n11126, n11121, n11116, n11111, n11106, n11101, n11096,
n11091, n11086, n11081, n11076, n11071, n11066, n11061, n11056,
n11051, n11046, n11041, n11036, n11031, n11026, n11021,
P2_P3_INSTQUEUEWR_ADDR_REG_4_, n11016, n10986, n10981, n10976, n10971,
n10966, n10961, n10956, n10951, n10946, n10941, n10936, n10931,
n10926, n10921, n10916, n10911, n10906, n10901, n10896, n10891,
n10886, n10881, n10876, n10871, n10866, n10861, n10856, n10851,
n10846, n10841, n10836, n10831, n10826, n10821, n10816, n10811,
n10806, n10801, n10796, n10791, n10786, n10781, n10776, n10771,
n10766, n10761, n10756, n10751, n10746, n10741, n10736, n10731,
n10726, n10721, n10716, n10711, n10706, n10701, n10696, n10691,
n10686, n10681, n10676, n10671, n10666, n10661, n10656, n10651,
n10646, n10641, n10636, n10631, n10626, n10621, n10616, n10611,
n10606, n10601, n10596, n10591, n10586, n10581, n10576, n10571,
n10566, n10561, n10556, n10551, n10546, n10541, n10536, n10531,
n10526, n10521, n10516, n10511, n10506, n10501, n10496, n10491,
n10486, n10481, n10476, n10471, n10466, n10461, n10456, n10451,
n10446, n10441, n10436, n10431, n10426, n10421, n10416, n10411,
n10406, n10401, n10396, n10391, n10386, n10381, n10376, n10371,
n10366, n10361, n10356, n10351, n10346, n10341, n10336, n10326,
n10321, n10316, n10311, n10306, n10301, n10296, n10291, n10286,
n10281, n10276, n10271, n10266, n10261, n10256, n10251, n10246,
n10241, n10236, n10231, n10226, n10221, n10216, n10211, n10206,
n10201, n10196, n10191, n10186, n10181, n10166, n10161, n10156,
n10151, n10146, n10141, n10136, n10131, n10126, n10121, n10116,
n10111, n10106, n10101, n10096, n10091, n10086, n10081, n10076,
n10071, n10066, n10061, P2_P3_REQUESTPENDING_REG, P2_P3_STATE_REG_1_,
P2_P3_STATE_REG_2_, P2_P3_REIP_REG_1_, P2_P3_STATE_REG_0_,
P2_P3_INSTQUEUEWR_ADDR_REG_1_, P2_P3_INSTQUEUEWR_ADDR_REG_3_,
P2_P3_FLUSH_REG, P2_P3_REIP_REG_0_, P2_P3_CODEFETCH_REG,
P2_P3_READREQUEST_REG, n9986, n9991, n9996, n10001, n10171, n10176,
n10331, n10991, n10996, n11001, n11006, n11011,
P2_P3_DATAWIDTH_REG_1_, n12161, n12171, n12176, n12186, n12196,
n12206, n12221, n12226, P2_P3_DATAWIDTH_REG_0_,
P2_P3_INSTADDRPOINTER_REG_31_, P2_P3_REIP_REG_31_, P2_P3_REIP_REG_30_,
P2_P3_REIP_REG_29_, P2_P3_REIP_REG_28_, P2_P3_REIP_REG_27_,
P2_P3_REIP_REG_26_, P2_P3_REIP_REG_25_, P2_P3_REIP_REG_24_,
P2_P3_REIP_REG_23_, P2_P3_REIP_REG_22_, P2_P3_REIP_REG_21_,
P2_P3_REIP_REG_20_, P2_P3_REIP_REG_19_, P2_P3_REIP_REG_18_,
P2_P3_REIP_REG_17_, P2_P3_REIP_REG_16_, P2_P3_REIP_REG_15_,
P2_P3_REIP_REG_14_, P2_P3_REIP_REG_13_, P2_P3_REIP_REG_11_,
P2_P3_REIP_REG_10_, P2_P3_REIP_REG_8_, P2_P3_REIP_REG_7_,
P2_P3_REIP_REG_5_, P2_P3_REIP_REG_4_, P2_P3_REIP_REG_3_,
P2_P3_REIP_REG_2_, P2_P3_INSTQUEUE_REG_0__0_,
P2_P3_INSTQUEUE_REG_1__0_, P2_P3_INSTQUEUE_REG_2__0_,
P2_P3_INSTQUEUE_REG_3__0_, P2_P3_INSTQUEUE_REG_4__0_,
P2_P3_INSTQUEUE_REG_5__0_, P2_P3_INSTQUEUE_REG_6__0_,
P2_P3_INSTQUEUE_REG_7__0_, P2_P3_INSTQUEUE_REG_8__0_,
P2_P3_INSTQUEUE_REG_9__0_, P2_P3_INSTQUEUE_REG_10__0_,
P2_P3_INSTQUEUE_REG_11__0_, P2_P3_INSTQUEUE_REG_12__0_,
P2_P3_INSTQUEUE_REG_13__0_, P2_P3_INSTQUEUE_REG_14__0_,
P2_P3_INSTQUEUE_REG_0__1_, P2_P3_INSTQUEUE_REG_1__1_,
P2_P3_INSTQUEUE_REG_2__1_, P2_P3_INSTQUEUE_REG_3__1_,
P2_P3_INSTQUEUE_REG_4__1_, P2_P3_INSTQUEUE_REG_5__1_,
P2_P3_INSTQUEUE_REG_6__1_, P2_P3_INSTQUEUE_REG_7__1_,
P2_P3_INSTQUEUE_REG_8__1_, P2_P3_INSTQUEUE_REG_9__1_,
P2_P3_INSTQUEUE_REG_10__1_, P2_P3_INSTQUEUE_REG_11__1_,
P2_P3_INSTQUEUE_REG_12__1_, P2_P3_INSTQUEUE_REG_13__1_,
P2_P3_INSTQUEUE_REG_14__1_, P2_P3_INSTQUEUE_REG_0__4_,
P2_P3_INSTQUEUE_REG_1__4_, P2_P3_INSTQUEUE_REG_2__4_,
P2_P3_INSTQUEUE_REG_3__4_, P2_P3_INSTQUEUE_REG_4__4_,
P2_P3_INSTQUEUE_REG_5__4_, P2_P3_INSTQUEUE_REG_6__4_,
P2_P3_INSTQUEUE_REG_7__4_, P2_P3_INSTQUEUE_REG_8__4_,
P2_P3_INSTQUEUE_REG_9__4_, P2_P3_INSTQUEUE_REG_10__4_,
P2_P3_INSTQUEUE_REG_11__4_, P2_P3_INSTQUEUE_REG_12__4_,
P2_P3_INSTQUEUE_REG_13__4_, P2_P3_INSTQUEUE_REG_14__4_,
P2_P3_INSTQUEUE_REG_0__2_, P2_P3_INSTQUEUE_REG_1__2_,
P2_P3_INSTQUEUE_REG_2__2_, P2_P3_INSTQUEUE_REG_3__2_,
P2_P3_INSTQUEUE_REG_4__2_, P2_P3_INSTQUEUE_REG_5__2_,
P2_P3_INSTQUEUE_REG_6__2_, P2_P3_INSTQUEUE_REG_7__2_,
P2_P3_INSTQUEUE_REG_8__2_, P2_P3_INSTQUEUE_REG_9__2_,
P2_P3_INSTQUEUE_REG_10__2_, P2_P3_INSTQUEUE_REG_11__2_,
P2_P3_INSTQUEUE_REG_12__2_, P2_P3_INSTQUEUE_REG_13__2_,
P2_P3_INSTQUEUE_REG_14__2_, P2_P3_INSTQUEUE_REG_0__3_,
P2_P3_INSTQUEUE_REG_1__3_, P2_P3_INSTQUEUE_REG_2__3_,
P2_P3_INSTQUEUE_REG_3__3_, P2_P3_INSTQUEUE_REG_4__3_,
P2_P3_INSTQUEUE_REG_5__3_, P2_P3_INSTQUEUE_REG_6__3_,
P2_P3_INSTQUEUE_REG_7__3_, P2_P3_INSTQUEUE_REG_8__3_,
P2_P3_INSTQUEUE_REG_9__3_, P2_P3_INSTQUEUE_REG_10__3_,
P2_P3_INSTQUEUE_REG_11__3_, P2_P3_INSTQUEUE_REG_12__3_,
P2_P3_INSTQUEUE_REG_13__3_, P2_P3_INSTQUEUE_REG_14__3_,
P2_P3_INSTQUEUE_REG_0__7_, P2_P3_INSTQUEUE_REG_1__7_,
P2_P3_INSTQUEUE_REG_2__7_, P2_P3_INSTQUEUE_REG_3__7_,
P2_P3_INSTQUEUE_REG_4__7_, P2_P3_INSTQUEUE_REG_5__7_,
P2_P3_INSTQUEUE_REG_6__7_, P2_P3_INSTQUEUE_REG_7__7_,
P2_P3_INSTQUEUE_REG_8__7_, P2_P3_INSTQUEUE_REG_9__7_,
P2_P3_INSTQUEUE_REG_10__7_, P2_P3_INSTQUEUE_REG_11__7_,
P2_P3_INSTQUEUE_REG_12__7_, P2_P3_INSTQUEUE_REG_13__7_,
P2_P3_INSTQUEUE_REG_14__7_, P2_P3_INSTQUEUE_REG_0__5_,
P2_P3_INSTQUEUE_REG_1__5_, P2_P3_INSTQUEUE_REG_2__5_,
P2_P3_INSTQUEUE_REG_3__5_, P2_P3_INSTQUEUE_REG_4__5_,
P2_P3_INSTQUEUE_REG_5__5_, P2_P3_INSTQUEUE_REG_6__5_,
P2_P3_INSTQUEUE_REG_7__5_, P2_P3_INSTQUEUE_REG_8__5_,
P2_P3_INSTQUEUE_REG_9__5_, P2_P3_INSTQUEUE_REG_10__5_,
P2_P3_INSTQUEUE_REG_11__5_, P2_P3_INSTQUEUE_REG_12__5_,
P2_P3_INSTQUEUE_REG_13__5_, P2_P3_INSTQUEUE_REG_14__5_,
P2_P3_INSTQUEUE_REG_0__6_, P2_P3_INSTQUEUE_REG_1__6_,
P2_P3_INSTQUEUE_REG_2__6_, P2_P3_INSTQUEUE_REG_3__6_,
P2_P3_INSTQUEUE_REG_4__6_, P2_P3_INSTQUEUE_REG_5__6_,
P2_P3_INSTQUEUE_REG_6__6_, P2_P3_INSTQUEUE_REG_7__6_,
P2_P3_INSTQUEUE_REG_8__6_, P2_P3_INSTQUEUE_REG_9__6_,
P2_P3_INSTQUEUE_REG_10__6_, P2_P3_INSTQUEUE_REG_11__6_,
P2_P3_INSTQUEUE_REG_12__6_, P2_P3_INSTQUEUE_REG_13__6_,
P2_P3_INSTQUEUE_REG_14__6_, P2_P3_MORE_REG,
P2_P3_INSTADDRPOINTER_REG_0_, P2_P3_INSTADDRPOINTER_REG_1_,
P2_P3_INSTADDRPOINTER_REG_2_, P2_P3_INSTADDRPOINTER_REG_3_,
P2_P3_INSTADDRPOINTER_REG_4_, P2_P3_INSTADDRPOINTER_REG_5_,
P2_P3_INSTADDRPOINTER_REG_6_, P2_P3_INSTADDRPOINTER_REG_7_,
P2_P3_INSTADDRPOINTER_REG_8_, P2_P3_INSTADDRPOINTER_REG_9_,
P2_P3_INSTADDRPOINTER_REG_10_, P2_P3_INSTADDRPOINTER_REG_11_,
P2_P3_INSTADDRPOINTER_REG_12_, P2_P3_INSTADDRPOINTER_REG_13_,
P2_P3_INSTADDRPOINTER_REG_14_, P2_P3_INSTADDRPOINTER_REG_15_,
P2_P3_INSTADDRPOINTER_REG_16_, P2_P3_INSTADDRPOINTER_REG_17_,
P2_P3_INSTADDRPOINTER_REG_18_, P2_P3_INSTADDRPOINTER_REG_19_,
P2_P3_INSTADDRPOINTER_REG_20_, P2_P3_INSTADDRPOINTER_REG_21_,
P2_P3_INSTADDRPOINTER_REG_22_, P2_P3_INSTADDRPOINTER_REG_23_,
P2_P3_INSTADDRPOINTER_REG_24_, P2_P3_INSTADDRPOINTER_REG_25_,
P2_P3_INSTADDRPOINTER_REG_26_, P2_P3_INSTADDRPOINTER_REG_27_,
P2_P3_INSTADDRPOINTER_REG_28_, P2_P3_INSTADDRPOINTER_REG_29_,
P2_P3_INSTADDRPOINTER_REG_30_, P2_P3_PHYADDRPOINTER_REG_0_,
P2_P3_PHYADDRPOINTER_REG_1_, P2_P3_PHYADDRPOINTER_REG_2_,
P2_P3_PHYADDRPOINTER_REG_3_, P2_P3_PHYADDRPOINTER_REG_4_,
P2_P3_PHYADDRPOINTER_REG_5_, P2_P3_PHYADDRPOINTER_REG_6_,
P2_P3_PHYADDRPOINTER_REG_7_, P2_P3_PHYADDRPOINTER_REG_8_,
P2_P3_PHYADDRPOINTER_REG_9_, P2_P3_PHYADDRPOINTER_REG_10_,
P2_P3_PHYADDRPOINTER_REG_11_, P2_P3_PHYADDRPOINTER_REG_12_,
P2_P3_PHYADDRPOINTER_REG_13_, P2_P3_PHYADDRPOINTER_REG_14_,
P2_P3_PHYADDRPOINTER_REG_15_, P2_P3_PHYADDRPOINTER_REG_16_,
P2_P3_PHYADDRPOINTER_REG_17_, P2_P3_PHYADDRPOINTER_REG_18_,
P2_P3_PHYADDRPOINTER_REG_19_, P2_P3_PHYADDRPOINTER_REG_20_,
P2_P3_PHYADDRPOINTER_REG_21_, P2_P3_PHYADDRPOINTER_REG_22_,
P2_P3_PHYADDRPOINTER_REG_23_, P2_P3_PHYADDRPOINTER_REG_24_,
P2_P3_PHYADDRPOINTER_REG_25_, P2_P3_PHYADDRPOINTER_REG_26_,
P2_P3_PHYADDRPOINTER_REG_27_, P2_P3_PHYADDRPOINTER_REG_28_,
P2_P3_PHYADDRPOINTER_REG_29_, P2_P3_PHYADDRPOINTER_REG_30_,
P2_P3_PHYADDRPOINTER_REG_31_, P2_P3_EAX_REG_15_, P2_P3_LWORD_REG_15_,
P2_P3_EAX_REG_14_, P2_P3_LWORD_REG_14_, P2_P3_EAX_REG_13_,
P2_P3_LWORD_REG_13_, P2_P3_EAX_REG_12_, P2_P3_LWORD_REG_12_,
P2_P3_EAX_REG_11_, P2_P3_LWORD_REG_11_, P2_P3_LWORD_REG_10_,
P2_P3_EAX_REG_9_, P2_P3_LWORD_REG_9_, P2_P3_EAX_REG_8_,
P2_P3_LWORD_REG_8_, P2_P3_EAX_REG_7_, P2_P3_LWORD_REG_7_,
P2_P3_EAX_REG_6_, P2_P3_LWORD_REG_6_, P2_P3_EAX_REG_5_,
P2_P3_LWORD_REG_5_, P2_P3_EAX_REG_4_, P2_P3_LWORD_REG_4_,
P2_P3_EAX_REG_3_, P2_P3_LWORD_REG_3_, P2_P3_EAX_REG_2_,
P2_P3_LWORD_REG_2_, P2_P3_EAX_REG_1_, P2_P3_LWORD_REG_1_,
P2_P3_EAX_REG_0_, P2_P3_LWORD_REG_0_, P2_P3_EAX_REG_30_,
P2_P3_UWORD_REG_14_, P2_P3_EAX_REG_29_, P2_P3_UWORD_REG_13_,
P2_P3_EAX_REG_28_, P2_P3_UWORD_REG_12_, P2_P3_EAX_REG_27_,
P2_P3_UWORD_REG_11_, P2_P3_EAX_REG_26_, P2_P3_UWORD_REG_10_,
P2_P3_EAX_REG_25_, P2_P3_UWORD_REG_9_, P2_P3_EAX_REG_24_,
P2_P3_UWORD_REG_8_, P2_P3_EAX_REG_23_, P2_P3_UWORD_REG_7_,
P2_P3_EAX_REG_22_, P2_P3_UWORD_REG_6_, P2_P3_EAX_REG_21_,
P2_P3_UWORD_REG_5_, P2_P3_EAX_REG_20_, P2_P3_UWORD_REG_4_,
P2_P3_EAX_REG_19_, P2_P3_UWORD_REG_3_, P2_P3_EAX_REG_18_,
P2_P3_UWORD_REG_2_, P2_P3_EAX_REG_17_, P2_P3_UWORD_REG_1_,
P2_P3_EAX_REG_16_, P2_P3_UWORD_REG_0_, P2_P3_EBX_REG_0_,
P2_P3_EBX_REG_1_, P2_P3_EBX_REG_2_, P2_P3_EBX_REG_3_,
P2_P3_EBX_REG_4_, P2_P3_EBX_REG_5_, P2_P3_EBX_REG_6_,
P2_P3_EBX_REG_7_, P2_P3_EBX_REG_8_, P2_P3_EBX_REG_9_,
P2_P3_EBX_REG_10_, P2_P3_EBX_REG_11_, P2_P3_EBX_REG_12_,
P2_P3_EBX_REG_13_, P2_P3_EBX_REG_14_, P2_P3_EBX_REG_15_,
P2_P3_EBX_REG_16_, P2_P3_EBX_REG_17_, P2_P3_EBX_REG_18_,
P2_P3_EBX_REG_19_, P2_P3_EBX_REG_20_, P2_P3_EBX_REG_21_,
P2_P3_EBX_REG_22_, P2_P3_EBX_REG_23_, P2_P3_EBX_REG_24_,
P2_P3_EBX_REG_25_, P2_P3_EBX_REG_26_, P2_P3_EBX_REG_27_,
P2_P3_EBX_REG_28_, P2_P3_EBX_REG_29_, P2_P3_EBX_REG_30_,
P2_P3_BYTEENABLE_REG_3_, P2_P3_BYTEENABLE_REG_2_,
P2_P3_BYTEENABLE_REG_1_, P2_P3_BYTEENABLE_REG_0_,
P2_P3_MEMORYFETCH_REG, P2_P1_INSTQUEUEWR_ADDR_REG_4_,
P2_P1_INSTQUEUEWR_ADDR_REG_0_, P2_P1_INSTQUEUERD_ADDR_REG_0_,
P2_P2_STATEBS16_REG, P2_P2_STATE2_REG_2_, P2_P2_STATE2_REG_3_,
P2_P2_STATE2_REG_1_, P2_P2_STATE2_REG_0_,
P2_P2_INSTQUEUERD_ADDR_REG_3_, P2_P2_INSTQUEUERD_ADDR_REG_2_,
P2_P2_INSTQUEUERD_ADDR_REG_1_, P2_P2_INSTQUEUERD_ADDR_REG_0_,
P2_P2_INSTQUEUEWR_ADDR_REG_0_, P2_P2_INSTQUEUEWR_ADDR_REG_2_,
P2_P2_EBX_REG_31_, P2_P2_INSTQUEUERD_ADDR_REG_4_, n14461, n14456,
n14446, n14436, n14426, n14411, n14401, n14396, n14391, n14386,
n14381, n14376, n14371, n14366, n14361, n14356, n14351, n14346,
n14341, n14336, n14331, n14326, n14321, n14316, n14311, n14306,
n14301, n14296, n14291, n14286, n14281, n14276, n14271, n14266,
n14261, n14256, n14251, n14246, n14241, n14236, n14231, n14226,
n14221, n14216, n14211, n14206, n14201, n14196, n14191, n14186,
n14181, n14176, n14171, n14166, n14161, n14156, n14151, n14146,
n14141, n14136, n14131, n14126, n14121, n14116, n14111, n14106,
n14101, n14096, n14091, n14086, n14081, n14071, n14066, n14061,
n14056, n14051, n14046, n14041, n14036, n14031, n14026, n14021,
n14016, n14011, n14006, n14001, n13996, n13991, n13986, n13981,
n13976, n13971, n13966, n13961, n13956, n13951, n13946, n13941,
n13936, n13931, n13926, n13921, n13916, n13911, n13906, n13901,
n13896, n13891, n13886, n13881, n13876, n13871, n13866, n13861,
n13856, n13851, n13846, n13841, n13836, n13831, n13826, n13821,
n13816, n13811, n13806, n13801, n13796, n13791, n13786, n13781,
n13776, n13771, n13766, n13761, n13756, n13751, n13746, n13741,
n13736, n13731, n13726, n13721, n13716, n13711, n13706, n13701,
n13696, n13691, n13686, n13681, n13676, n13671, n13666, n13661,
n13656, n13651, n13646, n13641, n13636, n13631, n13626, n13621,
n13616, n13611, n13606, n13601, n13596, n13591, n13586, n13581,
n13576, n13571, n13566, n13561, n13556, n13551, n13546, n13541,
n13536, n13531, n13526, n13521, n13516, n13511, n13506, n13501,
n13496, n13491, n13486, n13481, n13476, n13471, n13466, n13461,
n13456, n13451, n13446, n13441, n13436, n13431, n13426, n13421,
n13416, n13411, n13406, n13401, n13396, n13391, n13386, n13381,
n13376, n13371, n13366, n13361, n13356, n13351, n13346, n13341,
n13336, n13331, n13326, n13321, n13316, n13311, n13306, n13301,
n13296, n13291, n13286, n13281, n13276, n13271, n13266,
P2_P2_INSTQUEUEWR_ADDR_REG_4_, n13261, n13231, n13226, n13221, n13216,
n13211, n13206, n13201, n13196, n13191, n13186, n13181, n13176,
n13171, n13166, n13161, n13156, n13151, n13146, n13141, n13136,
n13131, n13126, n13121, n13116, n13111, n13106, n13101, n13096,
n13091, n13086, n13081, n13076, n13071, n13066, n13061, n13056,
n13051, n13046, n13041, n13036, n13031, n13026, n13021, n13016,
n13011, n13006, n13001, n12996, n12991, n12986, n12981, n12976,
n12971, n12966, n12961, n12956, n12951, n12946, n12941, n12936,
n12931, n12926, n12921, n12916, n12911, n12906, n12901, n12896,
n12891, n12886, n12881, n12876, n12871, n12866, n12861, n12856,
n12851, n12846, n12841, n12836, n12831, n12826, n12821, n12816,
n12811, n12806, n12801, n12796, n12791, n12786, n12781, n12776,
n12771, n12766, n12761, n12756, n12751, n12746, n12741, n12736,
n12731, n12726, n12721, n12716, n12711, n12706, n12701, n12696,
n12691, n12686, n12681, n12676, n12671, n12666, n12661, n12656,
n12651, n12646, n12641, n12636, n12631, n12626, n12621, n12616,
n12611, n12606, n12601, n12596, n12591, n12586, n12581, n12571,
n12566, n12561, n12556, n12551, n12546, n12541, n12536, n12531,
n12526, n12521, n12516, n12511, n12506, n12501, n12496, n12491,
n12486, n12481, n12476, n12471, n12466, n12461, n12456, n12451,
n12446, n12441, n12436, n12431, n12426, n12411, n12406, n12401,
n12396, n12391, n12386, n12381, n12376, n12371, n12366, n12361,
n12356, n12351, n12346, n12341, n12336, n12331, n12326, n12321,
n12316, n12311, n12306, n12301, n12296, n12291, n12286, n12281,
n12276, n12271, n12266, n12261, n12256, n12251,
P2_P2_REQUESTPENDING_REG, P2_P2_STATE_REG_1_, P2_P2_STATE_REG_2_,
P2_P2_REIP_REG_1_, P2_P2_STATE_REG_0_, P2_P2_INSTQUEUEWR_ADDR_REG_1_,
P2_P2_INSTQUEUEWR_ADDR_REG_3_, P2_P2_FLUSH_REG, P2_P2_REIP_REG_0_,
P2_P2_CODEFETCH_REG, P2_P2_READREQUEST_REG, n12231, n12236, n12241,
n12246, n12416, n12421, n12576, n13236, n13241, n13246, n13251,
n13256, P2_P2_DATAWIDTH_REG_1_, n14406, n14416, n14421, n14431,
n14441, n14451, n14466, n14471, P2_P2_DATAWIDTH_REG_0_,
P2_P2_INSTADDRPOINTER_REG_31_, P2_P2_REIP_REG_31_, P2_P2_REIP_REG_30_,
P2_P2_ADDRESS_REG_29_, P2_P2_REIP_REG_29_, P2_P2_ADDRESS_REG_28_,
P2_P2_REIP_REG_28_, P2_P2_ADDRESS_REG_27_, P2_P2_REIP_REG_27_,
P2_P2_ADDRESS_REG_26_, P2_P2_REIP_REG_26_, P2_P2_ADDRESS_REG_25_,
P2_P2_REIP_REG_25_, P2_P2_ADDRESS_REG_24_, P2_P2_REIP_REG_24_,
P2_P2_ADDRESS_REG_23_, P2_P2_REIP_REG_23_, P2_P2_ADDRESS_REG_22_,
P2_P2_REIP_REG_22_, P2_P2_ADDRESS_REG_21_, P2_P2_REIP_REG_21_,
P2_P2_ADDRESS_REG_20_, P2_P2_REIP_REG_20_, P2_P2_ADDRESS_REG_19_,
P2_P2_REIP_REG_19_, P2_P2_REIP_REG_18_, P2_P2_REIP_REG_17_,
P2_P2_REIP_REG_16_, P2_P2_REIP_REG_15_, P2_P2_REIP_REG_14_,
P2_P2_REIP_REG_13_, P2_P2_REIP_REG_11_, P2_P2_REIP_REG_10_,
P2_P2_REIP_REG_8_, P2_P2_REIP_REG_7_, P2_P2_REIP_REG_5_,
P2_P2_REIP_REG_4_, P2_P2_REIP_REG_3_, P2_P2_REIP_REG_2_,
P2_P2_INSTQUEUE_REG_0__0_, P2_P2_INSTQUEUE_REG_1__0_,
P2_P2_INSTQUEUE_REG_2__0_, P2_P2_INSTQUEUE_REG_3__0_,
P2_P2_INSTQUEUE_REG_4__0_, P2_P2_INSTQUEUE_REG_5__0_,
P2_P2_INSTQUEUE_REG_6__0_, P2_P2_INSTQUEUE_REG_7__0_,
P2_P2_INSTQUEUE_REG_8__0_, P2_P2_INSTQUEUE_REG_9__0_,
P2_P2_INSTQUEUE_REG_10__0_, P2_P2_INSTQUEUE_REG_11__0_,
P2_P2_INSTQUEUE_REG_12__0_, P2_P2_INSTQUEUE_REG_13__0_,
P2_P2_INSTQUEUE_REG_14__0_, P2_P2_INSTQUEUE_REG_0__1_,
P2_P2_INSTQUEUE_REG_1__1_, P2_P2_INSTQUEUE_REG_2__1_,
P2_P2_INSTQUEUE_REG_3__1_, P2_P2_INSTQUEUE_REG_4__1_,
P2_P2_INSTQUEUE_REG_5__1_, P2_P2_INSTQUEUE_REG_6__1_,
P2_P2_INSTQUEUE_REG_7__1_, P2_P2_INSTQUEUE_REG_8__1_,
P2_P2_INSTQUEUE_REG_9__1_, P2_P2_INSTQUEUE_REG_10__1_,
P2_P2_INSTQUEUE_REG_11__1_, P2_P2_INSTQUEUE_REG_12__1_,
P2_P2_INSTQUEUE_REG_13__1_, P2_P2_INSTQUEUE_REG_14__1_,
P2_P2_INSTQUEUE_REG_0__4_, P2_P2_INSTQUEUE_REG_1__4_,
P2_P2_INSTQUEUE_REG_2__4_, P2_P2_INSTQUEUE_REG_3__4_,
P2_P2_INSTQUEUE_REG_4__4_, P2_P2_INSTQUEUE_REG_5__4_,
P2_P2_INSTQUEUE_REG_6__4_, P2_P2_INSTQUEUE_REG_7__4_,
P2_P2_INSTQUEUE_REG_8__4_, P2_P2_INSTQUEUE_REG_9__4_,
P2_P2_INSTQUEUE_REG_10__4_, P2_P2_INSTQUEUE_REG_11__4_,
P2_P2_INSTQUEUE_REG_12__4_, P2_P2_INSTQUEUE_REG_13__4_,
P2_P2_INSTQUEUE_REG_14__4_, P2_P2_INSTQUEUE_REG_0__2_,
P2_P2_INSTQUEUE_REG_1__2_, P2_P2_INSTQUEUE_REG_2__2_,
P2_P2_INSTQUEUE_REG_3__2_, P2_P2_INSTQUEUE_REG_4__2_,
P2_P2_INSTQUEUE_REG_5__2_, P2_P2_INSTQUEUE_REG_6__2_,
P2_P2_INSTQUEUE_REG_7__2_, P2_P2_INSTQUEUE_REG_8__2_,
P2_P2_INSTQUEUE_REG_9__2_, P2_P2_INSTQUEUE_REG_10__2_,
P2_P2_INSTQUEUE_REG_11__2_, P2_P2_INSTQUEUE_REG_12__2_,
P2_P2_INSTQUEUE_REG_13__2_, P2_P2_INSTQUEUE_REG_14__2_,
P2_P2_INSTQUEUE_REG_0__3_, P2_P2_INSTQUEUE_REG_1__3_,
P2_P2_INSTQUEUE_REG_2__3_, P2_P2_INSTQUEUE_REG_3__3_,
P2_P2_INSTQUEUE_REG_4__3_, P2_P2_INSTQUEUE_REG_5__3_,
P2_P2_INSTQUEUE_REG_6__3_, P2_P2_INSTQUEUE_REG_7__3_,
P2_P2_INSTQUEUE_REG_8__3_, P2_P2_INSTQUEUE_REG_9__3_,
P2_P2_INSTQUEUE_REG_10__3_, P2_P2_INSTQUEUE_REG_11__3_,
P2_P2_INSTQUEUE_REG_12__3_, P2_P2_INSTQUEUE_REG_13__3_,
P2_P2_INSTQUEUE_REG_14__3_, P2_P2_INSTQUEUE_REG_0__7_,
P2_P2_INSTQUEUE_REG_1__7_, P2_P2_INSTQUEUE_REG_2__7_,
P2_P2_INSTQUEUE_REG_3__7_, P2_P2_INSTQUEUE_REG_4__7_,
P2_P2_INSTQUEUE_REG_5__7_, P2_P2_INSTQUEUE_REG_6__7_,
P2_P2_INSTQUEUE_REG_7__7_, P2_P2_INSTQUEUE_REG_8__7_,
P2_P2_INSTQUEUE_REG_9__7_, P2_P2_INSTQUEUE_REG_10__7_,
P2_P2_INSTQUEUE_REG_11__7_, P2_P2_INSTQUEUE_REG_12__7_,
P2_P2_INSTQUEUE_REG_13__7_, P2_P2_INSTQUEUE_REG_14__7_,
P2_P2_INSTQUEUE_REG_0__5_, P2_P2_INSTQUEUE_REG_1__5_,
P2_P2_INSTQUEUE_REG_2__5_, P2_P2_INSTQUEUE_REG_3__5_,
P2_P2_INSTQUEUE_REG_4__5_, P2_P2_INSTQUEUE_REG_5__5_,
P2_P2_INSTQUEUE_REG_6__5_, P2_P2_INSTQUEUE_REG_7__5_,
P2_P2_INSTQUEUE_REG_8__5_, P2_P2_INSTQUEUE_REG_9__5_,
P2_P2_INSTQUEUE_REG_10__5_, P2_P2_INSTQUEUE_REG_11__5_,
P2_P2_INSTQUEUE_REG_12__5_, P2_P2_INSTQUEUE_REG_13__5_,
P2_P2_INSTQUEUE_REG_14__5_, P2_P2_INSTQUEUE_REG_0__6_,
P2_P2_INSTQUEUE_REG_1__6_, P2_P2_INSTQUEUE_REG_2__6_,
P2_P2_INSTQUEUE_REG_3__6_, P2_P2_INSTQUEUE_REG_4__6_,
P2_P2_INSTQUEUE_REG_5__6_, P2_P2_INSTQUEUE_REG_6__6_,
P2_P2_INSTQUEUE_REG_7__6_, P2_P2_INSTQUEUE_REG_8__6_,
P2_P2_INSTQUEUE_REG_9__6_, P2_P2_INSTQUEUE_REG_10__6_,
P2_P2_INSTQUEUE_REG_11__6_, P2_P2_INSTQUEUE_REG_12__6_,
P2_P2_INSTQUEUE_REG_13__6_, P2_P2_INSTQUEUE_REG_14__6_,
P2_P2_MORE_REG, P2_P2_INSTADDRPOINTER_REG_0_,
P2_P2_INSTADDRPOINTER_REG_1_, P2_P2_INSTADDRPOINTER_REG_2_,
P2_P2_INSTADDRPOINTER_REG_3_, P2_P2_INSTADDRPOINTER_REG_4_,
P2_P2_INSTADDRPOINTER_REG_5_, P2_P2_INSTADDRPOINTER_REG_6_,
P2_P2_INSTADDRPOINTER_REG_7_, P2_P2_INSTADDRPOINTER_REG_8_,
P2_P2_INSTADDRPOINTER_REG_9_, P2_P2_INSTADDRPOINTER_REG_10_,
P2_P2_INSTADDRPOINTER_REG_11_, P2_P2_INSTADDRPOINTER_REG_12_,
P2_P2_INSTADDRPOINTER_REG_13_, P2_P2_INSTADDRPOINTER_REG_14_,
P2_P2_INSTADDRPOINTER_REG_15_, P2_P2_INSTADDRPOINTER_REG_16_,
P2_P2_INSTADDRPOINTER_REG_17_, P2_P2_INSTADDRPOINTER_REG_18_,
P2_P2_INSTADDRPOINTER_REG_19_, P2_P2_INSTADDRPOINTER_REG_20_,
P2_P2_INSTADDRPOINTER_REG_21_, P2_P2_INSTADDRPOINTER_REG_22_,
P2_P2_INSTADDRPOINTER_REG_23_, P2_P2_INSTADDRPOINTER_REG_24_,
P2_P2_INSTADDRPOINTER_REG_25_, P2_P2_INSTADDRPOINTER_REG_26_,
P2_P2_INSTADDRPOINTER_REG_27_, P2_P2_INSTADDRPOINTER_REG_28_,
P2_P2_INSTADDRPOINTER_REG_29_, P2_P2_INSTADDRPOINTER_REG_30_,
P2_P2_PHYADDRPOINTER_REG_0_, P2_P2_PHYADDRPOINTER_REG_1_,
P2_P2_PHYADDRPOINTER_REG_2_, P2_P2_PHYADDRPOINTER_REG_3_,
P2_P2_PHYADDRPOINTER_REG_4_, P2_P2_PHYADDRPOINTER_REG_5_,
P2_P2_PHYADDRPOINTER_REG_6_, P2_P2_PHYADDRPOINTER_REG_7_,
P2_P2_PHYADDRPOINTER_REG_8_, P2_P2_PHYADDRPOINTER_REG_9_,
P2_P2_PHYADDRPOINTER_REG_10_, P2_P2_PHYADDRPOINTER_REG_11_,
P2_P2_PHYADDRPOINTER_REG_12_, P2_P2_PHYADDRPOINTER_REG_13_,
P2_P2_PHYADDRPOINTER_REG_14_, P2_P2_PHYADDRPOINTER_REG_15_,
P2_P2_PHYADDRPOINTER_REG_16_, P2_P2_PHYADDRPOINTER_REG_17_,
P2_P2_PHYADDRPOINTER_REG_18_, P2_P2_PHYADDRPOINTER_REG_19_,
P2_P2_PHYADDRPOINTER_REG_20_, P2_P2_PHYADDRPOINTER_REG_21_,
P2_P2_PHYADDRPOINTER_REG_22_, P2_P2_PHYADDRPOINTER_REG_23_,
P2_P2_PHYADDRPOINTER_REG_24_, P2_P2_PHYADDRPOINTER_REG_25_,
P2_P2_PHYADDRPOINTER_REG_26_, P2_P2_PHYADDRPOINTER_REG_27_,
P2_P2_PHYADDRPOINTER_REG_28_, P2_P2_PHYADDRPOINTER_REG_29_,
P2_P2_PHYADDRPOINTER_REG_30_, P2_P2_PHYADDRPOINTER_REG_31_,
P2_P2_EAX_REG_15_, P2_P2_LWORD_REG_15_, P2_P2_EAX_REG_14_,
P2_P2_LWORD_REG_14_, P2_P2_EAX_REG_13_, P2_P2_LWORD_REG_13_,
P2_P2_EAX_REG_12_, P2_P2_LWORD_REG_12_, P2_P2_EAX_REG_11_,
P2_P2_LWORD_REG_11_, P2_P2_LWORD_REG_10_, P2_P2_EAX_REG_9_,
P2_P2_LWORD_REG_9_, P2_P2_EAX_REG_8_, P2_P2_LWORD_REG_8_,
P2_P2_EAX_REG_7_, P2_P2_LWORD_REG_7_, P2_P2_EAX_REG_6_,
P2_P2_LWORD_REG_6_, P2_P2_EAX_REG_5_, P2_P2_LWORD_REG_5_,
P2_P2_EAX_REG_4_, P2_P2_LWORD_REG_4_, P2_P2_EAX_REG_3_,
P2_P2_LWORD_REG_3_, P2_P2_EAX_REG_2_, P2_P2_LWORD_REG_2_,
P2_P2_EAX_REG_1_, P2_P2_LWORD_REG_1_, P2_P2_EAX_REG_0_,
P2_P2_LWORD_REG_0_, P2_P2_EAX_REG_30_, P2_P2_UWORD_REG_14_,
P2_P2_EAX_REG_29_, P2_P2_UWORD_REG_13_, P2_P2_EAX_REG_28_,
P2_P2_UWORD_REG_12_, P2_P2_EAX_REG_27_, P2_P2_UWORD_REG_11_,
P2_P2_EAX_REG_26_, P2_P2_UWORD_REG_10_, P2_P2_EAX_REG_25_,
P2_P2_UWORD_REG_9_, P2_P2_EAX_REG_24_, P2_P2_UWORD_REG_8_,
P2_P2_EAX_REG_23_, P2_P2_UWORD_REG_7_, P2_P2_EAX_REG_22_,
P2_P2_UWORD_REG_6_, P2_P2_EAX_REG_21_, P2_P2_UWORD_REG_5_,
P2_P2_EAX_REG_20_, P2_P2_UWORD_REG_4_, P2_P2_EAX_REG_19_,
P2_P2_UWORD_REG_3_, P2_P2_EAX_REG_18_, P2_P2_UWORD_REG_2_,
P2_P2_EAX_REG_17_, P2_P2_UWORD_REG_1_, P2_P2_EAX_REG_16_,
P2_P2_UWORD_REG_0_, P2_P2_EBX_REG_0_, P2_P2_EBX_REG_1_,
P2_P2_EBX_REG_2_, P2_P2_EBX_REG_3_, P2_P2_EBX_REG_4_,
P2_P2_EBX_REG_5_, P2_P2_EBX_REG_6_, P2_P2_EBX_REG_7_,
P2_P2_EBX_REG_8_, P2_P2_EBX_REG_9_, P2_P2_EBX_REG_10_,
P2_P2_EBX_REG_11_, P2_P2_EBX_REG_12_, P2_P2_EBX_REG_13_,
P2_P2_EBX_REG_14_, P2_P2_EBX_REG_15_, P2_P2_EBX_REG_16_,
P2_P2_EBX_REG_17_, P2_P2_EBX_REG_18_, P2_P2_EBX_REG_19_,
P2_P2_EBX_REG_20_, P2_P2_EBX_REG_21_, P2_P2_EBX_REG_22_,
P2_P2_EBX_REG_23_, P2_P2_EBX_REG_24_, P2_P2_EBX_REG_25_,
P2_P2_EBX_REG_26_, P2_P2_EBX_REG_27_, P2_P2_EBX_REG_28_,
P2_P2_EBX_REG_29_, P2_P2_EBX_REG_30_, P2_P2_BYTEENABLE_REG_3_,
P2_P2_BYTEENABLE_REG_2_, P2_P2_BYTEENABLE_REG_1_,
P2_P2_BYTEENABLE_REG_0_, P2_P2_MEMORYFETCH_REG, P2_P1_STATEBS16_REG,
P2_P1_STATE2_REG_2_, P2_P1_STATE2_REG_3_, P2_P1_STATE2_REG_1_,
P2_P1_STATE2_REG_0_, P2_P1_EBX_REG_31_, n16706, n16701, n16691,
n16681, n16671, n16656, n16646, n16641, n16636, n16631, n16626,
n16621, n16616, n16611, n16606, n16601, n16596, n16591, n16586,
n16581, n16576, n16571, n16566, n16561, n16556, n16551, n16546,
n16541, n16536, n16531, n16526, n16521, n16516, n16511, n16506,
n16501, n16496, n16491, n16486, n16481, n16476, n16471, n16466,
n16461, n16456, n16451, n16446, n16441, n16436, n16431, n16426,
n16421, n16416, n16411, n16406, n16401, n16396, n16391, n16386,
n16381, n16376, n16371, n16366, n16361, n16356, n16351, n16346,
n16341, n16336, n16331, n16326, n16316, n16311, n16306, n16301,
n16296, n16291, n16286, n16281, n16276, n16271, n16266, n16261,
n16256, n16251, n16246, n16241, n16236, n16231, n16226, n16221,
n16216, n16211, n16206, n16201, n16196, n16191, n16186, n16181,
n16176, n16171, n16166, n16161, n16156, n16151, n16146, n16141,
n16136, n16131, n16126, n16121, n16116, n16111, n16106, n16101,
n16096, n16091, n16086, n16081, n16076, n16071, n16066, n16061,
n16056, n16051, n16046, n16041, n16036, n16031, n16026, n16021,
n16016, n16011, n16006, n16001, n15996, n15991, n15986, n15981,
n15976, n15971, n15966, n15961, n15956, n15951, n15946, n15941,
n15936, n15931, n15926, n15921, n15916, n15911, n15906, n15901,
n15896, n15891, n15886, n15881, n15876, n15871, n15866, n15861,
n15856, n15851, n15846, n15841, n15836, n15831, n15826, n15821,
n15816, n15811, n15806, n15801, n15796, n15791, n15786, n15781,
n15776, n15771, n15766, n15761, n15756, n15751, n15746, n15741,
n15736, n15731, n15726, n15721, n15716, n15711, n15706, n15701,
n15696, n15691, n15686, n15681, n15676, n15671, n15666, n15661,
n15656, n15651, n15646, n15641, n15636, n15631, n15626, n15621,
n15616, n15611, n15606, n15601, n15596, n15591, n15586, n15581,
n15576, n15571, n15566, n15561, n15556, n15551, n15546, n15541,
n15536, n15531, n15526, n15521, n15516, n15511, n15506, n15476,
n15471, n15466, n15461, n15456, n15451, n15446, n15441, n15436,
n15431, n15426, n15421, n15416, n15411, n15406, n15401, n15396,
n15391, n15386, n15381, n15376, n15371, n15366, n15361, n15356,
n15351, n15346, n15341, n15336, n15331, n15326, n15321, n15316,
n15311, n15306, n15301, n15296, n15291, n15286, n15281, n15276,
n15271, n15266, n15261, n15256, n15251, n15246, n15241, n15236,
n15231, n15226, n15221, n15216, n15211, n15206, n15201, n15196,
n15191, n15186, n15181, n15176, n15171, n15166, n15161, n15156,
n15151, n15146, n15141, n15136, n15131, n15126, n15121, n15116,
n15111, n15106, n15101, n15096, n15091, n15086, n15081, n15076,
n15071, n15066, n15061, n15056, n15051, n15046, n15041, n15036,
n15031, n15026, n15021, n15016, n15011, n15006, n15001, n14996,
n14991, n14986, n14981, n14976, n14971, n14966, n14961, n14956,
n14951, n14946, n14941, n14936, n14931, n14926, n14921, n14916,
n14911, n14906, n14901, n14896, n14891, n14886, n14881, n14876,
n14871, n14866, n14861, n14856, n14851, n14846, n14841, n14836,
n14831, n14826, n14816, n14811, n14806, n14801, n14796, n14791,
n14786, n14781, n14776, n14771, n14766, n14761, n14756, n14751,
n14746, n14741, n14736, n14731, n14726, n14721, n14716, n14711,
n14706, n14701, n14696, n14691, n14686, n14681, n14676, n14671,
n14656, n14651, n14646, n14641, n14636, n14631, n14626, n14621,
n14616, n14611, n14606, n14601, n14596, n14591, n14586, n14581,
n14576, n14571, n14566, n14561, n14556, n14551, n14546, n14541,
n14536, n14531, n14526, n14521, n14516, n14511, n14506, n14501,
n14496, P2_P1_REQUESTPENDING_REG, P2_P1_STATE_REG_1_,
P2_P1_STATE_REG_2_, P2_P1_REIP_REG_1_, P2_P1_STATE_REG_0_,
P2_P1_FLUSH_REG, P2_P1_REIP_REG_0_, P2_P1_CODEFETCH_REG,
P2_P1_READREQUEST_REG, n14476, n14481, n14486, n14491, n14661, n14666,
n14821, n15481, n15486, n15491, n15496, n15501,
P2_P1_DATAWIDTH_REG_1_, n16651, n16661, n16666, n16676, n16686,
n16696, n16711, n16716, P2_P1_DATAWIDTH_REG_0_, P2_P1_REIP_REG_31_,
P2_P1_REIP_REG_30_, P2_P1_ADDRESS_REG_29_, P2_P1_REIP_REG_29_,
P2_P1_ADDRESS_REG_28_, P2_P1_REIP_REG_28_, P2_P1_ADDRESS_REG_27_,
P2_P1_REIP_REG_27_, P2_P1_ADDRESS_REG_26_, P2_P1_REIP_REG_26_,
P2_P1_ADDRESS_REG_25_, P2_P1_REIP_REG_25_, P2_P1_ADDRESS_REG_24_,
P2_P1_REIP_REG_24_, P2_P1_ADDRESS_REG_23_, P2_P1_REIP_REG_23_,
P2_P1_ADDRESS_REG_22_, P2_P1_REIP_REG_22_, P2_P1_ADDRESS_REG_21_,
P2_P1_REIP_REG_21_, P2_P1_ADDRESS_REG_20_, P2_P1_REIP_REG_20_,
P2_P1_ADDRESS_REG_19_, P2_P1_REIP_REG_19_, P2_P1_REIP_REG_18_,
P2_P1_REIP_REG_17_, P2_P1_REIP_REG_16_, P2_P1_REIP_REG_15_,
P2_P1_REIP_REG_14_, P2_P1_REIP_REG_13_, P2_P1_REIP_REG_11_,
P2_P1_REIP_REG_10_, P2_P1_REIP_REG_8_, P2_P1_REIP_REG_7_,
P2_P1_REIP_REG_5_, P2_P1_REIP_REG_4_, P2_P1_REIP_REG_3_,
P2_P1_REIP_REG_2_, P2_P1_INSTQUEUE_REG_0__0_,
P2_P1_INSTQUEUE_REG_1__0_, P2_P1_INSTQUEUE_REG_2__0_,
P2_P1_INSTQUEUE_REG_3__0_, P2_P1_INSTQUEUE_REG_4__0_,
P2_P1_INSTQUEUE_REG_5__0_, P2_P1_INSTQUEUE_REG_6__0_,
P2_P1_INSTQUEUE_REG_7__0_, P2_P1_INSTQUEUE_REG_8__0_,
P2_P1_INSTQUEUE_REG_9__0_, P2_P1_INSTQUEUE_REG_10__0_,
P2_P1_INSTQUEUE_REG_11__0_, P2_P1_INSTQUEUE_REG_12__0_,
P2_P1_INSTQUEUE_REG_13__0_, P2_P1_INSTQUEUE_REG_14__0_,
P2_P1_INSTQUEUE_REG_0__1_, P2_P1_INSTQUEUE_REG_1__1_,
P2_P1_INSTQUEUE_REG_2__1_, P2_P1_INSTQUEUE_REG_3__1_,
P2_P1_INSTQUEUE_REG_4__1_, P2_P1_INSTQUEUE_REG_5__1_,
P2_P1_INSTQUEUE_REG_6__1_, P2_P1_INSTQUEUE_REG_7__1_,
P2_P1_INSTQUEUE_REG_8__1_, P2_P1_INSTQUEUE_REG_9__1_,
P2_P1_INSTQUEUE_REG_10__1_, P2_P1_INSTQUEUE_REG_11__1_,
P2_P1_INSTQUEUE_REG_12__1_, P2_P1_INSTQUEUE_REG_13__1_,
P2_P1_INSTQUEUE_REG_14__1_, P2_P1_INSTQUEUE_REG_0__4_,
P2_P1_INSTQUEUE_REG_1__4_, P2_P1_INSTQUEUE_REG_2__4_,
P2_P1_INSTQUEUE_REG_3__4_, P2_P1_INSTQUEUE_REG_4__4_,
P2_P1_INSTQUEUE_REG_5__4_, P2_P1_INSTQUEUE_REG_6__4_,
P2_P1_INSTQUEUE_REG_7__4_, P2_P1_INSTQUEUE_REG_8__4_,
P2_P1_INSTQUEUE_REG_9__4_, P2_P1_INSTQUEUE_REG_10__4_,
P2_P1_INSTQUEUE_REG_11__4_, P2_P1_INSTQUEUE_REG_12__4_,
P2_P1_INSTQUEUE_REG_13__4_, P2_P1_INSTQUEUE_REG_14__4_,
P2_P1_INSTQUEUE_REG_0__2_, P2_P1_INSTQUEUE_REG_1__2_,
P2_P1_INSTQUEUE_REG_2__2_, P2_P1_INSTQUEUE_REG_3__2_,
P2_P1_INSTQUEUE_REG_4__2_, P2_P1_INSTQUEUE_REG_5__2_,
P2_P1_INSTQUEUE_REG_6__2_, P2_P1_INSTQUEUE_REG_7__2_,
P2_P1_INSTQUEUE_REG_8__2_, P2_P1_INSTQUEUE_REG_9__2_,
P2_P1_INSTQUEUE_REG_10__2_, P2_P1_INSTQUEUE_REG_11__2_,
P2_P1_INSTQUEUE_REG_12__2_, P2_P1_INSTQUEUE_REG_13__2_,
P2_P1_INSTQUEUE_REG_14__2_, P2_P1_INSTQUEUE_REG_0__3_,
P2_P1_INSTQUEUE_REG_1__3_, P2_P1_INSTQUEUE_REG_2__3_,
P2_P1_INSTQUEUE_REG_3__3_, P2_P1_INSTQUEUE_REG_4__3_,
P2_P1_INSTQUEUE_REG_5__3_, P2_P1_INSTQUEUE_REG_6__3_,
P2_P1_INSTQUEUE_REG_7__3_, P2_P1_INSTQUEUE_REG_8__3_,
P2_P1_INSTQUEUE_REG_9__3_, P2_P1_INSTQUEUE_REG_10__3_,
P2_P1_INSTQUEUE_REG_11__3_, P2_P1_INSTQUEUE_REG_12__3_,
P2_P1_INSTQUEUE_REG_13__3_, P2_P1_INSTQUEUE_REG_14__3_,
P2_P1_INSTQUEUE_REG_0__7_, P2_P1_INSTQUEUE_REG_1__7_,
P2_P1_INSTQUEUE_REG_2__7_, P2_P1_INSTQUEUE_REG_3__7_,
P2_P1_INSTQUEUE_REG_4__7_, P2_P1_INSTQUEUE_REG_5__7_,
P2_P1_INSTQUEUE_REG_6__7_, P2_P1_INSTQUEUE_REG_7__7_,
P2_P1_INSTQUEUE_REG_8__7_, P2_P1_INSTQUEUE_REG_9__7_,
P2_P1_INSTQUEUE_REG_10__7_, P2_P1_INSTQUEUE_REG_11__7_,
P2_P1_INSTQUEUE_REG_12__7_, P2_P1_INSTQUEUE_REG_13__7_,
P2_P1_INSTQUEUE_REG_14__7_, P2_P1_INSTQUEUE_REG_0__5_,
P2_P1_INSTQUEUE_REG_1__5_, P2_P1_INSTQUEUE_REG_2__5_,
P2_P1_INSTQUEUE_REG_3__5_, P2_P1_INSTQUEUE_REG_4__5_,
P2_P1_INSTQUEUE_REG_5__5_, P2_P1_INSTQUEUE_REG_6__5_,
P2_P1_INSTQUEUE_REG_7__5_, P2_P1_INSTQUEUE_REG_8__5_,
P2_P1_INSTQUEUE_REG_9__5_, P2_P1_INSTQUEUE_REG_10__5_,
P2_P1_INSTQUEUE_REG_11__5_, P2_P1_INSTQUEUE_REG_12__5_,
P2_P1_INSTQUEUE_REG_13__5_, P2_P1_INSTQUEUE_REG_14__5_,
P2_P1_INSTQUEUE_REG_0__6_, P2_P1_INSTQUEUE_REG_1__6_,
P2_P1_INSTQUEUE_REG_2__6_, P2_P1_INSTQUEUE_REG_3__6_,
P2_P1_INSTQUEUE_REG_4__6_, P2_P1_INSTQUEUE_REG_5__6_,
P2_P1_INSTQUEUE_REG_6__6_, P2_P1_INSTQUEUE_REG_7__6_,
P2_P1_INSTQUEUE_REG_8__6_, P2_P1_INSTQUEUE_REG_9__6_,
P2_P1_INSTQUEUE_REG_10__6_, P2_P1_INSTQUEUE_REG_11__6_,
P2_P1_INSTQUEUE_REG_12__6_, P2_P1_INSTQUEUE_REG_13__6_,
P2_P1_INSTQUEUE_REG_14__6_, P2_P1_MORE_REG,
P2_P1_PHYADDRPOINTER_REG_0_, P2_P1_PHYADDRPOINTER_REG_1_,
P2_P1_PHYADDRPOINTER_REG_2_, P2_P1_PHYADDRPOINTER_REG_3_,
P2_P1_PHYADDRPOINTER_REG_4_, P2_P1_PHYADDRPOINTER_REG_5_,
P2_P1_PHYADDRPOINTER_REG_6_, P2_P1_PHYADDRPOINTER_REG_7_,
P2_P1_PHYADDRPOINTER_REG_8_, P2_P1_PHYADDRPOINTER_REG_9_,
P2_P1_PHYADDRPOINTER_REG_10_, P2_P1_PHYADDRPOINTER_REG_11_,
P2_P1_PHYADDRPOINTER_REG_12_, P2_P1_PHYADDRPOINTER_REG_13_,
P2_P1_PHYADDRPOINTER_REG_14_, P2_P1_PHYADDRPOINTER_REG_15_,
P2_P1_PHYADDRPOINTER_REG_16_, P2_P1_PHYADDRPOINTER_REG_17_,
P2_P1_PHYADDRPOINTER_REG_18_, P2_P1_PHYADDRPOINTER_REG_19_,
P2_P1_PHYADDRPOINTER_REG_20_, P2_P1_PHYADDRPOINTER_REG_21_,
P2_P1_PHYADDRPOINTER_REG_22_, P2_P1_PHYADDRPOINTER_REG_23_,
P2_P1_PHYADDRPOINTER_REG_24_, P2_P1_PHYADDRPOINTER_REG_25_,
P2_P1_PHYADDRPOINTER_REG_26_, P2_P1_PHYADDRPOINTER_REG_27_,
P2_P1_PHYADDRPOINTER_REG_28_, P2_P1_PHYADDRPOINTER_REG_29_,
P2_P1_PHYADDRPOINTER_REG_30_, P2_P1_PHYADDRPOINTER_REG_31_,
P2_P1_LWORD_REG_15_, P2_P1_EAX_REG_14_, P2_P1_LWORD_REG_14_,
P2_P1_EAX_REG_13_, P2_P1_LWORD_REG_13_, P2_P1_LWORD_REG_12_,
P2_P1_EAX_REG_11_, P2_P1_LWORD_REG_11_, P2_P1_EAX_REG_10_,
P2_P1_LWORD_REG_10_, P2_P1_LWORD_REG_9_, P2_P1_EAX_REG_8_,
P2_P1_LWORD_REG_8_, P2_P1_EAX_REG_7_, P2_P1_LWORD_REG_7_,
P2_P1_LWORD_REG_6_, P2_P1_EAX_REG_5_, P2_P1_LWORD_REG_5_,
P2_P1_EAX_REG_4_, P2_P1_LWORD_REG_4_, P2_P1_LWORD_REG_3_,
P2_P1_EAX_REG_2_, P2_P1_LWORD_REG_2_, P2_P1_LWORD_REG_1_,
P2_P1_EAX_REG_0_, P2_P1_LWORD_REG_0_, P2_P1_EAX_REG_30_,
P2_P1_UWORD_REG_14_, P2_P1_EAX_REG_29_, P2_P1_UWORD_REG_13_,
P2_P1_EAX_REG_28_, P2_P1_UWORD_REG_12_, P2_P1_EAX_REG_27_,
P2_P1_UWORD_REG_11_, P2_P1_UWORD_REG_10_, P2_P1_EAX_REG_25_,
P2_P1_UWORD_REG_9_, P2_P1_EAX_REG_24_, P2_P1_UWORD_REG_8_,
P2_P1_UWORD_REG_7_, P2_P1_EAX_REG_22_, P2_P1_UWORD_REG_6_,
P2_P1_EAX_REG_21_, P2_P1_UWORD_REG_5_, P2_P1_UWORD_REG_4_,
P2_P1_EAX_REG_19_, P2_P1_UWORD_REG_3_, P2_P1_EAX_REG_18_,
P2_P1_UWORD_REG_2_, P2_P1_UWORD_REG_1_, P2_P1_EAX_REG_16_,
P2_P1_UWORD_REG_0_, P2_P1_EBX_REG_0_, P2_P1_EBX_REG_1_,
P2_P1_EBX_REG_2_, P2_P1_EBX_REG_3_, P2_P1_EBX_REG_4_,
P2_P1_EBX_REG_5_, P2_P1_EBX_REG_6_, P2_P1_EBX_REG_7_,
P2_P1_EBX_REG_8_, P2_P1_EBX_REG_9_, P2_P1_EBX_REG_10_,
P2_P1_EBX_REG_11_, P2_P1_EBX_REG_12_, P2_P1_EBX_REG_13_,
P2_P1_EBX_REG_14_, P2_P1_EBX_REG_15_, P2_P1_EBX_REG_16_,
P2_P1_EBX_REG_17_, P2_P1_EBX_REG_18_, P2_P1_EBX_REG_19_,
P2_P1_EBX_REG_20_, P2_P1_EBX_REG_21_, P2_P1_EBX_REG_22_,
P2_P1_EBX_REG_23_, P2_P1_EBX_REG_24_, P2_P1_EBX_REG_25_,
P2_P1_EBX_REG_26_, P2_P1_EBX_REG_27_, P2_P1_EBX_REG_28_,
P2_P1_EBX_REG_29_, P2_P1_EBX_REG_30_, P2_P1_BYTEENABLE_REG_3_,
P2_P1_BYTEENABLE_REG_2_, P2_P1_BYTEENABLE_REG_1_,
P2_P1_BYTEENABLE_REG_0_, P2_P1_MEMORYFETCH_REG, n1, n2, n3, n4, n6,
n7, n8, n9, n11, n12, n13, n14, n16, n17, n18, n19, n21, n22, n23,
n24, n26, n27, n28, n29, n31, n32, n33, n34, n36, n37, n38, n48, n50,
n52, n54, n56, n58, n60, n62, n64, n65, n67, n68, n70, n71, n73, n74,
n76, n77, n79, n80, n82, n83, n85, n88, n90, n92, n94, n96, n98, n100,
n102, n112, n114, n116, n118, n120, n123, n125, n128, n130, n133,
n135, n138, n140, n143, n145, n147, n148, n149, n150, n152, n153,
n154, n155, n157, n158, n162, n163, n164, n165, n167, n168, n169,
n170, n172, n173, n174, n175, n177, n178, n179, n180, n182, n184,
n185, n187, n188, n189, n190, n192, n193, n194, n195, n199, n200,
n202, n203, n204, n205, n207, n208, n209, n210, n212, n213, n214,
n215, n217, n218, n219, n220, n222, n223, n224, n225, n227, n228,
n229, n230, n232, n233, n234, n237, n238, n239, n240, n243, n245,
n247, n248, n249, n252, n253, n254, n255, n258, n259, n260, n262,
n264, n265, n267, n268, n270, n272, n273, n274, n277, n278, n279,
n280, n283, n284, n285, n287, n289, n290, n292, n304, n307, n309,
n312, n314, n317, n319, n322, n324, n325, n327, n329, n330, n333,
n335, n337, n339, n340, n342, n344, n347, n348, n350, n353, n355,
n358, n360, n363, n365, n368, n370, n383, n385, n388, n390, n393,
n395, n398, n400, n403, n405, n408, n410, n413, n415, n418, n419,
n420, n422, n423, n424, n425, n427, n428, n429, n430, n434, n435,
n437, n438, n439, n440, n442, n443, n444, n445, n446, n447, n448,
n449, n450, n452, n453, n455, n457, n458, n459, n460, n462, n463,
n464, n465, n467, n470, n472, n473, n474, n475, n477, n478, n479,
n480, n482, n483, n484, n485, n487, n489, n490, n492, n493, n494,
n495, n497, n498, n499, n500, n502, n503, n504, n505, n508, n509,
n510, n512, n514, n515, n517, n518, n519, n520, n522, n523, n524,
n527, n528, n529, n530, n532, n533, n534, n535, n537, n538, n539,
n540, n542, n543, n544, n545, n547, n548, n549, n550, n552, n553,
n555, n559, n563, n564, n565, n568, n569, n570, n573, n574, n575,
n577, n578, n579, n583, n584, n585, n587, n588, n589, n590, n592,
n593, n594, n595, n597, n598, n599, n600, n602, n603, n604, n607,
n608, n609, n610, n612, n613, n615, n617, n618, n619, n620, n622,
n623, n624, n625, n627, n628, n629, n630, n632, n633, n634, n635,
n637, n638, n639, n640, n642, n643, n644, n645, n647, n648, n649,
n650, n652, n653, n654, n655, n657, n659, n660, n662, n664, n665,
n667, n668, n669, n670, n672, n673, n674, n675, n677, n678, n679,
n680, n682, n683, n684, n685, n687, n688, n689, n690, n692, n693,
n694, n695, n697, n698, n699, n700, n702, n703, n704, n707, n708,
n709, n710, n712, n713, n714, n715, n717, n718, n719, n720, n722,
n723, n724, n725, n727, n728, n729, n730, n732, n733, n734, n735,
n737, n738, n739, n740, n742, n743, n744, n745, n747, n748, n749,
n750, n752, n753, n754, n757, n758, n759, n760, n762, n763, n764,
n765, n767, n768, n769, n770, n772, n773, n774, n775, n777, n778,
n779, n780, n782, n783, n784, n785, n786, n787, n788, n789, n790,
n792, n793, n794, n795, n797, n798, n799, n800, n802, n803, n804,
n805, n807, n810, n812, n813, n814, n815, n817, n818, n819, n820,
n822, n823, n824, n825, n827, n829, n830, n832, n833, n834, n835,
n837, n838, n839, n840, n842, n843, n844, n845, n847, n848, n849,
n850, n852, n853, n854, n855, n857, n858, n859, n860, n862, n863,
n864, n865, n867, n868, n869, n870, n872, n873, n874, n875, n877,
n878, n879, n880, n882, n883, n884, n885, n887, n888, n889, n890,
n892, n893, n894, n895, n897, n898, n899, n900, n902, n903, n904,
n905, n907, n908, n909, n910, n912, n913, n914, n915, n917, n933,
n934, n1018, n1019, n1022, n1024, n1027, n1028, n1030, n1032, n1033,
n1034, n1037, n1038, n1039, n1040, n1043, n1044, n1047, n1048, n1052,
n1053, n1054, n1057, n1059, n1060, n1062, n1063, n1064, n1065, n1067,
n1068, n1069, n1072, n1073, n1074, n1075, n1077, n1078, n1079, n1082,
n1083, n1084, n1085, n1087, n1088, n1089, n1090, n1092, n1093, n1095,
n1097, n1098, n1099, n1100, n1102, n1103, n1104, n1107, n1108, n1109,
n1110, n1112, n1113, n1114, n1115, n1117, n1118, n1119, n1120, n1122,
n1124, n1125, n1127, n1128, n1129, n1130, n1132, n1133, n1134, n1135,
n1137, n1140, n1142, n1143, n1144, n1145, n1147, n1148, n1149, n1150,
n1152, n1153, n1154, n1155, n1157, n1158, n1159, n1160, n1162, n1163,
n1165, n1167, n1168, n1169, n1170, n1173, n1174, n1175, n1177, n1179,
n1180, n1182, n1183, n1184, n1185, n1187, n1188, n1189, n1190, n1192,
n1193, n1194, n1195, n1197, n1198, n1199, n1200, n1202, n1203, n1204,
n1205, n1207, n1208, n1209, n1210, n1212, n1213, n1214, n1215, n1217,
n1218, n1220, n1222, n1223, n1224, n1225, n1227, n1228, n1229, n1230,
n1232, n1233, n1234, n1235, n1237, n1238, n1239, n1240, n1242, n1243,
n1244, n1245, n1247, n1248, n1249, n1250, n1252, n1253, n1254, n1255,
n1257, n1258, n1259, n1260, n1262, n1263, n1264, n1265, n1267, n1268,
n1269, n1270, n1272, n1273, n1274, n1277, n1278, n1279, n1280, n1282,
n1283, n1284, n1285, n1287, n1288, n1289, n1290, n1292, n1293, n1294,
n1295, n1297, n1298, n1299, n1300, n1302, n1303, n1304, n1305, n1307,
n1308, n1309, n1310, n1312, n1313, n1314, n1315, n1319, n1320, n1322,
n1324, n1325, n1327, n1328, n1329, n1330, n1332, n1333, n1334, n1335,
n1337, n1338, n1339, n1340, n1342, n1343, n1344, n1345, n1347, n1348,
n1349, n1350, n1352, n1353, n1354, n1355, n1357, n1358, n1360, n1362,
n1363, n1364, n1365, n1367, n1368, n1369, n1370, n1372, n1373, n1374,
n1375, n1377, n1378, n1379, n1380, n1382, n1383, n1384, n1385, n1387,
n1388, n1389, n1390, n1392, n1393, n1395, n1397, n1398, n1399, n1400,
n1402, n1403, n1404, n1405, n1407, n1408, n1409, n1410, n1412, n1413,
n1414, n1415, n1417, n1418, n1419, n1420, n1422, n1423, n1424, n1425,
n1428, n1429, n1430, n1432, n1433, n1434, n1435, n1437, n1438, n1439,
n1440, n1442, n1443, n1444, n1445, n1447, n1448, n1449, n1452, n1454,
n1455, n1457, n1458, n1459, n1460, n1462, n1463, n1464, n1465, n1467,
n1468, n1469, n1470, n1472, n1473, n1474, n1475, n1477, n1478, n1479,
n1482, n1484, n1485, n1487, n1488, n1489, n1490, n1492, n1493, n1494,
n1495, n1497, n1498, n1499, n1500, n1502, n1504, n1505, n1507, n1508,
n1509, n1510, n1512, n1513, n1514, n1515, n1517, n1518, n1519, n1520,
n1522, n1523, n1524, n1525, n1527, n1528, n1530, n1532, n1533, n1534,
n1535, n1537, n1538, n1539, n1540, n1542, n1543, n1544, n1547, n1548,
n1549, n1550, n1552, n1555, n1557, n1559, n1560, n1562, n1563, n1564,
n1565, n1567, n1568, n1569, n1570, n1572, n1573, n1575, n1577, n1578,
n1579, n1580, n1583, n1584, n1585, n1587, n1588, n1589, n1590, n1592,
n1594, n1595, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
n1607, n1608, n1609, n1610, n1613, n1614, n1615, n1618, n1619, n1620,
n1622, n1623, n1624, n1625, n1627, n1628, n1629, n1630, n1632, n1633,
n1634, n1635, n1637, n1639, n1640, n1642, n1643, n1644, n1645, n1647,
n1648, n1649, n1650, n1652, n1654, n1655, n1657, n1658, n1659, n1660,
n1662, n1663, n1664, n1665, n1667, n1668, n1669, n1670, n1673, n1674,
n1675, n1677, n1678, n1679, n1680, n1682, n1683, n1684, n1687, n1688,
n1689, n1690, n1693, n1694, n1695, n1697, n1698, n1699, n1700, n1703,
n1704, n1705, n1707, n1708, n1709, n1710, n1712, n1714, n1715, n1717,
n1718, n1719, n1720, n1722, n1724, n1725, n1727, n1728, n1729, n1730,
n1732, n1734, n1735, n1737, n1738, n1739, n1740, n1742, n1743, n1745,
n1747, n1748, n1749, n1750, n1752, n1754, n1755, n1757, n1758, n1760,
n1762, n1764, n1767, n1769, n1773, n1774, n1775, n1777, n1778, n1779,
n1780, n1782, n1783, n1784, n1785, n1787, n1788, n1790, n1792, n1793,
n1794, n1795, n1797, n1798, n1799, n1800, n1802, n1812, n1813, n1834,
n1838, n1843, n1844, n1845, n1847, n1848, n1849, n1850, n1852, n1853,
n1854, n1855, n1858, n1860, n1862, n1863, n1864, n1865, n1867, n1868,
n1869, n1870, n1872, n1873, n1874, n1875, n1877, n1878, n1879, n1880,
n1882, n1883, n1884, n1885, n1887, n1888, n1889, n1890, n1892, n1893,
n1894, n1900, n1902, n1903, n1904, n1905, n1907, n1908, n1909, n1910,
n1912, n1913, n1914, n1915, n1917, n1918, n1919, n1920, n1922, n1923,
n1924, n1925, n1927, n1928, n1929, n1930, n1932, n1933, n1934, n1935,
n1937, n1938, n1939, n1940, n1942, n1943, n1944, n1945, n1947, n1948,
n1949, n1950, n1952, n1953, n1954, n1955, n1957, n1958, n1959, n1960,
n1962, n1963, n1964, n1965, n1967, n1968, n1969, n1970, n1972, n1973,
n1974, n1975, n1977, n1978, n1979, n1980, n1982, n1983, n1984, n1985,
n1987, n1988, n1989, n1990, n1992, n1993, n1994, n1995, n1997, n2000,
n2002, n2003, n2004, n2005, n2007, n2008, n2009, n2010, n2011, n2012,
n2013, n2014, n2015, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
n2024, n2025, n2027, n2028, n2029, n2030, n2032, n2033, n2034, n2035,
n2037, n2038, n2039, n2040, n2042, n2043, n2044, n2045, n2047, n2048,
n2049, n2050, n2052, n2053, n2054, n2055, n2057, n2058, n2059, n2060,
n2062, n2064, n2065, n2067, n2068, n2069, n2070, n2072, n2073, n2074,
n2075, n2077, n2078, n2079, n2080, n2082, n2083, n2084, n2087, n2088,
n2090, n2092, n2093, n2094, n2095, n2097, n2098, n2100, n2102, n2103,
n2104, n2105, n2107, n2108, n2109, n2110, n2112, n2113, n2114, n2115,
n2117, n2118, n2119, n2120, n2122, n2123, n2124, n2125, n2127, n2128,
n2129, n2130, n2132, n2133, n2134, n2135, n2137, n2138, n2139, n2140,
n2142, n2143, n2144, n2145, n2147, n2148, n2149, n2150, n2152, n2153,
n2154, n2155, n2157, n2158, n2159, n2160, n2162, n2163, n2164, n2165,
n2167, n2168, n2169, n2170, n2172, n2173, n2174, n2175, n2177, n2178,
n2179, n2180, n2182, n2183, n2184, n2185, n2187, n2188, n2189, n2190,
n2192, n2193, n2194, n2195, n2197, n2198, n2199, n2200, n2202, n2203,
n2204, n2205, n2207, n2208, n2209, n2212, n2250, n2353, n2354, n2355,
n2357, n2358, n2359, n2360, n2362, n2363, n2364, n2365, n2367, n2368,
n2369, n2370, n2372, n2373, n2374, n2375, n2377, n2378, n2379, n2380,
n2382, n2383, n2384, n2385, n2387, n2388, n2389, n2392, n2393, n2394,
n2395, n2397, n2398, n2399, n2400, n2402, n2403, n2404, n2405, n2407,
n2408, n2409, n2410, n2412, n2413, n2414, n2415, n2417, n2418, n2419,
n2420, n2422, n2423, n2424, n2425, n2427, n2428, n2429, n2430, n2432,
n2433, n2437, n2438, n2439, n2442, n2443, n2444, n2445, n2447, n2448,
n2449, n2450, n2452, n2453, n2454, n2455, n2457, n2458, n2459, n2460,
n2462, n2463, n2464, n2465, n2467, n2468, n2469, n2470, n2472, n2473,
n2474, n2475, n2478, n2479, n2480, n2482, n2483, n2484, n2485, n2487,
n2488, n2489, n2490, n2492, n2493, n2494, n2495, n2497, n2498, n2499,
n2500, n2502, n2503, n2504, n2505, n2507, n2508, n2509, n2510, n2512,
n2514, n2515, n2517, n2518, n2519, n2520, n2522, n2523, n2524, n2525,
n2527, n2528, n2529, n2530, n2532, n2533, n2534, n2535, n2537, n2538,
n2539, n2540, n2542, n2543, n2544, n2545, n2547, n2549, n2550, n2552,
n2553, n2554, n2555, n2557, n2558, n2559, n2560, n2562, n2563, n2564,
n2565, n2567, n2568, n2569, n2570, n2572, n2574, n2575, n2577, n2578,
n2579, n2580, n2582, n2583, n2584, n2585, n2587, n2588, n2589, n2590,
n2592, n2593, n2594, n2595, n2597, n2598, n2599, n2600, n2602, n2603,
n2605, n2607, n2608, n2609, n2610, n2612, n2613, n2614, n2615, n2617,
n2618, n2619, n2620, n2622, n2623, n2624, n2625, n2628, n2629, n2630,
n2632, n2633, n2634, n2635, n2637, n2638, n2639, n2640, n2642, n2643,
n2644, n2645, n2647, n2648, n2649, n2652, n2653, n2654, n2655, n2657,
n2658, n2659, n2660, n2662, n2663, n2664, n2665, n2667, n2668, n2669,
n2670, n2672, n2673, n2675, n2677, n2678, n2679, n2680, n2682, n2683,
n2684, n2685, n2687, n2688, n2689, n2690, n2692, n2693, n2694, n2697,
n2698, n2699, n2700, n2702, n2703, n2704, n2705, n2707, n2708, n2709,
n2712, n2713, n2714, n2715, n2717, n2718, n2719, n2720, n2722, n2723,
n2724, n2725, n2728, n2729, n2730, n2732, n2733, n2734, n2735, n2738,
n2740, n2742, n2743, n2744, n2745, n2747, n2748, n2749, n2750, n2752,
n2753, n2754, n2755, n2757, n2758, n2759, n2760, n2763, n2764, n2765,
n2767, n2768, n2769, n2770, n2772, n2773, n2774, n2775, n2778, n2779,
n2780, n2782, n2783, n2784, n2785, n2787, n2788, n2789, n2790, n2793,
n2794, n2795, n2797, n2798, n2799, n2800, n2802, n2803, n2805, n2807,
n2808, n2809, n2812, n2813, n2814, n2815, n2817, n2818, n2820, n2822,
n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2832, n2833, n2834,
n2835, n2837, n2838, n2839, n2840, n2842, n2844, n2845, n2847, n2848,
n2849, n2850, n2853, n2854, n2855, n2857, n2858, n2859, n2860, n2863,
n2864, n2865, n2867, n2868, n2870, n2872, n2873, n2874, n2877, n2878,
n2882, n2884, n2889, n2890, n2892, n2893, n2894, n2895, n2897, n2898,
n2899, n2900, n2902, n2903, n2904, n2905, n2908, n2909, n2910, n2912,
n2913, n2914, n2915, n2917, n2918, n2919, n2929, n2930, n2978, n2979,
n2980, n2988, n2989, n3028, n3029, n3030, n3032, n3033, n3034, n3035,
n3037, n3038, n3039, n3040, n3042, n3044, n3045, n3048, n3052, n3053,
n3054, n3055, n3057, n3058, n3059, n3060, n3062, n3063, n3064, n3065,
n3067, n3068, n3069, n3072, n3073, n3075, n3077, n3078, n3083, n3084,
n3085, n3087, n3088, n3090, n3094, n3095, n3097, n3098, n3099, n3100,
n3102, n3103, n3104, n3105, n3107, n3108, n3109, n3110, n3112, n3113,
n3114, n3115, n3117, n3118, n3119, n3120, n3122, n3123, n3124, n3125,
n3127, n3128, n3129, n3130, n3132, n3133, n3134, n3135, n3137, n3138,
n3139, n3140, n3142, n3143, n3144, n3145, n3147, n3148, n3149, n3150,
n3152, n3153, n3155, n3158, n3159, n3160, n3162, n3163, n3165, n3167,
n3168, n3169, n3170, n3172, n3173, n3174, n3175, n3177, n3178, n3179,
n3180, n3183, n3184, n3185, n3187, n3188, n3189, n3192, n3193, n3195,
n3197, n3198, n3199, n3200, n3203, n3204, n3205, n3207, n3208, n3209,
n3210, n3212, n3213, n3215, n3217, n3218, n3219, n3220, n3222, n3223,
n3224, n3225, n3227, n3229, n3230, n3232, n3233, n3234, n3235, n3236,
n3237, n3238, n3239, n3242, n3243, n3244, n3245, n3246, n3384, n3387,
n3389, n3390, n3392, n3393, n3394, n3395, n3397, n3399, n3400, n3403,
n3404, n3405, n3407, n3408, n3409, n3410, n3412, n3413, n3414, n3418,
n3420, n3422, n3423, n3424, n3425, n3427, n3428, n3429, n3430, n3432,
n3433, n3434, n3435, n3437, n3438, n3439, n3440, n3442, n3443, n3444,
n3445, n3447, n3449, n3450, n3453, n3454, n3455, n3457, n3458, n3460,
n3463, n3464, n3465, n3467, n3468, n3469, n3470, n3473, n3474, n3475,
n3487, n3497, n3503, n3509, n3514, n3522, n3523, n3524, n3525, n3527,
n3528, n3529, n3530, n3532, n3533, n3534, n3535, n3537, n3538, n3540,
n3542, n3543, n3544, n3545, n3547, n3548, n3549, n3550, n3553, n3557,
n3558, n3559, n3560, n3562, n3563, n3565, n3567, n3568, n3569, n3570,
n3572, n3632, n3634, n3635, n3637, n3638, n3639, n3640, n3674, n3675,
n3677, n3678, n3679, n3680, n3682, n3683, n3684, n3685, n3687, n3688,
n3689, n3690, n3692, n3693, n3694, n3695, n3697, n3698, n3699, n3700,
n3702, n3703, n3704, n3744, n3745, n3747, n3749, n3794, n3797, n3822,
n3823, n3832, n3833, n3872, n3873, n3874, n3875, n3877, n3878, n3879,
n3880, n3882, n3883, n3884, n3885, n3888, n3889, n3892, n3895, n3897,
n3898, n3899, n3900, n3902, n3903, n3904, n3905, n3907, n3908, n3909,
n3910, n3912, n3913, n3915, n3917, n3919, n3920, n3922, n3927, n3928,
n3929, n3930, n3932, n3934, n3938, n3939, n3940, n3942, n3943, n3944,
n3945, n3947, n3948, n3949, n3950, n3952, n3953, n3954, n3955, n3957,
n3958, n3959, n3960, n3962, n3963, n3964, n3965, n3967, n3968, n3969,
n3970, n3972, n3973, n3974, n3975, n3977, n3978, n3979, n3980, n3982,
n3983, n3984, n3985, n3987, n3989, n3990, n3992, n3993, n3994, n3995,
n3997, n3999, n4000, n4002, n4003, n4005, n4007, n4008, n4009, n4010,
n4012, n4013, n4014, n4015, n4017, n4018, n4020, n4022, n4023, n4024,
n4027, n4028, n4030, n4032, n4033, n4035, n4037, n4038, n4039, n4040,
n4042, n4043, n4045, n4047, n4048, n4049, n4050, n4052, n4053, n4054,
n4057, n4058, n4059, n4060, n4062, n4063, n4064, n4067, n4068, n4069,
n4222, n4224, n4227, n4228, n4229, n4230, n4232, n4233, n4234, n4237,
n4238, n4240, n4242, n4243, n4244, n4245, n4247, n4248, n4249, n4250,
n4252, n4255, n4258, n4259, n4260, n4262, n4263, n4264, n4265, n4267,
n4268, n4269, n4270, n4272, n4273, n4274, n4275, n4277, n4278, n4279,
n4280, n4282, n4283, n4284, n4287, n4288, n4290, n4292, n4293, n4294,
n4295, n4298, n4300, n4302, n4303, n4304, n4305, n4307, n4308, n4310,
n4312, n4313, n4324, n4334, n4340, n4347, n4352, n4359, n4360, n4362,
n4363, n4364, n4365, n4367, n4368, n4369, n4370, n4372, n4373, n4374,
n4375, n4378, n4379, n4380, n4382, n4383, n4384, n4385, n4387, n4388,
n4390, n4394, n4395, n4397, n4398, n4399, n4400, n4403, n4404, n4405,
n4407, n4408, n4409, n4522, n4523, n4524, n4525, n4527, n4528, n4568,
n4569, n4570, n4572, n4573, n4574, n4575, n4577, n4578, n4579, n4580,
n4582, n4583, n4584, n4585, n4587, n4588, n4589, n4590, n4592, n4593,
n4594, n4595, n4597, n4598, n4638, n4639, n4640, n4643, n4687, n4711,
n4712, n4719, n4720, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
n4758, n4759, n4760, n4762, n4763, n4764, n4765, n4767, n4768, n4769,
n4770, n4772, n4773, n4774, n4777, n4778, n4780, n4782, n4784, n4785,
n4787, n4788, n4789, n4790, n4792, n4793, n4794, n4795, n4797, n4798,
n4799, n4800, n4802, n4803, n4804, n4805, n4807, n4808, n4809, n4810,
n4812, n4813, n4814, n4815, n4818, n4819, n4820, n4825, n4827, n4828,
n4829, n4832, n4833, n4834, n4835, n4838, n4839, n4842, n4843, n4844,
n4845, n4847, n4848, n4849, n4850, n4852, n4853, n4854, n4855, n4857,
n4858, n4859, n4860, n4862, n4863, n4864, n4865, n4867, n4868, n4869,
n4870, n4872, n4873, n4874, n4875, n4877, n4878, n4879, n4880, n4881,
n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
n4892, n4893, n4895, n4896, n4898, n4899, n4900, n4902, n4903, n4904,
n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
n4915, n4916, n4918, n4919, n4920, n4921, n4922, n4923, n4925, n4926,
n4928, n4929, n4930, n4932, n4933, n4935, n4937, n4938, n4939, n4940,
n4942, n4943, n4944, n4945, n4948, n4949, n4950, n4952, n4953, n4954,
n4955, n4957, n4958, n4959, n4962, n4963, n4964, n4965, n4967, n4968,
n4969, n4970, n4972, n4973, n4975, n4977, n4978, n4979, n4980, n5132,
n5134, n5137, n5138, n5139, n5140, n5142, n5143, n5144, n5147, n5148,
n5150, n5152, n5153, n5154, n5155, n5157, n5158, n5159, n5160, n5162,
n5165, n5168, n5169, n5170, n5172, n5173, n5174, n5175, n5177, n5178,
n5179, n5180, n5182, n5183, n5184, n5185, n5187, n5188, n5189, n5190,
n5192, n5193, n5194, n5195, n5197, n5198, n5200, n5202, n5204, n5205,
n5207, n5208, n5209, n5210, n5214, n5215, n5217, n5218, n5219, n5220,
n5223, n5224, n5225, n5237, n5247, n5253, n5269, n5270, n5272, n5273,
n5274, n5275, n5277, n5278, n5279, n5280, n5282, n5283, n5284, n5285,
n5288, n5289, n5290, n5292, n5293, n5294, n5295, n5297, n5298, n5299,
n5300, n5302, n5303, n5304, n5305, n5307, n5308, n5309, n5310, n5312,
n5314, n5315, n5317, n5318, n5319, n5320, n5434, n5435, n5437, n5438,
n5439, n5440, n5442, n5443, n5444, n5445, n5447, n5448, n5449, n5450,
n5452, n5453, n5454, n5455, n5457, n5458, n5459, n5460, n5462, n5463,
n5464, n5465, n5507, n5508, n5509, n5510, n5579, n5580, n5582, n5589,
n5590, n5629, n5630, n5632, n5633, n5634, n5635, n5637, n5638, n5639,
n5640, n5642, n5643, n5645, n5647, n5649, n5653, n5654, n5655, n5657,
n5658, n5659, n5660, n5662, n5663, n5664, n5665, n5667, n5668, n5669,
n5670, n5673, n5674, n5677, n5678, n5679, n5684, n5685, n5687, n5688,
n5689, n5692, n5695, n5697, n5698, n5699, n5700, n5702, n5703, n5704,
n5705, n5707, n5708, n5709, n5710, n5712, n5713, n5714, n5715, n5717,
n5718, n5719, n5720, n5722, n5723, n5724, n5725, n5727, n5728, n5729,
n5730, n5732, n5733, n5734, n5735, n5737, n5738, n5739, n5740, n5742,
n5743, n5744, n5747, n5748, n5749, n5750, n5752, n5753, n5754, n5757,
n5758, n5759, n5760, n5762, n5764, n5765, n5767, n5768, n5769, n5770,
n5772, n5773, n5774, n5775, n5777, n5778, n5779, n5782, n5783, n5784,
n5785, n5787, n5788, n5790, n5792, n5794, n5795, n5797, n5798, n5799,
n5802, n5803, n5804, n5805, n5807, n5808, n5809, n5810, n5812, n5814,
n5815, n5817, n5818, n5819, n5820, n5822, n5823, n5824, n5825, n5828,
n5829, n5830, n5832, n5833, n5834, n5835, n5837, n5838, n5839, n5842,
n5843, n5844, n5845, n5847, n5999, n6002, n6004, n6005, n6007, n6008,
n6009, n6010, n6012, n6014, n6015, n6018, n6019, n6020, n6022, n6023,
n6024, n6025, n6027, n6028, n6029, n6033, n6035, n6037, n6038, n6039,
n6040, n6042, n6043, n6044, n6045, n6047, n6048, n6049, n6050, n6052,
n6053, n6054, n6055, n6057, n6058, n6059, n6060, n6062, n6064, n6065,
n6068, n6069, n6070, n6072, n6073, n6075, n6078, n6079, n6080, n6082,
n6083, n6084, n6085, n6088, n6089, n6090, n6102, n6112, n6118, n6124,
n6129, n6137, n6138, n6139, n6140, n6142, n6143, n6144, n6145, n6147,
n6148, n6149, n6150, n6152, n6153, n6155, n6157, n6158, n6159, n6160,
n6162, n6163, n6164, n6165, n6168, n6172, n6173, n6174, n6175, n6177,
n6178, n6180, n6182, n6183, n6184, n6185, n6187, n6259, n6262, n6263,
n6264, n6265, n6267, n6268, n6308, n6309, n6310, n6312, n6313, n6314,
n6315, n6317, n6318, n6319, n6320, n6322, n6323, n6324, n6325, n6327,
n6328, n6329, n6330, n6332, n6333, n6334, n6335, n6337, n6338, n6378,
n6379, n6380, n6383, n6429, n6454, n6455, n6464, n6465, n6504, n6505,
n6507, n6508, n6509, n6510, n6512, n6513, n6514, n6515, n6517, n6518,
n6520, n6522, n6524, n6528, n6529, n6530, n6532, n6533, n6534, n6535,
n6537, n6538, n6539, n6540, n6542, n6543, n6544, n6545, n6548, n6549,
n6552, n6553, n6554, n6559, n6560, n6562, n6563, n6564, n6567, n6570,
n6572, n6573, n6574, n6575, n6577, n6578, n6579, n6580, n6582, n6583,
n6584, n6585, n6587, n6588, n6589, n6590, n6592, n6593, n6594, n6595,
n6597, n6598, n6599, n6600, n6602, n6603, n6604, n6605, n6607, n6608,
n6609, n6610, n6612, n6613, n6614, n6615, n6617, n6618, n6619, n6622,
n6623, n6624, n6625, n6627, n6628, n6629, n6632, n6633, n6634, n6635,
n6638, n6639, n6640, n6642, n6643, n6644, n6645, n6647, n6648, n6649,
n6650, n6653, n6654, n6655, n6657, n6659, n6660, n6663, n6664, n6665,
n6668, n6669, n6670, n6672, n6673, n6674, n6675, n6678, n6679, n6680,
n6682, n6683, n6684, n6685, n6687, n6689, n6690, n6692, n6693, n6694,
n6695, n6697, n6699, n6700, n6702, n6854, n6857, n6859, n6860, n6862,
n6863, n6864, n6865, n6867, n6869, n6870, n6873, n6874, n6875, n6877,
n6878, n6879, n6880, n6882, n6883, n6884, n6888, n6890, n6892, n6893,
n6894, n6895, n6897, n6898, n6899, n6900, n6902, n6903, n6904, n6905,
n6907, n6908, n6909, n6910, n6912, n6913, n6914, n6915, n6917, n6919,
n6920, n6923, n6924, n6925, n6927, n6928, n6930, n6933, n6934, n6935,
n6937, n6938, n6939, n6940, n6943, n6944, n6945, n6957, n6967, n6973,
n6979, n6984, n6992, n6993, n6994, n6995, n6997, n6998, n6999, n7000,
n7002, n7003, n7004, n7005, n7007, n7008, n7010, n7012, n7013, n7014,
n7015, n7017, n7018, n7019, n7020, n7023, n7027, n7028, n7029, n7030,
n7032, n7033, n7035, n7037, n7038, n7039, n7040, n7042, n7154, n7155,
n7157, n7158, n7159, n7160, n7200, n7202, n7203, n7204, n7205, n7207,
n7208, n7209, n7210, n7212, n7213, n7214, n7215, n7217, n7218, n7219,
n7220, n7222, n7223, n7224, n7225, n7227, n7228, n7229, n7230, n7270,
n7272, n7273, n7275, n7319, n7343, n7344, n7353, n7354, n7393, n7394,
n7395, n7397, n7398, n7399, n7400, n7402, n7403, n7404, n7405, n7407,
n7408, n7409, n7410, n7412, n7413, n7414, n7415, n7417, n7418, n7420,
n7422, n7424, n7428, n7429, n7430, n7432, n7433, n7434, n7435, n7437,
n7438, n7439, n7440, n7442, n7443, n7444, n7445, n7447, n7448, n7449,
n7450, n7452, n7453, n7454, n7455, n7457, n7458, n7459, n7462, n7463,
n7464, n7469, n7470, n7472, n7473, n7474, n7477, n7480, n7482, n7483,
n7484, n7485, n7487, n7488, n7489, n7490, n7492, n7493, n7494, n7495,
n7497, n7498, n7499, n7500, n7502, n7503, n7504, n7505, n7507, n7508,
n7509, n7510, n7512, n7513, n7514, n7515, n7517, n7518, n7519, n7520,
n7522, n7523, n7524, n7525, n7527, n7528, n7529, n7530, n7533, n7534,
n7535, n7537, n7538, n7539, n7540, n7543, n7544, n7545, n7547, n7548,
n7550, n7552, n7553, n7554, n7555, n7557, n7558, n7559, n7560, n7562,
n7563, n7564, n7565, n7567, n7569, n7570, n7572, n7573, n7574, n7575,
n7578, n7579, n7582, n7583, n7584, n7585, n7587, n7589, n7590, n7592,
n7593, n7594, n7595, n7597, n7598, n7599, n7602, n7603, n7604, n7605,
n7607, n7608, n7609, n7610, n7612, n7613, n7615, n7617, n7618, n7619,
n7620, n7622, n7623, n7624, n7625, n7627, n7629, n7630, n7632, n7633,
n7634, n7787, n7789, n7792, n7793, n7794, n7795, n7797, n7798, n7799,
n7802, n7803, n7805, n7807, n7808, n7809, n7810, n7812, n7813, n7814,
n7815, n7817, n7820, n7823, n7824, n7825, n7827, n7828, n7829, n7830,
n7832, n7833, n7834, n7835, n7837, n7838, n7839, n7840, n7842, n7843,
n7844, n7845, n7847, n7848, n7849, n7850, n7852, n7853, n7855, n7857,
n7859, n7860, n7862, n7863, n7865, n7868, n7869, n7870, n7872, n7873,
n7874, n7877, n7878, n7879, n7890, n7900, n7907, n7917, n7924, n7925,
n7927, n7928, n7929, n7930, n7932, n7933, n7934, n7935, n7937, n7938,
n7939, n7940, n7943, n7944, n7945, n7947, n7948, n7949, n7950, n7952,
n7953, n7954, n7955, n7957, n7958, n7959, n7960, n7962, n7963, n7964,
n7965, n7967, n7969, n7970, n7972, n7973, n7974, n7975, n8089, n8090,
n8092, n8093, n8094, n8095, n8097, n8098, n8099, n8100, n8102, n8103,
n8104, n8105, n8107, n8108, n8109, n8110, n8112, n8113, n8114, n8115,
n8117, n8118, n8119, n8160, n8162, n8163, n8164, n8208, n8209, n8210,
n8212, n8213, n8214, n8215, n8217, n8218, n8219, n8220, n8222, n8224,
n8225, n8227, n8229, n8230, n8232, n8233, n8234, n8235, n8237, n8238,
n8239, n8240, n8243, n8244, n8245, n8247, n8248, n8249, n8250, n8252,
n8253, n8254, n8255, n8257, n8258, n8259, n8260, n8262, n8263, n8264,
n8265, n8267, n8268, n8269, n8270, n8272, n8273, n8275, n8277, n8278,
n8279, n8280, n8282, n8283, n8284, n8285, n8287, n8288, n8289, n8290,
n8292, n8293, n8294, n8295, n8297, n8298, n8299, n8300, n8302, n8303,
n8304, n8305, n8307, n8309, n8310, n8312, n8313, n8314, n8315, n8317,
n8318, n8319, n8320, n8322, n8323, n8324, n8325, n8327, n8328, n8329,
n8330, n8332, n8333, n8334, n8335, n8337, n8338, n8339, n8340, n8342,
n8343, n8344, n8345, n8347, n8348, n8349, n8350, n8352, n8353, n8354,
n8355, n8357, n8358, n8359, n8360, n8362, n8363, n8364, n8365, n8367,
n8368, n8369, n8370, n8372, n8373, n8374, n8375, n8377, n8378, n8379,
n8380, n8382, n8383, n8384, n8385, n8387, n8388, n8389, n8392, n8393,
n8394, n8395, n8397, n8398, n8399, n8400, n8402, n8403, n8404, n8405,
n8407, n8408, n8409, n8410, n8412, n8413, n8414, n8415, n8417, n8418,
n8419, n8420, n8422, n8423, n8424, n8425, n8427, n8428, n8429, n8430,
n8432, n8433, n8434, n8435, n8437, n8438, n8439, n8440, n8442, n8443,
n8444, n8445, n8448, n8449, n8450, n8452, n8453, n8454, n8455, n8457,
n8458, n8459, n8460, n8462, n8463, n8464, n8465, n8467, n8468, n8469,
n8470, n8472, n8473, n8474, n8475, n8477, n8478, n8479, n8480, n8482,
n8483, n8484, n8485, n8487, n8488, n8489, n8490, n8492, n8493, n8494,
n8495, n8497, n8498, n8499, n8500, n8502, n8503, n8504, n8505, n8507,
n8508, n8509, n8510, n8512, n8513, n8514, n8515, n8517, n8518, n8519,
n8520, n8522, n8523, n8524, n8525, n8527, n8528, n8529, n8530, n8532,
n8533, n8534, n8535, n8537, n8538, n8539, n8540, n8542, n8543, n8544,
n8545, n8547, n8548, n8549, n8550, n8552, n8553, n8554, n8555, n8557,
n8558, n8559, n8560, n8562, n8563, n8564, n8565, n8567, n8568, n8569,
n8570, n8572, n8573, n8574, n8575, n8577, n8578, n8579, n8580, n8582,
n8583, n8584, n8585, n8587, n8588, n8589, n8590, n8592, n8593, n8594,
n8595, n8597, n8598, n8599, n8600, n8602, n8603, n8604, n8605, n8607,
n8608, n8609, n8610, n8612, n8613, n8614, n8615, n8617, n8618, n8619,
n8620, n8622, n8623, n8624, n8625, n8627, n8628, n8629, n8630, n8632,
n8633, n8634, n8635, n8637, n8638, n8639, n8640, n8642, n8643, n8644,
n8645, n8647, n8648, n8649, n8650, n8652, n8653, n8654, n8655, n8657,
n8658, n8659, n8660, n8662, n8663, n8664, n8665, n8667, n8668, n8669,
n8670, n8672, n8673, n8674, n8675, n8677, n8678, n8679, n8680, n8682,
n8683, n8684, n8685, n8687, n8688, n8689, n8690, n8692, n8693, n8694,
n8695, n8697, n8698, n8699, n8700, n8702, n8703, n8704, n8705, n8707,
n8708, n8709, n8710, n8712, n8713, n8714, n8715, n8717, n8718, n8719,
n8720, n8722, n8723, n8724, n8725, n8727, n8728, n8729, n8730, n8732,
n8733, n8734, n8735, n8737, n8738, n8739, n8740, n8742, n8743, n8744,
n8745, n8747, n8748, n8749, n8750, n8752, n8753, n8754, n8755, n8757,
n8758, n8759, n8760, n8762, n8763, n8764, n8765, n8767, n8768, n8769,
n8770, n8772, n8773, n8774, n8775, n8777, n8778, n8779, n8780, n8782,
n8783, n8784, n8785, n8787, n8788, n8789, n8790, n8792, n8793, n8794,
n8795, n8797, n8798, n8799, n8800, n8802, n8803, n8804, n8805, n8807,
n8808, n8809, n8810, n8812, n8813, n8814, n8815, n8817, n8818, n8819,
n8820, n8822, n8823, n8824, n8825, n8827, n8828, n8829, n8830, n8832,
n8833, n8834, n8835, n8837, n8838, n8839, n8840, n8842, n8843, n8844,
n8845, n8847, n8848, n8849, n8850, n8852, n8853, n8854, n8855, n8857,
n8858, n8859, n8860, n8862, n8863, n8864, n8865, n8867, n8868, n8869,
n8870, n8872, n8873, n8874, n8875, n8877, n8878, n8879, n8880, n8882,
n8883, n8884, n8885, n8887, n8888, n8889, n8890, n8892, n8893, n8894,
n8895, n8897, n8898, n8899, n8900, n8902, n8903, n8904, n8905, n8907,
n8908, n8909, n8910, n8912, n8913, n8914, n8915, n8917, n8918, n8919,
n8920, n8922, n8923, n8924, n8925, n8927, n8928, n8929, n8930, n8932,
n8933, n8934, n8935, n8937, n8938, n8939, n8940, n8942, n8943, n8944,
n8945, n8947, n8948, n8949, n8950, n8952, n8953, n8954, n8955, n8957,
n8958, n8959, n8960, n8962, n8963, n8964, n8965, n8967, n8968, n8969,
n8970, n8972, n8973, n8974, n8975, n8977, n8978, n8979, n8980, n8982,
n8983, n8984, n8985, n8987, n8988, n8989, n8990, n8992, n8993, n8994,
n8995, n8997, n8998, n8999, n9000, n9002, n9003, n9004, n9005, n9007,
n9008, n9009, n9010, n9012, n9013, n9014, n9015, n9017, n9018, n9019,
n9020, n9022, n9023, n9024, n9025, n9027, n9028, n9029, n9030, n9032,
n9033, n9034, n9035, n9037, n9038, n9039, n9040, n9042, n9043, n9044,
n9045, n9047, n9048, n9049, n9050, n9052, n9053, n9054, n9055, n9057,
n9058, n9059, n9060, n9062, n9063, n9064, n9065, n9067, n9068, n9069,
n9070, n9072, n9073, n9074, n9075, n9077, n9078, n9079, n9080, n9082,
n9083, n9084, n9085, n9087, n9088, n9089, n9090, n9092, n9093, n9094,
n9095, n9097, n9098, n9099, n9100, n9102, n9103, n9104, n9105, n9107,
n9108, n9109, n9110, n9112, n9113, n9114, n9115, n9117, n9118, n9119,
n9120, n9122, n9123, n9124, n9125, n9127, n9128, n9129, n9130, n9133,
n9134, n9135, n9137, n9138, n9139, n9140, n9142, n9143, n9144, n9145,
n9147, n9148, n9149, n9150, n9152, n9153, n9154, n9155, n9157, n9158,
n9159, n9160, n9162, n9163, n9164, n9165, n9167, n9168, n9169, n9170,
n9172, n9173, n9174, n9175, n9177, n9178, n9179, n9180, n9182, n9183,
n9184, n9185, n9187, n9188, n9189, n9190, n9192, n9193, n9194, n9195,
n9197, n9198, n9199, n9200, n9202, n9203, n9204, n9205, n9207, n9208,
n9209, n9210, n9212, n9213, n9214, n9215, n9217, n9218, n9219, n9220,
n9222, n9223, n9224, n9225, n9227, n9228, n9229, n9230, n9232, n9233,
n9234, n9235, n9237, n9238, n9239, n9240, n9242, n9243, n9244, n9245,
n9247, n9248, n9249, n9250, n9252, n9253, n9254, n9255, n9257, n9258,
n9259, n9260, n9262, n9263, n9264, n9265, n9267, n9268, n9269, n9270,
n9272, n9273, n9274, n9275, n9277, n9278, n9279, n9280, n9282, n9283,
n9284, n9285, n9287, n9288, n9289, n9290, n9292, n9293, n9294, n9295,
n9297, n9298, n9299, n9300, n9302, n9303, n9304, n9305, n9307, n9308,
n9309, n9310, n9312, n9313, n9314, n9315, n9317, n9318, n9319, n9320,
n9322, n9323, n9324, n9325, n9327, n9330, n9332, n9333, n9334, n9335,
n9337, n9338, n9339, n9340, n9342, n9343, n9344, n9345, n9347, n9348,
n9349, n9350, n9352, n9353, n9354, n9355, n9357, n9358, n9359, n9360,
n9362, n9363, n9364, n9365, n9367, n9368, n9369, n9370, n9372, n9373,
n9374, n9375, n9377, n9378, n9379, n9380, n9382, n9383, n9384, n9385,
n9387, n9388, n9389, n9390, n9392, n9393, n9394, n9395, n9397, n9398,
n9399, n9400, n9402, n9403, n9404, n9405, n9407, n9408, n9409, n9410,
n9412, n9413, n9414, n9415, n9417, n9418, n9419, n9420, n9422, n9423,
n9424, n9425, n9427, n9428, n9429, n9430, n9432, n9433, n9434, n9435,
n9437, n9438, n9439, n9440, n9442, n9443, n9445, n9447, n9448, n9449,
n9450, n9452, n9453, n9454, n9455, n9457, n9458, n9459, n9460, n9462,
n9463, n9464, n9465, n9467, n9468, n9469, n9470, n9472, n9473, n9474,
n9475, n9477, n9478, n9479, n9480, n9482, n9483, n9484, n9485, n9487,
n9488, n9489, n9490, n9492, n9493, n9494, n9495, n9497, n9498, n9499,
n9500, n9502, n9503, n9504, n9505, n9507, n9508, n9509, n9510, n9512,
n9513, n9514, n9515, n9517, n9518, n9519, n9520, n9522, n9523, n9524,
n9525, n9527, n9528, n9529, n9530, n9532, n9533, n9534, n9535, n9537,
n9538, n9539, n9540, n9542, n9543, n9544, n9545, n9547, n9548, n9549,
n9550, n9552, n9553, n9554, n9555, n9557, n9558, n9559, n9560, n9562,
n9563, n9564, n9565, n9567, n9568, n9569, n9570, n9572, n9573, n9574,
n9575, n9577, n9578, n9579, n9580, n9582, n9583, n9584, n9585, n9586,
n9587, n9588, n9589, n9590, n9592, n9593, n9594, n9595, n9597, n9598,
n9599, n9600, n9602, n9603, n9604, n9605, n9607, n9608, n9609, n9610,
n9612, n9613, n9614, n9615, n9617, n9618, n9619, n9620, n9622, n9623,
n9624, n9625, n9627, n9628, n9629, n9630, n9632, n9633, n9634, n9635,
n9637, n9638, n9639, n9640, n9642, n9643, n9644, n9645, n9647, n9648,
n9649, n9650, n9652, n9653, n9654, n9655, n9657, n9658, n9659, n9660,
n9662, n9663, n9664, n9665, n9667, n9668, n9669, n9670, n9672, n9673,
n9674, n9675, n9677, n9678, n9679, n9680, n9682, n9683, n9684, n9685,
n9687, n9688, n9689, n9690, n9692, n9693, n9694, n9695, n9697, n9698,
n9699, n9700, n9702, n9703, n9704, n9705, n9707, n9708, n9709, n9710,
n9712, n9713, n9714, n9715, n9717, n9718, n9719, n9720, n9722, n9723,
n9724, n9725, n9727, n9728, n9729, n9730, n9732, n9733, n9734, n9735,
n9737, n9738, n9739, n9740, n9742, n9743, n9744, n9745, n9747, n9748,
n9749, n9750, n9752, n9753, n9754, n9755, n9757, n9758, n9759, n9760,
n9762, n9763, n9764, n9765, n9767, n9768, n9769, n9770, n9772, n9773,
n9774, n9775, n9777, n9778, n9779, n9780, n9782, n9783, n9784, n9785,
n9787, n9788, n9789, n9790, n9792, n9793, n9794, n9795, n9797, n9798,
n9799, n9800, n9802, n9803, n9804, n9805, n9807, n9808, n9809, n9810,
n9812, n9813, n9814, n9815, n9817, n9818, n9819, n9820, n9822, n9823,
n9824, n9825, n9827, n9828, n9829, n9830, n9832, n9833, n9834, n9835,
n9837, n9838, n9839, n9840, n9842, n9843, n9844, n9845, n9847, n9848,
n9849, n9850, n9852, n9853, n9854, n9855, n9857, n9858, n9859, n9860,
n9862, n9863, n9864, n9868, n9869, n9873, n9874, n9875, n9877, n9880,
n9882, n9883, n9884, n9885, n9887, n9888, n9889, n9890, n9892, n9893,
n9894, n9895, n9897, n9898, n9899, n9900, n9902, n9905, n9907, n9908,
n9909, n9910, n9912, n9913, n9914, n9915, n9917, n9918, n9919, n9920,
n9922, n9923, n9924, n9925, n9927, n9928, n9929, n9930, n9932, n9933,
n9934, n9935, n9937, n9938, n9939, n9940, n9942, n9943, n9944, n9945,
n9947, n9948, n9949, n9950, n9952, n9953, n9954, n9955, n9957, n9958,
n9959, n9960, n9962, n9963, n9964, n9965, n9967, n9968, n9969, n9970,
n9972, n9973, n9974, n9975, n9977, n9978, n9979, n9980, n9982, n9983,
n9984, n9985, n9987, n9988, n9989, n9990, n9992, n9993, n9994, n9995,
n9997, n9998, n9999, n10000, n10002, n10003, n10004, n10005, n10006,
n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
n10055, n10056, n10057, n10058, n10059, n10060, n10062, n10063,
n10064, n10065, n10067, n10068, n10069, n10070, n10072, n10073,
n10074, n10075, n10077, n10078, n10079, n10080, n10082, n10083,
n10084, n10085, n10087, n10088, n10089, n10090, n10092, n10093,
n10094, n10095, n10097, n10098, n10099, n10100, n10102, n10103,
n10104, n10105, n10107, n10108, n10109, n10110, n10112, n10113,
n10114, n10115, n10117, n10118, n10119, n10120, n10122, n10123,
n10124, n10125, n10127, n10128, n10129, n10130, n10132, n10133,
n10134, n10135, n10137, n10138, n10139, n10140, n10142, n10143,
n10144, n10145, n10147, n10148, n10149, n10150, n10152, n10153,
n10154, n10155, n10157, n10158, n10159, n10160, n10162, n10163,
n10164, n10165, n10167, n10168, n10169, n10170, n10172, n10173,
n10174, n10175, n10177, n10178, n10179, n10180, n10182, n10183,
n10184, n10185, n10187, n10188, n10189, n10190, n10192, n10193,
n10194, n10195, n10197, n10198, n10199, n10200, n10202, n10203,
n10204, n10205, n10207, n10208, n10209, n10210, n10212, n10213,
n10214, n10215, n10217, n10218, n10219, n10220, n10222, n10223,
n10224, n10225, n10227, n10228, n10229, n10230, n10232, n10233,
n10234, n10235, n10237, n10238, n10239, n10240, n10242, n10243,
n10244, n10245, n10247, n10248, n10249, n10250, n10252, n10253,
n10254, n10255, n10257, n10258, n10259, n10260, n10262, n10263,
n10264, n10265, n10267, n10268, n10269, n10270, n10272, n10273,
n10274, n10275, n10277, n10278, n10279, n10280, n10282, n10283,
n10284, n10285, n10287, n10288, n10289, n10290, n10292, n10293,
n10294, n10295, n10297, n10298, n10299, n10300, n10302, n10303,
n10304, n10305, n10307, n10308, n10309, n10310, n10312, n10313,
n10314, n10315, n10317, n10318, n10319, n10320, n10322, n10323,
n10324, n10325, n10327, n10328, n10329, n10330, n10332, n10333,
n10334, n10335, n10337, n10338, n10339, n10340, n10342, n10343,
n10344, n10345, n10347, n10348, n10349, n10350, n10352, n10353,
n10354, n10355, n10357, n10358, n10359, n10360, n10362, n10363,
n10364, n10365, n10367, n10368, n10369, n10370, n10372, n10373,
n10374, n10375, n10377, n10378, n10379, n10380, n10382, n10383,
n10384, n10385, n10387, n10388, n10389, n10390, n10392, n10393,
n10394, n10395, n10397, n10398, n10399, n10400, n10402, n10403,
n10404, n10405, n10407, n10408, n10409, n10410, n10412, n10413,
n10414, n10415, n10417, n10418, n10419, n10420, n10422, n10423,
n10424, n10425, n10427, n10428, n10429, n10430, n10432, n10433,
n10434, n10435, n10437, n10438, n10439, n10440, n10442, n10443,
n10444, n10445, n10447, n10448, n10449, n10450, n10452, n10453,
n10454, n10455, n10457, n10458, n10459, n10460, n10462, n10463,
n10464, n10465, n10467, n10468, n10469, n10470, n10472, n10473,
n10474, n10475, n10477, n10478, n10479, n10480, n10482, n10483,
n10484, n10485, n10487, n10488, n10489, n10490, n10492, n10493,
n10494, n10495, n10497, n10498, n10499, n10500, n10502, n10503,
n10504, n10505, n10507, n10508, n10509, n10510, n10512, n10513,
n10514, n10515, n10517, n10518, n10519, n10520, n10522, n10523,
n10524, n10525, n10527, n10528, n10529, n10530, n10532, n10533,
n10534, n10535, n10537, n10538, n10539, n10540, n10542, n10543,
n10544, n10545, n10547, n10548, n10549, n10550, n10552, n10553,
n10554, n10555, n10557, n10558, n10559, n10560, n10562, n10563,
n10564, n10565, n10567, n10568, n10569, n10570, n10572, n10573,
n10574, n10575, n10577, n10578, n10579, n10580, n10582, n10583,
n10584, n10585, n10587, n10588, n10589, n10590, n10592, n10593,
n10594, n10595, n10597, n10598, n10599, n10600, n10602, n10603,
n10604, n10605, n10607, n10608, n10609, n10610, n10612, n10613,
n10614, n10615, n10617, n10618, n10619, n10620, n10622, n10623,
n10624, n10625, n10627, n10628, n10629, n10630, n10632, n10633,
n10634, n10635, n10637, n10638, n10639, n10640, n10642, n10643,
n10644, n10645, n10647, n10648, n10649, n10650, n10652, n10653,
n10654, n10655, n10657, n10658, n10659, n10660, n10662, n10663,
n10664, n10665, n10667, n10668, n10669, n10670, n10672, n10673,
n10674, n10675, n10677, n10678, n10679, n10680, n10682, n10683,
n10684, n10685, n10687, n10688, n10689, n10690, n10692, n10693,
n10694, n10695, n10697, n10698, n10699, n10700, n10702, n10703,
n10704, n10705, n10707, n10708, n10709, n10710, n10712, n10713,
n10714, n10715, n10717, n10718, n10719, n10720, n10722, n10723,
n10724, n10725, n10727, n10728, n10729, n10730, n10732, n10733,
n10734, n10735, n10737, n10738, n10739, n10740, n10742, n10743,
n10744, n10745, n10747, n10748, n10749, n10750, n10752, n10753,
n10754, n10755, n10757, n10758, n10759, n10760, n10762, n10763,
n10764, n10765, n10767, n10769, n10770, n10772, n10773, n10774,
n10775, n10777, n10778, n10779, n10780, n10782, n10783, n10784,
n10785, n10787, n10788, n10789, n10790, n10792, n10793, n10794,
n10795, n10797, n10798, n10799, n10800, n10802, n10803, n10804,
n10805, n10807, n10808, n10809, n10810, n10812, n10813, n10814,
n10815, n10817, n10818, n10819, n10820, n10822, n10823, n10824,
n10825, n10827, n10828, n10829, n10830, n10832, n10833, n10834,
n10835, n10837, n10838, n10839, n10840, n10842, n10843, n10844,
n10845, n10847, n10848, n10849, n10850, n10852, n10853, n10854,
n10855, n10857, n10858, n10859, n10860, n10862, n10863, n10864,
n10865, n10867, n10868, n10869, n10870, n10872, n10873, n10874,
n10875, n10877, n10878, n10879, n10880, n10882, n10883, n10884,
n10885, n10887, n10888, n10889, n10890, n10892, n10893, n10894,
n10895, n10897, n10898, n10899, n10900, n10902, n10903, n10904,
n10905, n10907, n10908, n10909, n10910, n10912, n10913, n10914,
n10915, n10917, n10918, n10919, n10920, n10922, n10923, n10924,
n10925, n10927, n10928, n10929, n10930, n10932, n10933, n10934,
n10935, n10937, n10938, n10939, n10940, n10942, n10943, n10944,
n10945, n10947, n10948, n10949, n10950, n10952, n10953, n10954,
n10955, n10957, n10958, n10959, n10960, n10962, n10963, n10964,
n10965, n10967, n10968, n10969, n10970, n10972, n10973, n10974,
n10975, n10977, n10978, n10979, n10980, n10982, n10983, n10984,
n10985, n10987, n10988, n10989, n10990, n10992, n10993, n10994,
n10995, n10997, n10998, n10999, n11000, n11002, n11003, n11004,
n11005, n11007, n11008, n11009, n11010, n11012, n11013, n11014,
n11015, n11017, n11018, n11019, n11020, n11022, n11023, n11024,
n11025, n11027, n11028, n11029, n11030, n11032, n11033, n11034,
n11035, n11037, n11038, n11039, n11040, n11042, n11043, n11044,
n11045, n11047, n11048, n11049, n11050, n11052, n11053, n11054,
n11055, n11057, n11058, n11059, n11060, n11062, n11063, n11064,
n11065, n11067, n11068, n11069, n11070, n11072, n11073, n11074,
n11075, n11077, n11078, n11079, n11080, n11082, n11083, n11084,
n11085, n11087, n11088, n11089, n11090, n11092, n11093, n11094,
n11095, n11097, n11098, n11099, n11100, n11102, n11103, n11104,
n11105, n11107, n11108, n11109, n11110, n11112, n11113, n11114,
n11115, n11117, n11118, n11119, n11120, n11122, n11123, n11124,
n11125, n11127, n11128, n11129, n11130, n11132, n11133, n11134,
n11135, n11137, n11138, n11139, n11140, n11142, n11143, n11144,
n11145, n11147, n11148, n11149, n11150, n11152, n11153, n11154,
n11155, n11157, n11158, n11159, n11160, n11162, n11163, n11164,
n11165, n11167, n11168, n11169, n11170, n11172, n11173, n11174,
n11175, n11177, n11178, n11179, n11180, n11182, n11183, n11184,
n11185, n11187, n11188, n11189, n11190, n11192, n11193, n11194,
n11195, n11197, n11198, n11199, n11200, n11202, n11203, n11204,
n11205, n11207, n11208, n11209, n11210, n11212, n11213, n11214,
n11215, n11217, n11218, n11219, n11220, n11222, n11223, n11224,
n11225, n11227, n11228, n11229, n11230, n11232, n11233, n11234,
n11235, n11237, n11238, n11239, n11240, n11242, n11243, n11244,
n11245, n11247, n11248, n11249, n11250, n11252, n11253, n11254,
n11255, n11257, n11258, n11259, n11260, n11262, n11263, n11264,
n11265, n11267, n11268, n11269, n11270, n11272, n11273, n11274,
n11275, n11277, n11278, n11279, n11280, n11282, n11283, n11284,
n11285, n11287, n11288, n11289, n11290, n11292, n11293, n11294,
n11295, n11297, n11298, n11299, n11300, n11302, n11303, n11304,
n11305, n11307, n11308, n11309, n11310, n11312, n11313, n11314,
n11315, n11317, n11318, n11319, n11320, n11322, n11323, n11324,
n11325, n11327, n11328, n11329, n11330, n11332, n11333, n11334,
n11335, n11337, n11338, n11339, n11340, n11342, n11343, n11344,
n11345, n11347, n11348, n11349, n11350, n11352, n11353, n11354,
n11355, n11357, n11358, n11359, n11360, n11362, n11363, n11364,
n11365, n11367, n11368, n11369, n11370, n11372, n11373, n11374,
n11375, n11377, n11378, n11379, n11380, n11382, n11383, n11384,
n11385, n11387, n11388, n11389, n11390, n11392, n11393, n11394,
n11395, n11397, n11398, n11399, n11400, n11402, n11403, n11404,
n11405, n11407, n11408, n11409, n11410, n11412, n11413, n11414,
n11415, n11417, n11418, n11419, n11420, n11422, n11423, n11424,
n11425, n11427, n11428, n11429, n11430, n11432, n11433, n11434,
n11435, n11437, n11438, n11439, n11440, n11442, n11443, n11444,
n11445, n11447, n11448, n11449, n11450, n11452, n11453, n11454,
n11455, n11457, n11458, n11459, n11460, n11462, n11463, n11464,
n11465, n11467, n11468, n11469, n11470, n11472, n11473, n11474,
n11475, n11477, n11478, n11479, n11480, n11482, n11483, n11484,
n11485, n11487, n11488, n11489, n11490, n11492, n11493, n11494,
n11495, n11497, n11498, n11499, n11500, n11502, n11503, n11504,
n11505, n11507, n11508, n11509, n11510, n11512, n11513, n11514,
n11515, n11517, n11518, n11519, n11520, n11522, n11523, n11524,
n11525, n11527, n11528, n11529, n11530, n11532, n11533, n11534,
n11535, n11537, n11538, n11539, n11540, n11542, n11543, n11544,
n11545, n11547, n11548, n11549, n11550, n11552, n11553, n11554,
n11555, n11557, n11558, n11559, n11560, n11562, n11563, n11564,
n11565, n11567, n11568, n11569, n11570, n11572, n11573, n11574,
n11575, n11577, n11578, n11579, n11580, n11582, n11583, n11584,
n11585, n11587, n11588, n11589, n11590, n11592, n11593, n11594,
n11595, n11597, n11598, n11599, n11600, n11602, n11603, n11604,
n11605, n11607, n11608, n11609, n11610, n11612, n11613, n11614,
n11615, n11617, n11618, n11619, n11620, n11622, n11623, n11624,
n11625, n11627, n11628, n11629, n11630, n11632, n11633, n11634,
n11635, n11637, n11638, n11639, n11640, n11642, n11643, n11644,
n11645, n11647, n11648, n11649, n11650, n11652, n11653, n11654,
n11655, n11657, n11658, n11659, n11660, n11662, n11663, n11664,
n11665, n11667, n11668, n11669, n11670, n11672, n11673, n11674,
n11675, n11677, n11678, n11679, n11680, n11682, n11683, n11684,
n11685, n11687, n11688, n11689, n11690, n11692, n11693, n11694,
n11695, n11697, n11698, n11699, n11700, n11702, n11703, n11704,
n11705, n11707, n11708, n11709, n11710, n11712, n11713, n11714,
n11715, n11717, n11718, n11719, n11720, n11722, n11723, n11724,
n11725, n11727, n11728, n11729, n11730, n11732, n11733, n11734,
n11735, n11737, n11738, n11739, n11740, n11742, n11743, n11744,
n11745, n11747, n11748, n11749, n11750, n11752, n11753, n11754,
n11755, n11757, n11758, n11759, n11760, n11762, n11763, n11764,
n11765, n11767, n11768, n11769, n11770, n11772, n11773, n11774,
n11775, n11777, n11778, n11779, n11780, n11782, n11783, n11784,
n11785, n11787, n11788, n11789, n11790, n11792, n11793, n11794,
n11795, n11797, n11798, n11799, n11800, n11802, n11803, n11804,
n11805, n11807, n11808, n11809, n11810, n11812, n11813, n11814,
n11815, n11817, n11818, n11819, n11820, n11822, n11823, n11824,
n11825, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
n11834, n11835, n11837, n11838, n11839, n11840, n11842, n11843,
n11844, n11845, n11847, n11848, n11849, n11850, n11852, n11853,
n11854, n11855, n11857, n11858, n11859, n11860, n11862, n11863,
n11864, n11865, n11867, n11868, n11869, n11870, n11872, n11873,
n11874, n11875, n11877, n11878, n11879, n11880, n11882, n11883,
n11884, n11885, n11887, n11888, n11889, n11890, n11892, n11893,
n11894, n11895, n11897, n11898, n11899, n11900, n11902, n11903,
n11904, n11905, n11907, n11908, n11909, n11910, n11912, n11913,
n11914, n11915, n11917, n11918, n11919, n11920, n11922, n11923,
n11924, n11925, n11927, n11928, n11929, n11930, n11932, n11933,
n11934, n11935, n11937, n11938, n11939, n11940, n11942, n11943,
n11944, n11945, n11947, n11948, n11949, n11950, n11952, n11953,
n11954, n11955, n11957, n11958, n11959, n11960, n11962, n11963,
n11964, n11965, n11967, n11968, n11969, n11970, n11972, n11973,
n11974, n11975, n11977, n11978, n11979, n11980, n11982, n11983,
n11984, n11985, n11987, n11988, n11989, n11990, n11992, n11993,
n11994, n11995, n11997, n11998, n11999, n12000, n12002, n12003,
n12004, n12005, n12007, n12008, n12009, n12010, n12012, n12013,
n12014, n12015, n12017, n12018, n12019, n12020, n12022, n12023,
n12024, n12025, n12027, n12028, n12029, n12030, n12032, n12033,
n12034, n12035, n12037, n12038, n12039, n12040, n12042, n12043,
n12044, n12045, n12047, n12048, n12049, n12050, n12052, n12053,
n12054, n12055, n12057, n12058, n12059, n12060, n12062, n12064,
n12065, n12067, n12068, n12069, n12070, n12072, n12073, n12074,
n12075, n12077, n12078, n12079, n12080, n12082, n12083, n12084,
n12085, n12087, n12088, n12089, n12090, n12092, n12093, n12094,
n12095, n12097, n12098, n12099, n12100, n12102, n12103, n12104,
n12105, n12107, n12108, n12109, n12110, n12112, n12113, n12114,
n12115, n12117, n12118, n12119, n12120, n12122, n12123, n12124,
n12125, n12127, n12128, n12129, n12130, n12132, n12133, n12134,
n12135, n12137, n12138, n12139, n12140, n12142, n12143, n12144,
n12145, n12147, n12148, n12149, n12150, n12152, n12153, n12154,
n12155, n12157, n12158, n12159, n12160, n12162, n12163, n12164,
n12165, n12167, n12168, n12169, n12170, n12172, n12173, n12174,
n12175, n12177, n12178, n12179, n12180, n12182, n12183, n12184,
n12185, n12187, n12188, n12189, n12190, n12192, n12193, n12194,
n12195, n12197, n12198, n12199, n12200, n12202, n12203, n12204,
n12205, n12207, n12208, n12209, n12210, n12212, n12213, n12214,
n12215, n12217, n12218, n12219, n12220, n12222, n12223, n12224,
n12225, n12227, n12228, n12229, n12230, n12232, n12233, n12234,
n12235, n12237, n12238, n12239, n12240, n12242, n12243, n12244,
n12245, n12247, n12248, n12249, n12250, n12252, n12253, n12254,
n12257, n12258, n12259, n12260, n12262, n12263, n12264, n12265,
n12267, n12268, n12269, n12270, n12272, n12273, n12274, n12275,
n12277, n12278, n12279, n12280, n12282, n12283, n12284, n12285,
n12287, n12288, n12289, n12290, n12292, n12293, n12294, n12295,
n12297, n12298, n12299, n12300, n12302, n12303, n12304, n12305,
n12307, n12308, n12309, n12310, n12312, n12313, n12314, n12315,
n12317, n12318, n12319, n12320, n12322, n12323, n12324, n12325,
n12327, n12328, n12329, n12330, n12332, n12333, n12334, n12335,
n12338, n12339, n12340, n12342, n12343, n12344, n12345, n12347,
n12348, n12349, n12350, n12352, n12353, n12354, n12355, n12357,
n12358, n12359, n12360, n12362, n12363, n12364, n12365, n12367,
n12368, n12369, n12370, n12372, n12373, n12374, n12375, n12377,
n12378, n12379, n12380, n12382, n12383, n12384, n12385, n12387,
n12388, n12389, n12390, n12392, n12393, n12394, n12395, n12397,
n12398, n12399, n12400, n12402, n12403, n12404, n12405, n12407,
n12408, n12409, n12410, n12412, n12413, n12414, n12415, n12417,
n12418, n12419, n12420, n12422, n12423, n12424, n12425, n12427,
n12428, n12429, n12430, n12432, n12433, n12434, n12435, n12437,
n12438, n12439, n12440, n12442, n12443, n12444, n12445, n12447,
n12448, n12449, n12450, n12452, n12453, n12454, n12455, n12457,
n12458, n12459, n12460, n12462, n12463, n12464, n12465, n12467,
n12468, n12469, n12470, n12472, n12473, n12474, n12475, n12477,
n12478, n12479, n12480, n12482, n12483, n12484, n12485, n12487,
n12488, n12489, n12490, n12492, n12493, n12494, n12495, n12497,
n12498, n12499, n12500, n12502, n12503, n12504, n12505, n12507,
n12508, n12509, n12510, n12512, n12513, n12514, n12515, n12517,
n12518, n12519, n12520, n12522, n12523, n12524, n12525, n12527,
n12528, n12529, n12530, n12532, n12533, n12534, n12535, n12537,
n12538, n12539, n12540, n12542, n12543, n12544, n12545, n12547,
n12548, n12549, n12550, n12552, n12553, n12554, n12555, n12557,
n12558, n12559, n12560, n12562, n12563, n12564, n12565, n12567,
n12568, n12569, n12570, n12572, n12573, n12574, n12575, n12577,
n12578, n12579, n12580, n12582, n12583, n12584, n12585, n12587,
n12588, n12589, n12590, n12592, n12593, n12594, n12595, n12597,
n12598, n12599, n12600, n12602, n12603, n12604, n12605, n12607,
n12608, n12609, n12610, n12612, n12613, n12614, n12615, n12617,
n12618, n12619, n12620, n12622, n12623, n12624, n12625, n12627,
n12628, n12629, n12630, n12632, n12633, n12634, n12635, n12637,
n12638, n12639, n12640, n12642, n12643, n12644, n12645, n12647,
n12648, n12649, n12650, n12652, n12653, n12654, n12655, n12657,
n12658, n12659, n12660, n12662, n12663, n12664, n12665, n12667,
n12668, n12669, n12670, n12672, n12673, n12674, n12675, n12677,
n12678, n12679, n12680, n12682, n12683, n12684, n12685, n12687,
n12688, n12689, n12690, n12692, n12693, n12694, n12695, n12697,
n12698, n12699, n12700, n12702, n12703, n12704, n12705, n12707,
n12708, n12709, n12710, n12712, n12713, n12714, n12715, n12717,
n12718, n12719, n12720, n12722, n12723, n12724, n12725, n12727,
n12728, n12729, n12730, n12732, n12733, n12734, n12735, n12737,
n12738, n12739, n12740, n12742, n12743, n12744, n12745, n12747,
n12748, n12749, n12750, n12752, n12753, n12754, n12755, n12757,
n12758, n12759, n12760, n12762, n12763, n12764, n12768, n12769,
n12770, n12772, n12773, n12774, n12775, n12777, n12778, n12779,
n12780, n12782, n12783, n12784, n12785, n12787, n12788, n12789,
n12790, n12792, n12793, n12794, n12795, n12797, n12798, n12799,
n12800, n12802, n12803, n12804, n12805, n12807, n12808, n12809,
n12810, n12812, n12813, n12814, n12815, n12817, n12818, n12819,
n12820, n12822, n12823, n12824, n12825, n12827, n12828, n12829,
n12830, n12832, n12833, n12834, n12835, n12837, n12838, n12839,
n12840, n12842, n12843, n12844, n12845, n12847, n12848, n12849,
n12850, n12852, n12853, n12854, n12855, n12857, n12858, n12859,
n12860, n12862, n12863, n12864, n12865, n12867, n12868, n12869,
n12870, n12872, n12873, n12874, n12875, n12877, n12878, n12879,
n12880, n12882, n12883, n12884, n12885, n12887, n12888, n12889,
n12890, n12892, n12893, n12894, n12895, n12897, n12898, n12899,
n12900, n12902, n12903, n12904, n12905, n12907, n12908, n12909,
n12910, n12912, n12913, n12914, n12915, n12919, n12920, n12922,
n12923, n12924, n12925, n12927, n12928, n12929, n12930, n12932,
n12933, n12934, n12935, n12937, n12938, n12939, n12940, n12942,
n12943, n12944, n12945, n12947, n12948, n12949, n12950, n12952,
n12953, n12954, n12955, n12957, n12958, n12959, n12960, n12962,
n12963, n12964, n12965, n12967, n12968, n12969, n12970, n12972,
n12973, n12974, n12975, n12977, n12978, n12979, n12980, n12982,
n12983, n12984, n12985, n12987, n12988, n12990, n12992, n12993,
n12994, n12997, n12998, n12999, n13000, n13002, n13003, n13004,
n13005, n13007, n13008, n13009, n13010, n13012, n13013, n13014,
n13015, n13017, n13018, n13019, n13020, n13022, n13023, n13024,
n13025, n13027, n13028, n13029, n13030, n13032, n13033, n13034,
n13035, n13037, n13038, n13039, n13040, n13042, n13043, n13044,
n13045, n13047, n13048, n13049, n13050, n13052, n13053, n13054,
n13055, n13057, n13058, n13059, n13060, n13062, n13063, n13064,
n13065, n13067, n13068, n13069, n13070, n13072, n13073, n13074,
n13075, n13077, n13078, n13079, n13080, n13082, n13083, n13084,
n13085, n13087, n13088, n13089, n13090, n13092, n13093, n13094,
n13095, n13097, n13098, n13099, n13100, n13102, n13103, n13104,
n13105, n13107, n13108, n13109, n13110, n13112, n13113, n13114,
n13115, n13117, n13118, n13119, n13120, n13122, n13123, n13124,
n13125, n13127, n13128, n13129, n13130, n13132, n13133, n13134,
n13135, n13137, n13138, n13139, n13140, n13142, n13143, n13144,
n13145, n13147, n13148, n13149, n13150, n13152, n13153, n13154,
n13155, n13157, n13158, n13159, n13160, n13162, n13163, n13164,
n13165, n13167, n13168, n13169, n13170, n13172, n13173, n13174,
n13175, n13177, n13178, n13179, n13180, n13182, n13183, n13184,
n13185, n13187, n13188, n13189, n13190, n13192, n13193, n13194,
n13195, n13197, n13198, n13199, n13200, n13202, n13203, n13204,
n13205, n13207, n13208, n13209, n13210, n13212, n13213, n13214,
n13215, n13217, n13218, n13219, n13220, n13222, n13223, n13224,
n13225, n13227, n13228, n13229, n13230, n13232, n13233, n13234,
n13235, n13237, n13238, n13239, n13240, n13242, n13243, n13244,
n13245, n13247, n13248, n13249, n13250, n13252, n13253, n13254,
n13255, n13257, n13258, n13259, n13260, n13262, n13263, n13264,
n13265, n13267, n13268, n13269, n13270, n13272, n13273, n13274,
n13275, n13277, n13278, n13279, n13280, n13282, n13283, n13284,
n13285, n13287, n13288, n13289, n13290, n13292, n13293, n13294,
n13295, n13297, n13298, n13299, n13300, n13302, n13303, n13304,
n13305, n13307, n13308, n13309, n13310, n13312, n13313, n13314,
n13315, n13317, n13318, n13319, n13320, n13322, n13323, n13324,
n13325, n13327, n13328, n13329, n13330, n13332, n13333, n13334,
n13335, n13337, n13338, n13339, n13340, n13342, n13343, n13344,
n13345, n13347, n13348, n13349, n13350, n13352, n13353, n13354,
n13355, n13357, n13358, n13359, n13360, n13362, n13363, n13364,
n13365, n13367, n13368, n13369, n13370, n13372, n13373, n13374,
n13375, n13377, n13378, n13379, n13380, n13382, n13383, n13384,
n13385, n13387, n13388, n13389, n13390, n13392, n13393, n13394,
n13395, n13397, n13398, n13399, n13400, n13402, n13403, n13404,
n13405, n13407, n13408, n13409, n13410, n13412, n13413, n13414,
n13415, n13417, n13418, n13419, n13420, n13422, n13423, n13424,
n13425, n13427, n13428, n13429, n13430, n13432, n13433, n13434,
n13435, n13437, n13438, n13439, n13440, n13442, n13443, n13444,
n13445, n13447, n13448, n13449, n13450, n13452, n13453, n13454,
n13455, n13457, n13458, n13459, n13460, n13462, n13463, n13464,
n13465, n13467, n13468, n13469, n13470, n13472, n13473, n13474,
n13475, n13477, n13478, n13479, n13480, n13482, n13483, n13484,
n13485, n13487, n13488, n13489, n13490, n13492, n13493, n13494,
n13495, n13497, n13498, n13499, n13500, n13502, n13503, n13504,
n13505, n13507, n13508, n13509, n13510, n13512, n13513, n13514,
n13515, n13517, n13518, n13519, n13520, n13522, n13523, n13524,
n13525, n13527, n13528, n13529, n13530, n13532, n13534, n13535,
n13537, n13538, n13539, n13540, n13542, n13543, n13544, n13545,
n13547, n13548, n13549, n13550, n13552, n13553, n13554, n13555,
n13557, n13558, n13559, n13560, n13562, n13563, n13564, n13565,
n13567, n13568, n13569, n13570, n13572, n13573, n13574, n13575,
n13577, n13578, n13579, n13580, n13584, n13585, n13587, n13588,
n13589, n13590, n13592, n13593, n13594, n13595, n13597, n13598,
n13599, n13600, n13602, n13603, n13604, n13605, n13607, n13608,
n13609, n13610, n13612, n13613, n13614, n13615, n13617, n13618,
n13620, n13622, n13623, n13624, n13625, n13627, n13628, n13629,
n13630, n13632, n13633, n13634, n13635, n13637, n13638, n13639,
n13640, n13642, n13643, n13644, n13645, n13647, n13648, n13649,
n13650, n13652, n13653, n13654, n13655, n13657, n13658, n13659,
n13660, n13662, n13663, n13664, n13665, n13667, n13668, n13669,
n13670, n13672, n13673, n13674, n13675, n13677, n13678, n13679,
n13680, n13682, n13683, n13684, n13685, n13687, n13688, n13689,
n13690, n13692, n13693, n13694, n13695, n13697, n13698, n13699,
n13700, n13702, n13703, n13704, n13705, n13707, n13708, n13709,
n13710, n13712, n13713, n13714, n13715, n13717, n13718, n13719,
n13720, n13722, n13723, n13724, n13725, n13727, n13728, n13729,
n13730, n13732, n13733, n13734, n13735, n13737, n13738, n13739,
n13740, n13742, n13743, n13744, n13745, n13747, n13748, n13749,
n13750, n13752, n13753, n13754, n13755, n13757, n13758, n13759,
n13760, n13762, n13763, n13764, n13765, n13767, n13768, n13769,
n13770, n13772, n13773, n13774, n13775, n13777, n13778, n13779,
n13780, n13782, n13783, n13784, n13785, n13787, n13788, n13789,
n13790, n13792, n13793, n13794, n13795, n13797, n13798, n13799,
n13800, n13802, n13803, n13804, n13805, n13807, n13808, n13809,
n13810, n13812, n13813, n13814, n13815, n13817, n13818, n13819,
n13820, n13822, n13823, n13824, n13825, n13827, n13828, n13829,
n13830, n13832, n13833, n13834, n13835, n13837, n13838, n13839,
n13840, n13842, n13843, n13844, n13845, n13847, n13848, n13849,
n13850, n13852, n13853, n13854, n13855, n13857, n13858, n13859,
n13860, n13862, n13863, n13864, n13865, n13867, n13868, n13869,
n13870, n13872, n13873, n13874, n13875, n13877, n13878, n13879,
n13880, n13882, n13883, n13884, n13885, n13887, n13888, n13889,
n13890, n13892, n13893, n13894, n13895, n13897, n13898, n13899,
n13900, n13902, n13903, n13904, n13905, n13907, n13908, n13909,
n13910, n13912, n13913, n13914, n13915, n13917, n13918, n13919,
n13920, n13922, n13923, n13924, n13925, n13927, n13928, n13929,
n13930, n13932, n13933, n13934, n13935, n13937, n13938, n13939,
n13940, n13942, n13943, n13944, n13945, n13947, n13948, n13949,
n13950, n13952, n13953, n13954, n13955, n13957, n13958, n13959,
n13960, n13962, n13963, n13964, n13965, n13967, n13968, n13969,
n13970, n13972, n13973, n13974, n13975, n13977, n13978, n13979,
n13980, n13982, n13983, n13984, n13985, n13987, n13988, n13989,
n13990, n13992, n13993, n13994, n13995, n13997, n13998, n13999,
n14000, n14002, n14003, n14004, n14005, n14007, n14008, n14009,
n14010, n14012, n14013, n14014, n14015, n14017, n14018, n14019,
n14020, n14022, n14023, n14024, n14025, n14027, n14028, n14029,
n14030, n14032, n14033, n14034, n14035, n14037, n14038, n14039,
n14040, n14042, n14043, n14044, n14045, n14047, n14048, n14049,
n14050, n14052, n14053, n14054, n14055, n14057, n14058, n14059,
n14060, n14062, n14063, n14064, n14065, n14067, n14068, n14069,
n14070, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
n14079, n14080, n14082, n14083, n14084, n14085, n14087, n14088,
n14089, n14090, n14092, n14093, n14094, n14095, n14097, n14098,
n14099, n14100, n14102, n14103, n14104, n14105, n14107, n14108,
n14109, n14110, n14112, n14113, n14114, n14115, n14117, n14118,
n14119, n14120, n14122, n14123, n14124, n14125, n14127, n14128,
n14129, n14130, n14132, n14133, n14134, n14135, n14137, n14138,
n14139, n14140, n14142, n14143, n14144, n14145, n14147, n14148,
n14149, n14150, n14152, n14153, n14154, n14155, n14157, n14158,
n14159, n14160, n14162, n14163, n14164, n14165, n14167, n14168,
n14169, n14170, n14172, n14173, n14174, n14175, n14177, n14178,
n14179, n14180, n14182, n14183, n14184, n14185, n14187, n14188,
n14189, n14190, n14192, n14193, n14194, n14195, n14197, n14198,
n14199, n14200, n14202, n14203, n14204, n14205, n14207, n14208,
n14209, n14210, n14212, n14213, n14214, n14215, n14217, n14218,
n14219, n14220, n14222, n14223, n14224, n14225, n14227, n14228,
n14229, n14230, n14232, n14233, n14234, n14235, n14237, n14238,
n14239, n14240, n14242, n14243, n14244, n14245, n14247, n14248,
n14249, n14250, n14252, n14253, n14254, n14255, n14257, n14258,
n14259, n14260, n14262, n14263, n14264, n14265, n14267, n14268,
n14269, n14270, n14272, n14273, n14274, n14275, n14277, n14278,
n14279, n14280, n14282, n14283, n14284, n14285, n14287, n14288,
n14289, n14290, n14292, n14293, n14294, n14295, n14297, n14298,
n14299, n14300, n14302, n14303, n14304, n14305, n14307, n14308,
n14309, n14310, n14312, n14313, n14314, n14315, n14317, n14318,
n14319, n14320, n14322, n14323, n14324, n14325, n14327, n14328,
n14329, n14330, n14332, n14333, n14334, n14335, n14337, n14338,
n14339, n14340, n14342, n14343, n14344, n14345, n14347, n14348,
n14349, n14350, n14352, n14353, n14354, n14355, n14357, n14358,
n14359, n14360, n14362, n14363, n14364, n14365, n14367, n14368,
n14369, n14370, n14372, n14373, n14374, n14375, n14377, n14378,
n14379, n14380, n14382, n14383, n14384, n14385, n14387, n14388,
n14389, n14390, n14392, n14393, n14397, n14398, n14399, n14400,
n14402, n14403, n14404, n14405, n14407, n14408, n14409, n14410,
n14412, n14413, n14414, n14415, n14417, n14418, n14419, n14420,
n14422, n14423, n14424, n14425, n14427, n14428, n14429, n14430,
n14432, n14433, n14434, n14435, n14437, n14438, n14439, n14440,
n14442, n14443, n14444, n14445, n14447, n14448, n14449, n14450,
n14452, n14453, n14454, n14455, n14457, n14458, n14459, n14460,
n14462, n14463, n14464, n14465, n14467, n14468, n14469, n14470,
n14472, n14473, n14474, n14475, n14477, n14478, n14479, n14480,
n14482, n14483, n14484, n14485, n14487, n14488, n14489, n14490,
n14492, n14493, n14494, n14495, n14497, n14498, n14499, n14500,
n14502, n14503, n14504, n14505, n14507, n14508, n14509, n14510,
n14512, n14513, n14514, n14515, n14517, n14518, n14519, n14520,
n14522, n14523, n14524, n14525, n14527, n14528, n14529, n14530,
n14532, n14533, n14534, n14535, n14537, n14538, n14539, n14540,
n14542, n14543, n14544, n14545, n14547, n14548, n14549, n14550,
n14552, n14553, n14554, n14555, n14557, n14558, n14559, n14560,
n14562, n14563, n14564, n14565, n14567, n14568, n14569, n14570,
n14572, n14573, n14574, n14575, n14577, n14578, n14579, n14580,
n14582, n14583, n14584, n14585, n14587, n14588, n14589, n14590,
n14592, n14593, n14594, n14595, n14597, n14598, n14599, n14600,
n14602, n14603, n14604, n14605, n14607, n14608, n14609, n14610,
n14612, n14613, n14614, n14615, n14617, n14618, n14619, n14620,
n14622, n14623, n14624, n14625, n14627, n14628, n14629, n14630,
n14632, n14633, n14634, n14635, n14637, n14638, n14639, n14640,
n14642, n14643, n14644, n14645, n14647, n14648, n14649, n14650,
n14652, n14653, n14654, n14655, n14657, n14658, n14659, n14660,
n14662, n14663, n14664, n14665, n14667, n14668, n14669, n14670,
n14672, n14673, n14674, n14675, n14677, n14678, n14679, n14680,
n14682, n14683, n14684, n14685, n14687, n14688, n14689, n14690,
n14692, n14693, n14694, n14695, n14697, n14698, n14699, n14700,
n14702, n14703, n14704, n14705, n14707, n14708, n14709, n14710,
n14712, n14713, n14714, n14715, n14717, n14718, n14719, n14720,
n14722, n14723, n14724, n14725, n14727, n14728, n14729, n14730,
n14732, n14733, n14734, n14735, n14737, n14738, n14739, n14740,
n14742, n14743, n14744, n14745, n14747, n14748, n14749, n14750,
n14752, n14753, n14754, n14755, n14757, n14758, n14759, n14760,
n14762, n14763, n14764, n14765, n14767, n14768, n14769, n14770,
n14772, n14773, n14774, n14775, n14777, n14778, n14779, n14780,
n14782, n14783, n14784, n14785, n14787, n14788, n14789, n14790,
n14792, n14793, n14794, n14795, n14797, n14798, n14799, n14800,
n14802, n14803, n14804, n14805, n14807, n14808, n14809, n14810,
n14812, n14813, n14814, n14815, n14817, n14818, n14819, n14820,
n14822, n14823, n14824, n14825, n14827, n14828, n14829, n14830,
n14832, n14833, n14834, n14835, n14837, n14838, n14839, n14840,
n14842, n14843, n14844, n14845, n14847, n14848, n14849, n14850,
n14852, n14853, n14854, n14855, n14857, n14858, n14859, n14860,
n14862, n14863, n14864, n14865, n14867, n14868, n14869, n14870,
n14872, n14873, n14874, n14875, n14877, n14878, n14879, n14880,
n14882, n14883, n14884, n14885, n14887, n14888, n14889, n14890,
n14892, n14893, n14894, n14895, n14897, n14898, n14899, n14900,
n14902, n14903, n14904, n14905, n14907, n14908, n14909, n14910,
n14912, n14913, n14914, n14915, n14917, n14918, n14919, n14920,
n14922, n14923, n14924, n14925, n14927, n14928, n14929, n14930,
n14932, n14933, n14934, n14935, n14937, n14938, n14939, n14940,
n14942, n14943, n14944, n14945, n14947, n14948, n14949, n14950,
n14952, n14953, n14954, n14955, n14957, n14958, n14959, n14960,
n14962, n14963, n14964, n14965, n14967, n14968, n14969, n14970,
n14972, n14973, n14974, n14975, n14977, n14978, n14979, n14980,
n14982, n14983, n14984, n14985, n14987, n14988, n14989, n14990,
n14992, n14993, n14994, n14995, n14997, n14998, n14999, n15000,
n15002, n15003, n15004, n15005, n15007, n15008, n15009, n15010,
n15012, n15013, n15014, n15015, n15017, n15018, n15019, n15020,
n15022, n15023, n15024, n15025, n15027, n15028, n15029, n15030,
n15032, n15033, n15034, n15035, n15037, n15038, n15039, n15040,
n15042, n15043, n15044, n15045, n15047, n15048, n15049, n15050,
n15052, n15053, n15054, n15055, n15057, n15058, n15059, n15060,
n15062, n15063, n15064, n15065, n15067, n15068, n15069, n15070,
n15072, n15073, n15074, n15075, n15077, n15078, n15079, n15080,
n15082, n15083, n15084, n15085, n15087, n15088, n15089, n15090,
n15092, n15093, n15094, n15095, n15097, n15098, n15099, n15100,
n15102, n15103, n15104, n15105, n15107, n15108, n15109, n15110,
n15112, n15113, n15114, n15115, n15117, n15118, n15119, n15120,
n15122, n15123, n15124, n15125, n15127, n15128, n15129, n15130,
n15132, n15133, n15134, n15135, n15137, n15138, n15139, n15140,
n15142, n15143, n15144, n15145, n15147, n15148, n15149, n15150,
n15152, n15153, n15154, n15155, n15157, n15158, n15159, n15160,
n15162, n15163, n15164, n15165, n15167, n15168, n15169, n15170,
n15172, n15173, n15174, n15175, n15177, n15178, n15179, n15180,
n15182, n15183, n15184, n15185, n15187, n15188, n15189, n15190,
n15192, n15193, n15194, n15195, n15197, n15198, n15199, n15200,
n15202, n15203, n15204, n15205, n15207, n15208, n15209, n15210,
n15212, n15213, n15214, n15215, n15217, n15218, n15219, n15220,
n15222, n15223, n15224, n15225, n15227, n15228, n15229, n15230,
n15232, n15233, n15234, n15235, n15237, n15238, n15239, n15240,
n15242, n15243, n15244, n15245, n15247, n15248, n15249, n15250,
n15252, n15253, n15254, n15255, n15257, n15258, n15259, n15260,
n15262, n15263, n15264, n15265, n15267, n15268, n15269, n15270,
n15272, n15273, n15274, n15275, n15277, n15278, n15279, n15280,
n15282, n15283, n15284, n15285, n15287, n15288, n15289, n15290,
n15292, n15293, n15294, n15295, n15297, n15298, n15299, n15300,
n15302, n15303, n15304, n15305, n15307, n15308, n15309, n15310,
n15312, n15313, n15314, n15315, n15317, n15318, n15319, n15320,
n15322, n15323, n15324, n15325, n15327, n15328, n15329, n15330,
n15332, n15333, n15334, n15335, n15337, n15338, n15339, n15340,
n15342, n15343, n15344, n15345, n15347, n15348, n15349, n15350,
n15352, n15353, n15354, n15355, n15357, n15358, n15359, n15360,
n15362, n15363, n15364, n15365, n15367, n15368, n15369, n15370,
n15372, n15373, n15374, n15375, n15377, n15378, n15379, n15380,
n15382, n15383, n15384, n15385, n15387, n15388, n15389, n15390,
n15392, n15393, n15394, n15395, n15397, n15398, n15399, n15400,
n15402, n15403, n15404, n15405, n15407, n15408, n15409, n15410,
n15412, n15413, n15414, n15415, n15417, n15418, n15419, n15420,
n15422, n15423, n15424, n15425, n15427, n15428, n15429, n15430,
n15432, n15433, n15434, n15435, n15437, n15438, n15439, n15440,
n15442, n15443, n15444, n15445, n15447, n15448, n15449, n15450,
n15452, n15453, n15454, n15455, n15457, n15458, n15459, n15460,
n15462, n15463, n15464, n15465, n15467, n15468, n15469, n15470,
n15472, n15473, n15474, n15475, n15477, n15478, n15479, n15480,
n15482, n15483, n15484, n15485, n15487, n15488, n15489, n15490,
n15492, n15493, n15494, n15495, n15497, n15498, n15499, n15500,
n15502, n15503, n15504, n15505, n15507, n15508, n15509, n15510,
n15512, n15513, n15514, n15515, n15517, n15518, n15519, n15520,
n15522, n15523, n15524, n15525, n15527, n15528, n15529, n15530,
n15532, n15533, n15534, n15535, n15537, n15538, n15539, n15540,
n15542, n15543, n15544, n15545, n15547, n15548, n15549, n15550,
n15552, n15553, n15554, n15555, n15557, n15558, n15559, n15560,
n15562, n15563, n15564, n15565, n15567, n15568, n15569, n15570,
n15572, n15573, n15574, n15575, n15577, n15578, n15579, n15580,
n15582, n15583, n15584, n15585, n15587, n15588, n15589, n15590,
n15592, n15593, n15594, n15595, n15597, n15598, n15599, n15600,
n15602, n15603, n15604, n15605, n15607, n15608, n15609, n15610,
n15612, n15613, n15614, n15615, n15617, n15618, n15619, n15620,
n15622, n15623, n15624, n15625, n15627, n15628, n15629, n15630,
n15632, n15633, n15634, n15635, n15637, n15638, n15639, n15640,
n15642, n15643, n15644, n15645, n15647, n15648, n15649, n15650,
n15652, n15653, n15654, n15655, n15657, n15658, n15659, n15660,
n15662, n15663, n15664, n15665, n15667, n15668, n15669, n15670,
n15672, n15673, n15674, n15675, n15677, n15678, n15679, n15680,
n15682, n15683, n15684, n15685, n15687, n15688, n15689, n15690,
n15692, n15693, n15694, n15695, n15697, n15698, n15699, n15700,
n15702, n15703, n15704, n15705, n15707, n15708, n15709, n15710,
n15712, n15713, n15714, n15715, n15717, n15718, n15719, n15720,
n15722, n15723, n15724, n15725, n15727, n15728, n15729, n15730,
n15732, n15733, n15734, n15735, n15737, n15738, n15739, n15740,
n15742, n15743, n15744, n15745, n15747, n15748, n15749, n15750,
n15752, n15753, n15754, n15755, n15757, n15758, n15759, n15760,
n15762, n15763, n15764, n15765, n15767, n15768, n15769, n15770,
n15772, n15773, n15774, n15775, n15777, n15778, n15779, n15780,
n15782, n15783, n15784, n15785, n15787, n15788, n15789, n15790,
n15792, n15793, n15794, n15795, n15797, n15798, n15799, n15800,
n15802, n15803, n15804, n15805, n15807, n15808, n15809, n15810,
n15812, n15813, n15814, n15815, n15817, n15818, n15819, n15820,
n15822, n15823, n15824, n15825, n15827, n15828, n15829, n15830,
n15832, n15833, n15834, n15835, n15837, n15838, n15839, n15840,
n15842, n15843, n15844, n15845, n15847, n15848, n15849, n15850,
n15852, n15853, n15854, n15855, n15857, n15858, n15859, n15860,
n15862, n15863, n15864, n15865, n15867, n15868, n15869, n15870,
n15872, n15873, n15874, n15875, n15877, n15878, n15879, n15880,
n15882, n15883, n15884, n15885, n15887, n15888, n15889, n15890,
n15892, n15893, n15894, n15895, n15897, n15898, n15899, n15900,
n15902, n15903, n15904, n15905, n15907, n15908, n15909, n15910,
n15912, n15913, n15914, n15915, n15917, n15918, n15919, n15920,
n15922, n15923, n15924, n15925, n15927, n15928, n15929, n15930,
n15932, n15933, n15934, n15935, n15937, n15938, n15939, n15940,
n15942, n15943, n15944, n15945, n15947, n15948, n15949, n15950,
n15952, n15953, n15954, n15955, n15957, n15958, n15959, n15960,
n15962, n15963, n15964, n15965, n15967, n15968, n15969, n15970,
n15972, n15973, n15974, n15975, n15977, n15978, n15979, n15980,
n15982, n15983, n15984, n15985, n15987, n15988, n15989, n15990,
n15992, n15993, n15994, n15995, n15997, n15998, n15999, n16000,
n16002, n16003, n16004, n16005, n16007, n16008, n16009, n16010,
n16012, n16013, n16014, n16015, n16017, n16018, n16019, n16020,
n16022, n16023, n16024, n16025, n16027, n16028, n16029, n16030,
n16032, n16033, n16034, n16035, n16037, n16038, n16039, n16040,
n16042, n16043, n16044, n16045, n16047, n16048, n16049, n16050,
n16052, n16053, n16054, n16055, n16057, n16058, n16059, n16060,
n16062, n16063, n16064, n16065, n16067, n16068, n16069, n16070,
n16072, n16073, n16074, n16075, n16077, n16078, n16079, n16080,
n16082, n16083, n16084, n16085, n16087, n16088, n16089, n16090,
n16092, n16093, n16094, n16095, n16097, n16098, n16099, n16100,
n16102, n16103, n16104, n16105, n16107, n16108, n16109, n16110,
n16112, n16113, n16114, n16115, n16117, n16118, n16119, n16120,
n16122, n16123, n16124, n16125, n16127, n16128, n16129, n16130,
n16132, n16133, n16134, n16135, n16137, n16138, n16139, n16140,
n16142, n16143, n16144, n16145, n16147, n16148, n16149, n16150,
n16152, n16153, n16154, n16155, n16157, n16158, n16159, n16160,
n16162, n16163, n16164, n16165, n16167, n16168, n16169, n16170,
n16172, n16173, n16174, n16175, n16177, n16178, n16179, n16180,
n16182, n16183, n16184, n16185, n16187, n16188, n16189, n16190,
n16192, n16193, n16194, n16195, n16197, n16198, n16199, n16200,
n16202, n16203, n16204, n16205, n16207, n16208, n16209, n16210,
n16212, n16213, n16214, n16215, n16217, n16218, n16219, n16220,
n16222, n16223, n16224, n16225, n16227, n16228, n16229, n16230,
n16232, n16233, n16234, n16235, n16237, n16238, n16239, n16240,
n16242, n16243, n16244, n16245, n16247, n16248, n16249, n16250,
n16252, n16253, n16254, n16255, n16257, n16258, n16259, n16260,
n16262, n16263, n16264, n16265, n16267, n16268, n16269, n16270,
n16272, n16273, n16274, n16275, n16277, n16278, n16279, n16280,
n16282, n16283, n16284, n16285, n16287, n16288, n16289, n16290,
n16292, n16293, n16294, n16295, n16297, n16298, n16299, n16300,
n16302, n16303, n16304, n16305, n16307, n16308, n16309, n16310,
n16312, n16313, n16314, n16315, n16317, n16318, n16319, n16320,
n16321, n16322, n16323, n16324, n16325, n16327, n16328, n16329,
n16330, n16332, n16333, n16334, n16335, n16337, n16338, n16339,
n16340, n16342, n16343, n16344, n16345, n16347, n16348, n16349,
n16350, n16352, n16353, n16354, n16355, n16357, n16358, n16359,
n16360, n16362, n16363, n16364, n16365, n16367, n16368, n16369,
n16370, n16372, n16373, n16374, n16375, n16377, n16378, n16379,
n16380, n16382, n16383, n16384, n16385, n16387, n16388, n16389,
n16390, n16392, n16393, n16394, n16395, n16397, n16398, n16399,
n16400, n16402, n16403, n16404, n16405, n16407, n16408, n16409,
n16410, n16412, n16413, n16414, n16415, n16417, n16418, n16419,
n16420, n16422, n16423, n16424, n16425, n16427, n16428, n16429,
n16430, n16432, n16433, n16434, n16435, n16437, n16438, n16439,
n16440, n16442, n16443, n16444, n16445, n16447, n16448, n16449,
n16450, n16452, n16453, n16454, n16455, n16457, n16458, n16459,
n16460, n16462, n16463, n16464, n16465, n16467, n16468, n16469,
n16470, n16472, n16473, n16474, n16475, n16477, n16478, n16479,
n16480, n16482, n16483, n16484, n16485, n16487, n16488, n16489,
n16490, n16493, n16494, n16495, n16497, n16498, n16499, n16500,
n16502, n16503, n16504, n16505, n16507, n16508, n16509, n16510,
n16512, n16513, n16514, n16515, n16517, n16518, n16519, n16520,
n16522, n16523, n16524, n16525, n16527, n16528, n16529, n16530,
n16532, n16533, n16534, n16535, n16537, n16538, n16539, n16540,
n16542, n16543, n16544, n16545, n16547, n16548, n16549, n16550,
n16552, n16553, n16554, n16555, n16557, n16558, n16559, n16560,
n16562, n16563, n16564, n16565, n16567, n16568, n16569, n16570,
n16572, n16573, n16574, n16575, n16577, n16578, n16579, n16580,
n16582, n16583, n16584, n16585, n16587, n16588, n16589, n16590,
n16592, n16593, n16594, n16595, n16597, n16598, n16599, n16600,
n16602, n16603, n16604, n16605, n16607, n16608, n16609, n16610,
n16612, n16613, n16614, n16615, n16617, n16618, n16619, n16620,
n16622, n16623, n16624, n16625, n16627, n16628, n16629, n16630,
n16632, n16633, n16634, n16635, n16637, n16638, n16639, n16640,
n16642, n16643, n16644, n16645, n16647, n16648, n16649, n16650,
n16652, n16653, n16654, n16655, n16657, n16658, n16659, n16660,
n16662, n16663, n16664, n16665, n16667, n16668, n16669, n16670,
n16672, n16673, n16674, n16675, n16677, n16678, n16679, n16680,
n16682, n16683, n16684, n16685, n16687, n16688, n16689, n16690,
n16692, n16693, n16694, n16695, n16697, n16698, n16699, n16700,
n16702, n16703, n16704, n16705, n16707, n16708, n16709, n16710,
n16712, n16713, n16714, n16715, n16717, n16718, n16719, n16720,
n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
n17393, n17394, n17395, n17398, n17399, n17400, n17401, n17402,
n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
n17956, n17957, n17959, n17960, n17961, n17962, n17963, n17964,
n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
n18333, n18334, n18335, n18336, n18337, n18338, n18340, n18341,
n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19295,
n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
n20649, n20650, n20651, n20652, n20653, n20655, n20656, n20657,
n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
n21090, n21091, n21093, n21094, n21095, n21096, n21097, n21098,
n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21107,
n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
n21596, n21597, n21598, n21599, n21600, n21601, n21603, n21604,
n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
n21677, n21678, n21679, n21681, n21682, n21683, n21684, n21685,
n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813,
n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
n21863, n21864, n21865, n21866, n21868, n21869, n21870, n21871,
n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
n22080, n22081, n22082, n22083, n22085, n22086, n22087, n22088,
n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
n22129, n22130, n22131, n22132, n22133, n22134, n22136, n22137,
n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
n22234, n22235, n22236, n22237, n22239, n22240, n22241, n22242,
n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
n22691, n22692, n22693, n22696, n22697, n22698, n22699, n22700,
n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764,
n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22789,
n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797,
n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813,
n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837,
n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845,
n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853,
n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861,
n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877,
n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885,
n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893,
n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909,
n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917,
n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941,
n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965,
n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989,
n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037,
n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053,
n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061,
n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077,
n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085,
n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093,
n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102,
n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110,
n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118,
n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
n23129, n23130, n23133, n23134, n23135, n23136, n23139, n23140,
n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148,
n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156,
n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164,
n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172,
n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196,
n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
n23205, n23206, n23207, n23209, n23210, n23211, n23212, n23213,
n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229,
n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237,
n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245,
n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261,
n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277,
n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301,
n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309,
n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325,
n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333,
n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357,
n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373,
n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381,
n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389,
n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397,
n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405,
n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429,
n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445,
n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461,
n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501,
n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517,
n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533,
n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549,
n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589,
n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621,
n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661,
n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733,
n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805,
n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853,
n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877,
n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901,
n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909,
n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949,
n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021,
n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045,
n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053,
n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069,
n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093,
n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117,
n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125,
n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141,
n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165,
n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173,
n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189,
n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213,
n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221,
n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229,
n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237,
n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253,
n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261,
n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285,
n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293,
n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301,
n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309,
n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325,
n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333,
n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341,
n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357,
n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365,
n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373,
n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381,
n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405,
n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429,
n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437,
n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477,
n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501,
n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509,
n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525,
n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549,
n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573,
n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581,
n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597,
n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613,
n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621,
n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629,
n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645,
n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653,
n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669,
n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685,
n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693,
n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701,
n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
n24710, n24711, n24712, n24713, n24714, n24716, n24717, n24718,
n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726,
n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734,
n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758,
n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766,
n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774,
n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782,
n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798,
n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806,
n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846,
n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870,
n24871, n24872, n24873, n24875, n24876, n24877, n24878, n24879,
n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
n24936, n24937, n24938, n24939, n24940, n24942, n24943, n24944,
n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960,
n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
n25411, n25412, n25413, n25414, n25415, n25418, n25419, n25420,
n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428,
n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436,
n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452,
n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468,
n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476,
n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484,
n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500,
n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508,
n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524,
n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540,
n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548,
n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556,
n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572,
n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580,
n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612,
n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620,
n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644,
n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652,
n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660,
n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668,
n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684,
n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692,
n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716,
n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724,
n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740,
n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756,
n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764,
n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780,
n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788,
n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796,
n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812,
n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828,
n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836,
n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844,
n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860,
n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876,
n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884,
n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900,
n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908,
n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916,
n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924,
n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932,
n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956,
n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980,
n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988,
n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004,
n26005, n26006, n26008, n26009, n26010, n26011, n26012, n26013,
n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021,
n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037,
n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055,
n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079,
n26080, n26081, n26082, n26083, n26084, n26085, n26087, n26088,
n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
n26233, n26234, n26235, n26236, n26237, n26239, n26240, n26241,
n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
n26330, n26331, n26332, n26333, n26334, n26335, n26337, n26338,
n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
n26699, n26700, n26701, n26702, n26703, n26704, n26707, n26708,
n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732,
n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804,
n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820,
n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836,
n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844,
n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852,
n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916,
n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940,
n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948,
n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964,
n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980,
n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988,
n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012,
n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020,
n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036,
n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084,
n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092,
n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108,
n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124,
n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156,
n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204,
n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220,
n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228,
n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236,
n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252,
n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268,
n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276,
n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292,
n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308,
n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324,
n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340,
n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348,
n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380,
n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412,
n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420,
n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452,
n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468,
n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508,
n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540,
n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572,
n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588,
n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660,
n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668,
n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684,
n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708,
n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732,
n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740,
n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756,
n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780,
n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788,
n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804,
n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812,
n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852,
n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868,
n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876,
n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884,
n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916,
n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020,
n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028,
n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068,
n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092,
n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100,
n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156,
n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164,
n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172,
n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228,
n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244,
n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292,
n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300,
n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308,
n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316,
n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332,
n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340,
n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356,
n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364,
n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372,
n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380,
n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388,
n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404,
n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428,
n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436,
n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444,
n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452,
n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460,
n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468,
n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476,
n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500,
n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508,
n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516,
n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524,
n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532,
n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540,
n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548,
n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572,
n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580,
n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596,
n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604,
n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620,
n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644,
n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668,
n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684,
n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692,
n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708,
n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716,
n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724,
n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732,
n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740,
n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748,
n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764,
n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780,
n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788,
n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796,
n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804,
n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812,
n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820,
n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828,
n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852,
n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860,
n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868,
n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876,
n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884,
n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892,
n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900,
n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28909,
n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917,
n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925,
n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933,
n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941,
n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949,
n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957,
n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965,
n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973,
n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981,
n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
n28990, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006,
n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014,
n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022,
n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030,
n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038,
n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046,
n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054,
n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086,
n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094,
n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102,
n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118,
n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126,
n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142,
n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150,
n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158,
n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166,
n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182,
n29183, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247,
n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263,
n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271,
n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279,
n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327,
n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343,
n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383,
n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391,
n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399,
n29400, n29401, n29402, n29404, n29405, n29406, n29407, n29408,
n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416,
n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424,
n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432,
n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448,
n29449, n29450, n29451, n29452, n29453, n29455, n29456, n29457,
n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
n29554, n29556, n29557, n29558, n29559, n29560, n29561, n29562,
n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578,
n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610,
n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642,
n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666,
n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682,
n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706,
n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722,
n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730,
n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738,
n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754,
n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802,
n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810,
n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826,
n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842,
n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850,
n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858,
n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874,
n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882,
n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898,
n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914,
n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922,
n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930,
n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938,
n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946,
n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954,
n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970,
n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986,
n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994,
n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002,
n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
n30011, n30012, n30013, n30014, n30015, n30016, n30019, n30020,
n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028,
n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036,
n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044,
n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052,
n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060,
n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068,
n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076,
n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084,
n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092,
n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100,
n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108,
n30109, n30110, n30111, n30112, n30114, n30115, n30116, n30117,
n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125,
n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141,
n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149,
n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157,
n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165,
n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173,
n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181,
n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189,
n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197,
n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205,
n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213,
n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221,
n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229,
n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237,
n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245,
n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253,
n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261,
n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269,
n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285,
n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293,
n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301,
n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309,
n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317,
n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325,
n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333,
n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341,
n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349,
n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357,
n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365,
n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373,
n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381,
n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389,
n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397,
n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405,
n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413,
n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421,
n30422, n30423, n30424, n30426, n30427, n30428, n30429, n30430,
n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438,
n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
n30455, n30456, n30457, n30460, n30461, n30464, n30465, n30466,
n30467, n30470, n30471, n30472, n30473, n30474, n30475, n30476,
n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492,
n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500,
n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508,
n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516,
n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524,
n30525, n30526, n30527, n30528, n30531, n30532, n30534, n30535,
n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543,
n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551,
n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559,
n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567,
n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575,
n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591,
n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599,
n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607,
n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615,
n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623,
n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639,
n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647,
n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663,
n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671,
n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679,
n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687,
n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695,
n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711,
n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719,
n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735,
n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743,
n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751,
n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759,
n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775,
n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783,
n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791,
n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807,
n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823,
n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831,
n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839,
n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855,
n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863,
n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879,
n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887,
n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895,
n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903,
n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911,
n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919,
n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927,
n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935,
n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951,
n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959,
n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967,
n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975,
n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983,
n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991,
n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999,
n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007,
n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015,
n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023,
n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031,
n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039,
n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047,
n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055,
n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063,
n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071,
n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079,
n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087,
n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095,
n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103,
n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119,
n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127,
n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143,
n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151,
n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159,
n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167,
n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175,
n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183,
n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191,
n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199,
n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207,
n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215,
n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223,
n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231,
n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239,
n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263,
n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271,
n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287,
n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295,
n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303,
n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311,
n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327,
n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335,
n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343,
n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351,
n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359,
n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367,
n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383,
n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399,
n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407,
n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415,
n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423,
n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431,
n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439,
n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455,
n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471,
n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479,
n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487,
n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503,
n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511,
n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527,
n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543,
n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551,
n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559,
n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567,
n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575,
n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583,
n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599,
n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615,
n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623,
n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631,
n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639,
n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647,
n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655,
n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663,
n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671,
n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687,
n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695,
n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711,
n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727,
n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735,
n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743,
n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759,
n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767,
n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775,
n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791,
n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799,
n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807,
n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815,
n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823,
n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831,
n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855,
n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863,
n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871,
n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887,
n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895,
n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903,
n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911,
n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
n31920, n31921, n31922, n31923, n31924, n31926, n31927, n31928,
n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936,
n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944,
n31945, n31946, n31948, n31949, n31950, n31951, n31952, n31953,
n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130,
n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162,
n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170,
n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187,
n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195,
n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211,
n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227,
n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
n32252, n32253, n32255, n32256, n32257, n32258, n32259, n32260,
n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268,
n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276,
n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292,
n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300,
n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316,
n32317, n32318, n32320, n32321, n32322, n32323, n32324, n32325,
n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333,
n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341,
n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349,
n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357,
n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365,
n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373,
n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381,
n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389,
n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397,
n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405,
n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413,
n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421,
n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429,
n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437,
n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445,
n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453,
n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461,
n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469,
n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477,
n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485,
n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493,
n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501,
n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509,
n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517,
n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525,
n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533,
n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541,
n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549,
n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557,
n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565,
n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573,
n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581,
n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589,
n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597,
n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605,
n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613,
n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621,
n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629,
n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637,
n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645,
n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653,
n32654, n32655, n32658, n32659, n32660, n32661, n32662, n32663,
n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671,
n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679,
n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687,
n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695,
n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703,
n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711,
n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719,
n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727,
n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735,
n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743,
n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751,
n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759,
n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767,
n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775,
n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783,
n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791,
n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799,
n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807,
n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815,
n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823,
n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831,
n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839,
n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847,
n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855,
n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863,
n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871,
n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879,
n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887,
n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895,
n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911,
n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919,
n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927,
n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935,
n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943,
n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951,
n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959,
n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967,
n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975,
n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983,
n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991,
n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999,
n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007,
n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015,
n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023,
n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031,
n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039,
n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055,
n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063,
n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071,
n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079,
n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087,
n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095,
n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103,
n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111,
n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119,
n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127,
n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135,
n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143,
n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151,
n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159,
n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167,
n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175,
n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183,
n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199,
n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207,
n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215,
n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223,
n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231,
n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239,
n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
n33248, n33249, n33250, n33252, n33253, n33254, n33255, n33256,
n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264,
n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272,
n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280,
n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288,
n33289, n33292, n33293, n33294, n33295, n33296, n33297, n33298,
n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306,
n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314,
n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
n33323, n33324, n33326, n33327, n33328, n33329, n33330, n33331,
n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348,
n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372,
n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388,
n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396,
n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412,
n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420,
n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428,
n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444,
n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460,
n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468,
n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476,
n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484,
n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492,
n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500,
n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508,
n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516,
n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532,
n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540,
n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548,
n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556,
n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564,
n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572,
n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580,
n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589,
n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597,
n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605,
n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613,
n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621,
n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629,
n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637,
n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645,
n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653,
n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661,
n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669,
n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677,
n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685,
n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693,
n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701,
n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709,
n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717,
n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725,
n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733,
n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741,
n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749,
n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757,
n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765,
n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773,
n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781,
n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789,
n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797,
n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805,
n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813,
n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821,
n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829,
n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837,
n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845,
n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853,
n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861,
n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869,
n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877,
n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885,
n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893,
n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901,
n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909,
n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917,
n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925,
n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933,
n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941,
n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949,
n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959,
n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967,
n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975,
n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983,
n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991,
n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999,
n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007,
n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015,
n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023,
n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031,
n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039,
n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047,
n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055,
n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063,
n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071,
n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079,
n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087,
n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095,
n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103,
n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111,
n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119,
n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127,
n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135,
n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143,
n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151,
n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159,
n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167,
n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175,
n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183,
n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191,
n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199,
n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207,
n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215,
n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223,
n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231,
n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239,
n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247,
n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255,
n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263,
n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271,
n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279,
n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287,
n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295,
n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303,
n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311,
n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319,
n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335,
n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343,
n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351,
n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359,
n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367,
n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375,
n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383,
n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391,
n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399,
n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407,
n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415,
n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423,
n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431,
n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439,
n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447,
n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455,
n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463,
n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471,
n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479,
n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487,
n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495,
n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503,
n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511,
n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519,
n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527,
n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535,
n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543,
n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551,
n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567,
n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575,
n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583,
n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591,
n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599,
n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607,
n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615,
n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623,
n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639,
n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647,
n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655,
n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663,
n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671,
n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679,
n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687,
n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695,
n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711,
n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719,
n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727,
n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735,
n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743,
n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751,
n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759,
n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767,
n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775,
n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783,
n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791,
n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799,
n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807,
n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815,
n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823,
n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831,
n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839,
n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855,
n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863,
n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871,
n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879,
n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887,
n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895,
n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903,
n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911,
n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919,
n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927,
n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935,
n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943,
n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951,
n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959,
n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967,
n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975,
n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983,
n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991,
n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999,
n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007,
n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015,
n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023,
n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031,
n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039,
n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047,
n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055,
n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063,
n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071,
n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079,
n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087,
n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095,
n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103,
n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111,
n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119,
n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127,
n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135,
n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143,
n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151,
n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159,
n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167,
n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175,
n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183,
n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191,
n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199,
n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207,
n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215,
n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223,
n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231,
n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239,
n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247,
n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255,
n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263,
n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271,
n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279,
n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287,
n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295,
n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303,
n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311,
n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319,
n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327,
n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335,
n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343,
n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351,
n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359,
n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367,
n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375,
n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383,
n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391,
n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399,
n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407,
n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415,
n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423,
n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431,
n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439,
n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447,
n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455,
n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463,
n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471,
n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479,
n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487,
n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495,
n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503,
n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511,
n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519,
n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527,
n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535,
n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543,
n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551,
n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559,
n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567,
n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575,
n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583,
n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591,
n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599,
n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607,
n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615,
n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623,
n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631,
n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639,
n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647,
n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655,
n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663,
n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671,
n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679,
n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687,
n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695,
n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703,
n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711,
n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719,
n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727,
n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735,
n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743,
n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751,
n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759,
n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775,
n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783,
n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791,
n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799,
n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807,
n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815,
n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823,
n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831,
n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839,
n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847,
n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855,
n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863,
n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871,
n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879,
n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887,
n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895,
n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911,
n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919,
n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927,
n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935,
n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943,
n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951,
n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959,
n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967,
n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975,
n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983,
n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991,
n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999,
n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007,
n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015,
n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023,
n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031,
n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039,
n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047,
n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055,
n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063,
n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071,
n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079,
n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36088,
n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096,
n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104,
n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112,
n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120,
n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128,
n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144,
n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160,
n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168,
n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176,
n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184,
n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192,
n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200,
n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208,
n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216,
n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232,
n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240,
n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248,
n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256,
n36257, n36258, n36259, n36260, n36261, n36263, n36264, n36265,
n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
n36546, n36548, n36549, n36550, n36551, n36552, n36553, n36554,
n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562,
n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570,
n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578,
n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594,
n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602,
n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618,
n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626,
n36627, n36629, n36630, n36631, n36632, n36633, n36634, n36635,
n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651,
n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659,
n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691,
n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699,
n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707,
n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715,
n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723,
n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731,
n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763,
n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771,
n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787,
n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795,
n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803,
n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835,
n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843,
n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852,
n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860,
n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868,
n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876,
n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884,
n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892,
n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900,
n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908,
n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916,
n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924,
n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932,
n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940,
n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948,
n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956,
n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964,
n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972,
n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980,
n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988,
n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996,
n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004,
n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012,
n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020,
n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028,
n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036,
n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044,
n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052,
n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060,
n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068,
n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076,
n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084,
n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092,
n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100,
n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108,
n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116,
n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124,
n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132,
n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140,
n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148,
n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156,
n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164,
n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172,
n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180,
n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188,
n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196,
n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204,
n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212,
n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220,
n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228,
n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236,
n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244,
n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252,
n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260,
n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268,
n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276,
n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284,
n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292,
n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300,
n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308,
n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316,
n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324,
n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332,
n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340,
n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348,
n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356,
n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364,
n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372,
n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380,
n37381, n37382, n37383, n37384, n37385, n37386, n37387, n37388,
n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396,
n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404,
n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412,
n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420,
n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428,
n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436,
n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444,
n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452,
n37453, n37454, n37455, n37456, n37457, n37458, n37459, n37460,
n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468,
n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476,
n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484,
n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492,
n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500,
n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508,
n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516,
n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524,
n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532,
n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540,
n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548,
n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556,
n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564,
n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572,
n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580,
n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588,
n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596,
n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604,
n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612,
n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620,
n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628,
n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636,
n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644,
n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652,
n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660,
n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668,
n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676,
n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684,
n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692,
n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700,
n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708,
n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716,
n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724,
n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732,
n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740,
n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748,
n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756,
n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764,
n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772,
n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780,
n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788,
n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796,
n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804,
n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812,
n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820,
n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828,
n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836,
n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844,
n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852,
n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860,
n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868,
n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876,
n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884,
n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892,
n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900,
n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908,
n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916,
n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924,
n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932,
n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940,
n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948,
n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956,
n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964,
n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972,
n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980,
n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988,
n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996,
n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004,
n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012,
n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020,
n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028,
n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036,
n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044,
n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052,
n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060,
n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068,
n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076,
n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084,
n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092,
n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100,
n38101, n38102, n38103, n38104, n38105, n38106, n38107, n38108,
n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116,
n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124,
n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132,
n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140,
n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148,
n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156,
n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164,
n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172,
n38173, n38174, n38175, n38176, n38177, n38178, n38179, n38180,
n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188,
n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196,
n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204,
n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212,
n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220,
n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228,
n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236,
n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244,
n38245, n38246, n38247, n38248, n38249, n38250, n38251, n38252,
n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260,
n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268,
n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276,
n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284,
n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292,
n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300,
n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308,
n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316,
n38317, n38318, n38319, n38320, n38321, n38322, n38323, n38324,
n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332,
n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340,
n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348,
n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356,
n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364,
n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372,
n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380,
n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388,
n38389, n38390, n38391, n38392, n38393, n38394, n38395, n38396,
n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404,
n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412,
n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420,
n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428,
n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436,
n38437, n38438, n38439, n38440, n38441, n38442, n38443, n38444,
n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452,
n38453, n38454, n38455, n38456, n38457, n38458, n38459, n38460,
n38461, n38462, n38463, n38464, n38465, n38466, n38467, n38468,
n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476,
n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484,
n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492,
n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500,
n38501, n38502, n38503, n38504, n38505, n38506, n38507, n38508,
n38509, n38510, n38511, n38512, n38513, n38514, n38515, n38516,
n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524,
n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532,
n38533, n38534, n38535, n38536, n38537, n38538, n38539, n38540,
n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548,
n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556,
n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564,
n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572,
n38573, n38574, n38575, n38576, n38577, n38578, n38579, n38580,
n38581, n38582, n38583, n38584, n38585, n38586, n38587, n38588,
n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596,
n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604,
n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612,
n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620,
n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628,
n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636,
n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644,
n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652,
n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660,
n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668,
n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676,
n38677, n38678, n38679, n38680, n38681, n38682, n38683, n38684,
n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692,
n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700,
n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708,
n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716,
n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724,
n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732,
n38733, n38734, n38735, n38736, n38737, n38739, n38740, n38741,
n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749,
n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757,
n38758, n38759, n38760, n38761, n38762, n38763, n38764, n38765,
n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773,
n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781,
n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789,
n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797,
n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805,
n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813,
n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821,
n38822, n38824, n38825, n38826, n38827, n38828, n38829, n38830,
n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838,
n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846,
n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862,
n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878,
n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886,
n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894,
n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902,
n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910,
n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918,
n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934,
n38935, n38936, n38937, n38938, n38941, n38942, n38943, n38944,
n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952,
n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960,
n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976,
n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984,
n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992,
n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000,
n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008,
n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024,
n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040,
n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048,
n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056,
n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064,
n39065, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082,
n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090,
n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114,
n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138,
n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154,
n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162,
n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170,
n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188,
n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196,
n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204,
n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212,
n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220,
n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39229,
n39230, n39231, n39232, n39233, n39234, n39235, n39236, n39237,
n39238, n39239, n39240, n39241, n39242, n39243, n39244, n39245,
n39246, n39247, n39248, n39249, n39250, n39251, n39252, n39253,
n39254, n39255, n39256, n39257, n39258, n39259, n39260, n39261,
n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269,
n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277,
n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285,
n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293,
n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301,
n39302, n39303, n39304, n39305, n39306, n39307, n39308, n39309,
n39310, n39311, n39312, n39313, n39314, n39315, n39316, n39317,
n39318, n39319, n39320, n39321, n39322, n39323, n39324, n39325,
n39326, n39327, n39328, n39329, n39330, n39331, n39332, n39333,
n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341,
n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349,
n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357,
n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365,
n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373,
n39374, n39375, n39376, n39377, n39378, n39379, n39380, n39381,
n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389,
n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397,
n39398, n39399, n39400, n39401, n39402, n39403, n39404, n39405,
n39406, n39407, n39408, n39409, n39410, n39411, n39412, n39413,
n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39423,
n39424, n39425, n39426, n39429, n39430, n39431, n39432, n39433,
n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
n39466, n39467, n39470, n39471, n39472, n39473, n39474, n39475,
n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483,
n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491,
n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499,
n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507,
n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523,
n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531,
n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539,
n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547,
n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555,
n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571,
n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579,
n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595,
n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603,
n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611,
n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619,
n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627,
n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635,
n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643,
n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39652,
n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660,
n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668,
n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676,
n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684,
n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692,
n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700,
n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708,
n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716,
n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724,
n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39734,
n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750,
n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758,
n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766,
n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774,
n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782,
n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790,
n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798,
n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806,
n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814,
n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822,
n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830,
n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838,
n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846,
n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854,
n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862,
n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870,
n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878,
n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886,
n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894,
n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910,
n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918,
n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926,
n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
n39935, n39936, n39937, n39938, n39940, n39941, n39942, n39943,
n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951,
n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959,
n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967,
n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975,
n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983,
n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991,
n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999,
n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007,
n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015,
n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023,
n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031,
n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039,
n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047,
n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055,
n40056, n40057, n40058, n40059, n40061, n40062, n40063, n40064,
n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072,
n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080,
n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088,
n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128,
n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136,
n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144,
n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152,
n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160,
n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192,
n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200,
n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208,
n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216,
n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224,
n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232,
n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248,
n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264,
n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272,
n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288,
n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296,
n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304,
n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320,
n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336,
n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344,
n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352,
n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360,
n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368,
n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376,
n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392,
n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408,
n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
n40417, n40418, n40419, n40420, n40421, n40423, n40424, n40425,
n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
n40458, n40459, n40460, n40461, n40464, n40465, n40466, n40467,
n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475,
n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491,
n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499,
n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507,
n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515,
n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523,
n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531,
n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539,
n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547,
n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563,
n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587,
n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595,
n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603,
n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611,
n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619,
n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635,
n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659,
n40660, n40661, n40663, n40664, n40665, n40666, n40667, n40668,
n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676,
n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684,
n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40692,
n40693, n40694, n40695, n40696, n40697, n40698, n40699, n40700,
n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708,
n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716,
n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724,
n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732,
n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740,
n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748,
n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756,
n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764,
n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772,
n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780,
n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788,
n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796,
n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804,
n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812,
n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820,
n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40829,
n40830, n40831, n40832, n40833, n40834, n40835, n40836, n40837,
n40838, n40839, n40840, n40841, n40842, n40843, n40844, n40845,
n40846, n40847, n40848, n40849, n40850, n40851, n40852, n40853,
n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861,
n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869,
n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877,
n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885,
n40886, n40887, n40888, n40889, n40890, n40891, n40892, n40893,
n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901,
n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909,
n40910, n40911, n40912, n40913, n40914, n40915, n40916, n40917,
n40918, n40919, n40920, n40921, n40922, n40923, n40924, n40925,
n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933,
n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941,
n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949,
n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957,
n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965,
n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973,
n40974, n40975, n40976, n40977, n40978, n40979, n40980, n40981,
n40982, n40983, n40984, n40985, n40986, n40987, n40988, n40989,
n40990, n40991, n40992, n40993, n40994, n40995, n40996, n40997,
n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005,
n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013,
n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021,
n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029,
n41030, n41031, n41032, n41033, n41034, n41035, n41036, n41037,
n41038, n41039, n41040, n41041, n41042, n41043, n41044, n41045,
n41046, n41047, n41048, n41049, n41050, n41051, n41052, n41053,
n41054, n41055, n41056, n41057, n41058, n41059, n41060, n41061,
n41062, n41063, n41064, n41065, n41066, n41067, n41068, n41069,
n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077,
n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085,
n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093,
n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101,
n41102, n41103, n41104, n41105, n41106, n41107, n41108, n41109,
n41110, n41111, n41112, n41113, n41114, n41115, n41116, n41117,
n41118, n41119, n41120, n41121, n41122, n41123, n41124, n41125,
n41126, n41127, n41128, n41129, n41130, n41131, n41132, n41133,
n41134, n41135, n41136, n41137, n41138, n41139, n41140, n41141,
n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149,
n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157,
n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165,
n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173,
n41174, n41175, n41176, n41177, n41178, n41179, n41180, n41181,
n41182, n41183, n41184, n41185, n41186, n41187, n41188, n41189,
n41190, n41191, n41192, n41193, n41194, n41195, n41196, n41197,
n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205,
n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213,
n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221,
n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229,
n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237,
n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245,
n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253,
n41254, n41255, n41256, n41257, n41258, n41259, n41260, n41261,
n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269,
n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277,
n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285,
n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293,
n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301,
n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309,
n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317,
n41318, n41319, n41320, n41321, n41322, n41323, n41324, n41325,
n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333,
n41334, n41335, n41336, n41337, n41338, n41339, n41340, n41341,
n41342, n41343, n41344, n41345, n41346, n41347, n41348, n41349,
n41350, n41351, n41352, n41353, n41354, n41355, n41356, n41357,
n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365,
n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373,
n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381,
n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389,
n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397,
n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405,
n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413,
n41414, n41415, n41416, n41417, n41418, n41419, n41420, n41421,
n41422, n41423, n41424, n41425, n41426, n41427, n41428, n41429,
n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437,
n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445,
n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453,
n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461,
n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469,
n41470, n41471, n41472, n41473, n41474, n41475, n41476, n41477,
n41478, n41479, n41480, n41481, n41482, n41483, n41484, n41485,
n41486, n41487, n41488, n41489, n41490, n41491, n41492, n41493,
n41494, n41495, n41496, n41497, n41498, n41499, n41500, n41501,
n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509,
n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517,
n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525,
n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533,
n41534, n41535, n41536, n41537, n41538, n41539, n41540, n41541,
n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549,
n41550, n41551, n41552, n41553, n41554, n41555, n41556, n41557,
n41558, n41559, n41560, n41561, n41562, n41563, n41564, n41565,
n41566, n41567, n41568, n41569, n41570, n41571, n41572, n41573,
n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581,
n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589,
n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597,
n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605,
n41606, n41607, n41608, n41609, n41610, n41611, n41612, n41613,
n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621,
n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629,
n41630, n41631, n41632, n41634, n41635, n41636, n41637, n41638,
n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646,
n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654,
n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662,
n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670,
n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678,
n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686,
n41687, n41689, n41690, n41691, n41692, n41693, n41694, n41695,
n41696, n41697, n41698, n41699, n41701, n41702, n41703, n41704,
n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712,
n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720,
n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728,
n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736,
n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744,
n41745, n41746, n41747, n41750, n41751, n41752, n41753, n41754,
n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762,
n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778,
n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794,
n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802,
n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818,
n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826,
n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850,
n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890,
n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898,
n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906,
n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922,
n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938,
n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946,
n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962,
n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970,
n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978,
n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994,
n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018,
n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026,
n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034,
n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042,
n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050,
n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066,
n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090,
n42091, n42092, n42093, n42095, n42096, n42097, n42098, n42099,
n42100, n42102, n42103, n42104, n42105, n42106, n42107, n42108,
n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116,
n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124,
n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132,
n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140,
n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148,
n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156,
n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164,
n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172,
n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180,
n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188,
n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196,
n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204,
n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212,
n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220,
n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228,
n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236,
n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244,
n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252,
n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260,
n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268,
n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276,
n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284,
n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292,
n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300,
n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308,
n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316,
n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324,
n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332,
n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340,
n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348,
n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356,
n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364,
n42365, n42367, n42368, n42369, n42370, n42371, n42372, n42373,
n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381,
n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389,
n42390, n42391, n42392, n42394, n42395, n42396, n42397, n42398,
n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406,
n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414,
n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422,
n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430,
n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438,
n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446,
n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454,
n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462,
n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478,
n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486,
n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494,
n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502,
n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510,
n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518,
n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42527,
n42528, n42529, n42530, n42531, n42532, n42533, n42534, n42535,
n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543,
n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551,
n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559,
n42560, n42561, n42562, n42563, n42564, n42565, n42566, n42567,
n42568, n42569, n42570, n42571, n42572, n42573, n42574, n42575,
n42576, n42577, n42578, n42579, n42580, n42581, n42582, n42583,
n42584, n42585, n42586, n42587, n42588, n42589, n42590, n42591,
n42592, n42593, n42594, n42595, n42596, n42597, n42598, n42599,
n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607,
n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615,
n42616, n42617, n42618, n42619, n42620, n42621, n42622, n42623,
n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631,
n42632, n42633, n42634, n42635, n42636, n42637, n42638, n42639,
n42640, n42641, n42642, n42643, n42644, n42645, n42646, n42647,
n42648, n42649, n42650, n42651, n42652, n42653, n42654, n42655,
n42656, n42657, n42658, n42659, n42660, n42661, n42662, n42663,
n42664, n42665, n42666, n42667, n42668, n42669, n42670, n42671,
n42672, n42673, n42674, n42675, n42676, n42677, n42678, n42679,
n42680, n42681, n42682, n42683, n42684, n42685, n42686, n42687,
n42688, n42689, n42690, n42691, n42692, n42693, n42694, n42695,
n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703,
n42704, n42705, n42706, n42707, n42708, n42709, n42710, n42711,
n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719,
n42720, n42721, n42722, n42723, n42724, n42725, n42726, n42727,
n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735,
n42736, n42737, n42738, n42739, n42740, n42741, n42742, n42743,
n42744, n42745, n42746, n42747, n42748, n42749, n42750, n42751,
n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759,
n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767,
n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775,
n42776, n42777, n42778, n42779, n42780, n42781, n42782, n42783,
n42784, n42785, n42786, n42787, n42788, n42789, n42790, n42791,
n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799,
n42800, n42801, n42802, n42803, n42804, n42805, n42806, n42807,
n42808, n42809, n42810, n42811, n42812, n42813, n42814, n42815,
n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823,
n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831,
n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42839,
n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847,
n42848, n42849, n42850, n42851, n42852, n42853, n42854, n42855,
n42856, n42857, n42858, n42859, n42860, n42861, n42862, n42863,
n42864, n42865, n42866, n42867, n42868, n42869, n42870, n42871,
n42872, n42873, n42874, n42875, n42876, n42877, n42878, n42879,
n42880, n42881, n42882, n42883, n42884, n42885, n42886, n42887,
n42888, n42889, n42890, n42891, n42892, n42893, n42894, n42895,
n42896, n42897, n42898, n42899, n42900, n42901, n42902, n42903,
n42904, n42905, n42906, n42907, n42908, n42909, n42910, n42911,
n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919,
n42920, n42921, n42922, n42923, n42924, n42925, n42926, n42927,
n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935,
n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943,
n42944, n42945, n42946, n42947, n42948, n42949, n42950, n42951,
n42952, n42953, n42954, n42955, n42956, n42957, n42958, n42959,
n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967,
n42968, n42969, n42970, n42971, n42972, n42973, n42974, n42975,
n42976, n42977, n42978, n42979, n42980, n42981, n42982, n42983,
n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991,
n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999,
n43000, n43001, n43002, n43003, n43004, n43005, n43006, n43007,
n43008, n43009, n43010, n43011, n43012, n43013, n43014, n43015,
n43016, n43017, n43018, n43019, n43020, n43021, n43022, n43023,
n43024, n43025, n43026, n43027, n43028, n43029, n43030, n43031,
n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43039,
n43040, n43041, n43042, n43043, n43044, n43045, n43046, n43047,
n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055,
n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063,
n43064, n43065, n43066, n43067, n43068, n43069, n43070, n43071,
n43072, n43073, n43074, n43075, n43076, n43077, n43078, n43079,
n43080, n43081, n43082, n43083, n43084, n43085, n43086, n43087,
n43088, n43089, n43090, n43091, n43092, n43093, n43094, n43095,
n43096, n43097, n43098, n43099, n43100, n43101, n43102, n43103,
n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111,
n43112, n43113, n43114, n43115, n43116, n43118, n43119, n43120,
n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128,
n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136,
n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144,
n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152,
n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160,
n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168,
n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176,
n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184,
n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192,
n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200,
n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208,
n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216,
n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224,
n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232,
n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240,
n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248,
n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256,
n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264,
n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272,
n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280,
n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43290,
n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306,
n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314,
n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330,
n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338,
n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346,
n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362,
n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378,
n43379, n43380, n43381, n43383, n43384, n43385, n43386, n43387,
n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395,
n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403,
n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411,
n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419,
n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427,
n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443,
n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459,
n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467,
n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475,
n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483,
n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491,
n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499,
n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515,
n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531,
n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539,
n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547,
n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555,
n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563,
n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571,
n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587,
n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603,
n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611,
n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619,
n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627,
n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635,
n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643,
n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659,
n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675,
n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683,
n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691,
n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699,
n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707,
n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715,
n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731,
n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747,
n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755,
n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763,
n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771,
n43772, n43773, n43776, n43777, n43780, n43781, n43782, n43783,
n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793,
n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801,
n43802, n43803, n43806, n43807, n43808, n43809, n43810, n43811,
n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819,
n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827,
n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835,
n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843,
n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851,
n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859,
n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875,
n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883,
n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891,
n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899,
n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907,
n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915,
n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923,
n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931,
n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947,
n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955,
n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963,
n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971,
n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979,
n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987,
n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995,
n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003,
n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011,
n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019,
n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027,
n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035,
n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043,
n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051,
n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059,
n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067,
n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075,
n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083,
n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091,
n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099,
n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107,
n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115,
n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123,
n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131,
n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139,
n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147,
n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163,
n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171,
n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179,
n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187,
n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195,
n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203,
n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211,
n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219,
n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227,
n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235,
n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243,
n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251,
n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259,
n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275,
n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283,
n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291,
n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299,
n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307,
n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315,
n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323,
n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331,
n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339,
n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347,
n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355,
n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363,
n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379,
n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395,
n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403,
n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411,
n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419,
n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427,
n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435,
n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443,
n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451,
n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459,
n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467,
n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475,
n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483,
n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491,
n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499,
n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507,
n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523,
n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531,
n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539,
n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547,
n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555,
n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563,
n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571,
n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579,
n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587,
n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595,
n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603,
n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611,
n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619,
n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627,
n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635,
n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643,
n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651,
n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659,
n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667,
n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683,
n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691,
n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707,
n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715,
n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723,
n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731,
n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739,
n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747,
n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755,
n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763,
n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771,
n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779,
n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787,
n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795,
n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803,
n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811,
n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819,
n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827,
n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835,
n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843,
n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851,
n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859,
n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867,
n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875,
n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883,
n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899,
n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907,
n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915,
n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923,
n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931,
n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939,
n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955,
n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963,
n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971,
n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979,
n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987,
n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995,
n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003,
n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011,
n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019,
n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027,
n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035,
n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043,
n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051,
n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059,
n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067,
n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075,
n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083,
n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091,
n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099,
n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107,
n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115,
n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123,
n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131,
n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139,
n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147,
n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155,
n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171,
n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179,
n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187,
n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195,
n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211,
n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219,
n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227,
n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235,
n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243,
n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251,
n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259,
n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267,
n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275,
n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283,
n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291,
n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299,
n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307,
n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315,
n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323,
n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331,
n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339,
n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347,
n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355,
n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363,
n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371,
n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379,
n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387,
n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395,
n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403,
n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411,
n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419,
n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427,
n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435,
n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443,
n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451,
n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459,
n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467,
n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475,
n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483,
n45484, n45485, n45486, n45487, n45488, n45491, n45492, n45493,
n45494, n45495, n45496, n45497, n45498, n45499, n45500, n45501,
n45502, n45503, n45504, n45505, n45506, n45507, n45508, n45509,
n45510, n45511, n45512, n45513, n45514, n45515, n45516, n45517,
n45518, n45519, n45520, n45521, n45522, n45523, n45524, n45525,
n45526, n45527, n45528, n45529, n45530, n45531, n45532, n45533,
n45534, n45535, n45536, n45537, n45538, n45539, n45540, n45541,
n45542, n45543, n45544, n45545, n45546, n45547, n45548, n45549,
n45550, n45551, n45552, n45553, n45554, n45555, n45556, n45557,
n45558, n45559, n45560, n45561, n45562, n45563, n45564, n45565,
n45566, n45567, n45568, n45569, n45570, n45571, n45572, n45573,
n45574, n45575, n45576, n45577, n45578, n45579, n45580, n45581,
n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589,
n45590, n45591, n45592, n45593, n45594, n45595, n45596, n45597,
n45598, n45599, n45600, n45601, n45602, n45603, n45604, n45605,
n45606, n45607, n45608, n45609, n45610, n45611, n45612, n45613,
n45614, n45615, n45616, n45617, n45618, n45619, n45620, n45621,
n45622, n45623, n45624, n45626, n45627, n45628, n45629, n45630,
n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638,
n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646,
n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654,
n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662,
n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670,
n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678,
n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686,
n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702,
n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710,
n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718,
n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726,
n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734,
n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742,
n45743, n45744, n45745, n45746, n45747, n45748, n45750, n45751,
n45752, n45753, n45754, n45755, n45756, n45757, n45758, n45759,
n45760, n45761, n45762, n45763, n45764, n45765, n45766, n45767,
n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775,
n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783,
n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791,
n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799,
n45800, n45802, n45803, n45804, n45805, n45806, n45807, n45808,
n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816,
n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824,
n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832,
n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840,
n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848,
n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856,
n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864,
n45865, n45867, n45868, n45869, n45870, n45871, n45872, n45873,
n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881,
n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889,
n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897,
n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905,
n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913,
n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921,
n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929,
n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937,
n45938, n45939, n45940, n45941, n45943, n45944, n45945, n45946,
n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954,
n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970,
n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978,
n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994,
n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002,
n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010,
n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46019,
n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027,
n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035,
n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043,
n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051,
n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059,
n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067,
n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075,
n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083,
n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091,
n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099,
n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107,
n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115,
n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123,
n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131,
n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139,
n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147,
n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155,
n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163,
n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171,
n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179,
n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195,
n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203,
n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211,
n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219,
n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227,
n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235,
n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243,
n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251,
n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259,
n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267,
n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275,
n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283,
n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291,
n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299,
n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307,
n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315,
n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323,
n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339,
n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347,
n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
n46356, n46359, n46360, n46361, n46362, n46363, n46364, n46365,
n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373,
n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381,
n46382, n46383, n46384, n46385, n46386, n46387, n46388, n46389,
n46390, n46391, n46392, n46393, n46394, n46395, n46396, n46397,
n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405,
n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413,
n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421,
n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429,
n46430, n46431, n46432, n46433, n46434, n46435, n46436, n46437,
n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445,
n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453,
n46454, n46455, n46456, n46457, n46458, n46459, n46460, n46461,
n46462, n46463, n46464, n46465, n46466, n46467, n46468, n46469,
n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477,
n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485,
n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493,
n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501,
n46502, n46503, n46504, n46505, n46506, n46507, n46508, n46509,
n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517,
n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525,
n46526, n46527, n46528, n46529, n46530, n46531, n46532, n46533,
n46534, n46535, n46536, n46537, n46538, n46539, n46540, n46541,
n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549,
n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557,
n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565,
n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573,
n46574, n46575, n46576, n46577, n46578, n46579, n46580, n46581,
n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589,
n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597,
n46598, n46599, n46600, n46601, n46602, n46603, n46604, n46605,
n46606, n46607, n46608, n46609, n46610, n46611, n46612, n46613,
n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621,
n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629,
n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637,
n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645,
n46646, n46647, n46648, n46649, n46650, n46651, n46652, n46653,
n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661,
n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669,
n46670, n46671, n46672, n46673, n46674, n46675, n46676, n46677,
n46678, n46679, n46680, n46681, n46682, n46683, n46684, n46685,
n46686, n46687, n46688, n46689, n46690, n46691, n46692, n46693,
n46694, n46695, n46696, n46697, n46698, n46699, n46700, n46701,
n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709,
n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717,
n46718, n46719, n46720, n46721, n46722, n46723, n46724, n46725,
n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733,
n46734, n46735, n46736, n46737, n46738, n46739, n46740, n46741,
n46742, n46743, n46744, n46745, n46746, n46747, n46748, n46749,
n46750, n46751, n46752, n46753, n46754, n46755, n46756, n46757,
n46758, n46759, n46760, n46761, n46762, n46763, n46764, n46765,
n46766, n46767, n46768, n46769, n46770, n46771, n46772, n46773,
n46774, n46775, n46776, n46777, n46778, n46779, n46780, n46781,
n46782, n46783, n46784, n46785, n46786, n46787, n46788, n46789,
n46790, n46791, n46792, n46793, n46794, n46795, n46796, n46797,
n46798, n46799, n46800, n46801, n46802, n46803, n46804, n46805,
n46806, n46807, n46808, n46809, n46810, n46811, n46812, n46813,
n46814, n46815, n46816, n46817, n46818, n46819, n46820, n46821,
n46822, n46823, n46824, n46825, n46826, n46827, n46828, n46829,
n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837,
n46838, n46839, n46840, n46841, n46842, n46843, n46844, n46845,
n46846, n46847, n46848, n46849, n46850, n46851, n46852, n46853,
n46854, n46855, n46856, n46857, n46858, n46859, n46860, n46861,
n46862, n46863, n46864, n46865, n46866, n46867, n46868, n46869,
n46870, n46871, n46872, n46873, n46874, n46875, n46876, n46877,
n46878, n46879, n46880, n46881, n46882, n46883, n46884, n46885,
n46886, n46887, n46888, n46889, n46890, n46891, n46892, n46893,
n46894, n46895, n46896, n46897, n46898, n46899, n46900, n46901,
n46902, n46903, n46904, n46905, n46906, n46907, n46908, n46909,
n46910, n46911, n46912, n46913, n46914, n46915, n46916, n46917,
n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925,
n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933,
n46934, n46935, n46936, n46937, n46938, n46939, n46940, n46941,
n46942, n46943, n46944, n46945, n46946, n46947, n46948, n46949,
n46950, n46951, n46952, n46953, n46954, n46955, n46956, n46957,
n46958, n46959, n46960, n46961, n46962, n46963, n46964, n46965,
n46966, n46967, n46968, n46969, n46970, n46971, n46972, n46973,
n46974, n46976, n46977, n46978, n46979, n46980, n46981, n46982,
n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990,
n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998,
n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006,
n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47016,
n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024,
n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032,
n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040,
n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048,
n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056,
n47057, n47059, n47060, n47061, n47062, n47063, n47064, n47065,
n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073,
n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081,
n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089,
n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097,
n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105,
n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113,
n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121,
n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129,
n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137,
n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145,
n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153,
n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161,
n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169,
n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177,
n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185,
n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193,
n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201,
n47202, n47203, n47204, n47205, n47206, n47207, n47209, n47210,
n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218,
n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226,
n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234,
n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250,
n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266,
n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274,
n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290,
n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298,
n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47307,
n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315,
n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323,
n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331,
n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339,
n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347,
n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355,
n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363,
n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371,
n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379,
n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387,
n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395,
n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403,
n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411,
n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419,
n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427,
n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435,
n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443,
n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451,
n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459,
n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467,
n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475,
n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483,
n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491,
n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499,
n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507,
n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515,
n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523,
n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531,
n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539,
n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547,
n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555,
n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563,
n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571,
n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579,
n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587,
n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595,
n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603,
n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611,
n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619,
n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627,
n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635,
n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643,
n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651,
n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659,
n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667,
n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675,
n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683,
n47684, n47687, n47688, n47689, n47690, n47691, n47692, n47693,
n47694, n47695, n47696, n47697, n47698, n47699, n47700, n47701,
n47702, n47703, n47704, n47705, n47706, n47707, n47708, n47709,
n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717,
n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725,
n47726, n47727, n47728, n47729, n47730, n47731, n47732, n47733,
n47734, n47735, n47736, n47737, n47738, n47739, n47740, n47741,
n47742, n47743, n47744, n47745, n47746, n47747, n47748, n47749,
n47750, n47751, n47752, n47753, n47754, n47755, n47756, n47757,
n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765,
n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773,
n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781,
n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789,
n47790, n47791, n47792, n47793, n47794, n47795, n47796, n47797,
n47798, n47799, n47800, n47801, n47802, n47803, n47804, n47805,
n47806, n47807, n47808, n47809, n47810, n47811, n47812, n47813,
n47814, n47815, n47816, n47817, n47818, n47819, n47820, n47821,
n47822, n47823, n47824, n47825, n47826, n47827, n47828, n47829,
n47830, n47831, n47832, n47833, n47834, n47835, n47836, n47837,
n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845,
n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853,
n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861,
n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869,
n47870, n47871, n47872, n47873, n47874, n47875, n47876, n47877,
n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885,
n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47893,
n47894, n47895, n47896, n47897, n47898, n47899, n47900, n47901,
n47902, n47903, n47904, n47905, n47906, n47907, n47908, n47909,
n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917,
n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925,
n47926, n47927, n47928, n47929, n47930, n47931, n47932, n47933,
n47934, n47935, n47936, n47937, n47938, n47939, n47940, n47941,
n47942, n47943, n47944, n47945, n47946, n47947, n47948, n47949,
n47950, n47951, n47952, n47953, n47954, n47955, n47956, n47957,
n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965,
n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973,
n47974, n47975, n47976, n47977, n47978, n47979, n47980, n47981,
n47982, n47983, n47984, n47985, n47986, n47987, n47988, n47989,
n47990, n47991, n47992, n47993, n47994, n47995, n47996, n47997,
n47998, n47999, n48000, n48001, n48002, n48003, n48004, n48005,
n48006, n48007, n48008, n48009, n48010, n48011, n48012, n48013,
n48014, n48015, n48016, n48017, n48018, n48019, n48020, n48021,
n48022, n48023, n48024, n48025, n48026, n48027, n48028, n48029,
n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037,
n48038, n48039, n48040, n48041, n48042, n48043, n48044, n48045,
n48046, n48047, n48048, n48049, n48050, n48051, n48052, n48053,
n48054, n48055, n48056, n48057, n48058, n48059, n48060, n48061,
n48062, n48063, n48064, n48065, n48066, n48067, n48068, n48069,
n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077,
n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085,
n48086, n48087, n48088, n48089, n48090, n48091, n48092, n48093,
n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101,
n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48109,
n48110, n48111, n48112, n48113, n48114, n48115, n48116, n48117,
n48118, n48119, n48120, n48121, n48122, n48123, n48124, n48125,
n48126, n48127, n48128, n48129, n48130, n48131, n48132, n48133,
n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141,
n48142, n48143, n48144, n48145, n48146, n48147, n48148, n48149,
n48150, n48151, n48152, n48153, n48154, n48155, n48156, n48157,
n48158, n48159, n48160, n48161, n48162, n48163, n48164, n48165,
n48166, n48167, n48168, n48169, n48170, n48171, n48172, n48173,
n48174, n48175, n48176, n48177, n48178, n48179, n48180, n48181,
n48182, n48183, n48184, n48185, n48186, n48187, n48188, n48189,
n48190, n48191, n48192, n48193, n48194, n48195, n48196, n48197,
n48198, n48199, n48200, n48201, n48202, n48203, n48204, n48205,
n48206, n48207, n48208, n48209, n48210, n48211, n48212, n48213,
n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221,
n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229,
n48230, n48231, n48232, n48233, n48234, n48235, n48236, n48237,
n48238, n48239, n48240, n48241, n48242, n48243, n48244, n48245,
n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253,
n48254, n48255, n48256, n48257, n48258, n48259, n48260, n48261,
n48262, n48263, n48264, n48265, n48266, n48267, n48268, n48269,
n48270, n48271, n48272, n48273, n48274, n48275, n48276, n48277,
n48278, n48279, n48280, n48281, n48282, n48283, n48284, n48285,
n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293,
n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301,
n48302, n48303, n48304, n48305, n48306, n48307, n48308, n48309,
n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317,
n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325,
n48326, n48327, n48328, n48329, n48330, n48331, n48332, n48333,
n48334, n48335, n48336, n48337, n48338, n48339, n48340, n48341,
n48342, n48343, n48344, n48345, n48346, n48347, n48348, n48349,
n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357,
n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365,
n48366, n48367, n48368, n48369, n48370, n48371, n48372, n48373,
n48374, n48375, n48376, n48377, n48378, n48379, n48380, n48381,
n48382, n48383, n48384, n48385, n48386, n48387, n48388, n48389,
n48390, n48391, n48392, n48393, n48394, n48395, n48396, n48397,
n48398, n48399, n48400, n48401, n48402, n48403, n48404, n48405,
n48406, n48407, n48408, n48409, n48410, n48411, n48412, n48413,
n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421,
n48422, n48423, n48424, n48425, n48426, n48427, n48428, n48429,
n48430, n48431, n48432, n48433, n48434, n48435, n48436, n48437,
n48438, n48439, n48440, n48441, n48442, n48443, n48444, n48445,
n48446, n48447, n48448, n48449, n48450, n48451, n48452, n48453,
n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461,
n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469,
n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477,
n48478, n48479, n48480, n48481, n48482, n48483, n48484, n48485,
n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493,
n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501,
n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509,
n48510, n48511, n48512, n48513, n48514, n48515, n48516, n48517,
n48518, n48519, n48520, n48521, n48522, n48523, n48524, n48525,
n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533,
n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541,
n48542, n48543, n48544, n48545, n48546, n48547, n48548, n48549,
n48550, n48551, n48552, n48553, n48554, n48555, n48556, n48557,
n48558, n48559, n48560, n48561, n48562, n48563, n48564, n48565,
n48566, n48567, n48568, n48569, n48570, n48571, n48572, n48573,
n48574, n48575, n48576, n48577, n48578, n48579, n48580, n48581,
n48582, n48583, n48584, n48585, n48586, n48587, n48588, n48589,
n48590, n48591, n48592, n48593, n48594, n48595, n48596, n48597,
n48598, n48599, n48600, n48601, n48602, n48603, n48604, n48605,
n48606, n48607, n48608, n48609, n48610, n48611, n48612, n48613,
n48614, n48615, n48616, n48617, n48618, n48619, n48620, n48621,
n48622, n48623, n48624, n48625, n48626, n48627, n48628, n48629,
n48630, n48631, n48632, n48633, n48634, n48635, n48636, n48637,
n48638, n48639, n48640, n48641, n48642, n48643, n48644, n48645,
n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653,
n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661,
n48662, n48663, n48664, n48665, n48666, n48667, n48668, n48669,
n48670, n48671, n48672, n48673, n48674, n48675, n48676, n48677,
n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685,
n48686, n48687, n48688, n48689, n48690, n48691, n48692, n48693,
n48694, n48695, n48696, n48697, n48698, n48699, n48700, n48701,
n48702, n48703, n48704, n48705, n48706, n48707, n48708, n48709,
n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717,
n48718, n48719, n48720, n48721, n48722, n48723, n48724, n48725,
n48726, n48727, n48728, n48729, n48730, n48731, n48732, n48733,
n48734, n48735, n48736, n48737, n48738, n48739, n48740, n48741,
n48742, n48743, n48744, n48745, n48746, n48747, n48748, n48749,
n48750, n48751, n48752, n48753, n48754, n48755, n48756, n48757,
n48758, n48759, n48760, n48761, n48762, n48763, n48764, n48765,
n48766, n48767, n48768, n48769, n48770, n48771, n48772, n48773,
n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781,
n48782, n48783, n48784, n48785, n48786, n48787, n48788, n48789,
n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797,
n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805,
n48806, n48807, n48808, n48809, n48810, n48811, n48812, n48813,
n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821,
n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829,
n48830, n48831, n48832, n48833, n48834, n48835, n48836, n48837,
n48838, n48839, n48840, n48841, n48842, n48843, n48844, n48845,
n48846, n48847, n48848, n48849, n48850, n48851, n48852, n48853,
n48854, n48855, n48856, n48857, n48858, n48859, n48860, n48861,
n48862, n48863, n48864, n48865, n48866, n48867, n48868, n48869,
n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877,
n48878, n48879, n48880, n48881, n48882, n48883, n48884, n48885,
n48886, n48887, n48888, n48889, n48890, n48891, n48892, n48893,
n48894, n48895, n48896, n48897, n48898, n48899, n48900, n48901,
n48902, n48903, n48904, n48905, n48906, n48907, n48908, n48909,
n48910, n48911, n48912, n48913, n48914, n48915, n48916, n48917,
n48918, n48919, n48920, n48921, n48922, n48923, n48924, n48925,
n48926, n48927, n48928, n48929, n48930, n48931, n48932, n48933,
n48934, n48935, n48936, n48937, n48938, n48939, n48940, n48941,
n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949,
n48950, n48951, n48952, n48953, n48954, n48955, n48956, n48957,
n48958, n48959, n48960, n48961, n48962, n48963, n48964, n48965,
n48966, n48967, n48968, n48969, n48970, n48971, n48972, n48973,
n48974, n48975, n48976, n48977, n48978, n48979, n48980, n48981,
n48982, n48983, n48984, n48985, n48986, n48987, n48988, n48989,
n48990, n48991, n48992, n48993, n48994, n48995, n48996, n48997,
n48998, n48999, n49000, n49001, n49002, n49003, n49004, n49005,
n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013,
n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021,
n49022, n49023, n49024, n49025, n49026, n49027, n49028, n49029,
n49030, n49031, n49032, n49033, n49034, n49035, n49036, n49037,
n49038, n49039, n49040, n49041, n49042, n49043, n49044, n49045,
n49046, n49047, n49048, n49049, n49050, n49051, n49052, n49053,
n49054, n49055, n49056, n49057, n49058, n49059, n49060, n49061,
n49062, n49063, n49064, n49065, n49066, n49067, n49068, n49069,
n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077,
n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085,
n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093,
n49094, n49095, n49096, n49097, n49098, n49099, n49100, n49101,
n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109,
n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117,
n49118, n49119, n49120, n49121, n49122, n49123, n49124, n49125,
n49126, n49127, n49128, n49129, n49130, n49131, n49132, n49133,
n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141,
n49142, n49143, n49144, n49145, n49146, n49147, n49148, n49149,
n49150, n49151, n49152, n49153, n49154, n49155, n49156, n49157,
n49158, n49159, n49160, n49161, n49162, n49163, n49164, n49165,
n49166, n49167, n49168, n49169, n49170, n49171, n49172, n49173,
n49174, n49175, n49176, n49177, n49178, n49179, n49180, n49181,
n49182, n49183, n49184, n49185, n49186, n49187, n49188, n49189,
n49190, n49191, n49192, n49193, n49194, n49195, n49196, n49197,
n49198, n49199, n49200, n49201, n49202, n49203, n49204, n49205,
n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213,
n49214, n49215, n49216, n49217, n49218, n49219, n49220, n49221,
n49222, n49223, n49224, n49225, n49226, n49227, n49228, n49229,
n49230, n49231, n49232, n49233, n49234, n49235, n49236, n49237,
n49238, n49239, n49240, n49241, n49242, n49243, n49244, n49245,
n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253,
n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261,
n49262, n49263, n49264, n49265, n49266, n49267, n49268, n49269,
n49270, n49271, n49272, n49273, n49274, n49275, n49276, n49277,
n49278, n49279, n49280, n49281, n49282, n49283, n49284, n49285,
n49286, n49287, n49288, n49289, n49290, n49291, n49292, n49293,
n49294, n49295, n49296, n49297, n49298, n49299, n49300, n49301,
n49302, n49303, n49304, n49305, n49306, n49307, n49308, n49309,
n49310, n49311, n49312, n49313, n49314, n49315, n49316, n49317,
n49318, n49319, n49320, n49321, n49322, n49323, n49324, n49325,
n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333,
n49334, n49335, n49336, n49337, n49338, n49339, n49340, n49341,
n49342, n49343, n49344, n49345, n49346, n49347, n49348, n49349,
n49350, n49351, n49352, n49353, n49354, n49355, n49356, n49357,
n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365,
n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373,
n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381,
n49382, n49383, n49384, n49385, n49386, n49387, n49388, n49389,
n49390, n49391, n49392, n49393, n49394, n49395, n49396, n49397,
n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405,
n49406, n49407, n49408, n49409, n49410, n49411, n49412, n49413,
n49414, n49415, n49416, n49417, n49418, n49419, n49420, n49421,
n49422, n49423, n49424, n49425, n49426, n49427, n49428, n49429,
n49430, n49431, n49432, n49433, n49434, n49435, n49436, n49437,
n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445,
n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453,
n49454, n49455, n49456, n49457, n49458, n49459, n49460, n49461,
n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469,
n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477,
n49478, n49479, n49480, n49481, n49482, n49483, n49484, n49486,
n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494,
n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502,
n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510,
n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518,
n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526,
n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534,
n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542,
n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550,
n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558,
n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566,
n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574,
n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582,
n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590,
n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598,
n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606,
n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614,
n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622,
n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630,
n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638,
n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646,
n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654,
n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662,
n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670,
n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678,
n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686,
n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694,
n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702,
n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710,
n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718,
n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726,
n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734,
n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742,
n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750,
n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758,
n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766,
n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774,
n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782,
n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790,
n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798,
n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806,
n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814,
n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822,
n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830,
n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838,
n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846,
n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854,
n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862,
n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870,
n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878,
n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886,
n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894,
n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902,
n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910,
n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918,
n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926,
n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934,
n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942,
n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950,
n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958,
n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966,
n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974,
n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982,
n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990,
n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998,
n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006,
n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014,
n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022,
n50023, n50024, n50025, n50026, n50027, n50030, n50031, n50032,
n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040,
n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056,
n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064,
n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072,
n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080,
n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088,
n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096,
n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104,
n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112,
n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120,
n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128,
n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136,
n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144,
n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152,
n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160,
n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168,
n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176,
n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184,
n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192,
n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200,
n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208,
n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216,
n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224,
n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232,
n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240,
n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248,
n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256,
n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264,
n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272,
n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280,
n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288,
n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296,
n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304,
n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312,
n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320,
n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328,
n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336,
n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344,
n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352,
n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360,
n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368,
n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376,
n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384,
n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392,
n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400,
n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408,
n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416,
n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424,
n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432,
n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440,
n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448,
n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456,
n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464,
n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472,
n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480,
n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488,
n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496,
n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504,
n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512,
n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520,
n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528,
n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536,
n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544,
n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552,
n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560,
n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568,
n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576,
n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584,
n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592,
n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600,
n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608,
n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616,
n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624,
n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632,
n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640,
n50641, n50642, n50643, n50644, n50645, n50647, n50648, n50649,
n50650, n50651, n50652, n50653, n50654, n50655, n50656, n50657,
n50658, n50659, n50660, n50661, n50662, n50663, n50664, n50665,
n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673,
n50674, n50675, n50676, n50677, n50678, n50679, n50680, n50681,
n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689,
n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697,
n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705,
n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713,
n50714, n50715, n50716, n50717, n50718, n50719, n50720, n50721,
n50722, n50723, n50724, n50725, n50726, n50727, n50728, n50729,
n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737,
n50738, n50739, n50740, n50741, n50742, n50743, n50744, n50745,
n50746, n50747, n50748, n50749, n50750, n50751, n50752, n50753,
n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761,
n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769,
n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777,
n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785,
n50786, n50787, n50788, n50789, n50790, n50791, n50792, n50793,
n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801,
n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809,
n50810, n50811, n50812, n50813, n50814, n50815, n50816, n50817,
n50818, n50819, n50820, n50821, n50822, n50823, n50824, n50825,
n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833,
n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841,
n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849,
n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857,
n50858, n50859, n50860, n50861, n50862, n50863, n50864, n50865,
n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873,
n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881,
n50882, n50883, n50884, n50885, n50886, n50887, n50888, n50889,
n50890, n50891, n50892, n50893, n50894, n50895, n50896, n50897,
n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905,
n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913,
n50914, n50915, n50917, n50918, n50919, n50920, n50921, n50922,
n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962,
n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970,
n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978,
n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994,
n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018,
n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034,
n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042,
n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050,
n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082,
n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090,
n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106,
n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114,
n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122,
n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138,
n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154,
n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162,
n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178,
n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194,
n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258,
n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266,
n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282,
n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298,
n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306,
n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322,
n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330,
n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338,
n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394,
n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410,
n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426,
n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442,
n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474,
n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498,
n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514,
n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522,
n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530,
n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538,
n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546,
n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554,
n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570,
n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586,
n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594,
n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602,
n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610,
n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618,
n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626,
n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642,
n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658,
n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666,
n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674,
n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682,
n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690,
n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698,
n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730,
n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738,
n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746,
n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754,
n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762,
n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770,
n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786,
n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794,
n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802,
n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810,
n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818,
n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826,
n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834,
n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842,
n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858,
n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866,
n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874,
n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882,
n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898,
n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906,
n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914,
n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930,
n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51947,
n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955,
n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963,
n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971,
n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979,
n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987,
n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995,
n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003,
n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011,
n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019,
n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027,
n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035,
n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043,
n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051,
n52052, n52053, n52054, n52055, n52056, n52057, n52058, n52059,
n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067,
n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075,
n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083,
n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091,
n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099,
n52100, n52101, n52102, n52103, n52104, n52105, n52106, n52107,
n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115,
n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123,
n52124, n52125, n52126, n52127, n52128, n52129, n52130, n52131,
n52132, n52133, n52134, n52135, n52136, n52137, n52138, n52139,
n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147,
n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155,
n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163,
n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171,
n52172, n52173, n52174, n52175, n52176, n52177, n52178, n52179,
n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187,
n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195,
n52196, n52197, n52198, n52199, n52200, n52201, n52202, n52203,
n52204, n52205, n52206, n52207, n52208, n52209, n52210, n52211,
n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219,
n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227,
n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235,
n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243,
n52244, n52245, n52246, n52247, n52248, n52249, n52250, n52251,
n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259,
n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267,
n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275,
n52276, n52277, n52278, n52279, n52280, n52281, n52282, n52283,
n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291,
n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299,
n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307,
n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315,
n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323,
n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331,
n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339,
n52340, n52341, n52342, n52343, n52344, n52345, n52346, n52347,
n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355,
n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363,
n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371,
n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379,
n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387,
n52388, n52389, n52390, n52391, n52392, n52393, n52394, n52395,
n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403,
n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411,
n52412, n52413, n52414, n52415, n52416, n52417, n52418, n52419,
n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427,
n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435,
n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443,
n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451,
n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459,
n52460, n52461, n52462, n52463, n52464, n52465, n52466, n52467,
n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475,
n52476, n52477, n52478, n52480, n52481, n52482, n52483, n52484,
n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492,
n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500,
n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508,
n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516,
n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524,
n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532,
n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540,
n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548,
n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556,
n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564,
n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572,
n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580,
n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588,
n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596,
n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604,
n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612,
n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620,
n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628,
n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636,
n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644,
n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652,
n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660,
n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668,
n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676,
n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684,
n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692,
n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700,
n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708,
n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716,
n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724,
n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732,
n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740,
n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748,
n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756,
n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764,
n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772,
n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780,
n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788,
n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796,
n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804,
n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812,
n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820,
n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828,
n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836,
n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844,
n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852,
n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860,
n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868,
n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876,
n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884,
n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892,
n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900,
n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908,
n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916,
n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924,
n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932,
n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940,
n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948,
n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956,
n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964,
n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972,
n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980,
n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988,
n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996,
n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004,
n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012,
n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020,
n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028,
n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036,
n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044,
n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052,
n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060,
n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068,
n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076,
n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084,
n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092,
n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100,
n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108,
n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116,
n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124,
n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132,
n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140,
n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148,
n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156,
n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164,
n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172,
n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180,
n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188,
n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196,
n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204,
n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212,
n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220,
n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228,
n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244,
n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252,
n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260,
n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268,
n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276,
n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284,
n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292,
n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300,
n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308,
n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316,
n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324,
n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332,
n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340,
n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348,
n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356,
n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364,
n53365, n53366, n53367, n53368, n53370, n53371, n53372, n53373,
n53374, n53375, n53376, n53377, n53378, n53379, n53380, n53381,
n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389,
n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397,
n53398, n53399, n53400, n53401, n53402, n53403, n53404, n53405,
n53406, n53407, n53408, n53409, n53410, n53411, n53412, n53413,
n53414, n53415, n53416, n53417, n53418, n53419, n53420, n53421,
n53422, n53423, n53424, n53425, n53426, n53427, n53428, n53429,
n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437,
n53438, n53439, n53440, n53441, n53442, n53443, n53444, n53445,
n53446, n53447, n53448, n53449, n53450, n53451, n53452, n53453,
n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461,
n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469,
n53470, n53471, n53472, n53473, n53474, n53475, n53476, n53477,
n53478, n53479, n53480, n53481, n53482, n53483, n53484, n53485,
n53486, n53487, n53488, n53489, n53490, n53491, n53492, n53493,
n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501,
n53502, n53503, n53504, n53505, n53506, n53507, n53508, n53509,
n53510, n53511, n53512, n53513, n53514, n53515, n53516, n53517,
n53518, n53519, n53520, n53521, n53522, n53523, n53524, n53525,
n53526, n53527, n53528, n53529, n53530, n53531, n53532, n53533,
n53534, n53535, n53536, n53537, n53538, n53539, n53540, n53541,
n53542, n53543, n53544, n53545, n53546, n53547, n53548, n53549,
n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557,
n53558, n53559, n53560, n53561, n53562, n53563, n53564, n53565,
n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573,
n53574, n53575, n53576, n53577, n53578, n53579, n53580, n53581,
n53582, n53583, n53584, n53585, n53586, n53587, n53588, n53589,
n53590, n53591, n53592, n53593, n53594, n53595, n53596, n53597,
n53598, n53599, n53600, n53601, n53602, n53603, n53604, n53605,
n53606, n53607, n53608, n53609, n53610, n53611, n53612, n53613,
n53614, n53615, n53616, n53617, n53618, n53619, n53620, n53621,
n53622, n53623, n53624, n53625, n53626, n53627, n53628, n53629,
n53630, n53631, n53632, n53633, n53634, n53635, n53636, n53637,
n53638, n53639, n53640, n53641, n53642, n53643, n53644, n53645,
n53646, n53647, n53648, n53649, n53650, n53651, n53652, n53653,
n53654, n53655, n53656, n53657, n53658, n53659, n53660, n53661,
n53662, n53663, n53664, n53665, n53666, n53667, n53668, n53669,
n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677,
n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685,
n53686, n53687, n53688, n53689, n53690, n53691, n53692, n53693,
n53694, n53695, n53696, n53697, n53698, n53699, n53700, n53701,
n53702, n53703, n53704, n53705, n53706, n53707, n53708, n53709,
n53710, n53711, n53712, n53713, n53714, n53715, n53716, n53717,
n53718, n53719, n53720, n53721, n53722, n53723, n53724, n53725,
n53726, n53727, n53728, n53729, n53730, n53731, n53732, n53733,
n53734, n53735, n53736, n53737, n53738, n53739, n53740, n53741,
n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749,
n53750, n53751, n53752, n53753, n53754, n53755, n53756, n53757,
n53758, n53759, n53760, n53761, n53762, n53763, n53764, n53765,
n53766, n53767, n53768, n53769, n53770, n53771, n53772, n53773,
n53774, n53775, n53776, n53777, n53778, n53779, n53780, n53781,
n53782, n53783, n53784, n53785, n53786, n53787, n53788, n53789,
n53790, n53791, n53792, n53793, n53794, n53795, n53796, n53797,
n53798, n53799, n53800, n53801, n53802, n53803, n53804, n53805,
n53806, n53807, n53808, n53809, n53810, n53811, n53812, n53813,
n53814, n53815, n53816, n53817, n53818, n53819, n53820, n53821,
n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829,
n53830, n53831, n53832, n53833, n53834, n53835, n53836, n53837,
n53838, n53839, n53840, n53841, n53842, n53843, n53844, n53845,
n53846, n53847, n53848, n53849, n53850, n53851, n53852, n53853,
n53854, n53855, n53856, n53857, n53858, n53859, n53860, n53861,
n53862, n53863, n53864, n53865, n53866, n53867, n53868, n53869,
n53870, n53871, n53872, n53873, n53874, n53875, n53876, n53877,
n53878, n53879, n53880, n53881, n53882, n53883, n53884, n53885,
n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893,
n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901,
n53902, n53903, n53904, n53905, n53906, n53907, n53908, n53909,
n53910, n53911, n53912, n53913, n53914, n53915, n53916, n53917,
n53918, n53919, n53920, n53921, n53922, n53923, n53924, n53925,
n53926, n53927, n53928, n53929, n53930, n53931, n53932, n53933,
n53934, n53935, n53936, n53937, n53938, n53939, n53940, n53941,
n53942, n53943, n53944, n53945, n53946, n53947, n53948, n53949,
n53950, n53951, n53952, n53953, n53954, n53955, n53956, n53957,
n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965,
n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973,
n53974, n53975, n53976, n53977, n53978, n53979, n53980, n53981,
n53982, n53983, n53984, n53985, n53986, n53987, n53988, n53989,
n53990, n53991, n53992, n53993, n53994, n53995, n53996, n53997,
n53998, n53999, n54000, n54001, n54002, n54003, n54004, n54005,
n54006, n54007, n54008, n54009, n54010, n54011, n54012, n54013,
n54014, n54015, n54016, n54017, n54018, n54019, n54020, n54021,
n54022, n54023, n54024, n54025, n54026, n54027, n54028, n54029,
n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037,
n54038, n54039, n54040, n54041, n54042, n54043, n54044, n54045,
n54046, n54047, n54048, n54049, n54050, n54051, n54052, n54053,
n54054, n54055, n54056, n54057, n54058, n54059, n54060, n54061,
n54062, n54063, n54064, n54065, n54066, n54067, n54068, n54069,
n54070, n54073, n54074, n54075, n54076, n54077, n54078, n54079,
n54080, n54081, n54082, n54083, n54084, n54085, n54086, n54087,
n54088, n54089, n54090, n54091, n54092, n54093, n54094, n54095,
n54096, n54097, n54098, n54099, n54100, n54101, n54102, n54103,
n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111,
n54112, n54113, n54114, n54115, n54116, n54117, n54118, n54119,
n54120, n54121, n54122, n54123, n54124, n54125, n54126, n54127,
n54128, n54129, n54130, n54131, n54132, n54133, n54134, n54135,
n54136, n54137, n54138, n54139, n54140, n54141, n54142, n54143,
n54144, n54145, n54146, n54147, n54148, n54149, n54150, n54151,
n54152, n54153, n54154, n54155, n54156, n54157, n54158, n54159,
n54160, n54161, n54162, n54163, n54164, n54165, n54166, n54167,
n54168, n54169, n54170, n54171, n54172, n54173, n54174, n54175,
n54176, n54177, n54178, n54179, n54180, n54181, n54182, n54183,
n54184, n54185, n54186, n54187, n54188, n54189, n54190, n54191,
n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199,
n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207,
n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215,
n54216, n54217, n54218, n54219, n54220, n54221, n54222, n54223,
n54224, n54225, n54226, n54227, n54228, n54229, n54230, n54231,
n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239,
n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54247,
n54248, n54249, n54250, n54251, n54252, n54253, n54254, n54255,
n54256, n54257, n54258, n54259, n54260, n54261, n54262, n54263,
n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271,
n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54279,
n54280, n54281, n54282, n54283, n54284, n54285, n54286, n54287,
n54288, n54289, n54290, n54291, n54292, n54293, n54294, n54295,
n54296, n54297, n54298, n54299, n54300, n54301, n54302, n54303,
n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311,
n54312, n54313, n54314, n54315, n54316, n54317, n54318, n54319,
n54320, n54321, n54322, n54323, n54324, n54325, n54326, n54327,
n54328, n54329, n54330, n54331, n54332, n54333, n54334, n54335,
n54336, n54337, n54338, n54339, n54340, n54341, n54342, n54343,
n54344, n54345, n54346, n54347, n54348, n54349, n54350, n54351,
n54352, n54353, n54354, n54355, n54356, n54357, n54358, n54359,
n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367,
n54368, n54369, n54370, n54371, n54372, n54373, n54374, n54375,
n54376, n54377, n54378, n54379, n54380, n54381, n54382, n54383,
n54384, n54385, n54386, n54387, n54388, n54389, n54390, n54391,
n54392, n54393, n54394, n54395, n54396, n54397, n54398, n54399,
n54400, n54401, n54402, n54403, n54404, n54405, n54406, n54407,
n54408, n54409, n54410, n54411, n54412, n54413, n54414, n54415,
n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423,
n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431,
n54432, n54433, n54434, n54435, n54436, n54437, n54438, n54439,
n54440, n54441, n54442, n54443, n54444, n54445, n54446, n54447,
n54448, n54449, n54450, n54451, n54452, n54453, n54454, n54455,
n54456, n54457, n54458, n54459, n54460, n54461, n54462, n54463,
n54464, n54465, n54466, n54467, n54468, n54469, n54470, n54471,
n54472, n54473, n54474, n54475, n54476, n54477, n54478, n54479,
n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487,
n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495,
n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503,
n54504, n54505, n54506, n54507, n54508, n54509, n54510, n54511,
n54512, n54513, n54514, n54515, n54516, n54517, n54518, n54519,
n54520, n54521, n54522, n54523, n54524, n54525, n54526, n54527,
n54528, n54529, n54530, n54531, n54532, n54533, n54534, n54535,
n54536, n54537, n54538, n54539, n54540, n54541, n54542, n54543,
n54544, n54545, n54546, n54547, n54548, n54549, n54550, n54551,
n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559,
n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567,
n54568, n54569, n54570, n54571, n54572, n54573, n54574, n54575,
n54576, n54577, n54578, n54579, n54580, n54581, n54582, n54583,
n54584, n54586, n54587, n54588, n54589, n54590, n54591, n54592,
n54593, n54594, n54595, n54596, n54597, n54598, n54599, n54600,
n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608,
n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616,
n54617, n54618, n54619, n54620, n54621, n54622, n54623, n54624,
n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632,
n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640,
n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648,
n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656,
n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664,
n54665, n54666, n54667, n54668, n54669, n54670, n54671, n54672,
n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680,
n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688,
n54689, n54690, n54691, n54692, n54693, n54694, n54695, n54696,
n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704,
n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712,
n54713, n54714, n54715, n54716, n54717, n54718, n54720, n54721,
n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729,
n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737,
n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745,
n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753,
n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761,
n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769,
n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777,
n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785,
n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793,
n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801,
n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809,
n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817,
n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825,
n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833,
n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841,
n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849,
n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857,
n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865,
n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873,
n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881,
n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889,
n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897,
n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905,
n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913,
n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921,
n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929,
n54930, n54932, n54933, n54934, n54935, n54936, n54937, n54938,
n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946,
n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954,
n54955, n54956, n54957, n54959, n54960, n54961, n54962, n54963,
n54964, n54965, n54966, n54967, n54968, n54969, n54970, n54971,
n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979,
n54980, n54981, n54982, n54983, n54984, n54985, n54986, n54987,
n54988, n54989, n54990, n54991, n54992, n54993, n54994, n54995,
n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003,
n55004, n55005, n55006, n55007, n55008, n55009, n55010, n55011,
n55012, n55013, n55014, n55015, n55016, n55017, n55018, n55019,
n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027,
n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035,
n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043,
n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051,
n55052, n55053, n55054, n55055, n55056, n55057, n55058, n55059,
n55060, n55061, n55062, n55063, n55064, n55065, n55066, n55067,
n55068, n55069, n55070, n55071, n55072, n55073, n55074, n55075,
n55076, n55077, n55078, n55079, n55080, n55081, n55082, n55083,
n55084, n55085, n55086, n55087, n55088, n55089, n55090, n55091,
n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099,
n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107,
n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115,
n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123,
n55124, n55125, n55126, n55127, n55128, n55129, n55130, n55131,
n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139,
n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147,
n55148, n55149, n55150, n55151, n55152, n55153, n55154, n55155,
n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163,
n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171,
n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179,
n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187,
n55188, n55189, n55190, n55191, n55192, n55193, n55195, n55196,
n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204,
n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212,
n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220,
n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228,
n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236,
n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244,
n55246, n55247, n55248, n55249, n55250, n55251, n55252, n55253,
n55254, n55255, n55256, n55257, n55258, n55259, n55260, n55261,
n55262, n55263, n55264, n55265, n55266, n55267, n55268, n55269,
n55270, n55271, n55272, n55273, n55274, n55275, n55276, n55277,
n55278, n55279, n55280, n55281, n55282, n55283, n55284, n55285,
n55286, n55287, n55288, n55289, n55290, n55291, n55292, n55293,
n55294, n55295, n55296, n55297, n55298, n55299, n55300, n55301,
n55302, n55303, n55304, n55305, n55306, n55307, n55308, n55309,
n55310, n55311, n55312, n55313, n55314, n55315, n55316, n55317,
n55318, n55319, n55320, n55321, n55322, n55323, n55324, n55325,
n55326, n55327, n55328, n55329, n55330, n55331, n55332, n55333,
n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341,
n55342, n55343, n55344, n55345, n55346, n55347, n55348, n55349,
n55351, n55352, n55353, n55354, n55355, n55356, n55357, n55358,
n55359, n55360, n55361, n55362, n55363, n55364, n55365, n55366,
n55367, n55368, n55369, n55370, n55371, n55372, n55373, n55374,
n55375, n55376, n55377, n55378, n55379, n55380, n55381, n55382,
n55383, n55384, n55385, n55386, n55387, n55388, n55389, n55390,
n55391, n55392, n55393, n55394, n55395, n55396, n55397, n55398,
n55399, n55400, n55401, n55402, n55403, n55404, n55405, n55406,
n55407, n55408, n55409, n55410, n55411, n55412, n55413, n55414,
n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55422,
n55423, n55424, n55425, n55426, n55427, n55428, n55429, n55430,
n55431, n55432, n55433, n55434, n55435, n55436, n55437, n55438,
n55439, n55440, n55441, n55442, n55443, n55444, n55445, n55446,
n55447, n55448, n55449, n55450, n55451, n55452, n55453, n55454,
n55455, n55456, n55457, n55458, n55459, n55460, n55461, n55462,
n55463, n55464, n55465, n55466, n55467, n55468, n55469, n55470,
n55471, n55472, n55473, n55474, n55475, n55476, n55477, n55478,
n55479, n55480, n55481, n55482, n55483, n55484, n55485, n55486,
n55487, n55488, n55489, n55490, n55491, n55492, n55493, n55494,
n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502,
n55503, n55504, n55505, n55506, n55507, n55508, n55509, n55510,
n55511, n55512, n55513, n55514, n55515, n55516, n55517, n55518,
n55519, n55520, n55521, n55522, n55523, n55524, n55525, n55526,
n55527, n55528, n55529, n55530, n55531, n55532, n55533, n55534,
n55535, n55536, n55537, n55538, n55539, n55540, n55541, n55542,
n55543, n55544, n55545, n55546, n55547, n55548, n55549, n55550,
n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558,
n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566,
n55567, n55568, n55569, n55570, n55571, n55572, n55573, n55574,
n55575, n55576, n55577, n55578, n55579, n55580, n55581, n55582,
n55583, n55584, n55585, n55586, n55587, n55588, n55589, n55590,
n55591, n55592, n55593, n55594, n55595, n55596, n55597, n55598,
n55599, n55600, n55601, n55602, n55603, n55604, n55605, n55606,
n55607, n55608, n55609, n55610, n55611, n55612, n55613, n55614,
n55615, n55616, n55617, n55618, n55619, n55620, n55621, n55622,
n55623, n55624, n55625, n55626, n55627, n55628, n55629, n55630,
n55631, n55632, n55633, n55634, n55635, n55636, n55637, n55638,
n55639, n55640, n55641, n55642, n55643, n55644, n55645, n55646,
n55647, n55648, n55649, n55650, n55651, n55652, n55653, n55654,
n55655, n55656, n55657, n55658, n55659, n55660, n55661, n55662,
n55663, n55664, n55665, n55666, n55667, n55668, n55669, n55670,
n55671, n55672, n55673, n55674, n55675, n55676, n55677, n55678,
n55679, n55680, n55681, n55682, n55683, n55684, n55685, n55686,
n55687, n55688, n55689, n55690, n55691, n55692, n55693, n55694,
n55695, n55696, n55697, n55698, n55699, n55700, n55701, n55702,
n55703, n55704, n55705, n55706, n55707, n55708, n55709, n55710,
n55711, n55712, n55713, n55714, n55715, n55716, n55717, n55718,
n55719, n55720, n55721, n55722, n55723, n55724, n55725, n55726,
n55727, n55728, n55729, n55730, n55731, n55732, n55733, n55734,
n55735, n55736, n55737, n55738, n55739, n55740, n55741, n55742,
n55743, n55744, n55745, n55746, n55747, n55748, n55749, n55750,
n55751, n55752, n55753, n55754, n55755, n55756, n55757, n55758,
n55759, n55760, n55761, n55762, n55763, n55764, n55765, n55766,
n55767, n55768, n55769, n55770, n55771, n55772, n55773, n55774,
n55775, n55776, n55777, n55778, n55779, n55780, n55781, n55782,
n55783, n55784, n55785, n55786, n55787, n55788, n55789, n55790,
n55791, n55792, n55793, n55794, n55795, n55796, n55797, n55798,
n55799, n55800, n55801, n55802, n55803, n55804, n55805, n55806,
n55807, n55808, n55809, n55812, n55813, n55814, n55815, n55816,
n55817, n55818, n55819, n55820, n55821, n55822, n55823, n55824,
n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832,
n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840,
n55841, n55842, n55843, n55844, n55845, n55846, n55847, n55848,
n55849, n55850, n55851, n55852, n55853, n55854, n55855, n55856,
n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864,
n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872,
n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880,
n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888,
n55889, n55890, n55891, n55892, n55893, n55894, n55895, n55896,
n55897, n55898, n55899, n55900, n55901, n55903, n55904, n55905,
n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913,
n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921,
n55922, n55923, n55924, n55925, n55926, n55927, n55928, n55929,
n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937,
n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945,
n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953,
n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961,
n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969,
n55970, n55971, n55972, n55973, n55974, n55975, n55976, n55977,
n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985,
n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993,
n55994, n55995, n55996, n55997, n55998, n55999, n56000, n56001,
n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009,
n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017,
n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025,
n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033,
n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041,
n56042, n56043, n56044, n56045, n56046, n56047, n56048, n56049,
n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057,
n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065,
n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073,
n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081,
n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089,
n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097,
n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105,
n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113,
n56114, n56115, n56116, n56117, n56118, n56119, n56120, n56121,
n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129,
n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137,
n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145,
n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153,
n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161,
n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169,
n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177,
n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185,
n56186, n56187, n56188, n56189, n56190, n56191, n56192, n56193,
n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201,
n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209,
n56210, n56211, n56212, n56213, n56214, n56216, n56217, n56218,
n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226,
n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234,
n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242,
n56243, n56244, n56245, n56246, n56247, n56250, n56251, n56254,
n56255, n56256, n56257, n56260, n56261, n56262, n56263, n56264,
n56265, n56266, n56267, n56268, n56269, n56270, n56271, n56272,
n56273, n56274, n56275, n56276, n56277, n56278, n56279, n56280,
n56281, n56282, n56283, n56284, n56285, n56286, n56287, n56288,
n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296,
n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304,
n56305, n56306, n56307, n56308, n56309, n56310, n56311, n56312,
n56313, n56314, n56315, n56316, n56317, n56318, n56319, n56320,
n56321, n56322, n56323, n56324, n56325, n56326, n56327, n56328,
n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337,
n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345,
n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353,
n56354, n56355, n56356, n56357, n56358, n56359, n56360, n56361,
n56362, n56363, n56364, n56365, n56366, n56367, n56368, n56369,
n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377,
n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385,
n56386, n56387, n56388, n56389, n56390, n56391, n56392, n56393,
n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401,
n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409,
n56410, n56411, n56412, n56413, n56414, n56415, n56416, n56417,
n56418, n56419, n56420, n56421, n56422, n56423, n56424, n56425,
n56426, n56427, n56428, n56429, n56430, n56431, n56432, n56433,
n56434, n56435, n56436, n56437, n56438, n56439, n56440, n56441,
n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449,
n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457,
n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56465,
n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473,
n56474, n56475, n56476, n56477, n56478, n56479, n56480, n56481,
n56482, n56483, n56484, n56485, n56486, n56487, n56488, n56489,
n56490, n56491, n56492, n56493, n56494, n56495, n56496, n56497,
n56498, n56499, n56500, n56501, n56502, n56503, n56504, n56505,
n56506, n56507, n56508, n56509, n56510, n56511, n56512, n56513,
n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521,
n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529,
n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537,
n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545,
n56546, n56547, n56548, n56549, n56550, n56551, n56552, n56553,
n56554, n56555, n56556, n56557, n56558, n56559, n56560, n56561,
n56562, n56563, n56564, n56565, n56566, n56567, n56568, n56569,
n56570, n56571, n56572, n56573, n56574, n56575, n56576, n56577,
n56578, n56579, n56580, n56581, n56582, n56583, n56584, n56585,
n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593,
n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601,
n56602, n56603, n56604, n56605, n56606, n56607, n56608, n56609,
n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56617,
n56618, n56619, n56620, n56621, n56622, n56623, n56624, n56625,
n56626, n56627, n56628, n56629, n56630, n56631, n56632, n56633,
n56634, n56635, n56636, n56637, n56638, n56639, n56640, n56641,
n56642, n56643, n56644, n56645, n56646, n56647, n56648, n56649,
n56650, n56651, n56652, n56653, n56654, n56655, n56656, n56657,
n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665,
n56666, n56667, n56668, n56669, n56670, n56671, n56672, n56673,
n56674, n56675, n56676, n56677, n56678, n56679, n56680, n56681,
n56682, n56683, n56684, n56685, n56686, n56687, n56688, n56689,
n56690, n56691, n56692, n56693, n56694, n56695, n56696, n56697,
n56698, n56699, n56700, n56701, n56702, n56703, n56704, n56705,
n56706, n56707, n56708, n56709, n56710, n56711, n56712, n56713,
n56714, n56715, n56716, n56717, n56718, n56719, n56720, n56721,
n56722, n56723, n56724, n56725, n56726, n56727, n56728, n56729,
n56730, n56731, n56732, n56733, n56734, n56735, n56736, n56737,
n56738, n56739, n56740, n56741, n56742, n56743, n56744, n56745,
n56746, n56747, n56748, n56749, n56750, n56751, n56752, n56753,
n56754, n56755, n56756, n56757, n56758, n56759, n56760, n56761,
n56762, n56763, n56764, n56765, n56766, n56767, n56768, n56769,
n56770, n56771, n56772, n56773, n56774, n56775, n56776, n56777,
n56778, n56779, n56780, n56781, n56782, n56783, n56784, n56785,
n56786, n56787, n56788, n56789, n56790, n56791, n56792, n56793,
n56794, n56795, n56796, n56797, n56798, n56799, n56800, n56801,
n56802, n56803, n56804, n56805, n56806, n56807, n56808, n56809,
n56810, n56811, n56812, n56813, n56814, n56815, n56816, n56817,
n56818, n56819, n56820, n56821, n56822, n56823, n56824, n56825,
n56826, n56827, n56828, n56829, n56830, n56831, n56832, n56833,
n56834, n56835, n56836, n56837, n56838, n56839, n56840, n56841,
n56842, n56843, n56844, n56845, n56846, n56847, n56848, n56849,
n56850, n56851, n56852, n56853, n56854, n56855, n56856, n56857,
n56858, n56859, n56860, n56861, n56862, n56863, n56864, n56865,
n56866, n56867, n56868, n56869, n56870, n56871, n56872, n56873,
n56874, n56875, n56876, n56877, n56878, n56879, n56880, n56881,
n56882, n56883, n56884, n56885, n56886, n56887, n56888, n56889,
n56890, n56891, n56892, n56893, n56894, n56895, n56896, n56897,
n56898, n56899, n56900, n56901, n56902, n56903, n56904, n56905,
n56906, n56907, n56908, n56909, n56910, n56911, n56912, n56913,
n56914, n56915, n56916, n56917, n56918, n56919, n56920, n56921,
n56922, n56923, n56924, n56925, n56926, n56927, n56928, n56929,
n56930, n56931, n56932, n56933, n56934, n56935, n56936, n56937,
n56938, n56939, n56940, n56941, n56942, n56943, n56944, n56945,
n56946, n56947, n56948, n56949, n56950, n56951, n56952, n56953,
n56954, n56955, n56956, n56957, n56958, n56959, n56960, n56961,
n56962, n56963, n56964, n56965, n56966, n56967, n56968, n56969,
n56970, n56971, n56972, n56973, n56974, n56975, n56976, n56977,
n56978, n56979, n56980, n56981, n56982, n56983, n56984, n56985,
n56986, n56987, n56988, n56989, n56990, n56991, n56992, n56993,
n56994, n56995, n56996, n56997, n56998, n56999, n57000, n57001,
n57002, n57003, n57004, n57005, n57006, n57007, n57008, n57009,
n57010, n57011, n57012, n57013, n57014, n57015, n57016, n57017,
n57018, n57019, n57020, n57021, n57022, n57023, n57024, n57025,
n57026, n57027, n57028, n57029, n57030, n57031, n57032, n57033,
n57034, n57035, n57036, n57037, n57038, n57039, n57040, n57041,
n57042, n57043, n57044, n57045, n57046, n57047, n57048, n57049,
n57050, n57051, n57052, n57053, n57054, n57055, n57056, n57057,
n57058, n57059, n57060, n57061, n57062, n57063, n57064, n57065,
n57066, n57067, n57068, n57069, n57070, n57071, n57072, n57073,
n57074, n57075, n57076, n57077, n57078, n57079, n57080, n57081,
n57082, n57083, n57084, n57085, n57086, n57087, n57088, n57089,
n57090, n57091, n57092, n57093, n57094, n57095, n57096, n57097,
n57098, n57099, n57100, n57101, n57102, n57103, n57104, n57105,
n57106, n57107, n57108, n57109, n57110, n57111, n57112, n57113,
n57114, n57115, n57116, n57117, n57118, n57119, n57120, n57121,
n57122, n57123, n57124, n57125, n57126, n57127, n57128, n57129,
n57130, n57131, n57132, n57133, n57134, n57135, n57136, n57137,
n57138, n57139, n57140, n57141, n57142, n57143, n57144, n57145,
n57146, n57147, n57148, n57149, n57150, n57151, n57152, n57153,
n57154, n57155, n57156, n57157, n57158, n57159, n57160, n57161,
n57162, n57163, n57164, n57165, n57166, n57167, n57168, n57169,
n57170, n57171, n57172, n57173, n57174, n57175, n57176, n57177,
n57178, n57179, n57180, n57181, n57182, n57183, n57184, n57185,
n57186, n57187, n57188, n57189, n57190, n57191, n57192, n57193,
n57194, n57195, n57196, n57197, n57198, n57199, n57200, n57201,
n57202, n57203, n57204, n57205, n57206, n57207, n57208, n57209,
n57210, n57211, n57212, n57213, n57214, n57215, n57216, n57217,
n57218, n57219, n57220, n57221, n57222, n57223, n57224, n57225,
n57226, n57227, n57228, n57229, n57230, n57231, n57232, n57233,
n57234, n57235, n57236, n57237, n57238, n57239, n57240, n57241,
n57242, n57243, n57244, n57245, n57246, n57247, n57248, n57249,
n57250, n57251, n57252, n57253, n57254, n57255, n57256, n57257,
n57258, n57259, n57260, n57261, n57262, n57263, n57264, n57265,
n57266, n57267, n57268, n57269, n57270, n57271, n57272, n57273,
n57274, n57275, n57276, n57277, n57278, n57279, n57280, n57281,
n57282, n57283, n57284, n57285, n57286, n57287, n57288, n57289,
n57290, n57291, n57292, n57293, n57294, n57295, n57296, n57297,
n57298, n57299, n57300, n57301, n57302, n57303, n57304, n57305,
n57306, n57307, n57308, n57309, n57310, n57311, n57312, n57313,
n57314, n57315, n57316, n57317, n57318, n57319, n57320, n57321,
n57322, n57323, n57324, n57325, n57326, n57327, n57328, n57329,
n57330, n57331, n57332, n57333, n57334, n57335, n57336, n57337,
n57338, n57339, n57340, n57341, n57342, n57343, n57344, n57345,
n57346, n57347, n57348, n57349, n57350, n57351, n57352, n57353,
n57354, n57355, n57356, n57357, n57358, n57359, n57360, n57361,
n57362, n57363, n57364, n57365, n57366, n57367, n57368, n57369,
n57370, n57371, n57372, n57373, n57374, n57375, n57376, n57377,
n57378, n57379, n57380, n57381, n57382, n57383, n57384, n57385,
n57386, n57387, n57388, n57389, n57390, n57391, n57392, n57393,
n57394, n57395, n57396, n57397, n57398, n57399, n57400, n57401,
n57402, n57403, n57404, n57405, n57406, n57407, n57408, n57409,
n57410, n57411, n57412, n57413, n57414, n57415, n57416, n57417,
n57418, n57419, n57420, n57421, n57422, n57423, n57424, n57425,
n57426, n57427, n57428, n57429, n57430, n57431, n57432, n57433,
n57434, n57435, n57436, n57437, n57438, n57439, n57440, n57441,
n57442, n57443, n57444, n57445, n57446, n57447, n57448, n57449,
n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457,
n57458, n57459, n57460, n57461, n57462, n57463, n57464, n57465,
n57466, n57467, n57468, n57469, n57470, n57471, n57472, n57473,
n57474, n57475, n57476, n57477, n57478, n57479, n57480, n57481,
n57482, n57483, n57484, n57485, n57486, n57487, n57488, n57489,
n57490, n57491, n57492, n57493, n57494, n57495, n57496, n57497,
n57498, n57499, n57500, n57501, n57502, n57503, n57504, n57505,
n57506, n57507, n57508, n57509, n57510, n57511, n57512, n57513,
n57514, n57515, n57516, n57517, n57518, n57519, n57520, n57521,
n57522, n57523, n57524, n57525, n57526, n57527, n57528, n57529,
n57530, n57531, n57532, n57533, n57534, n57535, n57536, n57537,
n57538, n57539, n57540, n57541, n57542, n57543, n57544, n57545,
n57546, n57547, n57548, n57549, n57550, n57551, n57552, n57553,
n57554, n57555, n57556, n57557, n57558, n57559, n57560, n57561,
n57562, n57563, n57564, n57565, n57566, n57567, n57568, n57569,
n57570, n57571, n57572, n57573, n57574, n57575, n57576, n57577,
n57578, n57579, n57580, n57581, n57582, n57583, n57584, n57585,
n57586, n57587, n57588, n57589, n57590, n57591, n57592, n57593,
n57594, n57595, n57596, n57597, n57598, n57599, n57600, n57601,
n57602, n57603, n57604, n57605, n57606, n57607, n57608, n57609,
n57610, n57611, n57612, n57613, n57614, n57615, n57616, n57617,
n57618, n57619, n57620, n57621, n57622, n57623, n57624, n57625,
n57626, n57627, n57628, n57629, n57630, n57631, n57632, n57633,
n57634, n57635, n57636, n57637, n57638, n57639, n57640, n57641,
n57642, n57643, n57644, n57645, n57646, n57647, n57648, n57649,
n57650, n57651, n57652, n57653, n57654, n57655, n57656, n57657,
n57658, n57659, n57660, n57661, n57662, n57663, n57664, n57665,
n57666, n57667, n57668, n57669, n57670, n57671, n57672, n57673,
n57674, n57675, n57676, n57677, n57678, n57679, n57680, n57681,
n57682, n57683, n57684, n57685, n57686, n57687, n57688, n57689,
n57690, n57691, n57692, n57693, n57694, n57695, n57696, n57697,
n57698, n57699, n57700, n57701, n57702, n57703, n57704, n57705,
n57706, n57707, n57708, n57709, n57710, n57711, n57712, n57713,
n57714, n57715, n57716, n57717, n57718, n57719, n57720, n57721,
n57722, n57723, n57724, n57725, n57726, n57727, n57728, n57729,
n57730, n57731, n57732, n57733, n57734, n57735, n57736, n57737,
n57738, n57739, n57740, n57741, n57742, n57743, n57744, n57745,
n57746, n57747, n57748, n57749, n57750, n57751, n57752, n57753,
n57754, n57755, n57756, n57757, n57758, n57759, n57760, n57761,
n57762, n57763, n57764, n57765, n57766, n57767, n57768, n57769,
n57770, n57771, n57772, n57773, n57774, n57775, n57776, n57777,
n57778, n57779, n57780, n57781, n57782, n57783, n57784, n57785,
n57786, n57787, n57788, n57789, n57790, n57791, n57792, n57793,
n57794, n57795, n57796, n57797, n57798, n57799, n57800, n57801,
n57802, n57803, n57804, n57805, n57806, n57807, n57808, n57809,
n57810, n57811, n57812, n57813, n57814, n57815, n57816, n57817,
n57818, n57819, n57820, n57821, n57822, n57823, n57824, n57825,
n57826, n57827, n57828, n57829, n57830, n57831, n57832, n57833,
n57834, n57835, n57836, n57837, n57838, n57839, n57840, n57841,
n57842, n57843, n57844, n57845, n57846, n57847, n57848, n57850,
n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858,
n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866,
n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874,
n57875, n57876, n57877, n57878, n57879, n57880, n57881, n57882,
n57883, n57884, n57885, n57886, n57887, n57888, n57889, n57890,
n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898,
n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906,
n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914,
n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922,
n57923, n57924, n57925, n57926, n57927, n57928, n57929, n57930,
n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938,
n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946,
n57947, n57948, n57949, n57950, n57951, n57952, n57953, n57954,
n57955, n57956, n57957, n57958, n57959, n57960, n57961, n57962,
n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978,
n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986,
n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994,
n57995, n57996, n57997, n57998, n57999, n58000, n58001, n58002,
n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010,
n58012, n58013, n58014, n58015, n58016, n58017, n58018, n58019,
n58020, n58021, n58022, n58023, n58024, n58025, n58026, n58027,
n58028, n58029, n58030, n58031, n58032, n58033, n58034, n58035,
n58036, n58037, n58038, n58039, n58040, n58041, n58042, n58043,
n58044, n58045, n58046, n58047, n58048, n58049, n58050, n58051,
n58052, n58053, n58054, n58055, n58056, n58057, n58058, n58059,
n58060, n58061, n58062, n58063, n58064, n58065, n58066, n58067,
n58068, n58069, n58070, n58071, n58072, n58073, n58074, n58075,
n58077, n58078, n58079, n58080, n58081, n58082, n58083, n58084,
n58085, n58086, n58087, n58088, n58089, n58090, n58091, n58092,
n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100,
n58101, n58102, n58103, n58104, n58105, n58106, n58107, n58108,
n58109, n58110, n58111, n58112, n58113, n58114, n58115, n58116,
n58117, n58118, n58119, n58120, n58121, n58122, n58123, n58124,
n58125, n58126, n58127, n58128, n58129, n58130, n58131, n58132,
n58133, n58134, n58135, n58136, n58137, n58138, n58139, n58140,
n58141, n58142, n58143, n58144, n58145, n58146, n58147, n58148,
n58149, n58150, n58151, n58153, n58154, n58155, n58156, n58157,
n58158, n58159, n58160, n58161, n58162, n58163, n58164, n58165,
n58166, n58167, n58168, n58169, n58170, n58171, n58172, n58173,
n58174, n58175, n58176, n58177, n58178, n58179, n58180, n58181,
n58182, n58183, n58184, n58185, n58186, n58187, n58188, n58189,
n58190, n58191, n58192, n58193, n58194, n58195, n58196, n58197,
n58198, n58199, n58200, n58201, n58202, n58203, n58204, n58205,
n58206, n58207, n58208, n58209, n58210, n58211, n58212, n58213,
n58214, n58215, n58216, n58218, n58219, n58220, n58221, n58222,
n58223, n58224, n58225, n58226, n58227, n58228, n58229, n58230,
n58231, n58232, n58233, n58234, n58235, n58236, n58237, n58238,
n58239, n58240, n58241, n58242, n58243, n58244, n58245, n58246,
n58247, n58248, n58249, n58250, n58251, n58252, n58253, n58254,
n58255, n58256, n58257, n58258, n58259, n58260, n58261, n58262,
n58263, n58264, n58265, n58266, n58267, n58268, n58269, n58270,
n58271, n58272, n58273, n58274, n58275, n58276, n58277, n58278,
n58279, n58280, n58281, n58282, n58283, n58284, n58285, n58286,
n58287, n58288, n58289, n58290, n58291, n58292, n58293, n58294,
n58295, n58296, n58297, n58298, n58299, n58300, n58301, n58302,
n58303, n58304, n58305, n58306, n58307, n58308, n58309, n58310,
n58311, n58312, n58313, n58314, n58315, n58316, n58317, n58318,
n58319, n58320, n58321, n58322, n58323, n58324, n58325, n58326,
n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334,
n58335, n58336, n58337, n58338, n58339, n58340, n58341, n58342,
n58343, n58344, n58345, n58346, n58347, n58348, n58349, n58350,
n58351, n58352, n58353, n58354, n58355, n58356, n58357, n58358,
n58359, n58360, n58361, n58362, n58363, n58364, n58365, n58366,
n58367, n58368, n58369, n58370, n58371, n58372, n58373, n58374,
n58375, n58376, n58377, n58378, n58379, n58380, n58381, n58382,
n58383, n58384, n58385, n58386, n58387, n58388, n58389, n58390,
n58391, n58392, n58393, n58394, n58395, n58396, n58397, n58398,
n58399, n58400, n58401, n58402, n58403, n58404, n58405, n58406,
n58407, n58408, n58409, n58410, n58411, n58412, n58413, n58414,
n58415, n58416, n58417, n58418, n58419, n58420, n58421, n58422,
n58423, n58424, n58425, n58426, n58427, n58428, n58429, n58430,
n58431, n58432, n58433, n58434, n58435, n58436, n58437, n58438,
n58439, n58440, n58441, n58442, n58443, n58444, n58445, n58446,
n58447, n58448, n58449, n58450, n58451, n58452, n58453, n58454,
n58455, n58456, n58457, n58458, n58459, n58460, n58461, n58462,
n58463, n58464, n58465, n58466, n58467, n58468, n58469, n58470,
n58471, n58472, n58473, n58474, n58475, n58476, n58477, n58478,
n58479, n58480, n58481, n58482, n58483, n58484, n58485, n58486,
n58487, n58488, n58489, n58490, n58491, n58492, n58493, n58494,
n58495, n58496, n58497, n58498, n58499, n58500, n58501, n58502,
n58503, n58504, n58505, n58506, n58507, n58508, n58509, n58510,
n58511, n58512, n58513, n58514, n58515, n58516, n58517, n58518,
n58519, n58520, n58521, n58522, n58523, n58524, n58525, n58526,
n58527, n58528, n58529, n58530, n58531, n58532, n58533, n58534,
n58535, n58536, n58537, n58538, n58539, n58540, n58541, n58542,
n58543, n58544, n58545, n58546, n58547, n58548, n58549, n58550,
n58551, n58552, n58555, n58556, n58557, n58558, n58559, n58560,
n58561, n58562, n58563, n58564, n58565, n58566, n58567, n58568,
n58569, n58570, n58571, n58572, n58573, n58574, n58575, n58576,
n58577, n58578, n58579, n58580, n58581, n58582, n58583, n58584,
n58585, n58586, n58587, n58588, n58589, n58590, n58591, n58592,
n58593, n58594, n58595, n58596, n58597, n58598, n58599, n58600,
n58601, n58602, n58603, n58604, n58605, n58606, n58607, n58608,
n58609, n58610, n58611, n58612, n58613, n58614, n58615, n58616,
n58617, n58618, n58619, n58620, n58621, n58622, n58623, n58624,
n58625, n58626, n58627, n58628, n58629, n58630, n58631, n58632,
n58633, n58634, n58635, n58636, n58637, n58638, n58639, n58640,
n58641, n58642, n58643, n58644, n58645, n58646, n58647, n58648,
n58649, n58650, n58651, n58652, n58653, n58654, n58655, n58656,
n58657, n58658, n58659, n58660, n58661, n58662, n58663, n58664,
n58665, n58666, n58667, n58668, n58669, n58670, n58671, n58672,
n58673, n58674, n58675, n58676, n58677, n58678, n58679, n58680,
n58681, n58682, n58683, n58684, n58685, n58686, n58687, n58688,
n58689, n58690, n58691, n58692, n58693, n58694, n58695, n58696,
n58697, n58698, n58699, n58700, n58701, n58702, n58703, n58704,
n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712,
n58713, n58714, n58715, n58716, n58717, n58718, n58719, n58720,
n58721, n58722, n58723, n58724, n58725, n58726, n58727, n58728,
n58729, n58730, n58731, n58732, n58733, n58734, n58735, n58736,
n58737, n58738, n58739, n58740, n58741, n58742, n58743, n58744,
n58745, n58746, n58747, n58748, n58749, n58750, n58751, n58752,
n58753, n58754, n58755, n58756, n58757, n58758, n58759, n58760,
n58761, n58762, n58763, n58764, n58765, n58766, n58767, n58768,
n58769, n58770, n58771, n58772, n58773, n58774, n58775, n58776,
n58777, n58778, n58779, n58780, n58781, n58782, n58783, n58784,
n58785, n58786, n58787, n58788, n58789, n58790, n58791, n58792,
n58793, n58794, n58795, n58796, n58797, n58798, n58799, n58800,
n58801, n58802, n58803, n58804, n58805, n58806, n58807, n58808,
n58809, n58810, n58811, n58812, n58813, n58814, n58815, n58816,
n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824,
n58825, n58826, n58827, n58828, n58829, n58830, n58831, n58832,
n58833, n58834, n58835, n58836, n58837, n58838, n58839, n58840,
n58841, n58842, n58843, n58844, n58845, n58846, n58847, n58848,
n58849, n58850, n58851, n58852, n58853, n58854, n58855, n58856,
n58857, n58858, n58859, n58860, n58861, n58862, n58863, n58864,
n58865, n58866, n58867, n58868, n58869, n58870, n58871, n58872,
n58873, n58874, n58875, n58876, n58877, n58878, n58879, n58880,
n58881, n58882, n58883, n58884, n58885, n58886, n58887, n58888,
n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896,
n58897, n58898, n58899, n58900, n58901, n58902, n58903, n58904,
n58905, n58906, n58907, n58908, n58909, n58910, n58911, n58912,
n58913, n58914, n58915, n58916, n58917, n58918, n58919, n58920,
n58921, n58922, n58923, n58924, n58925, n58926, n58927, n58928,
n58929, n58930, n58931, n58932, n58933, n58934, n58935, n58936,
n58937, n58938, n58939, n58940, n58941, n58942, n58943, n58944,
n58945, n58946, n58947, n58948, n58949, n58950, n58951, n58952,
n58953, n58954, n58955, n58956, n58957, n58958, n58959, n58960,
n58961, n58962, n58963, n58964, n58965, n58966, n58967, n58968,
n58969, n58970, n58971, n58972, n58973, n58974, n58975, n58976,
n58977, n58978, n58979, n58980, n58981, n58982, n58983, n58984,
n58985, n58986, n58987, n58988, n58989, n58990, n58991, n58992,
n58993, n58994, n58995, n58996, n58997, n58998, n58999, n59000,
n59001, n59002, n59003, n59004, n59005, n59006, n59007, n59008,
n59009, n59010, n59011, n59012, n59013, n59014, n59015, n59016,
n59017, n59018, n59019, n59020, n59021, n59022, n59023, n59024,
n59025, n59026, n59027, n59028, n59029, n59030, n59031, n59032,
n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040,
n59041, n59042, n59043, n59044, n59045, n59046, n59047, n59048,
n59049, n59050, n59051, n59052, n59053, n59054, n59055, n59056,
n59057, n59058, n59059, n59060, n59061, n59062, n59063, n59064,
n59065, n59066, n59067, n59068, n59069, n59070, n59071, n59072,
n59073, n59074, n59075, n59076, n59077, n59078, n59079, n59080,
n59081, n59082, n59083, n59084, n59085, n59086, n59087, n59088,
n59089, n59090, n59091, n59092, n59093, n59094, n59095, n59096,
n59097, n59098, n59099, n59100, n59101, n59102, n59103, n59104,
n59105, n59106, n59107, n59108, n59109, n59110, n59111, n59112,
n59113, n59114, n59115, n59116, n59117, n59118, n59119, n59120,
n59121, n59122, n59123, n59124, n59125, n59126, n59127, n59128,
n59129, n59130, n59131, n59132, n59133, n59134, n59135, n59136,
n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59144,
n59146, n59147, n59148, n59149, n59150, n59151, n59152, n59153,
n59154, n59155, n59156, n59157, n59158, n59159, n59160, n59161,
n59162, n59163, n59164, n59165, n59166, n59167, n59168, n59169,
n59170, n59171, n59172, n59173, n59174, n59175, n59176, n59177,
n59178, n59179, n59180, n59181, n59182, n59183, n59184, n59185,
n59186, n59189, n59190, n59191, n59192, n59193, n59194, n59195,
n59196, n59197, n59198, n59199, n59200, n59201, n59202, n59203,
n59204, n59205, n59206, n59207, n59208, n59209, n59210, n59211,
n59212, n59213, n59214, n59215, n59216, n59217, n59218, n59219,
n59220, n59221, n59222, n59223, n59224, n59225, n59226, n59228,
n59229, n59230, n59231, n59232, n59233, n59234, n59235, n59236,
n59237, n59238, n59239, n59240, n59241, n59242, n59243, n59244,
n59245, n59246, n59247, n59248, n59249, n59250, n59251, n59252,
n59253, n59254, n59255, n59256, n59257, n59258, n59259, n59260,
n59261, n59262, n59263, n59264, n59265, n59266, n59267, n59268,
n59269, n59270, n59271, n59272, n59273, n59274, n59275, n59276,
n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284,
n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292,
n59293, n59294, n59295, n59296, n59297, n59298, n59299, n59300,
n59301, n59302, n59303, n59304, n59305, n59306, n59307, n59308,
n59309, n59310, n59311, n59312, n59313, n59314, n59315, n59316,
n59317, n59318, n59319, n59320, n59321, n59322, n59323, n59324,
n59325, n59326, n59327, n59328, n59329, n59330, n59331, n59332,
n59333, n59334, n59335, n59336, n59337, n59338, n59339, n59340,
n59341, n59342, n59343, n59344, n59345, n59346, n59347, n59348,
n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356,
n59357, n59358, n59359, n59360, n59361, n59362, n59363, n59364,
n59365, n59366, n59367, n59368, n59369, n59370, n59371, n59372,
n59373, n59374, n59375, n59376, n59378, n59379, n59380, n59381,
n59382, n59383, n59384, n59385, n59386, n59387, n59388, n59389,
n59390, n59391, n59392, n59393, n59394, n59395, n59396, n59397,
n59398, n59399, n59400, n59401, n59402, n59403, n59404, n59405,
n59406, n59407, n59408, n59409, n59410, n59411, n59412, n59413,
n59414, n59415, n59416, n59417, n59418, n59419, n59420, n59421,
n59422, n59423, n59424, n59425, n59426, n59427, n59428, n59429,
n59430, n59431, n59432, n59433, n59434, n59435, n59436, n59437,
n59438, n59439, n59440, n59441, n59442, n59443, n59444, n59445,
n59446, n59447, n59448, n59449, n59450, n59451, n59452, n59453,
n59454, n59455, n59456, n59457, n59458, n59459, n59460, n59461,
n59462, n59463, n59464, n59465, n59466, n59467, n59468, n59469,
n59470, n59471, n59472, n59473, n59474, n59476, n59477, n59478,
n59479, n59480, n59481, n59482, n59483, n59484, n59485, n59486,
n59487, n59488, n59489, n59490, n59491, n59492, n59493, n59494,
n59495, n59496, n59497, n59498, n59499, n59500, n59501, n59502,
n59503, n59504, n59505, n59506, n59507, n59508, n59509, n59510,
n59511, n59512, n59513, n59514, n59515, n59516, n59517, n59518,
n59519, n59520, n59521, n59522, n59523, n59524, n59525, n59526,
n59527, n59528, n59529, n59530, n59531, n59532, n59533, n59534,
n59535, n59536, n59537, n59538, n59539, n59540, n59541, n59542,
n59543, n59544, n59545, n59546, n59547, n59548, n59549, n59550,
n59551, n59552, n59553, n59554, n59555, n59556, n59557, n59558,
n59559, n59560, n59561, n59562, n59563, n59564, n59565, n59566,
n59567, n59568, n59569, n59570, n59571, n59572, n59573, n59574,
n59575, n59576, n59577, n59578, n59579, n59580, n59581, n59582,
n59583, n59584, n59585, n59586, n59587, n59588, n59589, n59590,
n59591, n59592, n59593, n59594, n59595, n59596, n59597, n59598,
n59599, n59600, n59601, n59602, n59603, n59604, n59605, n59606,
n59607, n59608, n59609, n59610, n59611, n59612, n59613, n59614,
n59615, n59616, n59617, n59618, n59619, n59620, n59621, n59622,
n59623, n59624, n59625, n59626, n59627, n59628, n59629, n59630,
n59631, n59632, n59633, n59634, n59635, n59636, n59637, n59638,
n59639, n59640, n59641, n59642, n59643, n59644, n59645, n59646,
n59647, n59648, n59649, n59650, n59651, n59652, n59653, n59654,
n59655, n59656, n59657, n59658, n59659, n59660, n59661, n59662,
n59663, n59664, n59665, n59666, n59667, n59668, n59669, n59670,
n59671, n59672, n59673, n59674, n59675, n59676, n59677, n59678,
n59679, n59680, n59681, n59682, n59683, n59684, n59685, n59686,
n59687, n59688, n59689, n59690, n59691, n59692, n59693, n59694,
n59695, n59696, n59697, n59698, n59699, n59700, n59701, n59702,
n59703, n59704, n59705, n59706, n59707, n59708, n59709, n59710,
n59711, n59712, n59713, n59714, n59715, n59716, n59717, n59718,
n59719, n59720, n59721, n59722, n59723, n59724, n59725, n59726,
n59727, n59728, n59729, n59730, n59731, n59732, n59733, n59734,
n59735, n59736, n59737, n59738, n59739, n59740, n59741, n59742,
n59743, n59744, n59745, n59746, n59747, n59748, n59749, n59750,
n59751, n59752, n59753, n59754, n59755, n59756, n59757, n59758,
n59759, n59760, n59761, n59762, n59763, n59764, n59765, n59766,
n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774,
n59775, n59776, n59777, n59778, n59779, n59780, n59781, n59782,
n59783, n59784, n59785, n59786, n59787, n59788, n59789, n59790,
n59791, n59792, n59793, n59794, n59795, n59796, n59797, n59798,
n59799, n59800, n59801, n59802, n59803, n59804, n59805, n59806,
n59807, n59808, n59809, n59810, n59811, n59812, n59813, n59814,
n59815, n59816, n59817, n59818, n59819, n59820, n59821, n59822,
n59823, n59824, n59825, n59826, n59827, n59828, n59829, n59830,
n59831, n59832, n59833, n59834, n59835, n59836, n59837, n59838,
n59839, n59840, n59841, n59842, n59843, n59844, n59845, n59846,
n59849, n59850, n59851, n59852, n59853, n59854, n59855, n59856,
n59857, n59858, n59859, n59860, n59861, n59862, n59863, n59864,
n59865, n59866, n59867, n59868, n59869, n59870, n59871, n59872,
n59873, n59874, n59875, n59876, n59877, n59878, n59879, n59880,
n59881, n59882, n59883, n59884, n59885, n59886, n59887, n59888,
n59889, n59890, n59891, n59892, n59893, n59894, n59895, n59896,
n59897, n59898, n59899, n59900, n59901, n59902, n59903, n59904,
n59905, n59906, n59907, n59908, n59909, n59910, n59911, n59912,
n59913, n59914, n59915, n59916, n59917, n59918, n59919, n59920,
n59921, n59922, n59923, n59924, n59925, n59926, n59927, n59928,
n59929, n59930, n59931, n59932, n59933, n59934, n59935, n59936,
n59937, n59938, n59939, n59940, n59941, n59942, n59943, n59944,
n59945, n59946, n59947, n59948, n59949, n59950, n59951, n59952,
n59953, n59954, n59955, n59956, n59957, n59958, n59959, n59960,
n59961, n59962, n59963, n59964, n59965, n59966, n59967, n59968,
n59969, n59970, n59971, n59972, n59973, n59974, n59975, n59976,
n59977, n59978, n59979, n59980, n59981, n59982, n59983, n59984,
n59985, n59986, n59987, n59988, n59989, n59990, n59991, n59992,
n59993, n59994, n59995, n59996, n59997, n59998, n59999, n60000,
n60001, n60002, n60003, n60004, n60005, n60006, n60007, n60008,
n60009, n60010, n60011, n60012, n60013, n60014, n60015, n60016,
n60017, n60018, n60019, n60020, n60021, n60022, n60023, n60024,
n60025, n60026, n60027, n60028, n60029, n60030, n60031, n60032,
n60033, n60034, n60035, n60036, n60037, n60038, n60039, n60040,
n60041, n60042, n60043, n60044, n60045, n60046, n60047, n60048,
n60049, n60050, n60051, n60052, n60053, n60054, n60055, n60056,
n60057, n60058, n60059, n60060, n60061, n60062, n60063, n60064,
n60065, n60066, n60067, n60068, n60069, n60070, n60071, n60072,
n60073, n60074, n60075, n60076, n60077, n60078, n60079, n60080,
n60081, n60082, n60083, n60084, n60085, n60086, n60087, n60088,
n60089, n60090, n60091, n60092, n60093, n60094, n60095, n60096,
n60097, n60098, n60099, n60100, n60101, n60102, n60103, n60104,
n60105, n60106, n60107, n60108, n60109, n60110, n60111, n60112,
n60113, n60114, n60115, n60116, n60117, n60118, n60119, n60120,
n60121, n60122, n60123, n60124, n60125, n60126, n60127, n60128,
n60129, n60130, n60131, n60132, n60133, n60134, n60135, n60136,
n60137, n60138, n60139, n60140, n60141, n60142, n60143, n60144,
n60145, n60146, n60147, n60148, n60149, n60150, n60151, n60152,
n60153, n60154, n60155, n60156, n60157, n60158, n60159, n60160,
n60161, n60162, n60163, n60164, n60165, n60166, n60167, n60168,
n60169, n60170, n60171, n60172, n60173, n60174, n60175, n60176,
n60177, n60178, n60179, n60180, n60181, n60182, n60183, n60184,
n60185, n60186, n60187, n60188, n60189, n60190, n60191, n60192,
n60193, n60194, n60195, n60196, n60197, n60198, n60199, n60200,
n60201, n60202, n60203, n60204, n60205, n60206, n60207, n60208,
n60209, n60210, n60211, n60212, n60213, n60214, n60215, n60216,
n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224,
n60225, n60226, n60227, n60228, n60229, n60230, n60231, n60232,
n60233, n60234, n60235, n60236, n60237, n60238, n60239, n60240,
n60241, n60242, n60243, n60244, n60245, n60246, n60247, n60248,
n60249, n60250, n60251, n60252, n60253, n60254, n60255, n60256,
n60257, n60258, n60259, n60260, n60261, n60262, n60263, n60264,
n60265, n60266, n60267, n60268, n60269, n60270, n60271, n60272,
n60273, n60274, n60275, n60276, n60277, n60278, n60279, n60280,
n60281, n60282, n60283, n60284, n60285, n60286, n60287, n60288,
n60289, n60290, n60291, n60292, n60293, n60294, n60295, n60296,
n60297, n60298, n60299, n60300, n60301, n60302, n60303, n60304,
n60305, n60306, n60307, n60308, n60309, n60310, n60311, n60312,
n60313, n60314, n60315, n60316, n60317, n60318, n60319, n60320,
n60321, n60322, n60323, n60324, n60325, n60326, n60327, n60328,
n60329, n60330, n60331, n60332, n60333, n60334, n60335, n60336,
n60337, n60338, n60339, n60340, n60341, n60342, n60343, n60344,
n60345, n60346, n60347, n60348, n60349, n60350, n60351, n60352,
n60353, n60354, n60355, n60356, n60357, n60358, n60359, n60360,
n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368,
n60369, n60370, n60371, n60372, n60373, n60374, n60375, n60376,
n60377, n60378, n60379, n60380, n60381, n60382, n60383, n60384,
n60385, n60386, n60387, n60388, n60389, n60390, n60391, n60392,
n60393, n60394, n60395, n60396, n60397, n60398, n60399, n60400,
n60401, n60402, n60403, n60404, n60405, n60406, n60407, n60408,
n60409, n60410, n60411, n60412, n60413, n60414, n60415, n60416,
n60417, n60418, n60419, n60420, n60421, n60422, n60423, n60424,
n60425, n60426, n60427, n60428, n60429, n60430, n60431, n60432,
n60433, n60434, n60435, n60436, n60437, n60438, n60439, n60440,
n60441, n60442, n60443, n60444, n60445, n60446, n60447, n60448,
n60449, n60450, n60451, n60452, n60453, n60454, n60455, n60456,
n60457, n60458, n60459, n60460, n60461, n60462, n60463, n60464,
n60465, n60466, n60467, n60468, n60469, n60470, n60471, n60472,
n60473, n60474, n60475, n60476, n60477, n60478, n60479, n60480,
n60481, n60482, n60483, n60484, n60485, n60486, n60487, n60488,
n60489, n60490, n60491, n60492, n60493, n60494, n60495, n60496,
n60497, n60498, n60499, n60500, n60501, n60502, n60503, n60504,
n60505, n60506, n60507, n60508, n60509, n60510, n60511, n60512,
n60513, n60514, n60515, n60516, n60517, n60518, n60519, n60520,
n60521, n60522, n60523, n60524, n60525, n60526, n60527, n60528,
n60529, n60530, n60531, n60532, n60533, n60534, n60535, n60536,
n60537, n60538, n60539, n60540, n60541, n60542, n60543, n60544,
n60545, n60546, n60547, n60548, n60549, n60550, n60551, n60552,
n60553, n60554, n60555, n60556, n60557, n60558, n60559, n60560,
n60561, n60562, n60563, n60564, n60565, n60566, n60567, n60568,
n60569, n60570, n60571, n60572, n60573, n60574, n60575, n60576,
n60577, n60578, n60579, n60580, n60581, n60582, n60583, n60584,
n60585, n60586, n60587, n60588, n60589, n60590, n60591, n60592,
n60593, n60594, n60595, n60596, n60597, n60598, n60599, n60600,
n60601, n60602, n60603, n60604, n60605, n60606, n60607, n60608,
n60609, n60610, n60611, n60612, n60613, n60614, n60615, n60616,
n60617, n60618, n60619, n60620, n60621, n60622, n60623, n60624,
n60625, n60626, n60627, n60628, n60629, n60630, n60631, n60632,
n60633, n60634, n60635, n60636, n60637, n60638, n60639, n60640,
n60641, n60642, n60643, n60644, n60645, n60646, n60647, n60648,
n60649, n60650, n60651, n60652, n60653, n60654, n60655, n60656,
n60657, n60658, n60659, n60660, n60661, n60662, n60663, n60664,
n60665, n60666, n60667, n60668, n60669, n60670, n60671, n60672,
n60673, n60674, n60675, n60676, n60677, n60678, n60679, n60680,
n60681, n60682, n60683, n60684, n60685, n60686, n60687, n60688,
n60689, n60690, n60691, n60692, n60693, n60694, n60695, n60696,
n60697, n60698, n60699, n60700, n60701, n60702, n60703, n60704,
n60705, n60706, n60707, n60708, n60709, n60710, n60711, n60712,
n60713, n60714, n60715, n60716, n60717, n60718, n60719, n60720,
n60721, n60722, n60723, n60724, n60725, n60726, n60727, n60728,
n60729, n60730, n60731, n60732, n60733, n60734, n60735, n60736,
n60737, n60738, n60739, n60740, n60741, n60742, n60743, n60744,
n60745, n60746, n60747, n60748, n60749, n60750, n60751, n60752,
n60753, n60754, n60755, n60756, n60757, n60758, n60759, n60760,
n60761, n60762, n60763, n60764, n60765, n60766, n60767, n60768,
n60769, n60770, n60771, n60772, n60773, n60774, n60775, n60776,
n60777, n60778, n60779, n60780, n60781, n60782, n60783, n60784,
n60785, n60786, n60787, n60788, n60789, n60790, n60791, n60792,
n60793, n60794, n60795, n60796, n60797, n60798, n60799, n60800,
n60801, n60802, n60803, n60804, n60805, n60806, n60807, n60808,
n60809, n60810, n60811, n60812, n60813, n60814, n60815, n60816,
n60817, n60818, n60819, n60820, n60821, n60822, n60823, n60824,
n60825, n60826, n60827, n60828, n60829, n60830, n60831, n60832,
n60833, n60834, n60835, n60836, n60837, n60838, n60839, n60840,
n60841, n60842, n60843, n60844, n60845, n60846, n60847, n60848,
n60849, n60850, n60851, n60852, n60853, n60854, n60855, n60856,
n60857, n60858, n60859, n60860, n60861, n60862, n60863, n60864,
n60865, n60866, n60867, n60868, n60869, n60870, n60871, n60872,
n60873, n60874, n60875, n60876, n60877, n60878, n60879, n60880,
n60881, n60882, n60883, n60884, n60885, n60886, n60887, n60888,
n60889, n60890, n60891, n60892, n60893, n60894, n60895, n60896,
n60897, n60898, n60899, n60900, n60901, n60902, n60903, n60904,
n60905, n60906, n60907, n60908, n60909, n60910, n60911, n60912,
n60913, n60914, n60915, n60916, n60917, n60918, n60919, n60920,
n60921, n60922, n60923, n60924, n60925, n60926, n60927, n60928,
n60929, n60930, n60931, n60932, n60933, n60934, n60935, n60936,
n60937, n60938, n60939, n60940, n60941, n60942, n60943, n60944,
n60945, n60946, n60947, n60948, n60949, n60950, n60951, n60952,
n60953, n60954, n60955, n60956, n60957, n60958, n60959, n60960,
n60961, n60962, n60963, n60964, n60965, n60966, n60967, n60968,
n60969, n60970, n60971, n60972, n60973, n60974, n60975, n60976,
n60977, n60978, n60979, n60980, n60981, n60982, n60983, n60984,
n60985, n60986, n60987, n60988, n60989, n60990, n60991, n60992,
n60993, n60994, n60995, n60996, n60997, n60998, n60999, n61000,
n61001, n61002, n61003, n61004, n61005, n61006, n61007, n61008,
n61009, n61010, n61011, n61012, n61013, n61014, n61015, n61016,
n61017, n61018, n61019, n61020, n61021, n61022, n61023, n61024,
n61025, n61026, n61027, n61028, n61029, n61030, n61031, n61032,
n61033, n61034, n61035, n61036, n61037, n61038, n61039, n61040,
n61041, n61042, n61043, n61044, n61045, n61046, n61047, n61048,
n61049, n61050, n61051, n61052, n61053, n61054, n61055, n61056,
n61057, n61058, n61059, n61060, n61061, n61062, n61063, n61064,
n61065, n61066, n61067, n61068, n61069, n61070, n61071, n61072,
n61073, n61074, n61075, n61076, n61077, n61078, n61079, n61080,
n61081, n61082, n61083, n61084, n61085, n61086, n61087, n61088,
n61089, n61090, n61091, n61092, n61093, n61094, n61095, n61096,
n61097, n61098, n61099, n61100, n61101, n61102, n61103, n61104,
n61105, n61106, n61107, n61108, n61109, n61110, n61111, n61112,
n61113, n61114, n61115, n61116, n61117, n61118, n61119, n61120,
n61121, n61122, n61123, n61124, n61125, n61126, n61127, n61128,
n61129, n61130, n61131, n61132, n61133, n61134, n61135, n61136,
n61137, n61138, n61139, n61140, n61141, n61142, n61143, n61144,
n61145, n61146, n61147, n61148, n61149, n61150, n61151, n61152,
n61153, n61154, n61155, n61156, n61157, n61158, n61159, n61160,
n61161, n61162, n61163, n61164, n61165, n61166, n61167, n61168,
n61169, n61170, n61171, n61172, n61173, n61174, n61175, n61176,
n61177, n61178, n61179, n61180, n61181, n61182, n61183, n61184,
n61185, n61186, n61187, n61188, n61189, n61190, n61191, n61192,
n61193, n61194, n61195, n61196, n61197, n61198, n61199, n61200,
n61201, n61202, n61203, n61204, n61205, n61206, n61207, n61208,
n61209, n61210, n61211, n61212, n61213, n61214, n61215, n61216,
n61217, n61218, n61219, n61220, n61221, n61222, n61223, n61224,
n61225, n61226, n61227, n61228, n61229, n61230, n61231, n61232,
n61233, n61234, n61235, n61236, n61237, n61238, n61239, n61240,
n61241, n61242, n61243, n61244, n61245, n61246, n61247, n61248,
n61249, n61250, n61251, n61252, n61253, n61254, n61255, n61256,
n61257, n61258, n61259, n61260, n61261, n61262, n61263, n61264,
n61265, n61266, n61267, n61268, n61269, n61270, n61271, n61272,
n61273, n61274, n61275, n61276, n61277, n61278, n61279, n61280,
n61281, n61282, n61283, n61284, n61285, n61286, n61287, n61288,
n61289, n61290, n61291, n61292, n61293, n61294, n61295, n61296,
n61297, n61298, n61299, n61300, n61301, n61302, n61303, n61304,
n61305, n61306, n61307, n61308, n61309, n61310, n61311, n61312,
n61313, n61314, n61315, n61316, n61317, n61318, n61319, n61320,
n61321, n61322, n61323, n61324, n61325, n61326, n61327, n61328,
n61329, n61330, n61331, n61332, n61333, n61334, n61335, n61336,
n61337, n61338, n61339, n61340, n61341, n61342, n61343, n61344,
n61345, n61346, n61347, n61348, n61349, n61350, n61351, n61352,
n61353, n61354, n61355, n61356, n61357, n61358, n61359, n61360,
n61361, n61362, n61363, n61364, n61365, n61366, n61367, n61368,
n61369, n61370, n61371, n61372, n61373, n61374, n61375, n61376,
n61377, n61378, n61379, n61380, n61381, n61382, n61383, n61384,
n61385, n61386, n61387, n61388, n61389, n61390, n61391, n61392,
n61393, n61394, n61395, n61396, n61397, n61398, n61399, n61400,
n61401, n61402, n61403, n61404, n61405, n61406, n61407, n61408,
n61409, n61410, n61411, n61412, n61413, n61414, n61415, n61416,
n61417, n61418, n61419, n61420, n61421, n61422, n61423, n61424,
n61425, n61426, n61427, n61428, n61429, n61430, n61431, n61432,
n61433, n61434, n61435, n61436, n61437, n61438, n61439, n61440,
n61441, n61442, n61443, n61444, n61445, n61446, n61447, n61448,
n61449, n61450, n61451, n61452, n61453, n61454, n61455, n61456,
n61457, n61458, n61459, n61460, n61461, n61462, n61463, n61464,
n61465, n61466, n61467, n61468, n61469, n61470, n61471, n61472,
n61473, n61474, n61475, n61476, n61477, n61478, n61479, n61480,
n61481, n61482, n61483, n61484, n61485, n61486, n61487, n61488,
n61489, n61490, n61491, n61492, n61493, n61494, n61495, n61496,
n61497, n61498, n61499, n61500, n61501, n61502, n61503, n61504,
n61505, n61506, n61507, n61508, n61509, n61510, n61511, n61512,
n61513, n61514, n61515, n61516, n61517, n61518, n61519, n61520,
n61521, n61522, n61523, n61524, n61525, n61526, n61527, n61528,
n61529, n61530, n61531, n61532, n61533, n61534, n61535, n61536,
n61537, n61538, n61539, n61540, n61541, n61542, n61543, n61544,
n61545, n61546, n61547, n61548, n61549, n61550, n61551, n61552,
n61553, n61554, n61555, n61556, n61557, n61558, n61559, n61560,
n61561, n61562, n61563, n61564, n61565, n61566, n61567, n61568,
n61569, n61570, n61571, n61572, n61573, n61574, n61575, n61576,
n61577, n61578, n61579, n61580, n61581, n61582, n61583, n61584,
n61585, n61586, n61587, n61588, n61589, n61590, n61591, n61592,
n61593, n61594, n61595, n61596, n61597, n61598, n61599, n61600,
n61601, n61602, n61603, n61604, n61605, n61606, n61607, n61608,
n61609, n61610, n61611, n61612, n61613, n61614, n61615, n61616,
n61617, n61618, n61619, n61620, n61621, n61622, n61623, n61624,
n61625, n61626, n61627, n61628, n61629, n61630, n61631, n61632,
n61633, n61634, n61635, n61636, n61637, n61638, n61639, n61640,
n61641, n61642, n61643, n61644, n61645, n61646, n61647, n61648,
n61649, n61650, n61651, n61652, n61653, n61654, n61655, n61656,
n61657, n61658, n61659, n61660, n61661, n61662, n61663, n61664,
n61665, n61666, n61667, n61668, n61669, n61670, n61671, n61672,
n61673, n61674, n61675, n61676, n61677, n61678, n61679, n61680,
n61681, n61682, n61683, n61684, n61685, n61686, n61687, n61688,
n61689, n61690, n61691, n61692, n61693, n61694, n61695, n61696,
n61697, n61698, n61699, n61700, n61701, n61702, n61703, n61704,
n61705, n61706, n61707, n61708, n61709, n61710, n61711, n61712,
n61713, n61714, n61715, n61716, n61717, n61718, n61719, n61720,
n61721, n61722, n61723, n61724, n61725, n61726, n61727, n61728,
n61729, n61730, n61731, n61732, n61733, n61734, n61735, n61736,
n61737, n61738, n61739, n61740, n61741, n61742, n61743, n61744,
n61745, n61746, n61747, n61748, n61749, n61750, n61751, n61752,
n61753, n61754, n61755, n61756, n61757, n61758, n61759, n61760,
n61761, n61762, n61763, n61764, n61765, n61766, n61767, n61768,
n61769, n61770, n61771, n61772, n61773, n61774, n61775, n61776,
n61777, n61778, n61779, n61780, n61781, n61782, n61783, n61784,
n61785, n61786, n61787, n61788, n61789, n61790, n61791, n61792,
n61793, n61794, n61795, n61796, n61797, n61798, n61799, n61800,
n61801, n61802, n61803, n61804, n61805, n61806, n61807, n61808,
n61809, n61810, n61811, n61812, n61813, n61814, n61815, n61816,
n61817, n61818, n61819, n61820, n61821, n61822, n61823, n61824,
n61825, n61826, n61827, n61828, n61829, n61830, n61831, n61832,
n61833, n61834, n61835, n61836, n61837, n61838, n61839, n61840,
n61841, n61842, n61843, n61844, n61845, n61846, n61847, n61848,
n61849, n61850, n61851, n61852, n61853, n61854, n61855, n61856,
n61857, n61858, n61859, n61860, n61861, n61862, n61863, n61864,
n61865, n61866, n61867, n61868, n61869, n61870, n61871, n61872,
n61873, n61874, n61875, n61876, n61877, n61878, n61879, n61880,
n61881, n61882, n61883, n61884, n61885, n61886, n61887, n61888,
n61889, n61890, n61891, n61892, n61893, n61894, n61895, n61896,
n61897, n61898, n61899, n61900, n61901, n61902, n61903, n61904,
n61905, n61906, n61907, n61908, n61909, n61910, n61911, n61912,
n61913, n61914, n61915, n61916, n61917, n61918, n61919, n61920,
n61921, n61922, n61923, n61924, n61925, n61926, n61927, n61928,
n61929, n61930, n61931, n61932, n61933, n61934, n61935, n61936,
n61937, n61938, n61939, n61940, n61941, n61942, n61943, n61944,
n61945, n61946, n61947, n61948, n61949, n61950, n61951, n61952,
n61953, n61954, n61955, n61956, n61957, n61958, n61959, n61960,
n61961, n61962, n61963, n61964, n61965, n61966, n61967, n61968,
n61969, n61970, n61971, n61972, n61973, n61974, n61975, n61976,
n61977, n61978, n61979, n61980, n61981, n61982, n61983, n61984,
n61985, n61986, n61987, n61988, n61989, n61990, n61991, n61992,
n61993, n61994, n61995, n61996, n61997, n61998, n61999, n62000,
n62001, n62002, n62003, n62004, n62005, n62006, n62007, n62008,
n62009, n62010, n62011, n62012, n62013, n62014, n62015, n62016,
n62017, n62018, n62019, n62020, n62021, n62022, n62023, n62024,
n62025, n62026, n62027, n62028, n62029, n62030, n62031, n62032,
n62033, n62034, n62035, n62036, n62037, n62038, n62039, n62040,
n62041, n62042, n62043, n62044, n62045, n62046, n62047, n62048,
n62049, n62050, n62051, n62052, n62053, n62054, n62055, n62056,
n62057, n62058, n62059, n62060, n62061, n62062, n62063, n62064,
n62065, n62066, n62067, n62068, n62069, n62070, n62071, n62072,
n62073, n62074, n62075, n62076, n62077, n62078, n62079, n62080,
n62081, n62082, n62083, n62084, n62085, n62086, n62087, n62088,
n62089, n62090, n62091, n62092, n62093, n62094, n62095, n62096,
n62097, n62098, n62099, n62100, n62101, n62102, n62103, n62104,
n62105, n62106, n62107, n62108, n62109, n62110, n62111, n62112,
n62113, n62114, n62115, n62116, n62117, n62118, n62119, n62120,
n62121, n62122, n62123, n62124, n62125, n62126, n62127, n62128,
n62129, n62130, n62131, n62132, n62133, n62134, n62135, n62136,
n62137, n62138, n62139, n62140, n62141, n62142, n62143, n62144,
n62145, n62146, n62147, n62148, n62149, n62150, n62151, n62152,
n62153, n62154, n62155, n62156, n62157, n62158, n62159, n62160,
n62161, n62162, n62163, n62164, n62165, n62166, n62167, n62168,
n62169, n62170, n62171, n62172, n62173, n62174, n62175, n62176,
n62177, n62178, n62179, n62180, n62181, n62182, n62183, n62184,
n62185, n62186, n62187, n62188, n62189, n62190, n62191, n62192,
n62193, n62194, n62195, n62196, n62197, n62198, n62199, n62200,
n62201, n62202, n62203, n62204, n62205, n62206, n62207, n62208,
n62209, n62210, n62211, n62212, n62214, n62215, n62216, n62217,
n62218, n62219, n62220, n62221, n62222, n62223, n62224, n62225,
n62226, n62227, n62228, n62229, n62230, n62231, n62232, n62233,
n62234, n62235, n62236, n62237, n62238, n62239, n62240, n62241,
n62242, n62243, n62244, n62245, n62246, n62247, n62248, n62249,
n62250, n62251, n62252, n62253, n62254, n62255, n62256, n62257,
n62258, n62259, n62260, n62261, n62262, n62263, n62264, n62265,
n62266, n62267, n62268, n62269, n62270, n62271, n62272, n62273,
n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281,
n62282, n62283, n62284, n62285, n62286, n62287, n62288, n62289,
n62290, n62291, n62292, n62293, n62294, n62295, n62296, n62297,
n62298, n62299, n62300, n62301, n62302, n62303, n62304, n62305,
n62306, n62307, n62308, n62309, n62310, n62311, n62312, n62313,
n62314, n62315, n62316, n62317, n62318, n62319, n62320, n62321,
n62322, n62325, n62326, n62327, n62328, n62329, n62330, n62331,
n62332, n62333, n62334, n62335, n62336, n62337, n62338, n62339,
n62340, n62341, n62342, n62343, n62344, n62345, n62346, n62347,
n62348, n62349, n62350, n62351, n62352, n62353, n62354, n62355,
n62356, n62357, n62358, n62359, n62360, n62361, n62362, n62363,
n62364, n62365, n62366, n62367, n62368, n62369, n62370, n62371,
n62372, n62373, n62374, n62375, n62376, n62377, n62378, n62379,
n62380, n62381, n62382, n62383, n62384, n62385, n62386, n62387,
n62388, n62389, n62390, n62391, n62392, n62393, n62394, n62395,
n62396, n62397, n62398, n62399, n62400, n62401, n62402, n62403,
n62404, n62405, n62406, n62407, n62408, n62409, n62410, n62411,
n62412, n62413, n62414, n62415, n62416, n62417, n62418, n62419,
n62420, n62421, n62422, n62423, n62424, n62425, n62426, n62427,
n62428, n62429, n62430, n62431, n62432, n62433, n62434, n62435,
n62436, n62437, n62438, n62439, n62440, n62441, n62442, n62443,
n62444, n62445, n62446, n62447, n62448, n62449, n62450, n62451,
n62452, n62453, n62454, n62455, n62456, n62457, n62458, n62459,
n62460, n62461, n62462, n62463, n62464, n62465, n62466, n62467,
n62468, n62469, n62470, n62471, n62472, n62473, n62474, n62475,
n62476, n62477, n62478, n62479, n62480, n62481, n62482, n62483,
n62484, n62485, n62486, n62487, n62488, n62489, n62490, n62491,
n62492, n62493, n62494, n62496, n62497, n62498, n62499, n62500,
n62501, n62502, n62503, n62504, n62505, n62506, n62507, n62508,
n62509, n62510, n62511, n62512, n62513, n62514, n62515, n62516,
n62517, n62518, n62519, n62520, n62521, n62522, n62523, n62524,
n62525, n62526, n62527, n62528, n62529, n62530, n62531, n62532,
n62533, n62534, n62535, n62536, n62537, n62538, n62539, n62540,
n62541, n62542, n62543, n62544, n62545, n62546, n62547, n62548,
n62549, n62550, n62551, n62552, n62553, n62554, n62555, n62556,
n62557, n62558, n62559, n62560, n62561, n62562, n62563, n62564,
n62565, n62566, n62567, n62568, n62569, n62570, n62571, n62572,
n62575, n62576, n62577, n62578, n62579, n62580, n62581, n62582,
n62583, n62584, n62585, n62586, n62587, n62588, n62589, n62590,
n62591, n62592, n62593, n62594, n62595, n62596, n62597, n62598,
n62599, n62600, n62601, n62602, n62603, n62604, n62605, n62606,
n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614,
n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622,
n62623, n62624, n62625, n62626, n62627, n62628, n62629, n62630,
n62631, n62632, n62633, n62634, n62635, n62636, n62637, n62638,
n62639, n62640, n62641, n62642, n62643, n62644, n62645, n62646,
n62647, n62648, n62649, n62651, n62652, n62653, n62654, n62655,
n62656, n62657, n62658, n62659, n62660, n62661, n62662, n62663,
n62664, n62665, n62666, n62667, n62668, n62669, n62670, n62671,
n62672, n62673, n62674, n62675, n62676, n62677, n62678, n62679,
n62680, n62681, n62682, n62683, n62684, n62685, n62686, n62687,
n62688, n62689, n62690, n62691, n62692, n62693, n62694, n62695,
n62696, n62697, n62698, n62699, n62700, n62701, n62702, n62703,
n62704, n62705, n62706, n62707, n62708, n62709, n62710, n62711,
n62712, n62713, n62714, n62715, n62716, n62717, n62718, n62719,
n62720, n62721, n62722, n62723, n62724, n62725, n62726, n62727,
n62728, n62729, n62730, n62731, n62732, n62733, n62734, n62735,
n62736, n62737, n62738, n62739, n62740, n62741, n62742, n62743,
n62744, n62745, n62746, n62747, n62748, n62749, n62750, n62751,
n62752, n62753, n62754, n62755, n62756, n62757, n62758, n62759,
n62760, n62761, n62762, n62763, n62764, n62765, n62766, n62767,
n62768, n62769, n62770, n62771, n62772, n62773, n62774, n62775,
n62776, n62777, n62778, n62779, n62780, n62781, n62782, n62783,
n62784, n62785, n62786, n62787, n62788, n62789, n62790, n62791,
n62792, n62793, n62794, n62795, n62796, n62797, n62798, n62799,
n62800, n62801, n62802, n62803, n62804, n62805, n62806, n62807,
n62808, n62809, n62810, n62811, n62812, n62813, n62814, n62815,
n62816, n62817, n62818, n62819, n62820, n62821, n62822, n62823,
n62824, n62825, n62826, n62827, n62828, n62829, n62830, n62831,
n62832, n62833, n62834, n62835, n62836, n62837, n62838, n62839,
n62840, n62841, n62842, n62843, n62844, n62845, n62846, n62847,
n62848, n62849, n62850, n62851, n62852, n62853, n62854, n62855,
n62856, n62857, n62858, n62859, n62860, n62861, n62862, n62863,
n62864, n62865, n62866, n62867, n62868, n62869, n62870, n62871,
n62872, n62873, n62874, n62875, n62876, n62877, n62878, n62879,
n62880, n62881, n62882, n62883, n62884, n62885, n62886, n62887,
n62888, n62889, n62890, n62891, n62892, n62893, n62894, n62895,
n62896, n62897, n62898, n62899, n62900, n62901, n62903, n62904,
n62905, n62906, n62907, n62908, n62909, n62910, n62911, n62912,
n62913, n62914, n62915, n62916, n62917, n62918, n62919, n62920,
n62921, n62922, n62923, n62924, n62925, n62926, n62927, n62928,
n62929, n62930, n62931, n62932, n62933, n62934, n62935, n62936,
n62937, n62938, n62939, n62940, n62941, n62942, n62943, n62944,
n62945, n62946, n62947, n62948, n62949, n62950, n62951, n62952,
n62953, n62954, n62955, n62956, n62957, n62958, n62959, n62960,
n62961, n62962, n62963, n62964, n62965, n62966, n62967, n62968,
n62969, n62970, n62973, n62974, n62975, n62978, n62979, n62980,
n62981, n62982, n62983, n62984, n62985, n62986, n62987, n62988,
n62989, n62990, n62991, n62992, n62993, n62994, n62995, n62996,
n62997, n62998, n62999, n63000, n63001, n63002, n63003, n63004,
n63005, n63006, n63007, n63008, n63009, n63010, n63011, n63012,
n63013, n63014, n63015, n63016, n63017, n63018, n63019, n63020,
n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028,
n63029, n63030, n63031, n63032, n63033, n63034, n63035, n63036,
n63037, n63038, n63039, n63040, n63041, n63042, n63043, n63044,
n63045, n63046, n63047, n63048, n63049, n63050, n63051, n63052,
n63053, n63054, n63055, n63056, n63057, n63058, n63059, n63060,
n63061, n63062, n63063, n63064, n63065, n63066, n63067, n63068,
n63069, n63070, n63071, n63072, n63073, n63074, n63075, n63076,
n63077, n63078, n63079, n63080, n63081, n63082, n63083, n63084,
n63085, n63086, n63087, n63088, n63089, n63090, n63091, n63092,
n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100,
n63101, n63102, n63103, n63104, n63105, n63106, n63107, n63108,
n63109, n63110, n63111, n63112, n63113, n63114, n63115, n63116,
n63117, n63118, n63119, n63120, n63121, n63122, n63123, n63124,
n63125, n63126, n63127, n63128, n63129, n63130, n63131, n63132,
n63133, n63134, n63135, n63136, n63137, n63138, n63139, n63140,
n63141, n63142, n63143, n63144, n63145, n63146, n63147, n63148,
n63149, n63150, n63151, n63152, n63153, n63154, n63155, n63156,
n63157, n63158, n63159, n63160, n63161, n63162, n63163, n63164,
n63165, n63167, n63168, n63169, n63170, n63171, n63172, n63173,
n63174, n63175, n63176, n63177, n63178, n63179, n63180, n63181,
n63182, n63183, n63184, n63185, n63186, n63187, n63188, n63189,
n63190, n63191, n63192, n63193, n63194, n63195, n63196, n63197,
n63198, n63199, n63200, n63201, n63202, n63203, n63204, n63205,
n63206, n63207, n63208, n63209, n63210, n63211, n63212, n63213,
n63214, n63215, n63216, n63218, n63219, n63220, n63221, n63222,
n63223, n63224, n63225, n63226, n63227, n63228, n63229, n63230,
n63231, n63232, n63233, n63234, n63235, n63236, n63237, n63238,
n63239, n63240, n63241, n63242, n63243, n63244, n63245, n63246,
n63247, n63248, n63249, n63250, n63251, n63252, n63253, n63254,
n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262,
n63263, n63264, n63265, n63266, n63267, n63268, n63269, n63270,
n63271, n63272, n63273, n63274, n63275, n63276, n63277, n63278,
n63279, n63280, n63281, n63282, n63283, n63284, n63285, n63288,
n63289, n63290, n63291, n63292, n63293, n63294, n63295, n63296,
n63299, n63300, n63301, n63302, n63303, n63304, n63305, n63306,
n63307, n63308, n63309, n63310, n63311, n63312, n63313, n63314,
n63315, n63316, n63317, n63318, n63319, n63320, n63321, n63322,
n63323, n63324, n63325, n63326, n63327, n63328, n63329, n63330,
n63331, n63332, n63333, n63334, n63335, n63336, n63337, n63338,
n63339, n63340, n63341, n63342, n63343, n63344, n63345, n63346,
n63347, n63348, n63349, n63350, n63351, n63352, n63353, n63354,
n63355, n63356, n63357, n63358, n63359, n63360, n63361, n63362,
n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370,
n63371, n63372, n63373, n63374, n63375, n63376, n63377, n63378,
n63379, n63380, n63381, n63382, n63383, n63384, n63385, n63386,
n63387, n63388, n63389, n63390, n63391, n63392, n63393, n63394,
n63395, n63396, n63397, n63398, n63399, n63400, n63401, n63402,
n63403, n63404, n63405, n63406, n63407, n63408, n63409, n63410,
n63411, n63412, n63414, n63415, n63416, n63417, n63418, n63419,
n63420, n63421, n63422, n63423, n63424, n63425, n63426, n63427,
n63428, n63429, n63430, n63431, n63432, n63433, n63434, n63435,
n63436, n63437, n63438, n63439, n63440, n63441, n63442, n63443,
n63444, n63445, n63446, n63447, n63448, n63449, n63450, n63451,
n63452, n63453, n63454, n63455, n63456, n63457, n63459, n63460,
n63461, n63462, n63463, n63464, n63465, n63466, n63467, n63468,
n63469, n63470, n63471, n63472, n63473, n63474, n63475, n63476,
n63477, n63478, n63479, n63480, n63481, n63482, n63483, n63484,
n63485, n63486, n63487, n63488, n63489, n63490, n63491, n63492,
n63493, n63494, n63495, n63496, n63497, n63498, n63499, n63500,
n63501, n63502, n63503, n63504, n63505, n63506, n63507, n63508,
n63509, n63510, n63511, n63512, n63513, n63514, n63515, n63516,
n63517, n63518, n63519, n63520, n63521, n63522, n63523, n63524,
n63525, n63526, n63527, n63528, n63529, n63530, n63531, n63532,
n63533, n63534, n63535, n63536, n63537, n63538, n63539, n63540,
n63541, n63542, n63543, n63544, n63545, n63546, n63547, n63548,
n63549, n63550, n63551, n63552, n63553, n63554, n63555, n63556,
n63557, n63558, n63559, n63560, n63561, n63562, n63563, n63564,
n63565, n63566, n63567, n63568, n63569, n63570, n63571, n63572,
n63573, n63574, n63575, n63576, n63577, n63578, n63579, n63580,
n63581, n63582, n63583, n63584, n63585, n63586, n63587, n63588,
n63589, n63590, n63591, n63592, n63593, n63594, n63595, n63596,
n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604,
n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612,
n63613, n63614, n63615, n63616, n63617, n63618, n63619, n63620,
n63621, n63622, n63623, n63624, n63625, n63626, n63627, n63628,
n63629, n63630, n63631, n63632, n63633, n63634, n63635, n63636,
n63637, n63638, n63639, n63640, n63641, n63642, n63643, n63644,
n63645, n63646, n63647, n63648, n63649, n63650, n63651, n63652,
n63653, n63654, n63655, n63656, n63657, n63658, n63659, n63660,
n63661, n63662, n63663, n63664, n63665, n63666, n63667, n63668,
n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676,
n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684,
n63685, n63686, n63687, n63688, n63689, n63690, n63691, n63692,
n63693, n63694, n63695, n63696, n63697, n63698, n63699, n63700,
n63701, n63702, n63703, n63704, n63705, n63706, n63707, n63708,
n63709, n63710, n63711, n63712, n63713, n63714, n63715, n63716,
n63717, n63718, n63719, n63720, n63721, n63722, n63723, n63724,
n63725, n63726, n63727, n63728, n63729, n63730, n63731, n63732,
n63733, n63734, n63735, n63736, n63737, n63738, n63739, n63740,
n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748,
n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756,
n63757, n63758, n63759, n63760, n63761, n63762, n63763, n63764,
n63765, n63766, n63767, n63768, n63769, n63770, n63771, n63772,
n63773, n63774, n63775, n63776, n63777, n63778, n63779, n63780,
n63781, n63782, n63783, n63784, n63785, n63786, n63787, n63788,
n63789, n63790, n63791, n63792, n63793, n63794, n63795, n63796,
n63797, n63798, n63799, n63800, n63801, n63802, n63803, n63804,
n63805, n63806, n63807, n63808, n63809, n63810, n63811, n63812,
n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820,
n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828,
n63829, n63830, n63831, n63832, n63833, n63834, n63835, n63836,
n63837, n63838, n63839, n63840, n63841, n63842, n63843, n63844,
n63845, n63846, n63847, n63848, n63849, n63850, n63851, n63852,
n63853, n63854, n63855, n63856, n63857, n63858, n63859, n63860,
n63861, n63862, n63863, n63864, n63865, n63866, n63867, n63868,
n63869, n63870, n63871, n63872, n63873, n63874, n63875, n63876,
n63877, n63878, n63879, n63880, n63881, n63882, n63883, n63884,
n63885, n63886, n63887, n63888, n63889, n63890, n63891, n63892,
n63893, n63894, n63895, n63896, n63897, n63898, n63899, n63900,
n63901, n63902, n63903, n63904, n63905, n63906, n63907, n63908,
n63909, n63910, n63911, n63912, n63913, n63914, n63915, n63916,
n63917, n63918, n63919, n63920, n63921, n63922, n63923, n63924,
n63925, n63926, n63927, n63928, n63929, n63930, n63931, n63932,
n63933, n63934, n63935, n63936, n63937, n63938, n63939, n63940,
n63941, n63942, n63943, n63944, n63945, n63946, n63947, n63948,
n63949, n63950, n63951, n63952, n63953, n63954, n63955, n63956,
n63957, n63958, n63959, n63960, n63961, n63962, n63963, n63964,
n63965, n63966, n63967, n63968, n63969, n63970, n63971, n63972,
n63975, n63976, n63977, n63978, n63979, n63980, n63981, n63982,
n63983, n63984, n63985, n63986, n63987, n63988, n63989, n63990,
n63991, n63992, n63993, n63994, n63995, n63996, n63997, n63998,
n63999, n64000, n64001, n64002, n64003, n64004, n64005, n64006,
n64007, n64008, n64009, n64010, n64011, n64012, n64013, n64014,
n64015, n64016, n64017, n64018, n64019, n64020, n64021, n64022,
n64023, n64024, n64025, n64026, n64027, n64028, n64029, n64030,
n64031, n64032, n64033, n64034, n64035, n64036, n64037, n64038,
n64039, n64040, n64041, n64042, n64043, n64044, n64045, n64046,
n64047, n64048, n64049, n64050, n64051, n64052, n64053, n64054,
n64055, n64056, n64057, n64058, n64059, n64060, n64061, n64062,
n64063, n64064, n64065, n64066, n64067, n64068, n64069, n64070,
n64071, n64072, n64073, n64074, n64075, n64076, n64077, n64078,
n64079, n64080, n64081, n64082, n64083, n64084, n64085, n64086,
n64087, n64088, n64089, n64090, n64091, n64092, n64093, n64094,
n64095, n64096, n64097, n64098, n64099, n64100, n64101, n64102,
n64103, n64104, n64105, n64106, n64107, n64108, n64109, n64110,
n64111, n64112, n64113, n64114, n64115, n64116, n64117, n64118,
n64119, n64120, n64121, n64122, n64123, n64124, n64125, n64127,
n64128, n64129, n64130, n64131, n64132, n64133, n64134, n64135,
n64136, n64137, n64138, n64139, n64140, n64141, n64142, n64143,
n64144, n64145, n64146, n64147, n64148, n64149, n64150, n64151,
n64152, n64153, n64154, n64155, n64156, n64157, n64158, n64159,
n64160, n64161, n64162, n64163, n64164, n64165, n64166, n64167,
n64168, n64169, n64170, n64171, n64172, n64173, n64174, n64175,
n64176, n64177, n64178, n64179, n64180, n64181, n64182, n64183,
n64184, n64185, n64186, n64187, n64188, n64189, n64190, n64191,
n64192, n64193, n64194, n64195, n64196, n64197, n64198, n64199,
n64200, n64201, n64202, n64203, n64204, n64205, n64206, n64208,
n64209, n64210, n64211, n64212, n64213, n64214, n64215, n64216,
n64217, n64218, n64219, n64220, n64221, n64222, n64223, n64224,
n64225, n64226, n64227, n64228, n64229, n64230, n64231, n64232,
n64233, n64234, n64235, n64236, n64237, n64238, n64239, n64240,
n64241, n64242, n64243, n64244, n64245, n64246, n64247, n64248,
n64249, n64250, n64251, n64252, n64253, n64254, n64255, n64256,
n64257, n64258, n64259, n64260, n64261, n64262, n64263, n64264,
n64265, n64266, n64267, n64268, n64269, n64270, n64271, n64272,
n64273, n64274, n64275, n64276, n64277, n64278, n64279, n64280,
n64281, n64282, n64283, n64284, n64285, n64286, n64287, n64288,
n64289, n64290, n64291, n64292, n64293, n64294, n64295, n64296,
n64297, n64298, n64299, n64300, n64301, n64302, n64303, n64304,
n64305, n64306, n64307, n64308, n64309, n64310, n64311, n64312,
n64313, n64314, n64315, n64316, n64317, n64318, n64319, n64320,
n64321, n64322, n64323, n64324, n64325, n64326, n64327, n64328,
n64329, n64330, n64331, n64332, n64333, n64334, n64335, n64336,
n64337, n64338, n64339, n64340, n64341, n64342, n64343, n64344,
n64345, n64346, n64347, n64348, n64349, n64350, n64351, n64352,
n64353, n64354, n64355, n64356, n64357, n64358, n64359, n64360,
n64361, n64362, n64363, n64364, n64365, n64366, n64367, n64368,
n64369, n64370, n64371, n64372, n64373, n64374, n64375, n64376,
n64377, n64378, n64379, n64380, n64381, n64382, n64383, n64384,
n64385, n64386, n64387, n64388, n64389, n64390, n64391, n64392,
n64393, n64394, n64395, n64396, n64397, n64398, n64399, n64400,
n64401, n64402, n64403, n64404, n64405, n64406, n64407, n64408,
n64409, n64410, n64411, n64412, n64413, n64414, n64415, n64416,
n64417, n64418, n64419, n64420, n64421, n64422, n64423, n64424,
n64425, n64426, n64427, n64428, n64429, n64430, n64431, n64432,
n64433, n64434, n64435, n64436, n64437, n64438, n64439, n64440,
n64441, n64442, n64443, n64444, n64445, n64446, n64447, n64448,
n64449, n64450, n64451, n64452, n64453, n64454, n64455, n64456,
n64457, n64458, n64459, n64460, n64461, n64462, n64463, n64464,
n64465, n64466, n64467, n64468, n64469, n64470, n64471, n64472,
n64473, n64474, n64475, n64476, n64477, n64478, n64479, n64480,
n64481, n64482, n64483, n64484, n64485, n64486, n64487, n64488,
n64489, n64490, n64491, n64492, n64493, n64494, n64495, n64496,
n64497, n64498, n64499, n64500, n64501, n64502, n64503, n64504,
n64505, n64506, n64507, n64508, n64509, n64510, n64511, n64512,
n64513, n64514, n64515, n64516, n64517, n64518, n64519, n64520,
n64521, n64522, n64523, n64524, n64525, n64526, n64527, n64528,
n64529, n64530, n64531, n64532, n64533, n64534, n64535, n64536,
n64537, n64538, n64539, n64540, n64541, n64542, n64543, n64544,
n64545, n64546, n64547, n64548, n64549, n64550, n64551, n64552,
n64553, n64554, n64555, n64556, n64557, n64558, n64559, n64560,
n64561, n64562, n64563, n64564, n64565, n64566, n64567, n64568,
n64569, n64570, n64571, n64572, n64573, n64574, n64575, n64576,
n64577, n64578, n64579, n64580, n64581, n64582, n64583, n64585,
n64586, n64587, n64588, n64589, n64590, n64591, n64592, n64593,
n64594, n64595, n64596, n64597, n64598, n64599, n64600, n64601,
n64602, n64603, n64604, n64605, n64606, n64607, n64608, n64609,
n64610, n64611, n64612, n64613, n64614, n64615, n64616, n64619,
n64620, n64623, n64624, n64625, n64626, n64629, n64630, n64631,
n64632, n64633, n64634, n64635, n64636, n64637, n64638, n64639,
n64640, n64641, n64642, n64643, n64644, n64645, n64646, n64647,
n64648, n64649, n64650, n64651, n64652, n64653, n64654, n64655,
n64656, n64657, n64658, n64659, n64660, n64661, n64662, n64663,
n64664, n64665, n64666, n64667, n64668, n64669, n64670, n64671,
n64672, n64673, n64674, n64675, n64676, n64677, n64678, n64679,
n64680, n64681, n64682, n64683, n64684, n64685, n64686, n64687,
n64690, n64691, n64693, n64694, n64695, n64696, n64697, n64698,
n64699, n64700, n64701, n64702, n64703, n64704, n64705, n64706,
n64707, n64708, n64709, n64710, n64711, n64712, n64713, n64714,
n64715, n64716, n64717, n64718, n64719, n64720, n64721, n64722,
n64723, n64724, n64725, n64726, n64727, n64728, n64729, n64730,
n64731, n64732, n64733, n64734, n64735, n64736, n64737, n64738,
n64739, n64740, n64741, n64742, n64743, n64744, n64745, n64746,
n64747, n64748, n64749, n64750, n64751, n64752, n64753, n64754,
n64755, n64756, n64757, n64758, n64759, n64760, n64761, n64762,
n64763, n64764, n64765, n64766, n64767, n64768, n64769, n64770,
n64771, n64772, n64773, n64774, n64775, n64776, n64777, n64778,
n64779, n64780, n64781, n64782, n64783, n64784, n64785, n64786,
n64787, n64788, n64789, n64790, n64791, n64792, n64793, n64794,
n64795, n64796, n64797, n64798, n64799, n64800, n64801, n64802,
n64803, n64804, n64805, n64806, n64807, n64808, n64809, n64810,
n64811, n64812, n64813, n64814, n64815, n64816, n64817, n64818,
n64819, n64820, n64821, n64822, n64823, n64824, n64825, n64826,
n64827, n64828, n64829, n64830, n64831, n64832, n64833, n64834,
n64835, n64836, n64837, n64838, n64839, n64840, n64841, n64842,
n64843, n64844, n64845, n64846, n64847, n64848, n64849, n64850,
n64851, n64852, n64853, n64854, n64855, n64856, n64857, n64858,
n64859, n64860, n64861, n64862, n64863, n64864, n64865, n64866,
n64867, n64868, n64869, n64870, n64871, n64872, n64873, n64874,
n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882,
n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890,
n64891, n64892, n64893, n64894, n64895, n64896, n64897, n64898,
n64899, n64900, n64901, n64902, n64903, n64904, n64905, n64906,
n64907, n64908, n64909, n64910, n64911, n64912, n64913, n64914,
n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922,
n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930,
n64931, n64932, n64933, n64934, n64935, n64936, n64937, n64938,
n64939, n64940, n64941, n64942, n64943, n64944, n64945, n64946,
n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954,
n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962,
n64963, n64964, n64965, n64966, n64967, n64968, n64969, n64970,
n64971, n64972, n64973, n64974, n64975, n64976, n64977, n64978,
n64979, n64980, n64981, n64982, n64983, n64984, n64985, n64986,
n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994,
n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002,
n65003, n65004, n65005, n65006, n65007, n65008, n65009, n65010,
n65011, n65012, n65013, n65014, n65015, n65016, n65017, n65018,
n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026,
n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034,
n65035, n65036, n65037, n65038, n65039, n65040, n65041, n65042,
n65043, n65044, n65045, n65046, n65047, n65048, n65049, n65050,
n65051, n65052, n65053, n65054, n65055, n65056, n65057, n65058,
n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066,
n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074,
n65075, n65076, n65077, n65078, n65079, n65080, n65081, n65082,
n65083, n65084, n65085, n65086, n65087, n65088, n65089, n65090,
n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098,
n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106,
n65107, n65108, n65109, n65110, n65111, n65112, n65113, n65114,
n65115, n65116, n65117, n65118, n65119, n65120, n65121, n65122,
n65123, n65124, n65125, n65126, n65127, n65128, n65129, n65130,
n65131, n65132, n65133, n65134, n65135, n65136, n65137, n65138,
n65139, n65140, n65141, n65142, n65143, n65144, n65145, n65146,
n65147, n65148, n65149, n65150, n65151, n65152, n65153, n65154,
n65155, n65156, n65157, n65158, n65159, n65160, n65161, n65162,
n65163, n65164, n65165, n65166, n65167, n65168, n65169, n65170,
n65171, n65172, n65173, n65174, n65175, n65176, n65177, n65178,
n65179, n65180, n65181, n65182, n65183, n65184, n65185, n65186,
n65187, n65188, n65189, n65190, n65191, n65192, n65193, n65194,
n65195, n65196, n65197, n65198, n65199, n65200, n65201, n65202,
n65203, n65204, n65205, n65206, n65207, n65208, n65209, n65210,
n65211, n65212, n65213, n65214, n65215, n65216, n65217, n65218,
n65219, n65220, n65221, n65222, n65223, n65224, n65225, n65226,
n65227, n65228, n65229, n65230, n65231, n65232, n65233, n65234,
n65235, n65236, n65237, n65238, n65239, n65240, n65241, n65242,
n65243, n65244, n65245, n65246, n65247, n65248, n65249, n65250,
n65251, n65252, n65253, n65254, n65255, n65256, n65257, n65258,
n65259, n65260, n65261, n65262, n65263, n65264, n65265, n65266,
n65267, n65268, n65269, n65270, n65271, n65272, n65273, n65274,
n65275, n65276, n65277, n65278, n65279, n65280, n65281, n65282,
n65283, n65284, n65285, n65286, n65287, n65288, n65289, n65290,
n65291, n65292, n65293, n65294, n65295, n65296, n65297, n65298,
n65299, n65300, n65301, n65302, n65303, n65304, n65305, n65306,
n65307, n65308, n65309, n65310, n65311, n65312, n65313, n65314,
n65315, n65316, n65317, n65318, n65319, n65320, n65321, n65322,
n65323, n65324, n65325, n65326, n65327, n65328, n65329, n65330,
n65331, n65332, n65333, n65334, n65336, n65337, n65338, n65339,
n65340, n65341, n65342, n65343, n65344, n65345, n65346, n65347,
n65348, n65349, n65350, n65351, n65352, n65353, n65354, n65355,
n65356, n65357, n65358, n65359, n65360, n65361, n65362, n65363,
n65364, n65365, n65366, n65367, n65368, n65369, n65370, n65371,
n65372, n65373, n65374, n65375, n65376, n65377, n65378, n65379,
n65380, n65381, n65382, n65383, n65384, n65385, n65386, n65387,
n65388, n65389, n65390, n65391, n65392, n65393, n65394, n65395,
n65396, n65397, n65398, n65399, n65400, n65401, n65402, n65403,
n65404, n65405, n65406, n65407, n65408, n65409, n65410, n65411,
n65412, n65413, n65414, n65415, n65416, n65417, n65418, n65419,
n65420, n65421, n65422, n65423, n65424, n65425, n65426, n65427,
n65428, n65429, n65430, n65431, n65432, n65433, n65434, n65435,
n65436, n65437, n65438, n65439, n65440, n65441, n65442, n65443,
n65444, n65445, n65446, n65447, n65448, n65449, n65450, n65451,
n65452, n65453, n65454, n65455, n65456, n65457, n65458, n65459,
n65460, n65461, n65462, n65463, n65464, n65465, n65466, n65467,
n65468, n65469, n65470, n65471, n65472, n65473, n65474, n65475,
n65476, n65477, n65478, n65479, n65480, n65481, n65482, n65483,
n65484, n65485, n65486, n65487, n65488, n65489, n65490, n65491,
n65492, n65493, n65494, n65495, n65496, n65497, n65498, n65499,
n65500, n65501, n65502, n65503, n65504, n65505, n65506, n65507,
n65508, n65509, n65510, n65511, n65512, n65513, n65514, n65515,
n65516, n65517, n65518, n65519, n65520, n65521, n65522, n65523,
n65524, n65525, n65526, n65527, n65528, n65529, n65530, n65531,
n65532, n65533, n65534, n65535, n65536, n65537, n65538, n65539,
n65540, n65541, n65542, n65543, n65544, n65545, n65546, n65547,
n65548, n65549, n65550, n65551, n65552, n65553, n65554, n65555,
n65556, n65557, n65558, n65559, n65560, n65561, n65562, n65563,
n65564, n65565, n65566, n65567, n65568, n65569, n65570, n65571,
n65572, n65573, n65574, n65575, n65576, n65577, n65578, n65579,
n65580, n65581, n65582, n65583, n65584, n65585, n65586, n65587,
n65588, n65589, n65590, n65591, n65592, n65593, n65594, n65595,
n65596, n65597, n65598, n65599, n65600, n65601, n65602, n65603,
n65604, n65605, n65606, n65607, n65608, n65609, n65610, n65611,
n65612, n65613, n65614, n65615, n65616, n65617, n65618, n65619,
n65620, n65621, n65622, n65623, n65624, n65625, n65626, n65627,
n65628, n65629, n65630, n65631, n65632, n65633, n65634, n65635,
n65636, n65637, n65638, n65639, n65640, n65641, n65642, n65643,
n65644, n65645, n65646, n65647, n65648, n65649, n65650, n65651,
n65652, n65653, n65654, n65655, n65656, n65657, n65658, n65659,
n65660, n65661, n65662, n65663, n65664, n65665, n65666, n65667,
n65668, n65669, n65670, n65671, n65672, n65673, n65674, n65675,
n65676, n65677, n65678, n65679, n65680, n65681, n65682, n65683,
n65684, n65685, n65686, n65687, n65688, n65689, n65690, n65691,
n65692, n65693, n65694, n65695, n65696, n65697, n65698, n65699,
n65700, n65701, n65702, n65703, n65704, n65705, n65706, n65707,
n65708, n65709, n65710, n65711, n65712, n65713, n65714, n65715,
n65716, n65717, n65718, n65719, n65720, n65721, n65722, n65723,
n65724, n65725, n65726, n65727, n65728, n65729, n65730, n65731,
n65732, n65733, n65734, n65735, n65736, n65737, n65738, n65739,
n65740, n65741, n65742, n65743, n65744, n65745, n65746, n65747,
n65748, n65749, n65750, n65751, n65752, n65753, n65754, n65755,
n65756, n65757, n65758, n65759, n65760, n65761, n65762, n65763,
n65764, n65765, n65766, n65767, n65768, n65769, n65770, n65771,
n65772, n65773, n65774, n65775, n65776, n65777, n65778, n65779,
n65780, n65781, n65782, n65783, n65784, n65785, n65786, n65787,
n65788, n65789, n65790, n65791, n65792, n65793, n65794, n65795,
n65796, n65797, n65798, n65799, n65800, n65801, n65802, n65803,
n65804, n65805, n65806, n65807, n65808, n65809, n65810, n65811,
n65812, n65813, n65814, n65815, n65816, n65817, n65818, n65819,
n65820, n65821, n65822, n65823, n65824, n65825, n65826, n65827,
n65828, n65829, n65830, n65831, n65832, n65833, n65834, n65835,
n65836, n65837, n65838, n65839, n65840, n65841, n65842, n65843,
n65844, n65845, n65846, n65847, n65848, n65849, n65850, n65851,
n65852, n65853, n65854, n65855, n65856, n65857, n65858, n65859,
n65860, n65861, n65862, n65863, n65864, n65865, n65866, n65867,
n65868, n65869, n65870, n65871, n65872, n65873, n65874, n65875,
n65876, n65877, n65878, n65879, n65880, n65881, n65882, n65883,
n65884, n65885, n65886, n65887, n65888, n65889, n65890, n65891,
n65892, n65893, n65894, n65895, n65896, n65897, n65898, n65899,
n65900, n65901, n65902, n65903, n65904, n65905, n65906, n65907,
n65908, n65909, n65910, n65911, n65912, n65913, n65914, n65915,
n65916, n65917, n65918, n65919, n65920, n65921, n65922, n65923,
n65924, n65925, n65926, n65927, n65928, n65929, n65930, n65931,
n65932, n65933, n65934, n65935, n65936, n65937, n65938, n65939,
n65940, n65941, n65942, n65943, n65944, n65945, n65946, n65947,
n65948, n65949, n65950, n65951, n65952, n65953, n65954, n65955,
n65956, n65957, n65958, n65959, n65960, n65961, n65962, n65963,
n65964, n65965, n65966, n65967, n65968, n65969, n65970, n65971,
n65972, n65973, n65974, n65975, n65976, n65977, n65978, n65979,
n65980, n65981, n65982, n65983, n65984, n65985, n65986, n65987,
n65988, n65989, n65990, n65991, n65992, n65993, n65994, n65995,
n65996, n65997, n65998, n65999, n66000, n66001, n66002, n66003,
n66004, n66005, n66006, n66007, n66008, n66009, n66010, n66011,
n66012, n66013, n66014, n66015, n66016, n66017, n66018, n66019,
n66020, n66021, n66022, n66023, n66024, n66025, n66026, n66027,
n66028, n66029, n66030, n66031, n66032, n66033, n66034, n66035,
n66036, n66037, n66038, n66039, n66040, n66041, n66042, n66043,
n66044, n66045, n66046, n66047, n66048, n66049, n66050, n66051,
n66052, n66053, n66054, n66055, n66056, n66057, n66058, n66059,
n66060, n66061, n66062, n66063, n66064, n66065, n66066, n66067,
n66068, n66069, n66070, n66071, n66072, n66073, n66074, n66075,
n66076, n66077, n66078, n66079, n66080, n66081, n66082, n66083,
n66084, n66085, n66086, n66087, n66088, n66089, n66090, n66091,
n66092, n66093, n66094, n66095, n66096, n66097, n66098, n66099,
n66100, n66101, n66102, n66103, n66104, n66105, n66106, n66107,
n66108, n66109, n66110, n66111, n66112, n66113, n66114, n66115,
n66116, n66117, n66118, n66119, n66120, n66121, n66122, n66123,
n66124, n66125, n66126, n66127, n66128, n66129, n66130, n66131,
n66132, n66133, n66134, n66135, n66136, n66137, n66138, n66139,
n66140, n66141, n66142, n66143, n66144, n66145, n66146, n66147,
n66148, n66149, n66150, n66151, n66152, n66153, n66154, n66155,
n66156, n66157, n66158, n66159, n66160, n66161, n66162, n66163,
n66164, n66165, n66166, n66167, n66168, n66169, n66170, n66171,
n66172, n66173, n66174, n66175, n66176, n66177, n66178, n66179,
n66180, n66181, n66182, n66183, n66184, n66185, n66186, n66187,
n66188, n66189, n66190, n66191, n66192, n66193, n66194, n66195,
n66196, n66197, n66198, n66199, n66200, n66201, n66202, n66203,
n66204, n66205, n66206, n66207, n66208, n66209, n66210, n66211,
n66212, n66213, n66214, n66215, n66216, n66217, n66218, n66219,
n66220, n66221, n66222, n66223, n66224, n66225, n66226, n66227,
n66228, n66229, n66230, n66231, n66232, n66233, n66234, n66235,
n66236, n66237, n66238, n66239, n66240, n66241, n66242, n66243,
n66244, n66245, n66246, n66247, n66248, n66249, n66250, n66251,
n66252, n66253, n66254, n66255, n66256, n66257, n66258, n66259,
n66260, n66261, n66262, n66263, n66264, n66265, n66266, n66267,
n66268, n66269, n66270, n66271, n66272, n66273, n66274, n66275,
n66276, n66277, n66278, n66279, n66280, n66281, n66282, n66283,
n66284, n66285, n66286, n66287, n66288, n66290, n66291, n66292,
n66293, n66294, n66295, n66296, n66297, n66298, n66299, n66300,
n66301, n66302, n66303, n66304, n66305, n66306, n66307, n66308,
n66309, n66310, n66311, n66312, n66313, n66314, n66315, n66316,
n66317, n66318, n66319, n66320, n66321, n66322, n66323, n66324,
n66325, n66326, n66327, n66328, n66329, n66330, n66331, n66332,
n66333, n66334, n66335, n66336, n66337, n66338, n66339, n66340,
n66341, n66342, n66343, n66344, n66345, n66346, n66347, n66348,
n66349, n66350, n66351, n66352, n66353, n66354, n66355, n66356,
n66357, n66358, n66359, n66360, n66361, n66362, n66363, n66364,
n66365, n66366, n66367, n66368, n66369, n66370, n66371, n66372,
n66373, n66374, n66375, n66376, n66377, n66378, n66379, n66380,
n66381, n66382, n66383, n66384, n66385, n66386, n66387, n66388,
n66389, n66390, n66391, n66392, n66393, n66394, n66395, n66396,
n66397, n66398, n66399, n66400, n66401, n66402, n66403, n66404,
n66405, n66406, n66407, n66408, n66409, n66410, n66411, n66412,
n66413, n66414, n66415, n66416, n66417, n66418, n66419, n66420,
n66421, n66422, n66423, n66424, n66425, n66426, n66427, n66428,
n66429, n66430, n66431, n66432, n66433, n66434, n66435, n66436,
n66437, n66438, n66439, n66440, n66441, n66442, n66443, n66444,
n66445, n66446, n66447, n66448, n66449, n66450, n66451, n66452,
n66453, n66454, n66455, n66456, n66457, n66458, n66459, n66460,
n66461, n66462, n66463, n66464, n66465, n66466, n66467, n66468,
n66469, n66470, n66471, n66472, n66473, n66474, n66475, n66476,
n66477, n66478, n66479, n66480, n66481, n66482, n66483, n66484,
n66485, n66486, n66487, n66488, n66489, n66490, n66491, n66492,
n66493, n66494, n66495, n66496, n66497, n66498, n66499, n66500,
n66501, n66502, n66503, n66504, n66505, n66506, n66507, n66508,
n66509, n66510, n66511, n66512, n66513, n66514, n66515, n66516,
n66517, n66518, n66519, n66520, n66521, n66522, n66523, n66524,
n66525, n66526, n66527, n66528, n66529, n66530, n66531, n66532,
n66533, n66534, n66535, n66536, n66537, n66538, n66539, n66540,
n66541, n66542, n66543, n66544, n66545, n66546, n66547, n66548,
n66549, n66551, n66552, n66553, n66554, n66555, n66556, n66557,
n66558, n66559, n66560, n66561, n66562, n66563, n66564, n66565,
n66566, n66567, n66568, n66569, n66570, n66571, n66572, n66573,
n66574, n66575, n66576, n66577, n66578, n66579, n66580, n66581,
n66582, n66583, n66584, n66585, n66586, n66587, n66588, n66589,
n66590, n66591, n66592, n66593, n66594, n66595, n66596, n66597,
n66598, n66599, n66600, n66601, n66602, n66603, n66604, n66605,
n66606, n66607, n66608, n66609, n66610, n66611, n66612, n66613,
n66614, n66615, n66616, n66617, n66618, n66619, n66620, n66621,
n66622, n66623, n66624, n66625, n66626, n66627, n66628, n66629,
n66630, n66631, n66632, n66633, n66634, n66635, n66636, n66637,
n66638, n66639, n66640, n66641, n66642, n66643, n66644, n66645,
n66646, n66647, n66648, n66649, n66650, n66651, n66652, n66653,
n66654, n66655, n66656, n66657, n66658, n66659, n66660, n66661,
n66662, n66663, n66664, n66665, n66666, n66667, n66668, n66669,
n66670, n66671, n66672, n66673, n66674, n66675, n66676, n66677,
n66678, n66679, n66680, n66681, n66682, n66683, n66684, n66685,
n66686, n66687, n66688, n66689, n66690, n66691, n66692, n66693,
n66694, n66695, n66696, n66697, n66698, n66699, n66700, n66701,
n66702, n66703, n66704, n66705, n66706, n66707, n66708, n66710,
n66711, n66712, n66713, n66714, n66715, n66716, n66717, n66718,
n66719, n66720, n66721, n66722, n66723, n66724, n66725, n66726,
n66727, n66728, n66729, n66730, n66731, n66732, n66733, n66734,
n66735, n66736, n66737, n66738, n66739, n66740, n66741, n66742,
n66743, n66744, n66745, n66746, n66747, n66748, n66749, n66750,
n66751, n66752, n66753, n66754, n66755, n66756, n66757, n66758,
n66759, n66760, n66761, n66762, n66763, n66764, n66765, n66766,
n66767, n66768, n66769, n66770, n66771, n66772, n66773, n66774,
n66775, n66776, n66777, n66778, n66779, n66780, n66781, n66782,
n66783, n66784, n66785, n66786, n66787, n66788, n66789, n66790,
n66791, n66792, n66793, n66794, n66795, n66796, n66797, n66798,
n66799, n66800, n66801, n66802, n66803, n66804, n66805, n66806,
n66807, n66808, n66809, n66810, n66811, n66812, n66813, n66814,
n66815, n66816, n66818, n66819, n66820, n66821, n66822, n66823,
n66824, n66825, n66826, n66827, n66828, n66829, n66830, n66831,
n66832, n66833, n66834, n66835, n66836, n66837, n66838, n66839,
n66840, n66841, n66842, n66843, n66844, n66845, n66846, n66847,
n66848, n66849, n66850, n66851, n66852, n66853, n66854, n66855,
n66856, n66857, n66858, n66859, n66860, n66861, n66862, n66863,
n66864, n66865, n66866, n66867, n66868, n66869, n66870, n66871,
n66872, n66873, n66874, n66875, n66876, n66877, n66878, n66879,
n66880, n66881, n66882, n66883, n66884, n66885, n66886, n66887,
n66888, n66889, n66890, n66891, n66892, n66894, n66895, n66896,
n66897, n66898, n66899, n66900, n66901, n66902, n66903, n66904,
n66905, n66906, n66907, n66908, n66909, n66910, n66911, n66912,
n66913, n66914, n66915, n66916, n66917, n66918, n66919, n66920,
n66921, n66922, n66923, n66924, n66925, n66926, n66927, n66928,
n66929, n66930, n66931, n66932, n66933, n66934, n66935, n66936,
n66937, n66938, n66939, n66940, n66941, n66942, n66943, n66944,
n66945, n66946, n66947, n66948, n66949, n66950, n66951, n66952,
n66953, n66954, n66955, n66956, n66957, n66959, n66960, n66961,
n66962, n66963, n66964, n66965, n66966, n66967, n66968, n66969,
n66970, n66971, n66972, n66973, n66974, n66975, n66976, n66977,
n66978, n66979, n66980, n66981, n66982, n66983, n66984, n66985,
n66986, n66987, n66988, n66989, n66990, n66991, n66992, n66993,
n66994, n66995, n66996, n66997, n66998, n66999, n67000, n67001,
n67002, n67003, n67004, n67005, n67006, n67007, n67008, n67009,
n67010, n67011, n67012, n67013, n67014, n67015, n67016, n67017,
n67018, n67019, n67020, n67021, n67022, n67023, n67024, n67025,
n67026, n67027, n67028, n67029, n67030, n67031, n67032, n67033,
n67034, n67035, n67036, n67037, n67038, n67039, n67040, n67041,
n67042, n67043, n67044, n67045, n67046, n67047, n67048, n67049,
n67050, n67051, n67052, n67053, n67054, n67055, n67056, n67057,
n67058, n67059, n67060, n67061, n67062, n67063, n67064, n67065,
n67066, n67067, n67068, n67069, n67070, n67071, n67072, n67073,
n67074, n67075, n67076, n67077, n67078, n67079, n67080, n67081,
n67082, n67083, n67084, n67085, n67086, n67087, n67088, n67089,
n67090, n67091, n67092, n67093, n67094, n67095, n67096, n67097,
n67098, n67099, n67100, n67101, n67102, n67103, n67104, n67105,
n67106, n67107, n67108, n67109, n67110, n67111, n67112, n67113,
n67114, n67115, n67116, n67117, n67118, n67119, n67120, n67121,
n67122, n67123, n67124, n67125, n67126, n67127, n67128, n67129,
n67130, n67131, n67132, n67133, n67134, n67135, n67136, n67137,
n67138, n67139, n67140, n67141, n67142, n67143, n67144, n67145,
n67146, n67147, n67148, n67149, n67150, n67151, n67152, n67153,
n67154, n67155, n67156, n67157, n67158, n67159, n67160, n67161,
n67162, n67163, n67164, n67165, n67166, n67167, n67168, n67169,
n67170, n67171, n67172, n67173, n67174, n67175, n67176, n67177,
n67178, n67179, n67180, n67181, n67182, n67183, n67184, n67185,
n67186, n67187, n67188, n67189, n67190, n67191, n67192, n67193,
n67194, n67195, n67196, n67197, n67198, n67199, n67200, n67201,
n67202, n67203, n67204, n67205, n67206, n67207, n67208, n67209,
n67210, n67211, n67212, n67213, n67214, n67215, n67216, n67217,
n67218, n67219, n67220, n67221, n67222, n67223, n67224, n67225,
n67226, n67227, n67228, n67229, n67230, n67231, n67232, n67233,
n67234, n67235, n67236, n67237, n67238, n67239, n67240, n67241,
n67242, n67243, n67244, n67245, n67246, n67247, n67248, n67249,
n67250, n67251, n67252, n67253, n67254, n67255, n67256, n67257,
n67258, n67259, n67260, n67261, n67262, n67263, n67264, n67265,
n67266, n67267, n67268, n67269, n67270, n67271, n67272, n67273,
n67274, n67275, n67276, n67277, n67278, n67279, n67280, n67281,
n67282, n67283, n67284, n67285, n67286, n67287, n67288, n67289,
n67290, n67291, n67292, n67293, n67294, n67295, n67296, n67297,
n67298, n67299, n67300, n67301, n67302, n67303, n67304, n67305,
n67306, n67307, n67308, n67309, n67310, n67311, n67312, n67313,
n67314, n67315, n67316, n67317, n67318, n67319, n67320, n67321,
n67322, n67323, n67324, n67325, n67326, n67327, n67328, n67329,
n67330, n67331, n67332, n67333, n67334, n67335, n67336, n67337,
n67338, n67339, n67340, n67341, n67342, n67343, n67344, n67345,
n67346, n67347, n67348, n67349, n67350, n67351, n67352, n67353,
n67354, n67355, n67356, n67357, n67358, n67359, n67360, n67361,
n67362, n67363, n67364, n67365, n67366, n67367, n67368, n67369,
n67370, n67371, n67372, n67373, n67374, n67375, n67376, n67377,
n67378, n67379, n67380, n67381, n67382, n67383, n67384, n67385,
n67386, n67387, n67388, n67389, n67390, n67391, n67392, n67393,
n67394, n67395, n67396, n67397, n67398, n67399, n67400, n67401,
n67402, n67403, n67404, n67405, n67406, n67407, n67408, n67409,
n67410, n67411, n67412, n67413, n67414, n67415, n67416, n67417,
n67418, n67419, n67420, n67423, n67424, n67425, n67426, n67427,
n67428, n67429, n67430, n67431, n67432, n67433, n67434, n67435,
n67436, n67437, n67438, n67439, n67440, n67441, n67442, n67443,
n67444, n67445, n67446, n67447, n67448, n67449, n67450, n67451,
n67452, n67453, n67454, n67455, n67456, n67457, n67458, n67459,
n67460, n67461, n67462, n67463, n67464, n67465, n67466, n67467,
n67468, n67469, n67470, n67471, n67472, n67473, n67474, n67475,
n67476, n67477, n67478, n67479, n67480, n67481, n67482, n67483,
n67484, n67485, n67486, n67487, n67488, n67489, n67490, n67491,
n67492, n67493, n67494, n67495, n67496, n67497, n67498, n67499,
n67500, n67501, n67502, n67503, n67504, n67505, n67506, n67507,
n67508, n67509, n67510, n67511, n67512, n67513, n67514, n67515,
n67516, n67517, n67518, n67519, n67520, n67521, n67522, n67523,
n67524, n67525, n67526, n67527, n67528, n67529, n67530, n67531,
n67532, n67533, n67534, n67535, n67536, n67537, n67538, n67539,
n67540, n67541, n67542, n67543, n67544, n67545, n67546, n67547,
n67548, n67549, n67550, n67551, n67552, n67553, n67554, n67555,
n67556, n67557, n67558, n67559, n67560, n67561, n67562, n67563,
n67564, n67565, n67566, n67567, n67568, n67569, n67570, n67571,
n67572, n67573, n67574, n67575, n67576, n67577, n67578, n67579,
n67580, n67581, n67582, n67583, n67584, n67585, n67586, n67587,
n67588, n67589, n67590, n67591, n67592, n67593, n67594, n67595,
n67596, n67597, n67598, n67599, n67600, n67601, n67602, n67603,
n67604, n67605, n67606, n67607, n67608, n67609, n67610, n67611,
n67612, n67613, n67614, n67615, n67616, n67617, n67618, n67619,
n67620, n67621, n67622, n67623, n67624, n67625, n67626, n67627,
n67628, n67629, n67630, n67631, n67632, n67633, n67634, n67635,
n67636, n67637, n67638, n67639, n67640, n67641, n67642, n67643,
n67644, n67645, n67646, n67647, n67648, n67649, n67650, n67651,
n67652, n67653, n67654, n67655, n67656, n67657, n67658, n67659,
n67660, n67661, n67662, n67663, n67664, n67665, n67666, n67667,
n67668, n67669, n67670, n67671, n67672, n67673, n67674, n67675,
n67676, n67677, n67678, n67679, n67680, n67681, n67682, n67683,
n67684, n67685, n67686, n67687, n67688, n67689, n67690, n67691,
n67692, n67693, n67694, n67695, n67696, n67697, n67698, n67699,
n67700, n67701, n67702, n67703, n67704, n67705, n67706, n67707,
n67708, n67709, n67710, n67711, n67712, n67713, n67714, n67715,
n67716, n67717, n67718, n67719, n67720, n67721, n67722, n67723,
n67724, n67725, n67726, n67727, n67728, n67729, n67730, n67731,
n67732, n67733, n67734, n67735, n67736, n67737, n67738, n67739,
n67740, n67741, n67742, n67743, n67744, n67745, n67746, n67747,
n67748, n67749, n67750, n67751, n67752, n67753, n67754, n67755,
n67756, n67757, n67758, n67759, n67760, n67761, n67762, n67763,
n67764, n67765, n67766, n67767, n67768, n67769, n67770, n67771,
n67772, n67773, n67774, n67775, n67776, n67777, n67778, n67779,
n67780, n67781, n67782, n67783, n67784, n67785, n67786, n67787,
n67788, n67789, n67790, n67791, n67792, n67793, n67794, n67795,
n67796, n67797, n67798, n67799, n67800, n67801, n67802, n67803,
n67804, n67805, n67806, n67807, n67808, n67809, n67810, n67811,
n67812, n67813, n67814, n67815, n67816, n67817, n67818, n67819,
n67820, n67821, n67822, n67823, n67824, n67825, n67826, n67827,
n67828, n67829, n67830, n67831, n67832, n67833, n67834, n67835,
n67836, n67837, n67838, n67839, n67840, n67841, n67842, n67843,
n67844, n67845, n67846, n67847, n67848, n67849, n67850, n67851,
n67852, n67853, n67854, n67855, n67856, n67857, n67858, n67859,
n67860, n67861, n67862, n67863, n67864, n67865, n67866, n67867,
n67868, n67869, n67870, n67871, n67872, n67873, n67874, n67875,
n67876, n67877, n67878, n67879, n67880, n67881, n67882, n67883,
n67884, n67885, n67886, n67887, n67888, n67889, n67890, n67891,
n67892, n67893, n67894, n67895, n67896, n67897, n67898, n67899,
n67900, n67901, n67902, n67903, n67904, n67905, n67906, n67907,
n67908, n67909, n67910, n67911, n67912, n67913, n67914, n67915,
n67916, n67917, n67918, n67919, n67920, n67921, n67922, n67923,
n67924, n67925, n67926, n67927, n67928, n67929, n67930, n67931,
n67932, n67933, n67934, n67935, n67936, n67937, n67938, n67939,
n67940, n67941, n67942, n67943, n67944, n67945, n67946, n67947,
n67948, n67949, n67950, n67951, n67952, n67953, n67954, n67955,
n67956, n67957, n67958, n67959, n67960, n67961, n67962, n67963,
n67964, n67965, n67966, n67967, n67968, n67969, n67970, n67971,
n67972, n67973, n67974, n67975, n67976, n67977, n67978, n67979,
n67980, n67981, n67982, n67983, n67984, n67985, n67986, n67987,
n67988, n67989, n67990, n67991, n67992, n67993, n67994, n67995,
n67996, n67997, n67998, n67999, n68000, n68001, n68002, n68003,
n68004, n68005, n68006, n68007, n68008, n68009, n68011, n68012,
n68013, n68014, n68015, n68016, n68017, n68018, n68019, n68020,
n68021, n68022, n68023, n68024, n68025, n68026, n68027, n68028,
n68029, n68030, n68031, n68032, n68033, n68034, n68035, n68036,
n68037, n68038, n68039, n68040, n68041, n68042, n68043, n68044,
n68045, n68046, n68047, n68048, n68051, n68052, n68053, n68054,
n68055, n68056, n68057, n68058, n68059, n68060, n68061, n68062,
n68063, n68064, n68065, n68066, n68067, n68068, n68069, n68070,
n68071, n68072, n68073, n68074, n68075, n68076, n68077, n68078,
n68079, n68080, n68081, n68082, n68083, n68084, n68085, n68086,
n68087, n68088, n68090, n68091, n68092, n68093, n68094, n68095,
n68096, n68097, n68098, n68099, n68100, n68101, n68102, n68103,
n68104, n68105, n68106, n68107, n68108, n68109, n68110, n68111,
n68112, n68113, n68114, n68115, n68116, n68117, n68118, n68119,
n68120, n68121, n68122, n68123, n68124, n68125, n68126, n68127,
n68128, n68129, n68130, n68131, n68132, n68133, n68134, n68135,
n68136, n68137, n68138, n68139, n68140, n68141, n68142, n68143,
n68144, n68145, n68146, n68147, n68148, n68149, n68150, n68151,
n68152, n68153, n68154, n68155, n68156, n68157, n68158, n68159,
n68160, n68161, n68162, n68163, n68164, n68165, n68166, n68167,
n68168, n68169, n68170, n68171, n68172, n68173, n68174, n68175,
n68176, n68177, n68178, n68179, n68180, n68181, n68182, n68183,
n68184, n68185, n68186, n68187, n68188, n68189, n68190, n68191,
n68192, n68193, n68194, n68195, n68196, n68197, n68198, n68199,
n68200, n68201, n68202, n68203, n68204, n68205, n68206, n68207,
n68208, n68209, n68210, n68211, n68212, n68213, n68214, n68215,
n68216, n68217, n68218, n68219, n68220, n68221, n68222, n68223,
n68224, n68225, n68226, n68227, n68228, n68229, n68230, n68231,
n68232, n68233, n68234, n68235, n68236, n68237, n68238, n68240,
n68241, n68242, n68243, n68244, n68245, n68246, n68247, n68248,
n68249, n68250, n68251, n68252, n68253, n68254, n68255, n68256,
n68257, n68258, n68259, n68260, n68261, n68262, n68263, n68264,
n68265, n68266, n68267, n68268, n68269, n68270, n68271, n68272,
n68273, n68274, n68275, n68276, n68277, n68278, n68279, n68280,
n68281, n68282, n68283, n68284, n68285, n68286, n68287, n68288,
n68289, n68290, n68291, n68292, n68293, n68294, n68295, n68296,
n68297, n68298, n68299, n68300, n68301, n68302, n68303, n68304,
n68305, n68306, n68307, n68308, n68309, n68310, n68311, n68312,
n68313, n68314, n68315, n68316, n68317, n68318, n68319, n68320,
n68321, n68322, n68323, n68324, n68325, n68326, n68327, n68328,
n68329, n68330, n68331, n68332, n68333, n68334, n68335, n68336,
n68338, n68339, n68340, n68341, n68342, n68343, n68344, n68345,
n68346, n68347, n68348, n68349, n68350, n68351, n68352, n68353,
n68354, n68355, n68356, n68357, n68358, n68359, n68360, n68361,
n68362, n68363, n68364, n68365, n68366, n68367, n68368, n68369,
n68370, n68371, n68372, n68373, n68374, n68375, n68376, n68377,
n68378, n68379, n68380, n68381, n68382, n68383, n68384, n68385,
n68386, n68387, n68388, n68389, n68390, n68391, n68392, n68393,
n68394, n68395, n68396, n68397, n68398, n68399, n68400, n68401,
n68402, n68403, n68404, n68405, n68406, n68407, n68408, n68409,
n68410, n68411, n68412, n68413, n68414, n68415, n68416, n68417,
n68418, n68419, n68420, n68421, n68422, n68423, n68424, n68425,
n68426, n68427, n68428, n68429, n68430, n68431, n68432, n68433,
n68434, n68435, n68436, n68437, n68438, n68439, n68440, n68441,
n68442, n68443, n68444, n68445, n68446, n68447, n68448, n68449,
n68450, n68451, n68452, n68453, n68454, n68455, n68456, n68457,
n68458, n68459, n68460, n68461, n68462, n68463, n68464, n68465,
n68466, n68467, n68468, n68469, n68470, n68471, n68472, n68473,
n68474, n68475, n68476, n68477, n68478, n68479, n68480, n68481,
n68482, n68483, n68484, n68485, n68486, n68487, n68488, n68489,
n68490, n68491, n68492, n68493, n68494, n68495, n68496, n68497,
n68498, n68499, n68500, n68501, n68502, n68503, n68504, n68505,
n68506, n68507, n68508, n68509, n68510, n68511, n68512, n68513,
n68514, n68515, n68516, n68517, n68518, n68519, n68520, n68521,
n68522, n68523, n68524, n68525, n68526, n68527, n68528, n68529,
n68530, n68531, n68532, n68533, n68534, n68535, n68536, n68537,
n68538, n68539, n68540, n68541, n68542, n68543, n68544, n68545,
n68546, n68547, n68548, n68549, n68550, n68551, n68552, n68553,
n68554, n68555, n68556, n68557, n68558, n68559, n68560, n68561,
n68562, n68563, n68564, n68565, n68566, n68567, n68568, n68569,
n68570, n68571, n68572, n68573, n68574, n68575, n68576, n68577,
n68578, n68579, n68580, n68581, n68582, n68583, n68584, n68585,
n68586, n68587, n68588, n68589, n68590, n68591, n68592, n68593,
n68594, n68595, n68596, n68597, n68598, n68599, n68600, n68601,
n68602, n68603, n68604, n68605, n68606, n68607, n68608, n68609,
n68610, n68611, n68612, n68613, n68614, n68615, n68616, n68617,
n68618, n68619, n68620, n68621, n68622, n68623, n68624, n68625,
n68626, n68627, n68628, n68629, n68630, n68631, n68632, n68633,
n68634, n68635, n68636, n68637, n68638, n68639, n68640, n68641,
n68642, n68643, n68644, n68645, n68646, n68647, n68648, n68649,
n68650, n68651, n68652, n68653, n68654, n68655, n68656, n68657,
n68658, n68659, n68660, n68661, n68662, n68663, n68664, n68665,
n68666, n68667, n68668, n68669, n68670, n68671, n68672, n68673,
n68674, n68675, n68676, n68677, n68678, n68679, n68680, n68681,
n68682, n68683, n68684, n68685, n68686, n68687, n68688, n68689,
n68690, n68691, n68692, n68693, n68694, n68695, n68696, n68697,
n68698, n68699, n68700, n68701, n68702, n68703, n68704, n68705,
n68708, n68709, n68710, n68711, n68712, n68713, n68714, n68715,
n68716, n68717, n68718, n68719, n68720, n68721, n68722, n68723,
n68724, n68725, n68726, n68727, n68728, n68729, n68730, n68731,
n68732, n68733, n68734, n68735, n68736, n68737, n68738, n68739,
n68740, n68741, n68742, n68743, n68744, n68745, n68746, n68747,
n68748, n68749, n68750, n68751, n68752, n68753, n68754, n68755,
n68756, n68757, n68758, n68759, n68760, n68761, n68762, n68763,
n68764, n68765, n68766, n68767, n68768, n68769, n68770, n68771,
n68772, n68773, n68774, n68775, n68776, n68777, n68778, n68779,
n68780, n68781, n68782, n68783, n68784, n68785, n68786, n68787,
n68788, n68789, n68790, n68791, n68792, n68793, n68794, n68795,
n68796, n68797, n68798, n68799, n68800, n68801, n68802, n68803,
n68804, n68805, n68806, n68807, n68808, n68809, n68810, n68811,
n68812, n68813, n68814, n68815, n68816, n68817, n68818, n68819,
n68820, n68821, n68822, n68823, n68824, n68825, n68826, n68827,
n68828, n68829, n68830, n68831, n68832, n68833, n68834, n68835,
n68836, n68837, n68838, n68839, n68840, n68841, n68842, n68843,
n68844, n68845, n68846, n68847, n68848, n68849, n68850, n68851,
n68852, n68853, n68854, n68855, n68856, n68857, n68858, n68859,
n68860, n68861, n68862, n68863, n68864, n68865, n68866, n68867,
n68868, n68869, n68870, n68871, n68872, n68873, n68874, n68875,
n68876, n68877, n68878, n68879, n68880, n68881, n68882, n68883,
n68884, n68885, n68886, n68887, n68888, n68889, n68890, n68891,
n68892, n68893, n68894, n68895, n68896, n68897, n68898, n68899,
n68900, n68901, n68902, n68903, n68904, n68905, n68906, n68907,
n68908, n68909, n68910, n68911, n68912, n68913, n68914, n68915,
n68916, n68917, n68918, n68919, n68920, n68921, n68922, n68923,
n68924, n68925, n68926, n68927, n68928, n68929, n68930, n68931,
n68932, n68933, n68934, n68935, n68936, n68937, n68938, n68939,
n68940, n68941, n68942, n68943, n68944, n68945, n68946, n68947,
n68948, n68949, n68950, n68951, n68952, n68953, n68954, n68955,
n68956, n68957, n68958, n68959, n68960, n68961, n68962, n68963,
n68964, n68965, n68966, n68967, n68968, n68969, n68970, n68971,
n68972, n68973, n68974, n68975, n68976, n68977, n68978, n68979,
n68980, n68981, n68982, n68983, n68984, n68985, n68986, n68987,
n68988, n68989, n68990, n68991, n68992, n68993, n68994, n68995,
n68996, n68997, n68998, n68999, n69000, n69001, n69002, n69003,
n69004, n69005, n69006, n69007, n69008, n69009, n69010, n69011,
n69012, n69013, n69014, n69015, n69016, n69017, n69018, n69019,
n69020, n69021, n69022, n69023, n69024, n69025, n69026, n69027,
n69028, n69029, n69030, n69031, n69032, n69033, n69034, n69035,
n69036, n69037, n69038, n69039, n69040, n69041, n69042, n69043,
n69044, n69045, n69046, n69047, n69048, n69049, n69050, n69051,
n69052, n69053, n69054, n69055, n69056, n69057, n69058, n69059,
n69060, n69061, n69062, n69063, n69064, n69065, n69066, n69067,
n69068, n69069, n69070, n69071, n69072, n69073, n69074, n69075,
n69076, n69077, n69078, n69079, n69080, n69081, n69082, n69083,
n69084, n69085, n69086, n69087, n69088, n69089, n69090, n69091,
n69092, n69093, n69094, n69095, n69096, n69097, n69098, n69099,
n69100, n69101, n69102, n69103, n69104, n69105, n69106, n69107,
n69108, n69109, n69110, n69111, n69112, n69113, n69114, n69115,
n69116, n69117, n69118, n69119, n69120, n69121, n69122, n69123,
n69124, n69125, n69126, n69127, n69128, n69129, n69130, n69131,
n69132, n69133, n69134, n69135, n69136, n69137, n69138, n69139,
n69140, n69141, n69142, n69143, n69144, n69145, n69146, n69147,
n69148, n69149, n69150, n69151, n69152, n69153, n69154, n69155,
n69156, n69157, n69158, n69159, n69160, n69161, n69162, n69163,
n69164, n69165, n69166, n69167, n69168, n69169, n69170, n69171,
n69172, n69173, n69174, n69175, n69176, n69177, n69178, n69179,
n69180, n69181, n69182, n69183, n69184, n69185, n69186, n69187,
n69188, n69189, n69190, n69191, n69192, n69193, n69194, n69195,
n69196, n69197, n69198, n69199, n69200, n69201, n69202, n69203,
n69204, n69205, n69206, n69207, n69208, n69209, n69210, n69211,
n69212, n69213, n69214, n69215, n69216, n69217, n69218, n69219,
n69220, n69221, n69222, n69223, n69224, n69225, n69226, n69227,
n69228, n69229, n69230, n69231, n69232, n69233, n69234, n69235,
n69236, n69237, n69238, n69239, n69240, n69241, n69242, n69243,
n69244, n69245, n69246, n69247, n69248, n69249, n69250, n69251,
n69252, n69253, n69254, n69255, n69256, n69257, n69258, n69259,
n69260, n69261, n69262, n69263, n69264, n69265, n69266, n69267,
n69268, n69269, n69270, n69271, n69272, n69273, n69274, n69275,
n69276, n69277, n69278, n69279, n69280, n69281, n69282, n69283,
n69284, n69285, n69286, n69287, n69288, n69289, n69290, n69291,
n69292, n69293, n69294, n69295, n69296, n69297, n69298, n69299,
n69300, n69301, n69302, n69303, n69304, n69305, n69306, n69307,
n69308, n69309, n69310, n69311, n69312, n69313, n69314, n69315,
n69316, n69317, n69318, n69319, n69320, n69321, n69322, n69323,
n69324, n69325, n69326, n69327, n69328, n69329, n69330, n69331,
n69332, n69333, n69334, n69335, n69336, n69337, n69338, n69339,
n69340, n69341, n69342, n69343, n69344, n69345, n69346, n69347,
n69348, n69349, n69350, n69351, n69352, n69353, n69354, n69355,
n69356, n69357, n69358, n69359, n69360, n69361, n69362, n69363,
n69364, n69365, n69366, n69367, n69368, n69369, n69370, n69371,
n69372, n69373, n69374, n69375, n69376, n69377, n69378, n69379,
n69380, n69381, n69382, n69383, n69384, n69385, n69386, n69387,
n69388, n69389, n69390, n69391, n69392, n69393, n69394, n69395,
n69396, n69397, n69398, n69399, n69400, n69401, n69402, n69403,
n69404, n69405, n69406, n69407, n69408, n69409, n69410, n69411,
n69412, n69413, n69414, n69415, n69416, n69417, n69418, n69419,
n69420, n69421, n69422, n69423, n69424, n69425, n69426, n69427,
n69428, n69429, n69430, n69431, n69432, n69433, n69434, n69435,
n69436, n69437, n69438, n69439, n69440, n69441, n69442, n69443,
n69444, n69445, n69446, n69447, n69448, n69449, n69450, n69451,
n69452, n69453, n69454, n69455, n69456, n69457, n69458, n69459,
n69460, n69461, n69462, n69463, n69464, n69465, n69466, n69467,
n69468, n69469, n69470, n69471, n69472, n69473, n69474, n69475,
n69476, n69477, n69478, n69479, n69480, n69481, n69482, n69483,
n69484, n69485, n69486, n69487, n69488, n69489, n69490, n69491,
n69492, n69493, n69494, n69495, n69496, n69497, n69498, n69499,
n69500, n69501, n69502, n69503, n69504, n69505, n69506, n69507,
n69508, n69509, n69510, n69511, n69512, n69513, n69514, n69515,
n69516, n69517, n69518, n69519, n69520, n69521, n69522, n69523,
n69524, n69525, n69526, n69527, n69528, n69529, n69530, n69531,
n69532, n69533, n69534, n69535, n69536, n69537, n69538, n69539,
n69540, n69541, n69542, n69543, n69544, n69545, n69546, n69547,
n69548, n69549, n69550, n69551, n69552, n69553, n69554, n69555,
n69556, n69557, n69558, n69559, n69560, n69561, n69562, n69563,
n69564, n69565, n69566, n69567, n69568, n69569, n69570, n69571,
n69572, n69573, n69574, n69575, n69576, n69577, n69578, n69579,
n69580, n69581, n69582, n69583, n69584, n69585, n69586, n69587,
n69588, n69589, n69590, n69591, n69592, n69593, n69594, n69595,
n69596, n69597, n69598, n69599, n69600, n69601, n69602, n69603,
n69604, n69605, n69606, n69607, n69608, n69609, n69610, n69611,
n69612, n69613, n69614, n69615, n69616, n69617, n69618, n69619,
n69620, n69621, n69622, n69623, n69624, n69625, n69626, n69627,
n69628, n69629, n69630, n69631, n69632, n69633, n69634, n69635,
n69636, n69637, n69638, n69639, n69640, n69641, n69642, n69643,
n69644, n69645, n69646, n69647, n69648, n69649, n69650, n69651,
n69652, n69653, n69654, n69655, n69656, n69657, n69658, n69659,
n69660, n69661, n69662, n69663, n69664, n69665, n69666, n69667,
n69668, n69669, n69670, n69671, n69672, n69673, n69674, n69675,
n69676, n69677, n69678, n69679, n69680, n69681, n69682, n69683,
n69684, n69685, n69686, n69687, n69688, n69689, n69690, n69691,
n69692, n69693, n69694, n69695, n69696, n69697, n69698, n69699,
n69700, n69701, n69702, n69703, n69704, n69705, n69706, n69707,
n69708, n69709, n69710, n69711, n69712, n69713, n69714, n69715,
n69716, n69717, n69718, n69719, n69720, n69721, n69722, n69723,
n69724, n69725, n69726, n69727, n69728, n69729, n69730, n69731,
n69732, n69733, n69734, n69735, n69736, n69737, n69738, n69739,
n69740, n69741, n69742, n69743, n69744, n69745, n69746, n69747,
n69748, n69749, n69750, n69751, n69752, n69753, n69754, n69755,
n69756, n69757, n69758, n69759, n69760, n69761, n69762, n69763,
n69764, n69765, n69766, n69767, n69768, n69769, n69770, n69771,
n69772, n69773, n69774, n69775, n69776, n69777, n69778, n69779,
n69780, n69781, n69782, n69783, n69784, n69785, n69786, n69787,
n69788, n69789, n69790, n69791, n69792, n69793, n69794, n69795,
n69796, n69797, n69798, n69799, n69800, n69801, n69802, n69803,
n69804, n69805, n69806, n69807, n69808, n69809, n69810, n69811,
n69812, n69813, n69814, n69815, n69816, n69817, n69818, n69819,
n69820, n69821, n69822, n69823, n69824, n69825, n69826, n69827,
n69828, n69829, n69830, n69831, n69832, n69833, n69834, n69835,
n69836, n69837, n69838, n69839, n69840, n69841, n69842, n69843,
n69844, n69845, n69846, n69847, n69848, n69849, n69850, n69851,
n69852, n69853, n69854, n69855, n69856, n69857, n69858, n69859,
n69860, n69861, n69862, n69863, n69864, n69865, n69866, n69867,
n69868, n69869, n69870, n69871, n69872, n69873, n69874, n69875,
n69876, n69877, n69878, n69879, n69880, n69881, n69882, n69883,
n69884, n69885, n69886, n69887, n69888, n69889, n69890, n69891,
n69892, n69893, n69894, n69895, n69896, n69897, n69898, n69899,
n69900, n69901, n69902, n69903, n69904, n69905, n69906, n69907,
n69908, n69909, n69910, n69911, n69912, n69913, n69914, n69915,
n69916, n69917, n69918, n69919, n69920, n69921, n69922, n69923,
n69924, n69925, n69926, n69927, n69928, n69929, n69930, n69931,
n69932, n69933, n69934, n69935, n69936, n69937, n69938, n69939,
n69940, n69941, n69942, n69943, n69944, n69945, n69946, n69947,
n69948, n69949, n69950, n69951, n69952, n69953, n69954, n69955,
n69956, n69957, n69958, n69959, n69960, n69961, n69962, n69963,
n69964, n69965, n69966, n69967, n69968, n69969, n69970, n69971,
n69972, n69973, n69974, n69975, n69976, n69977, n69978, n69979,
n69980, n69981, n69982, n69983, n69984, n69985, n69986, n69987,
n69988, n69989, n69990, n69991, n69992, n69993, n69994, n69995,
n69996, n69997, n69998, n69999, n70000, n70001, n70002, n70003,
n70004, n70005, n70006, n70007, n70008, n70009, n70010, n70011,
n70012, n70013, n70014, n70015, n70016, n70017, n70018, n70019,
n70020, n70021, n70022, n70023, n70024, n70025, n70026, n70027,
n70028, n70029, n70030, n70031, n70032, n70033, n70034, n70035,
n70036, n70037, n70038, n70039, n70040, n70041, n70042, n70043,
n70044, n70045, n70046, n70047, n70048, n70049, n70050, n70051,
n70052, n70053, n70054, n70055, n70056, n70057, n70058, n70059,
n70060, n70061, n70062, n70063, n70064, n70065, n70066, n70067,
n70068, n70069, n70070, n70071, n70072, n70073, n70074, n70075,
n70076, n70077, n70078, n70079, n70080, n70081, n70082, n70083,
n70084, n70085, n70086, n70087, n70088, n70089, n70090, n70091,
n70092, n70093, n70094, n70095, n70096, n70097, n70098, n70099,
n70100, n70101, n70102, n70103, n70104, n70105, n70106, n70107,
n70108, n70109, n70110, n70111, n70112, n70113, n70114, n70115,
n70116, n70117, n70118, n70119, n70120, n70121, n70122, n70123,
n70124, n70125, n70126, n70127, n70128, n70129, n70130, n70131,
n70132, n70133, n70134, n70135, n70136, n70137, n70138, n70139,
n70140, n70141, n70142, n70143, n70144, n70145, n70146, n70147,
n70148, n70149, n70150, n70151, n70152, n70153, n70154, n70155,
n70156, n70157, n70158, n70159, n70160, n70161, n70162, n70163,
n70164, n70165, n70166, n70167, n70168, n70169, n70170, n70171,
n70172, n70173, n70174, n70175, n70176, n70177, n70178, n70179,
n70180, n70181, n70182, n70183, n70184, n70185, n70186, n70187,
n70188, n70189, n70190, n70191, n70192, n70193, n70194, n70195,
n70196, n70197, n70198, n70199, n70200, n70201, n70202, n70203,
n70204, n70205, n70206, n70207, n70208, n70209, n70210, n70211,
n70212, n70213, n70214, n70215, n70216, n70217, n70218, n70219,
n70220, n70221, n70222, n70223, n70224, n70225, n70226, n70227,
n70228, n70229, n70230, n70231, n70232, n70233, n70234, n70235,
n70236, n70237, n70238, n70239, n70240, n70241, n70242, n70243,
n70244, n70245, n70246, n70247, n70248, n70249, n70250, n70251,
n70252, n70253, n70254, n70255, n70256, n70257, n70258, n70259,
n70260, n70261, n70262, n70263, n70264, n70265, n70266, n70267,
n70268, n70269, n70270, n70271, n70272, n70273, n70274, n70275,
n70276, n70277, n70278, n70279, n70280, n70281, n70282, n70283,
n70284, n70285, n70286, n70287, n70288, n70289, n70290, n70291,
n70292, n70293, n70294, n70295, n70296, n70297, n70298, n70299,
n70300, n70301, n70302, n70303, n70304, n70305, n70306, n70307,
n70308, n70309, n70310, n70311, n70312, n70313, n70314, n70315,
n70316, n70317, n70318, n70319, n70320, n70321, n70322, n70323,
n70324, n70325, n70326, n70327, n70328, n70329, n70330, n70331,
n70332, n70333, n70334, n70335, n70336, n70337, n70338, n70339,
n70340, n70341, n70342, n70343, n70344, n70345, n70346, n70347,
n70348, n70349, n70350, n70351, n70352, n70353, n70354, n70355,
n70356, n70357, n70358, n70359, n70360, n70361, n70362, n70363,
n70364, n70365, n70366, n70367, n70368, n70369, n70370, n70371,
n70372, n70373, n70374, n70375, n70376, n70377, n70378, n70379,
n70380, n70381, n70382, n70383, n70384, n70385, n70386, n70387,
n70388, n70389, n70390, n70391, n70392, n70393, n70394, n70395,
n70396, n70397, n70398, n70399, n70400, n70401, n70402, n70403,
n70404, n70405, n70406, n70407, n70408, n70409, n70410, n70411,
n70412, n70413, n70414, n70415, n70416, n70417, n70418, n70419,
n70420, n70421, n70422, n70423, n70424, n70425, n70426, n70427,
n70428, n70429, n70430, n70431, n70432, n70433, n70434, n70435,
n70436, n70437, n70438, n70439, n70440, n70441, n70442, n70443,
n70444, n70445, n70446, n70447, n70448, n70449, n70450, n70451,
n70452, n70453, n70454, n70455, n70456, n70457, n70458, n70459,
n70460, n70461, n70462, n70463, n70464, n70465, n70466, n70467,
n70468, n70469, n70470, n70471, n70472, n70473, n70474, n70475,
n70476, n70477, n70478, n70479, n70480, n70481, n70482, n70483,
n70484, n70485, n70486, n70487, n70488, n70489, n70490, n70491,
n70492, n70493, n70494, n70495, n70496, n70497, n70498, n70499,
n70500, n70501, n70502, n70503, n70504, n70505, n70506, n70507,
n70508, n70509, n70510, n70511, n70512, n70513, n70514, n70515,
n70516, n70517, n70518, n70519, n70520, n70521, n70522, n70523,
n70524, n70525, n70526, n70527, n70528, n70529, n70530, n70531,
n70532, n70533, n70534, n70535, n70536, n70537, n70538, n70539,
n70540, n70541, n70542, n70543, n70544, n70545, n70546, n70547,
n70548, n70549, n70550, n70551, n70552, n70553, n70554, n70555,
n70556, n70557, n70558, n70559, n70560, n70561, n70562, n70563,
n70564, n70565, n70566, n70567, n70568, n70569, n70570, n70571,
n70572, n70573, n70574, n70575, n70576, n70577, n70578, n70579,
n70580, n70581, n70582, n70583, n70584, n70585, n70586, n70587,
n70588, n70589, n70590, n70591, n70592, n70593, n70594, n70595,
n70596, n70597, n70598, n70599, n70600, n70601, n70602, n70603,
n70604, n70605, n70606, n70607, n70608, n70609, n70610, n70611,
n70612, n70613, n70614, n70615, n70616, n70617, n70618, n70619,
n70620, n70621, n70622, n70623, n70624, n70625, n70626, n70627,
n70628, n70629, n70630, n70631, n70632, n70633, n70634, n70635,
n70636, n70637, n70638, n70639, n70640, n70641, n70642, n70643,
n70644, n70645, n70646, n70647, n70648, n70649, n70650, n70651,
n70652, n70653, n70654, n70655, n70656, n70657, n70658, n70659,
n70660, n70661, n70662, n70663, n70664, n70665, n70666, n70667,
n70668, n70669, n70670, n70671, n70672, n70673, n70674, n70675,
n70676, n70677, n70678, n70679, n70680, n70681, n70682, n70683,
n70684, n70685, n70686, n70687, n70688, n70689, n70690, n70691,
n70692, n70693, n70694, n70695, n70696, n70697, n70698, n70699,
n70700, n70701, n70702, n70703, n70704, n70705, n70706, n70707,
n70708, n70709, n70710, n70711, n70712, n70713, n70714, n70715,
n70716, n70717, n70718, n70719, n70720, n70721, n70722, n70723,
n70724, n70725, n70726, n70727, n70728, n70729, n70730, n70731,
n70732, n70733, n70734, n70735, n70736, n70737, n70738, n70739,
n70740, n70741, n70742, n70743, n70744, n70745, n70746, n70747,
n70748, n70749, n70750, n70751, n70752, n70753, n70754, n70755,
n70756, n70757, n70758, n70759, n70760, n70761, n70762, n70763,
n70764, n70765, n70766, n70767, n70768, n70769, n70770, n70771,
n70772, n70773, n70774, n70775, n70776, n70777, n70778, n70779,
n70780, n70781, n70782, n70783, n70784, n70785, n70786, n70787,
n70788, n70789, n70790, n70791, n70792, n70793, n70794, n70795,
n70796, n70797, n70798, n70799, n70800, n70801, n70802, n70803,
n70804, n70805, n70806, n70807, n70808, n70809, n70810, n70811,
n70812, n70814, n70815, n70816, n70817, n70818, n70819, n70820,
n70821, n70822, n70823, n70824, n70825, n70826, n70827, n70828,
n70829, n70830, n70831, n70832, n70833, n70834, n70835, n70836,
n70837, n70838, n70839, n70840, n70841, n70842, n70843, n70844,
n70845, n70846, n70847, n70848, n70849, n70850, n70851, n70852,
n70853, n70854, n70855, n70856, n70857, n70858, n70859, n70860,
n70861, n70862, n70863, n70864, n70865, n70866, n70867, n70868,
n70869, n70870, n70871, n70872, n70873, n70874, n70875, n70876,
n70877, n70878, n70879, n70880, n70881, n70882, n70883, n70884,
n70885, n70886, n70887, n70888, n70889, n70890, n70891, n70892,
n70893, n70894, n70895, n70896, n70897, n70898, n70899, n70900,
n70901, n70902, n70903, n70904, n70905, n70906, n70907, n70908,
n70909, n70910, n70911, n70912, n70913, n70914, n70915, n70916,
n70917, n70918, n70919, n70920, n70921, n70922, n70923, n70924,
n70925, n70926, n70927, n70928, n70929, n70930, n70931, n70932,
n70933, n70934, n70935, n70936, n70937, n70938, n70939, n70940,
n70941, n70942, n70943, n70944, n70945, n70946, n70947, n70948,
n70949, n70950, n70951, n70952, n70953, n70954, n70955, n70956,
n70957, n70958, n70959, n70960, n70961, n70962, n70963, n70964,
n70965, n70966, n70967, n70968, n70969, n70970, n70971, n70972,
n70973, n70974, n70975, n70976, n70979, n70980, n70981, n70982,
n70983, n70984, n70985, n70986, n70987, n70988, n70989, n70990,
n70991, n70992, n70993, n70994, n70995, n70996, n70997, n70998,
n70999, n71000, n71001, n71002, n71003, n71004, n71005, n71006,
n71007, n71008, n71009, n71010, n71011, n71012, n71013, n71014,
n71015, n71016, n71017, n71018, n71019, n71020, n71021, n71022,
n71023, n71024, n71025, n71026, n71027, n71028, n71029, n71030,
n71031, n71032, n71033, n71034, n71035, n71036, n71037, n71038,
n71039, n71040, n71041, n71042, n71043, n71044, n71045, n71046,
n71047, n71048, n71049, n71050, n71051, n71052, n71053, n71054,
n71055, n71056, n71057, n71058, n71059, n71060, n71061, n71062,
n71063, n71064, n71065, n71066, n71067, n71068, n71069, n71070,
n71071, n71072, n71073, n71074, n71075, n71076, n71077, n71078,
n71079, n71080, n71081, n71082, n71083, n71084, n71085, n71086,
n71087, n71088, n71089, n71090, n71091, n71092, n71093, n71094,
n71095, n71096, n71097, n71098, n71099, n71100, n71101, n71102,
n71103, n71104, n71105, n71106, n71107, n71108, n71109, n71110,
n71111, n71112, n71113, n71114, n71115, n71116, n71117, n71118,
n71119, n71120, n71121, n71122, n71123, n71124, n71125, n71126,
n71127, n71128, n71129, n71130, n71131, n71132, n71133, n71134,
n71135, n71136, n71137, n71138, n71139, n71140, n71141, n71142,
n71143, n71144, n71145, n71146, n71147, n71148, n71149, n71150,
n71151, n71152, n71153, n71154, n71155, n71156, n71157, n71158,
n71159, n71160, n71161, n71162, n71163, n71164, n71165, n71166,
n71167, n71168, n71169, n71170, n71171, n71172, n71173, n71174,
n71175, n71176, n71177, n71178, n71179, n71180, n71181, n71182,
n71183, n71184, n71185, n71186, n71187, n71188, n71189, n71190,
n71191, n71192, n71193, n71194, n71195, n71196, n71197, n71198,
n71199, n71200, n71201, n71202, n71203, n71204, n71205, n71206,
n71207, n71208, n71209, n71210, n71211, n71212, n71213, n71214,
n71215, n71216, n71217, n71218, n71219, n71220, n71221, n71222,
n71223, n71224, n71225, n71226, n71227, n71228, n71229, n71230,
n71231, n71232, n71233, n71234, n71235, n71236, n71237, n71238,
n71239, n71240, n71241, n71242, n71243, n71244, n71245, n71246,
n71247, n71248, n71249, n71250, n71251, n71252, n71253, n71254,
n71255, n71256, n71257, n71258, n71259, n71260, n71261, n71262,
n71263, n71264, n71265, n71266, n71267, n71268, n71269, n71270,
n71271, n71272, n71273, n71274, n71275, n71276, n71277, n71278,
n71279, n71280, n71281, n71282, n71283, n71284, n71285, n71286,
n71287, n71288, n71289, n71290, n71291, n71292, n71293, n71294,
n71295, n71296, n71297, n71298, n71299, n71300, n71301, n71302,
n71303, n71304, n71305, n71306, n71307, n71308, n71309, n71310,
n71311, n71312, n71313, n71314, n71315, n71316, n71317, n71318,
n71319, n71320, n71321, n71322, n71323, n71324, n71325, n71326,
n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334,
n71335, n71336, n71337, n71338, n71339, n71340, n71341, n71342,
n71343, n71344, n71345, n71346, n71347, n71348, n71349, n71350,
n71351, n71352, n71353, n71354, n71355, n71356, n71357, n71358,
n71359, n71360, n71361, n71362, n71363, n71364, n71365, n71366,
n71367, n71368, n71369, n71370, n71371, n71372, n71373, n71374,
n71375, n71376, n71377, n71378, n71379, n71380, n71381, n71382,
n71383, n71384, n71385, n71386, n71387, n71388, n71389, n71390,
n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398,
n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406,
n71407, n71408, n71409, n71410, n71411, n71412, n71413, n71414,
n71415, n71416, n71417, n71418, n71419, n71420, n71421, n71422,
n71423, n71424, n71425, n71426, n71427, n71428, n71429, n71430,
n71431, n71432, n71433, n71434, n71435, n71436, n71437, n71438,
n71439, n71440, n71441, n71442, n71443, n71444, n71445, n71446,
n71447, n71448, n71449, n71450, n71451, n71452, n71453, n71454,
n71455, n71456, n71457, n71458, n71459, n71460, n71461, n71462,
n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470,
n71471, n71472, n71473, n71474, n71475, n71476, n71477, n71478,
n71479, n71480, n71481, n71482, n71483, n71484, n71485, n71486,
n71487, n71488, n71489, n71490, n71491, n71492, n71493, n71494,
n71495, n71496, n71497, n71498, n71499, n71500, n71501, n71502,
n71503, n71504, n71505, n71506, n71507, n71508, n71509, n71510,
n71511, n71512, n71513, n71514, n71515, n71516, n71517, n71518,
n71519, n71520, n71521, n71522, n71523, n71524, n71525, n71526,
n71527, n71528, n71529, n71530, n71531, n71532, n71533, n71534,
n71535, n71536, n71537, n71538, n71539, n71540, n71541, n71542,
n71543, n71544, n71545, n71546, n71547, n71548, n71549, n71550,
n71551, n71552, n71553, n71554, n71555, n71556, n71557, n71558,
n71559, n71560, n71561, n71562, n71563, n71564, n71565, n71566,
n71567, n71568, n71569, n71570, n71571, n71572, n71573, n71574,
n71575, n71576, n71577, n71578, n71579, n71580, n71581, n71582,
n71583, n71584, n71585, n71586, n71587, n71588, n71589, n71590,
n71591, n71592, n71593, n71594, n71595, n71596, n71597, n71598,
n71599, n71600, n71601, n71602, n71603, n71604, n71605, n71606,
n71607, n71608, n71609, n71610, n71611, n71612, n71613, n71614,
n71615, n71616, n71617, n71618, n71619, n71620, n71621, n71622,
n71623, n71624, n71625, n71626, n71627, n71628, n71629, n71630,
n71631, n71632, n71633, n71634, n71635, n71636, n71637, n71638,
n71639, n71640, n71641, n71642, n71643, n71644, n71645, n71646,
n71647, n71648, n71649, n71650, n71651, n71652, n71653, n71654,
n71655, n71656, n71657, n71658, n71659, n71660, n71661, n71662,
n71663, n71664, n71665, n71666, n71667, n71668, n71669, n71670,
n71671, n71672, n71673, n71674, n71675, n71676, n71677, n71678,
n71679, n71680, n71681, n71682, n71683, n71684, n71685, n71686,
n71687, n71688, n71689, n71690, n71691, n71692, n71693, n71694,
n71695, n71696, n71697, n71698, n71699, n71700, n71701, n71702,
n71703, n71704, n71705, n71706, n71707, n71708, n71709, n71710,
n71711, n71712, n71713, n71714, n71715, n71716, n71717, n71718,
n71719, n71720, n71721, n71722, n71723, n71724, n71725, n71726,
n71727, n71728, n71729, n71730, n71731, n71732, n71733, n71734,
n71735, n71736, n71737, n71738, n71739, n71740, n71741, n71742,
n71743, n71744, n71745, n71746, n71747, n71748, n71749, n71750,
n71751, n71752, n71753, n71754, n71755, n71756, n71757, n71758,
n71759, n71760, n71761, n71762, n71763, n71764, n71765, n71766,
n71767, n71768, n71769, n71770, n71771, n71772, n71773, n71774,
n71775, n71776, n71777, n71778, n71779, n71780, n71781, n71782,
n71783, n71784, n71785, n71786, n71787, n71788, n71789, n71790,
n71791, n71792, n71793, n71794, n71795, n71796, n71797, n71798,
n71799, n71800, n71801, n71802, n71803, n71804, n71805, n71806,
n71807, n71808, n71809, n71810, n71811, n71813, n71814, n71815,
n71816, n71817, n71818, n71819, n71820, n71821, n71822, n71823,
n71824, n71825, n71826, n71827, n71828, n71829, n71830, n71831,
n71832, n71833, n71834, n71835, n71836, n71837, n71838, n71839,
n71840, n71841, n71842, n71843, n71844, n71845, n71846, n71847,
n71848, n71849, n71850, n71851, n71852, n71853, n71854, n71855,
n71856, n71857, n71858, n71859, n71860, n71861, n71862, n71863,
n71864, n71865, n71866, n71867, n71868, n71869, n71870, n71871,
n71872, n71873, n71874, n71875, n71876, n71877, n71878, n71879,
n71880, n71881, n71882, n71883, n71884, n71885, n71886, n71887,
n71888, n71889, n71890, n71891, n71892, n71893, n71894, n71895,
n71896, n71897, n71898, n71899, n71900, n71901, n71902, n71903,
n71904, n71905, n71906, n71907, n71908, n71909, n71910, n71911,
n71912, n71913, n71914, n71915, n71916, n71917, n71918, n71919,
n71920, n71921, n71922, n71923, n71924, n71925, n71926, n71927,
n71928, n71929, n71930, n71931, n71932, n71933, n71934, n71935,
n71936, n71937, n71938, n71939, n71940, n71941, n71942, n71943,
n71944, n71945, n71946, n71947, n71948, n71949, n71950, n71951,
n71952, n71953, n71954, n71955, n71956, n71957, n71958, n71959,
n71960, n71961, n71962, n71963, n71964, n71965, n71966, n71967,
n71968, n71969, n71970, n71971, n71972, n71973, n71974, n71975,
n71976, n71977, n71978, n71979, n71980, n71981, n71982, n71983,
n71984, n71985, n71986, n71987, n71988, n71989, n71990, n71991,
n71992, n71993, n71994, n71995, n71996, n71997, n71998, n71999,
n72000, n72001, n72002, n72003, n72004, n72005, n72006, n72007,
n72008, n72009, n72010, n72011, n72012, n72013, n72014, n72015,
n72016, n72017, n72018, n72019, n72020, n72021, n72022, n72023,
n72024, n72025, n72026, n72027, n72028, n72029, n72030, n72031,
n72032, n72033, n72034, n72035, n72036, n72037, n72038, n72039,
n72040, n72041, n72042, n72043, n72044, n72045, n72046, n72047,
n72048, n72049, n72050, n72051, n72052, n72053, n72054, n72055,
n72056, n72057, n72058, n72059, n72060, n72061, n72062, n72063,
n72064, n72065, n72066, n72067, n72068, n72069, n72070, n72071,
n72072, n72073, n72074, n72075, n72076, n72077, n72078, n72079,
n72080, n72081, n72082, n72083, n72084, n72085, n72086, n72087,
n72088, n72089, n72090, n72091, n72092, n72093, n72094, n72095,
n72096, n72097, n72098, n72099, n72100, n72101, n72102, n72103,
n72104, n72105, n72106, n72107, n72108, n72109, n72110, n72111,
n72112, n72113, n72114, n72115, n72116, n72117, n72118, n72119,
n72120, n72121, n72122, n72123, n72124, n72125, n72126, n72127,
n72128, n72129, n72130, n72131, n72132, n72133, n72134, n72135,
n72136, n72137, n72138, n72139, n72140, n72141, n72142, n72143,
n72144, n72145, n72146, n72147, n72148, n72149, n72150, n72151,
n72152, n72153, n72154, n72155, n72156, n72157, n72158, n72159,
n72160, n72161, n72162, n72163, n72164, n72165, n72166, n72167,
n72168, n72169, n72170, n72171, n72172, n72173, n72174, n72175,
n72176, n72177, n72178, n72179, n72180, n72181, n72182, n72183,
n72184, n72185, n72186, n72187, n72188, n72189, n72190, n72191,
n72192, n72193, n72194, n72195, n72196, n72197, n72198, n72199,
n72200, n72201, n72202, n72203, n72204, n72205, n72206, n72207,
n72208, n72209, n72210, n72211, n72212, n72213, n72214, n72215,
n72216, n72217, n72218, n72219, n72220, n72221, n72222, n72223,
n72224, n72225, n72226, n72227, n72228, n72229, n72230, n72231,
n72232, n72233, n72234, n72235, n72236, n72237, n72238, n72239,
n72240, n72241, n72242, n72243, n72244, n72245, n72246, n72247,
n72248, n72249, n72250, n72251, n72252, n72253, n72254, n72255,
n72256, n72257, n72258, n72259, n72260, n72261, n72262, n72263,
n72264, n72265, n72266, n72267, n72268, n72269, n72270, n72271,
n72272, n72273, n72274, n72275, n72276, n72277, n72278, n72279,
n72280, n72281, n72282, n72283, n72284, n72285, n72286, n72287,
n72288, n72289, n72290, n72291, n72292, n72293, n72294, n72295,
n72296, n72297, n72298, n72299, n72300, n72301, n72302, n72303,
n72304, n72305, n72306, n72307, n72308, n72309, n72310, n72311,
n72312, n72313, n72314, n72315, n72316, n72317, n72318, n72319,
n72320, n72321, n72322, n72323, n72324, n72325, n72326, n72327,
n72328, n72329, n72330, n72331, n72332, n72333, n72334, n72335,
n72336, n72337, n72338, n72339, n72340, n72341, n72342, n72343,
n72344, n72345, n72346, n72347, n72348, n72349, n72350, n72351,
n72352, n72353, n72354, n72355, n72356, n72357, n72358, n72359,
n72360, n72361, n72362, n72363, n72364, n72365, n72366, n72367,
n72368, n72369, n72370, n72371, n72372, n72373, n72374, n72375,
n72376, n72377, n72378, n72379, n72380, n72381, n72382, n72383,
n72384, n72385, n72386, n72387, n72388, n72389, n72390, n72391,
n72392, n72393, n72394, n72395, n72396, n72397, n72398, n72399,
n72400, n72401, n72402, n72403, n72404, n72405, n72406, n72407,
n72408, n72409, n72410, n72411, n72412, n72413, n72414, n72415,
n72416, n72417, n72418, n72419, n72420, n72421, n72422, n72423,
n72424, n72425, n72426, n72427, n72428, n72429, n72430, n72431,
n72432, n72433, n72434, n72435, n72436, n72437, n72438, n72439,
n72440, n72441, n72442, n72443, n72444, n72445, n72446, n72447,
n72448, n72449, n72450, n72451, n72452, n72453, n72454, n72455,
n72456, n72457, n72458, n72459, n72460, n72461, n72462, n72463,
n72464, n72465, n72466, n72467, n72468, n72469, n72470, n72471,
n72472, n72473, n72474, n72475, n72476, n72477, n72478, n72479,
n72480, n72481, n72482, n72483, n72484, n72485, n72486, n72487,
n72488, n72489, n72490, n72491, n72492, n72493, n72494, n72495,
n72496, n72497, n72498, n72499, n72500, n72501, n72502, n72503,
n72504, n72505, n72506, n72507, n72508, n72509, n72510, n72511,
n72512, n72513, n72514, n72515, n72516, n72517, n72518, n72519,
n72520, n72521, n72522, n72523, n72524, n72525, n72526, n72527,
n72528, n72529, n72530, n72531, n72532, n72533, n72534, n72535,
n72536, n72537, n72538, n72539, n72540, n72541, n72542, n72543,
n72544, n72545, n72546, n72547, n72548, n72549, n72550, n72551,
n72552, n72553, n72554, n72555, n72556, n72557, n72558, n72559,
n72560, n72561, n72562, n72563, n72564, n72565, n72566, n72567,
n72568, n72569, n72570, n72571, n72572, n72573, n72574, n72575,
n72576, n72577, n72578, n72579, n72580, n72581, n72582, n72583,
n72584, n72585, n72586, n72587, n72588, n72589, n72590, n72591,
n72592, n72593, n72594, n72595, n72596, n72597, n72598, n72599,
n72600, n72601, n72602, n72603, n72604, n72605, n72606, n72607,
n72608, n72609, n72610, n72611, n72612, n72613, n72614, n72615,
n72616, n72617, n72618, n72619, n72620, n72621, n72622, n72623,
n72624, n72625, n72626, n72627, n72628, n72629, n72630, n72631,
n72632, n72633, n72634, n72635, n72636, n72637, n72638, n72639,
n72640, n72641, n72642, n72643, n72644, n72645, n72646, n72647,
n72648, n72649, n72650, n72651, n72652, n72653, n72654, n72655,
n72656, n72657, n72658, n72659, n72660, n72661, n72662, n72663,
n72664, n72665, n72666, n72667, n72668, n72669, n72670, n72671,
n72672, n72673, n72674, n72675, n72676, n72677, n72678, n72679,
n72680, n72681, n72682, n72683, n72684, n72685, n72686, n72687,
n72688, n72689, n72690, n72691, n72692, n72693, n72694, n72695,
n72696, n72697, n72698, n72699, n72700, n72701, n72702, n72703,
n72704, n72705, n72706, n72707, n72708, n72709, n72710, n72711,
n72712, n72713, n72714, n72715, n72716, n72717, n72718, n72719,
n72720, n72721, n72722, n72723, n72724, n72725, n72726, n72727,
n72728, n72729, n72730, n72731, n72732, n72733, n72734, n72735,
n72736, n72737, n72738, n72739, n72740, n72741, n72742, n72743,
n72744, n72745, n72746, n72747, n72748, n72749, n72750, n72751,
n72752, n72753, n72754, n72755, n72756, n72757, n72758, n72759,
n72760, n72761, n72762, n72763, n72764, n72765, n72766, n72767,
n72768, n72769, n72770, n72771, n72772, n72773, n72774, n72775,
n72776, n72777, n72778, n72779, n72780, n72781, n72782, n72783,
n72784, n72785, n72786, n72787, n72788, n72789, n72790, n72791,
n72792, n72793, n72794, n72795, n72796, n72797, n72798, n72799,
n72800, n72801, n72802, n72803, n72804, n72805, n72806, n72807,
n72808, n72809, n72810, n72811, n72812, n72813, n72814, n72815,
n72816, n72817, n72818, n72819, n72820, n72821, n72822, n72823,
n72824, n72825, n72826, n72827, n72828, n72829, n72830, n72831,
n72832, n72833, n72834, n72835, n72836, n72837, n72838, n72839,
n72840, n72841, n72842, n72843, n72844, n72845, n72846, n72847,
n72848, n72849, n72850, n72851, n72852, n72853, n72854, n72855,
n72856, n72857, n72858, n72859, n72860, n72861, n72862, n72863,
n72864, n72865, n72866, n72867, n72868, n72869, n72870, n72871,
n72872, n72873, n72874, n72875, n72876, n72877, n72878, n72879,
n72880, n72881, n72882, n72883, n72884, n72885, n72886, n72887,
n72888, n72889, n72890, n72891, n72892, n72893, n72894, n72895,
n72896, n72897, n72898, n72899, n72900, n72901, n72902, n72903,
n72904, n72905, n72906, n72907, n72908, n72909, n72910, n72911,
n72912, n72913, n72914, n72915, n72916, n72917, n72918, n72919,
n72920, n72921, n72922, n72923, n72924, n72925, n72926, n72927,
n72928, n72929, n72930, n72931, n72932, n72933, n72934, n72935,
n72936, n72937, n72938, n72939, n72940, n72941, n72942, n72943,
n72944, n72945, n72946, n72947, n72948, n72949, n72950, n72951,
n72952, n72953, n72954, n72955, n72956, n72957, n72958, n72959,
n72960, n72961, n72962, n72963, n72964, n72965, n72966, n72967,
n72968, n72969, n72970, n72971, n72972, n72973, n72974, n72975,
n72976, n72977, n72978, n72979, n72980, n72981, n72982, n72983,
n72984, n72985, n72986, n72987, n72988, n72989, n72990, n72991,
n72992, n72993, n72994, n72995, n72996, n72997, n72998, n72999,
n73000, n73001, n73002, n73003, n73004, n73005, n73006, n73007,
n73008, n73009, n73010, n73011, n73012, n73013, n73014, n73015,
n73016, n73017, n73018, n73019, n73020, n73021, n73022, n73023,
n73024, n73025, n73026, n73027, n73028, n73029, n73030, n73031,
n73032, n73033, n73034, n73035, n73036, n73037, n73038, n73039,
n73040, n73041, n73042, n73043, n73044, n73045, n73046, n73047,
n73048, n73049, n73050, n73051, n73052, n73053, n73054, n73055,
n73056, n73057, n73058, n73059, n73060, n73061, n73062, n73063,
n73064, n73065, n73066, n73067, n73068, n73069, n73070, n73071,
n73072, n73073, n73074, n73075, n73076, n73077, n73078, n73079,
n73080, n73081, n73082, n73083, n73084, n73085, n73086, n73087,
n73088, n73089, n73090, n73091, n73092, n73093, n73094, n73095,
n73096, n73097, n73098, n73099, n73100, n73101, n73102, n73103,
n73104, n73105, n73106, n73107, n73108, n73109, n73110, n73111,
n73112, n73113, n73114, n73115, n73116, n73117, n73118, n73119,
n73120, n73121, n73122, n73123, n73124, n73125, n73126, n73127,
n73128, n73129, n73130, n73131, n73132, n73133, n73134, n73135,
n73136, n73137, n73138, n73139, n73140, n73141, n73142, n73143,
n73144, n73145, n73146, n73147, n73148, n73149, n73150, n73151,
n73152, n73153, n73154, n73155, n73156, n73157, n73158, n73159,
n73160, n73161, n73162, n73163, n73164, n73165, n73166, n73167,
n73168, n73169, n73170, n73171, n73172, n73173, n73174, n73175,
n73176, n73177, n73178, n73179, n73180, n73181, n73182, n73183,
n73184, n73185, n73186, n73187, n73188, n73189, n73190, n73191,
n73192, n73193, n73194, n73195, n73196, n73197, n73198, n73199,
n73200, n73201, n73202, n73203, n73204, n73205, n73206, n73207,
n73208, n73209, n73210, n73211, n73212, n73213, n73214, n73215,
n73216, n73217, n73218, n73219, n73220, n73221, n73222, n73223,
n73224, n73225, n73226, n73227, n73228, n73229, n73230, n73231,
n73232, n73233, n73234, n73235, n73236, n73237, n73238, n73239,
n73240, n73241, n73242, n73243, n73244, n73245, n73246, n73247,
n73248, n73249, n73250, n73251, n73252, n73253, n73254, n73255,
n73256, n73257, n73258, n73259, n73260, n73261, n73262, n73263,
n73264, n73265, n73266, n73267, n73268, n73269, n73270, n73271,
n73272, n73273, n73274, n73275, n73276, n73277, n73278, n73279,
n73280, n73281, n73282, n73283, n73284, n73285, n73286, n73287,
n73288, n73289, n73290, n73291, n73292, n73293, n73294, n73295,
n73296, n73297, n73298, n73299, n73300, n73301, n73302, n73303,
n73304, n73305, n73306, n73307, n73308, n73309, n73310, n73311,
n73312, n73313, n73314, n73315, n73316, n73317, n73318, n73319,
n73320, n73321, n73322, n73323, n73324, n73325, n73326, n73327,
n73328, n73329, n73330, n73331, n73332, n73333, n73334, n73335,
n73336, n73337, n73338, n73339, n73340, n73341, n73342, n73343,
n73344, n73345, n73346, n73347, n73348, n73349, n73350, n73351,
n73352, n73353, n73354, n73355, n73356, n73357, n73358, n73359,
n73360, n73361, n73362, n73363, n73364, n73365, n73366, n73367,
n73368, n73369, n73370, n73371, n73372, n73373, n73374, n73375,
n73376, n73377, n73378, n73379, n73380, n73381, n73382, n73383,
n73384, n73385, n73386, n73387, n73388, n73389, n73390, n73391,
n73392, n73393, n73394, n73395, n73396, n73397, n73398, n73399,
n73400, n73401, n73402, n73403, n73404, n73405, n73406, n73407,
n73408, n73409, n73410, n73411, n73412, n73413, n73414, n73415,
n73416, n73417, n73418, n73419, n73420, n73421, n73422, n73423,
n73424, n73425, n73426, n73427, n73428, n73429, n73430, n73431,
n73432, n73433, n73434, n73435, n73436, n73437, n73438, n73439,
n73440, n73441, n73442, n73443, n73444, n73445, n73446, n73447,
n73448, n73449, n73450, n73451, n73452, n73453, n73454, n73455,
n73456, n73457, n73458, n73459, n73460, n73461, n73462, n73463,
n73464, n73465, n73466, n73467, n73468, n73469, n73470, n73471,
n73472, n73473, n73474, n73475, n73476, n73477, n73478, n73479,
n73480, n73481, n73482, n73483, n73484, n73485, n73486, n73487,
n73488, n73489, n73490, n73491, n73492, n73493, n73494, n73495,
n73496, n73497, n73498, n73499, n73500, n73501, n73502, n73503,
n73504, n73505, n73506, n73507, n73508, n73509, n73510, n73511,
n73512, n73513, n73514, n73515, n73516, n73517, n73518, n73519,
n73520, n73521, n73522, n73523, n73524, n73525, n73526, n73527,
n73528, n73529, n73530, n73531, n73532, n73533, n73534, n73535,
n73536, n73537, n73538, n73539, n73540, n73541, n73542, n73543,
n73544, n73545, n73546, n73547, n73548, n73549, n73550, n73551,
n73552, n73553, n73554, n73555, n73556, n73557, n73558, n73559,
n73560, n73561, n73562, n73563, n73564, n73565, n73566, n73567,
n73568, n73569, n73570, n73571, n73572, n73573, n73574, n73575,
n73576, n73577, n73578, n73579, n73580, n73581, n73582, n73583,
n73584, n73585, n73586, n73587, n73588, n73589, n73590, n73591,
n73592, n73593, n73594, n73595, n73596, n73597, n73598, n73599,
n73600, n73601, n73602, n73603, n73604, n73605, n73606, n73607,
n73608, n73609, n73610, n73611, n73612, n73613, n73614, n73615,
n73616, n73617, n73618, n73619, n73620, n73621, n73622, n73623,
n73624, n73625, n73626, n73627, n73628, n73629, n73630, n73631,
n73632, n73633, n73634, n73635, n73636, n73637, n73638, n73639,
n73640, n73641, n73642, n73643, n73644, n73645, n73646, n73647,
n73648, n73649, n73650, n73651, n73652, n73653, n73654, n73655,
n73656, n73657, n73658, n73659, n73660, n73661, n73662, n73663,
n73664, n73665, n73666, n73667, n73668, n73669, n73670, n73671,
n73672, n73673, n73674, n73675, n73676, n73677, n73678, n73679,
n73680, n73681, n73682, n73683, n73684, n73685, n73686, n73687,
n73688, n73689, n73690, n73691, n73692, n73693, n73694, n73695,
n73696, n73697, n73698, n73699, n73700, n73701, n73702, n73703,
n73704, n73705, n73706, n73707, n73708, n73709, n73710, n73711,
n73712, n73713, n73714, n73715, n73716, n73717, n73718, n73719,
n73720, n73721, n73722, n73723, n73724, n73725, n73726, n73727,
n73728, n73729, n73730, n73731, n73732, n73733, n73734, n73735,
n73736, n73737, n73738, n73739, n73740, n73741, n73742, n73743,
n73744, n73745, n73746, n73747, n73748, n73749, n73750, n73751,
n73752, n73753, n73754, n73755, n73756, n73757, n73758, n73759,
n73760, n73761, n73762, n73763, n73764, n73765, n73766, n73767,
n73768, n73769, n73770, n73771, n73772, n73773, n73774, n73775,
n73776, n73777, n73778, n73779, n73780, n73781, n73782, n73783,
n73784, n73785, n73786, n73787, n73788, n73789, n73790, n73791,
n73792, n73793, n73794, n73795, n73796, n73797, n73798, n73799,
n73800, n73801, n73802, n73803, n73804, n73805, n73806, n73807,
n73808, n73809, n73810, n73811, n73812, n73813, n73814, n73815,
n73816, n73817, n73818, n73819, n73820, n73821, n73822, n73823,
n73824, n73825, n73826, n73827, n73828, n73829, n73830, n73831,
n73832, n73833, n73834, n73835, n73836, n73837, n73838, n73839,
n73840, n73841, n73842, n73843, n73844, n73845, n73846, n73847,
n73848, n73849, n73850, n73851, n73852, n73853, n73854, n73855,
n73856, n73857, n73858, n73859, n73860, n73861, n73862, n73863,
n73864, n73865, n73866, n73867, n73868, n73869, n73870, n73871,
n73872, n73873, n73874, n73875, n73876, n73877, n73878, n73879,
n73880, n73881, n73882, n73883, n73884, n73885, n73886, n73887,
n73888, n73889, n73890, n73891, n73892, n73893, n73894, n73895,
n73896, n73897, n73898, n73899, n73900, n73901, n73902, n73903,
n73904, n73905, n73906, n73907, n73908, n73909, n73910, n73911,
n73912, n73913, n73914, n73915, n73916, n73917, n73918, n73919,
n73920, n73921, n73922, n73923, n73924, n73925, n73926, n73927,
n73928, n73929, n73930, n73931, n73932, n73933, n73934, n73935,
n73936, n73937, n73938, n73939, n73940, n73941, n73942, n73943,
n73944, n73945, n73946, n73947, n73948, n73949, n73950, n73951,
n73952, n73953, n73954, n73955, n73956, n73957, n73958, n73959,
n73960, n73961, n73962, n73963, n73964, n73965, n73966, n73967,
n73968, n73969, n73970, n73971, n73972, n73973, n73974, n73975,
n73976, n73977, n73978, n73979, n73980, n73981, n73982, n73983,
n73984, n73985, n73986, n73987, n73988, n73989, n73990, n73991,
n73992, n73993, n73994, n73995, n73996, n73997, n73998, n73999,
n74000, n74001, n74002, n74003, n74004, n74005, n74006, n74007,
n74008, n74009, n74010, n74011, n74012, n74013, n74014, n74015,
n74016, n74017, n74018, n74019, n74020, n74021, n74022, n74023,
n74024, n74025, n74026, n74027, n74028, n74029, n74030, n74031,
n74032, n74033, n74034, n74035, n74036, n74037, n74038, n74039,
n74040, n74041, n74042, n74043, n74044, n74045, n74046, n74047,
n74048, n74049, n74050, n74051, n74052, n74053, n74054, n74055,
n74056, n74057, n74058, n74059, n74060, n74061, n74062, n74063,
n74064, n74065, n74066, n74067, n74068, n74069, n74070, n74071,
n74072, n74073, n74074, n74075, n74076, n74077, n74078, n74079,
n74080, n74081, n74082, n74083, n74084, n74085, n74086, n74087,
n74088, n74089, n74090, n74091, n74092, n74093, n74094, n74095,
n74096, n74097, n74098, n74099, n74100, n74101, n74102, n74103,
n74104, n74105, n74106, n74107, n74108, n74109, n74110, n74111,
n74112, n74113, n74114, n74115, n74116, n74117, n74118, n74119,
n74120, n74121, n74122, n74123, n74124, n74125, n74126, n74127,
n74128, n74129, n74130, n74131, n74132, n74133, n74134, n74135,
n74136, n74137, n74138, n74139, n74140, n74141, n74142, n74143,
n74144, n74145, n74146, n74147, n74148, n74149, n74150, n74151,
n74152, n74153, n74154, n74155, n74156, n74157, n74158, n74159,
n74160, n74161, n74162, n74163, n74164, n74165, n74166, n74167,
n74168, n74169, n74170, n74171, n74172, n74173, n74174, n74175,
n74176, n74177, n74178, n74179, n74180, n74181, n74182, n74183,
n74184, n74185, n74186, n74187, n74188, n74189, n74190, n74191,
n74192, n74193, n74194, n74195, n74196, n74197, n74198, n74199,
n74200, n74201, n74202, n74203, n74204, n74205, n74206, n74207,
n74208, n74209, n74210, n74211, n74212, n74213, n74214, n74215,
n74216, n74217, n74218, n74219, n74220, n74221, n74222, n74223,
n74224, n74225, n74226, n74227, n74228, n74229, n74230, n74231,
n74232, n74233, n74234, n74235, n74236, n74237, n74238, n74239,
n74240, n74241, n74242, n74243, n74244, n74245, n74246, n74247,
n74248, n74249, n74250, n74251, n74252, n74253, n74254, n74255,
n74256, n74257, n74258, n74259, n74260, n74261, n74262, n74263,
n74264, n74265, n74266, n74267, n74268, n74269, n74270, n74271,
n74272, n74273, n74274, n74275, n74276, n74277, n74278, n74279,
n74280, n74281, n74282, n74283, n74284, n74285, n74286, n74287,
n74288, n74289, n74290, n74291, n74292, n74293, n74294, n74295,
n74296, n74297, n74298, n74299, n74300, n74301, n74302, n74303,
n74304, n74305, n74306, n74307, n74308, n74309, n74310, n74311,
n74312, n74313, n74314, n74315, n74316, n74317, n74318, n74319,
n74320, n74321, n74322, n74323, n74324, n74325, n74326, n74327,
n74328, n74329, n74330, n74331, n74332, n74333, n74334, n74335,
n74336, n74337, n74338, n74339, n74340, n74341, n74342, n74343,
n74344, n74345, n74346, n74347, n74348, n74349, n74350, n74351,
n74352, n74353, n74354, n74355, n74356, n74357, n74358, n74359,
n74360, n74361, n74362, n74363, n74364, n74365, n74366, n74367,
n74368, n74369, n74370, n74371, n74372, n74373, n74374, n74375,
n74376, n74377, n74378, n74379, n74380, n74381, n74382, n74383,
n74384, n74385, n74386, n74387, n74388, n74389, n74390, n74391,
n74392, n74393, n74394, n74395, n74396, n74397, n74398, n74399,
n74400, n74401, n74402, n74403, n74404, n74405, n74406, n74407,
n74408, n74409, n74410, n74411, n74412, n74413, n74414, n74415,
n74416, n74417, n74418, n74419, n74420, n74421, n74422, n74423,
n74424, n74425, n74426, n74427, n74428, n74429, n74430, n74431,
n74432, n74433, n74434, n74435, n74436, n74437, n74438, n74439,
n74440, n74441, n74442, n74443, n74444, n74445, n74446, n74447,
n74448, n74449, n74450, n74451, n74452, n74453, n74454, n74455,
n74456, n74457, n74458, n74459, n74460, n74461, n74462, n74463,
n74464, n74465, n74466, n74467, n74468, n74469, n74470, n74471,
n74472, n74473, n74474, n74475, n74476, n74477, n74478, n74479,
n74480, n74481, n74482, n74483, n74484, n74485, n74486, n74487,
n74488, n74489, n74490, n74491, n74492, n74493, n74494, n74495,
n74496, n74497, n74498, n74499, n74500, n74501, n74502, n74503,
n74504, n74505, n74506, n74507, n74508, n74509, n74510, n74511,
n74512, n74513, n74514, n74515, n74516, n74517, n74518, n74519,
n74520, n74521, n74522, n74523, n74524, n74525, n74526, n74527,
n74528, n74529, n74530, n74531, n74532, n74533, n74534, n74535,
n74536, n74537, n74538, n74539, n74540, n74541, n74542, n74543,
n74544, n74545, n74546, n74547, n74548, n74549, n74550, n74551,
n74552, n74553, n74554, n74555, n74556, n74557, n74558, n74559,
n74560, n74561, n74562, n74563, n74564, n74565, n74566, n74567,
n74568, n74569, n74570, n74571, n74572, n74573, n74574, n74575,
n74576, n74577, n74578, n74579, n74580, n74581, n74582, n74583,
n74584, n74585, n74586, n74587, n74588, n74589, n74590, n74591,
n74592, n74593, n74594, n74595, n74596, n74597, n74598, n74599,
n74600, n74601, n74602, n74603, n74604, n74605, n74606, n74607,
n74608, n74609, n74610, n74611, n74612, n74613, n74614, n74615,
n74616, n74617, n74618, n74619, n74620, n74621, n74622, n74623,
n74624, n74625, n74626, n74627, n74628, n74629, n74630, n74631,
n74632, n74633, n74634, n74635, n74636, n74637, n74638, n74639,
n74640, n74641, n74642, n74643, n74644, n74645, n74646, n74647,
n74648, n74649, n74650, n74651, n74652, n74653, n74654, n74655,
n74656, n74657, n74658, n74659, n74660, n74661, n74662, n74663,
n74664, n74665, n74666, n74667, n74668, n74669, n74670, n74671,
n74672, n74673, n74674, n74675, n74676, n74677, n74678, n74679,
n74680, n74681, n74682, n74683, n74684, n74685, n74686, n74687,
n74688, n74689, n74690, n74691, n74692, n74693, n74694, n74695,
n74696, n74697, n74698, n74699, n74700, n74701, n74702, n74703,
n74704, n74705, n74706, n74707, n74708, n74709, n74710, n74711,
n74712, n74713, n74714, n74715, n74716, n74717, n74718, n74719,
n74720, n74721, n74722, n74723, n74724, n74725, n74726, n74727,
n74728, n74729, n74730, n74731, n74732, n74733, n74734, n74735,
n74736, n74737, n74738, n74739, n74740, n74741, n74742, n74743,
n74744, n74745, n74746, n74747, n74748, n74749, n74750, n74751,
n74752, n74753, n74754, n74755, n74756, n74757, n74758, n74759,
n74760, n74761, n74762, n74763, n74764, n74765, n74766, n74767,
n74768, n74769, n74770, n74771, n74772, n74773, n74774, n74775,
n74776, n74777, n74778, n74779, n74780, n74781, n74782, n74783,
n74784, n74785, n74786, n74787, n74788, n74789, n74790, n74791,
n74792, n74793, n74794, n74795, n74796, n74797, n74798, n74799,
n74800, n74801, n74802, n74803, n74804, n74805, n74806, n74807,
n74808, n74809, n74810, n74811, n74812, n74813, n74814, n74815,
n74816, n74817, n74818, n74819, n74820, n74821, n74822, n74823,
n74824, n74825, n74826, n74827, n74828, n74829, n74830, n74831,
n74832, n74833, n74834, n74835, n74836, n74837, n74838, n74839,
n74840, n74841, n74842, n74843, n74844, n74845, n74846, n74847,
n74848, n74849, n74850, n74851, n74852, n74853, n74854, n74855,
n74856, n74857, n74858, n74859, n74860, n74861, n74862, n74863,
n74864, n74865, n74866, n74867, n74868, n74869, n74870, n74871,
n74872, n74873, n74874, n74875, n74876, n74877, n74878, n74879,
n74880, n74881, n74882, n74883, n74884, n74885, n74886, n74887,
n74888, n74889, n74890, n74891, n74892, n74893, n74894, n74895,
n74896, n74897, n74898, n74899, n74900, n74901, n74902, n74903,
n74904, n74905, n74906, n74907, n74908, n74909, n74910, n74911,
n74912, n74913, n74914, n74915, n74916, n74917, n74918, n74919,
n74920, n74921, n74922, n74923, n74924, n74925, n74926, n74927,
n74928, n74929, n74930, n74931, n74932, n74933, n74934, n74935,
n74936, n74937, n74938, n74939, n74940, n74941, n74942, n74943,
n74944, n74945, n74946, n74947, n74948, n74949, n74950, n74951,
n74952, n74953, n74954, n74955, n74956, n74957, n74958, n74959,
n74960, n74961, n74962, n74963, n74964, n74965, n74966, n74967,
n74968, n74969, n74970, n74971, n74972, n74973, n74974, n74975,
n74976, n74977, n74978, n74979, n74980, n74981, n74982, n74983,
n74984, n74985, n74986, n74987, n74988, n74989, n74990, n74991,
n74992, n74993, n74994, n74995, n74996, n74997, n74998, n74999,
n75000, n75001, n75002, n75003, n75004, n75005, n75006, n75007,
n75008, n75009, n75010, n75011, n75012, n75013, n75014, n75015,
n75016, n75017, n75018, n75019, n75020, n75021, n75022, n75023,
n75024, n75025, n75026, n75027, n75028, n75029, n75030, n75031,
n75032, n75033, n75034, n75035, n75036, n75037, n75038, n75039,
n75040, n75041, n75042, n75043, n75044, n75045, n75046, n75047,
n75048, n75049, n75050, n75051, n75052, n75053, n75054, n75055,
n75056, n75057, n75058, n75059, n75060, n75061, n75062, n75063,
n75064, n75065, n75066, n75067, n75068, n75069, n75070, n75071,
n75072, n75073, n75074, n75075, n75076, n75077, n75078, n75079,
n75080, n75081, n75082, n75083, n75084, n75085, n75086, n75087,
n75088, n75089, n75090, n75091, n75092, n75093, n75094, n75095,
n75096, n75097, n75098, n75099, n75100, n75101, n75102, n75103,
n75104, n75105, n75106, n75107, n75108, n75109, n75110, n75111,
n75112, n75113, n75114, n75115, n75116, n75117, n75118, n75119,
n75120, n75121, n75122, n75123, n75124, n75125, n75126, n75127,
n75128, n75129, n75130, n75131, n75132, n75133, n75134, n75135,
n75136, n75137, n75138, n75139, n75140, n75141, n75142, n75143,
n75144, n75145, n75146, n75147, n75148, n75149, n75150, n75151,
n75152, n75153, n75154, n75155, n75156, n75157, n75158, n75159,
n75160, n75161, n75162, n75163, n75164, n75165, n75166, n75167,
n75168, n75169, n75170, n75171, n75172, n75173, n75174, n75175,
n75176, n75177, n75178, n75179, n75180, n75181, n75182, n75183,
n75184, n75185, n75186, n75187, n75188, n75189, n75190, n75191,
n75192, n75193, n75194, n75195, n75196, n75197, n75198, n75199,
n75200, n75201, n75202, n75203, n75204, n75205, n75206, n75207,
n75208, n75209, n75210, n75211, n75212, n75213, n75214, n75215,
n75216, n75217, n75218, n75219, n75220, n75221, n75222, n75223,
n75224, n75225, n75226, n75227, n75228, n75229, n75230, n75231,
n75232, n75233, n75234, n75235, n75236, n75237, n75238, n75239,
n75240, n75241, n75242, n75243, n75244, n75245, n75246, n75247,
n75248, n75249, n75250, n75251, n75252, n75253, n75254, n75255,
n75256, n75257, n75258, n75259, n75260, n75261, n75262, n75263,
n75264, n75265, n75266, n75267, n75268, n75269, n75270, n75271,
n75272, n75273, n75274, n75275, n75276, n75277, n75278, n75279,
n75280, n75281, n75282, n75283, n75284, n75285, n75286, n75287,
n75288, n75289, n75290, n75291, n75292, n75293, n75294, n75295,
n75296, n75297, n75298, n75299, n75300, n75301, n75302, n75303,
n75304, n75305, n75306, n75307, n75308, n75309, n75310, n75311,
n75312, n75313, n75314, n75315, n75316, n75317, n75318, n75319,
n75320, n75321, n75322, n75323, n75324, n75325, n75326, n75327,
n75328, n75329, n75330, n75331, n75332, n75333, n75334, n75335,
n75336, n75337, n75338, n75339, n75340, n75341, n75342, n75343,
n75344, n75345, n75346, n75347, n75348, n75349, n75350, n75351,
n75352, n75353, n75354, n75355, n75356, n75357, n75358, n75359,
n75360, n75361, n75362, n75363, n75364, n75365, n75366, n75367,
n75368, n75369, n75370, n75371, n75372, n75373, n75374, n75375,
n75376, n75377, n75378, n75379, n75380, n75381, n75382, n75383,
n75384, n75385, n75386, n75387, n75388, n75389, n75390, n75391,
n75392, n75393, n75394, n75395, n75396, n75397, n75398, n75399,
n75400, n75401, n75402, n75403, n75404, n75405, n75406, n75407,
n75408, n75409, n75410, n75411, n75412, n75413, n75414, n75415,
n75416, n75417, n75418, n75419, n75420, n75421, n75422, n75423,
n75424, n75425, n75426, n75427, n75428, n75429, n75430, n75431,
n75432, n75433, n75434, n75435, n75436, n75437, n75438, n75439,
n75440, n75441, n75442, n75443, n75444, n75445, n75446, n75447,
n75448, n75449, n75450, n75451, n75452, n75453, n75454, n75455,
n75456, n75457, n75458, n75459, n75460, n75461, n75462, n75463,
n75464, n75465, n75466, n75467, n75468, n75469, n75470, n75471,
n75472, n75473, n75474, n75475, n75476, n75477, n75478, n75479,
n75480, n75481, n75482, n75483, n75484, n75485, n75486, n75487,
n75488, n75489, n75490, n75491, n75492, n75493, n75494, n75495,
n75496, n75497, n75498, n75499, n75500, n75501, n75502, n75503,
n75504, n75505, n75506, n75507, n75508, n75509, n75510, n75511,
n75512, n75513, n75514, n75515, n75516, n75517, n75518, n75519,
n75520, n75521, n75522, n75523, n75524, n75525, n75526, n75527,
n75528, n75529, n75530, n75531, n75532, n75533, n75534, n75535,
n75536, n75537, n75538, n75539, n75540, n75541, n75542, n75543,
n75544, n75545, n75546, n75547, n75548, n75549, n75550, n75551,
n75552, n75553, n75554, n75555, n75556, n75557, n75558, n75559,
n75560, n75561, n75562, n75563, n75564, n75565, n75566, n75567,
n75568, n75569, n75570, n75571, n75572, n75573, n75574, n75575,
n75576, n75577, n75578, n75579, n75580, n75581, n75582, n75583,
n75584, n75585, n75586, n75587, n75588, n75589, n75590, n75591,
n75592, n75593, n75594, n75595, n75596, n75597, n75598, n75599,
n75600, n75601, n75602, n75603, n75604, n75605, n75606, n75607,
n75608, n75609, n75610, n75611, n75612, n75613, n75614, n75615,
n75616, n75617, n75618, n75619, n75620, n75621, n75622, n75623,
n75624, n75625, n75626, n75627, n75628, n75629, n75630, n75631,
n75632, n75633, n75634, n75635, n75636, n75637, n75638, n75639,
n75640, n75641, n75642, n75643, n75644, n75645, n75646, n75647,
n75648, n75649, n75650, n75651, n75652, n75653, n75654, n75655,
n75656, n75657, n75658, n75659, n75660, n75661, n75662, n75663,
n75664, n75665, n75666, n75667, n75668, n75669, n75670, n75671,
n75672, n75673, n75674, n75675, n75676, n75677, n75678, n75679,
n75680, n75681, n75682, n75683, n75684, n75685, n75686, n75687,
n75688, n75689, n75690, n75691, n75692, n75693, n75694, n75695,
n75696, n75697, n75698, n75699, n75700, n75701, n75702, n75703,
n75704, n75705, n75706, n75707, n75708, n75709, n75710, n75711,
n75712, n75713, n75714, n75715, n75716, n75717, n75718, n75719,
n75720, n75721, n75722, n75723, n75724, n75725, n75726, n75727,
n75728, n75729, n75730, n75731, n75732, n75733, n75734, n75735,
n75736, n75737, n75738, n75739, n75740, n75741, n75742, n75743,
n75744, n75745, n75746, n75747, n75748, n75749, n75750, n75751,
n75752, n75753, n75754, n75755, n75756, n75757, n75758, n75759,
n75760, n75761, n75762, n75763, n75764, n75765, n75766, n75767,
n75768, n75769, n75770, n75771, n75772, n75773, n75774, n75775,
n75776, n75777, n75778, n75779, n75780, n75781, n75782, n75783,
n75784, n75785, n75786, n75787, n75788, n75789, n75790, n75791,
n75792, n75793, n75794, n75795, n75796, n75797, n75798, n75799,
n75800, n75801, n75802, n75803, n75804, n75805, n75806, n75807,
n75808, n75809, n75810, n75811, n75812, n75813, n75814, n75815,
n75816, n75817, n75818, n75819, n75820, n75821, n75822, n75823,
n75824, n75825, n75826, n75827, n75828, n75829, n75830, n75831,
n75832, n75833, n75834, n75835, n75836, n75837, n75838, n75839,
n75840, n75841, n75842, n75843, n75844, n75845, n75846, n75847,
n75848, n75849, n75850, n75851, n75852, n75853, n75854, n75855,
n75856, n75857, n75858, n75859, n75860, n75861, n75862, n75863,
n75864, n75865, n75866, n75867, n75868, n75869, n75870, n75871,
n75872, n75873, n75874, n75875, n75876, n75877, n75878, n75879,
n75880, n75881, n75882, n75883, n75884, n75885, n75886, n75887,
n75888, n75889, n75890, n75891, n75892, n75893, n75894, n75895,
n75896, n75897, n75898, n75899, n75900, n75901, n75902, n75903,
n75904, n75905, n75906, n75907, n75908, n75909, n75910, n75911,
n75912, n75913, n75914, n75915, n75916, n75917, n75918, n75919,
n75920, n75921, n75922, n75923, n75924, n75925, n75926, n75927,
n75928, n75929, n75930, n75931, n75932, n75933, n75934, n75935,
n75936, n75937, n75938, n75939, n75940, n75941, n75942, n75943,
n75944, n75945, n75946, n75947, n75948, n75949, n75950, n75951,
n75952, n75953, n75954, n75955, n75956, n75957, n75958, n75959,
n75960, n75961, n75962, n75963, n75964, n75965, n75966, n75967,
n75968, n75969, n75970, n75971, n75972, n75973, n75974, n75975,
n75976, n75977, n75978, n75979, n75980, n75981, n75982, n75983,
n75984, n75985, n75986, n75987, n75988, n75989, n75990, n75991,
n75992, n75993, n75994, n75995, n75996, n75997, n75998, n75999,
n76000, n76001, n76002, n76003, n76004, n76005, n76006, n76007,
n76008, n76009, n76010, n76011, n76012, n76013, n76014, n76015,
n76016, n76017, n76018, n76019, n76020, n76021, n76022, n76023,
n76024, n76025, n76026, n76027, n76028, n76029, n76030, n76031,
n76032, n76033, n76034, n76035, n76036, n76037, n76038, n76039,
n76040, n76041, n76042, n76043, n76044, n76045, n76046, n76047,
n76048, n76049, n76050, n76051, n76052, n76053, n76054, n76055,
n76056, n76057, n76058, n76059, n76060, n76061, n76062, n76063,
n76064, n76065, n76066, n76067, n76068, n76069, n76070, n76071,
n76072, n76073, n76074, n76075, n76076, n76077, n76078, n76079,
n76080, n76081, n76082, n76083, n76084, n76085, n76086, n76087,
n76088, n76089, n76090, n76091, n76092, n76093, n76094, n76095,
n76096, n76097, n76098, n76099, n76100, n76101, n76102, n76103,
n76104, n76105, n76106, n76107, n76108, n76109, n76110, n76111,
n76112, n76113, n76114, n76115, n76116, n76117, n76118, n76119,
n76120, n76121, n76122, n76123, n76124, n76125, n76126, n76127,
n76128, n76129, n76130, n76131, n76132, n76133, n76134, n76135,
n76136, n76137, n76138, n76139, n76140, n76141, n76142, n76143,
n76144, n76145, n76146, n76147, n76148, n76149, n76150, n76151,
n76152, n76153, n76154, n76155, n76156, n76157, n76158, n76159,
n76160, n76161, n76162, n76163, n76164, n76165, n76166, n76167,
n76168, n76169, n76170, n76171, n76172, n76173, n76174, n76175,
n76176, n76177, n76178, n76179, n76180, n76181, n76182, n76183,
n76184, n76185, n76186, n76187, n76188, n76189, n76190, n76191,
n76192, n76193, n76194, n76195, n76196, n76197, n76198, n76199,
n76200, n76201, n76202, n76203, n76204, n76205, n76206, n76207,
n76208, n76209, n76210, n76211, n76212, n76213, n76214, n76215,
n76216, n76217, n76218, n76219, n76220, n76221, n76222, n76223,
n76224, n76225, n76226, n76227, n76228, n76229, n76230, n76231,
n76232, n76233, n76234, n76235, n76236, n76237, n76238, n76239,
n76240, n76241, n76242, n76243, n76244, n76245, n76246, n76247,
n76248, n76249, n76250, n76251, n76252, n76253, n76254, n76255,
n76256, n76257, n76258, n76259, n76260, n76261, n76262, n76263,
n76264, n76265, n76266, n76267, n76268, n76269, n76270, n76271,
n76272, n76273, n76274, n76275, n76276, n76277, n76278, n76279,
n76280, n76281, n76282, n76283, n76284, n76285, n76286, n76287,
n76288, n76289, n76290, n76291, n76292, n76293, n76294, n76295,
n76296, n76297, n76298, n76299, n76300, n76301, n76302, n76303,
n76304, n76305, n76306, n76307, n76308, n76309, n76310, n76311,
n76312, n76313, n76314, n76315, n76316, n76317, n76318, n76319,
n76320, n76321, n76322, n76323, n76324, n76325, n76326, n76327,
n76328, n76329, n76330, n76331, n76332, n76333, n76334, n76335,
n76336, n76337, n76338, n76339, n76340, n76341, n76342, n76343,
n76344, n76345, n76346, n76347, n76348, n76349, n76350, n76351,
n76352, n76353, n76354, n76355, n76356, n76357, n76358, n76359,
n76360, n76361, n76362, n76363, n76364, n76365, n76366, n76367,
n76368, n76369, n76370, n76371, n76372, n76373, n76374, n76375,
n76376, n76377, n76378, n76379, n76380, n76381, n76382, n76383,
n76384, n76385, n76386, n76387, n76388, n76389, n76390, n76391,
n76392, n76393, n76394, n76395, n76396, n76397, n76398, n76399,
n76400, n76401, n76402, n76403, n76404, n76405, n76406, n76407,
n76408, n76409, n76410, n76411, n76412, n76413, n76414, n76415,
n76416, n76417, n76418, n76419, n76420, n76421, n76422, n76423,
n76424, n76425, n76426, n76427, n76428, n76429, n76430, n76431,
n76432, n76433, n76434, n76435, n76436, n76437, n76438, n76439,
n76440, n76441, n76442, n76443, n76444, n76445, n76446, n76447,
n76448, n76449, n76450, n76451, n76452, n76453, n76454, n76455,
n76456, n76457, n76458, n76459, n76460, n76461, n76462, n76463,
n76464, n76465, n76466, n76467, n76468, n76469, n76470, n76471,
n76472, n76473, n76474, n76475, n76476, n76477, n76478, n76479,
n76480, n76481, n76482, n76483, n76484, n76485, n76486, n76487,
n76488, n76489, n76490, n76491, n76492, n76493, n76494, n76495,
n76496, n76497, n76498, n76499, n76500, n76501, n76502, n76503,
n76504, n76505, n76506, n76507, n76508, n76509, n76510, n76511,
n76512, n76513, n76514, n76515, n76516, n76517, n76518, n76519,
n76520, n76521, n76522, n76523, n76524, n76525, n76526, n76527,
n76528, n76529, n76530, n76531, n76532, n76533, n76534, n76535,
n76536, n76537, n76538, n76539, n76540, n76541, n76542, n76543,
n76544, n76545, n76546, n76547, n76548, n76549, n76550, n76551,
n76552, n76553, n76554, n76555, n76556, n76557, n76558, n76559,
n76560, n76561, n76562, n76563, n76564, n76565, n76566, n76567,
n76568, n76569, n76570, n76571, n76572, n76573, n76574, n76575,
n76576, n76577, n76578, n76579, n76580, n76581, n76582, n76583,
n76584, n76585, n76586, n76587, n76588, n76589, n76590, n76591,
n76592, n76593, n76594, n76595, n76596, n76597, n76598, n76599,
n76600, n76601, n76602, n76603, n76604, n76605, n76606, n76607,
n76608, n76609, n76610, n76611, n76612, n76613, n76614, n76615,
n76616, n76617, n76618, n76619, n76620, n76621, n76622, n76623,
n76624, n76625, n76626, n76627, n76628, n76629, n76630, n76631,
n76632, n76633, n76634, n76635, n76636, n76637, n76638, n76639,
n76640, n76641, n76642, n76643, n76644, n76645, n76646, n76647,
n76648, n76649, n76650, n76651, n76652, n76653, n76654, n76655,
n76656, n76657, n76658, n76659, n76660, n76661, n76662, n76663,
n76664, n76665, n76666, n76667, n76668, n76669, n76670, n76671,
n76672, n76673, n76674, n76675, n76676, n76677, n76678, n76679,
n76680, n76681, n76682, n76683, n76684, n76685, n76686, n76687,
n76688, n76689, n76690, n76691, n76692, n76693, n76694, n76695,
n76696, n76697, n76698, n76699, n76700, n76701, n76702, n76703,
n76704, n76705, n76706, n76707, n76708, n76709, n76710, n76711,
n76712, n76713, n76714, n76715, n76716, n76717, n76718, n76719,
n76720, n76721, n76722, n76723, n76724, n76725, n76726, n76727,
n76728, n76729, n76730, n76731, n76732, n76733, n76734, n76735,
n76736, n76737, n76738, n76739, n76740, n76741, n76742, n76743,
n76744, n76745, n76746, n76747, n76748, n76749, n76750, n76751,
n76752, n76753, n76754, n76755, n76756, n76757, n76758, n76759,
n76760, n76761, n76762, n76763, n76764, n76765, n76766, n76767,
n76768, n76769, n76770, n76771, n76772, n76773, n76774, n76775,
n76776, n76777, n76778, n76779, n76780, n76781, n76782, n76783,
n76784, n76785, n76786, n76787, n76788, n76789, n76790, n76791,
n76792, n76793, n76794, n76795, n76796, n76797, n76798, n76799,
n76800, n76801, n76802, n76803, n76804, n76805, n76806, n76807,
n76808, n76809, n76810, n76811, n76812, n76813, n76814, n76815,
n76816, n76817, n76818, n76819, n76820, n76821, n76822, n76823,
n76824, n76825, n76826, n76827, n76828, n76829, n76830, n76831,
n76832, n76833, n76834, n76835, n76836, n76837, n76838, n76839,
n76840, n76841, n76842, n76843, n76844, n76845, n76846, n76847,
n76848, n76849, n76850, n76851, n76852, n76853, n76854, n76855,
n76856, n76857, n76858, n76859, n76860, n76861, n76862, n76863,
n76864, n76865, n76866, n76867, n76868, n76869, n76870, n76871,
n76872, n76873, n76874, n76875, n76876, n76877, n76878, n76879,
n76880, n76881, n76882, n76883, n76884, n76885, n76886, n76887,
n76888, n76889, n76890, n76891, n76892, n76893, n76894, n76895,
n76896, n76897, n76898, n76899, n76900, n76901, n76902, n76903,
n76904, n76905, n76906, n76907, n76908, n76909, n76910, n76911,
n76912, n76913, n76914, n76915, n76916, n76917, n76918, n76919,
n76920, n76921, n76922, n76923, n76924, n76925, n76926, n76927,
n76928, n76929, n76930;

dff P3_STATE_REG_reg ( clk, reset, P3_STATE_REG, n76042 );
not U_inv0 ( n72968, P3_STATE_REG );
dff P4_STATE_REG_reg ( clk, reset, P4_STATE_REG, n76922 );
not U_inv1 ( n72969, P4_STATE_REG );
dff P2_P1_MEMORYFETCH_REG_reg ( clk, reset, P2_P1_MEMORYFETCH_REG, n16716 );
dff P2_P1_M_IO_N_REG_reg ( clk, reset, P2_P1_M_IO_N_REG, n16696 );
dff P2_READY11_REG_reg ( clk, reset, P2_READY11_REG, n796 );
dff P2_BUF1_REG_0__reg ( clk, reset, P2_BUF1_REG_0_, n461 );
not U_inv2 ( n75455, P2_BUF1_REG_0_ );
dff P2_P2_INSTQUEUE_REG_15__0__reg ( clk, reset, ex_wire0, n12631 );
not U_inv3 ( n73660, ex_wire0 );
dff P2_P2_PHYADDRPOINTER_REG_27__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_27_, n13581 );
not U_inv4 ( n74851, P2_P2_PHYADDRPOINTER_REG_27_ );
dff P2_P2_PHYADDRPOINTER_REG_28__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_28_, n13586 );
not U_inv5 ( n75245, P2_P2_PHYADDRPOINTER_REG_28_ );
dff P2_P2_REIP_REG_28__reg ( clk, reset, P2_P2_REIP_REG_28_, n14381 );
not U_inv6 ( n75300, P2_P2_REIP_REG_28_ );
dff P2_P2_REIP_REG_29__reg ( clk, reset, P2_P2_REIP_REG_29_, n14386 );
not U_inv7 ( n73316, P2_P2_REIP_REG_29_ );
dff P2_P2_REIP_REG_30__reg ( clk, reset, P2_P2_REIP_REG_30_, n14391 );
not U_inv8 ( n75063, P2_P2_REIP_REG_30_ );
dff P2_P2_ADDRESS_REG_29__reg ( clk, reset, P2_P2_ADDRESS_REG_29_, n12251 );
dff P2_P2_INSTQUEUE_REG_15__7__reg ( clk, reset, ex_wire1, n12596 );
not U_inv9 ( n74179, ex_wire1 );
dff P2_P2_STATE2_REG_3__reg ( clk, reset, P2_P2_STATE2_REG_3_, n12576 );
dff P2_P2_INSTQUEUE_REG_15__6__reg ( clk, reset, ex_wire2, n12601 );
not U_inv10 ( n74057, ex_wire2 );
dff P2_P2_FLUSH_REG_reg ( clk, reset, P2_P2_FLUSH_REG, n14426 );
not U_inv11 ( n75234, P2_P2_FLUSH_REG );
dff P2_P2_INSTQUEUERD_ADDR_REG_4__reg ( clk, reset, P2_P2_INSTQUEUERD_ADDR_REG_4_, n13236 );
not U_inv12 ( n74614, P2_P2_INSTQUEUERD_ADDR_REG_4_ );
dff P2_P2_INSTADDRPOINTER_REG_31__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_31_, n13441 );
not U_inv13 ( n75067, P2_P2_INSTADDRPOINTER_REG_31_ );
dff P2_P2_EAX_REG_16__reg ( clk, reset, P2_P2_EAX_REG_16_, n14001 );
not U_inv14 ( n75380, P2_P2_EAX_REG_16_ );
dff P2_P2_EAX_REG_17__reg ( clk, reset, P2_P2_EAX_REG_17_, n14006 );
not U_inv15 ( n74819, P2_P2_EAX_REG_17_ );
dff P2_P2_UWORD_REG_1__reg ( clk, reset, P2_P2_UWORD_REG_1_, n13751 );
not U_inv16 ( n75479, P2_P2_UWORD_REG_1_ );
dff P2_P2_DATAO_REG_17__reg ( clk, reset, P2_P2_DATAO_REG_17_, n13846 );
not U_inv17 ( n75518, P2_P2_DATAO_REG_17_ );
dff P2_BUF2_REG_17__reg ( clk, reset, P2_BUF2_REG_17_, n706 );
not U_inv18 ( n75360, P2_BUF2_REG_17_ );
dff P2_P3_INSTQUEUE_REG_15__1__reg ( clk, reset, ex_wire3, n10381 );
not U_inv19 ( n73628, ex_wire3 );
dff P2_P3_PHYADDRPOINTER_REG_27__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_27_, n11336 );
not U_inv20 ( n74848, P2_P3_PHYADDRPOINTER_REG_27_ );
dff P2_P3_PHYADDRPOINTER_REG_28__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_28_, n11341 );
not U_inv21 ( n75244, P2_P3_PHYADDRPOINTER_REG_28_ );
dff P2_P3_REIP_REG_28__reg ( clk, reset, P2_P3_REIP_REG_28_, n12136 );
not U_inv22 ( n75361, P2_P3_REIP_REG_28_ );
dff P2_P3_REIP_REG_29__reg ( clk, reset, P2_P3_REIP_REG_29_, n12141 );
not U_inv23 ( n73319, P2_P3_REIP_REG_29_ );
dff P2_P3_REIP_REG_30__reg ( clk, reset, P2_P3_REIP_REG_30_, n12146 );
not U_inv24 ( n75070, P2_P3_REIP_REG_30_ );
dff P2_P3_PHYADDRPOINTER_REG_30__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_30_, n11351 );
not U_inv25 ( n75188, P2_P3_PHYADDRPOINTER_REG_30_ );
dff P2_P3_PHYADDRPOINTER_REG_31__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_31_, n11356 );
dff P2_P3_REIP_REG_0__reg ( clk, reset, P2_P3_REIP_REG_0_, n11996 );
not U_inv26 ( n75257, P2_P3_REIP_REG_0_ );
dff P2_P3_BYTEENABLE_REG_3__reg ( clk, reset, P2_P3_BYTEENABLE_REG_3_, n12156 );
dff P2_P3_BE_N_REG_3__reg ( clk, reset, P2_P3_BE_N_REG_3_, n9986 );
dff P2_READY22_REG_reg ( clk, reset, P2_READY22_REG, n791 );
dff P2_P3_STATE_REG_2__reg ( clk, reset, P2_P3_STATE_REG_2_, n10156 );
not U_inv27 ( n72927, P2_P3_STATE_REG_2_ );
dff P2_P3_STATE_REG_0__reg ( clk, reset, P2_P3_STATE_REG_0_, n10166 );
not U_inv28 ( n73186, P2_P3_STATE_REG_0_ );
dff P2_P3_STATE_REG_1__reg ( clk, reset, P2_P3_STATE_REG_1_, n10161 );
not U_inv29 ( n74657, P2_P3_STATE_REG_1_ );
dff P2_P3_ADS_N_REG_reg ( clk, reset, P2_P3_ADS_N_REG, n12216 );
not U_inv30 ( n75969, P2_P3_ADS_N_REG );
dff P2_P3_DATAWIDTH_REG_0__reg ( clk, reset, P2_P3_DATAWIDTH_REG_0_, n10171 );
dff P2_P3_STATEBS16_REG_reg ( clk, reset, P2_P3_STATEBS16_REG, n12191 );
not U_inv31 ( n74889, P2_P3_STATEBS16_REG );
dff P2_P3_INSTQUEUE_REG_15__7__reg ( clk, reset, ex_wire4, n10351 );
not U_inv32 ( n74177, ex_wire4 );
dff P2_P3_STATE2_REG_3__reg ( clk, reset, P2_P3_STATE2_REG_3_, n10331 );
dff P2_P3_INSTQUEUERD_ADDR_REG_4__reg ( clk, reset, P2_P3_INSTQUEUERD_ADDR_REG_4_, n10991 );
not U_inv33 ( n74613, P2_P3_INSTQUEUERD_ADDR_REG_4_ );
dff P2_P3_FLUSH_REG_reg ( clk, reset, P2_P3_FLUSH_REG, n12181 );
not U_inv34 ( n75233, P2_P3_FLUSH_REG );
dff P2_P3_INSTQUEUEWR_ADDR_REG_4__reg ( clk, reset, P2_P3_INSTQUEUEWR_ADDR_REG_4_, n11016 );
not U_inv35 ( n75034, P2_P3_INSTQUEUEWR_ADDR_REG_4_ );
dff P2_P3_INSTADDRPOINTER_REG_31__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_31_, n11196 );
not U_inv36 ( n75068, P2_P3_INSTADDRPOINTER_REG_31_ );
dff P2_P3_DATAO_REG_31__reg ( clk, reset, P2_P3_DATAO_REG_31_, n11671 );
not U_inv37 ( n73429, P2_P3_DATAO_REG_31_ );
dff P2_P3_INSTQUEUEWR_ADDR_REG_1__reg ( clk, reset, P2_P3_INSTQUEUEWR_ADDR_REG_1_, n11031 );
not U_inv38 ( n74562, P2_P3_INSTQUEUEWR_ADDR_REG_1_ );
dff P2_P3_INSTQUEUEWR_ADDR_REG_3__reg ( clk, reset, P2_P3_INSTQUEUEWR_ADDR_REG_3_, n11021 );
not U_inv39 ( n73139, P2_P3_INSTQUEUEWR_ADDR_REG_3_ );
dff P2_P3_EAX_REG_0__reg ( clk, reset, P2_P3_EAX_REG_0_, n11676 );
not U_inv40 ( n74487, P2_P3_EAX_REG_0_ );
dff P2_P3_EAX_REG_1__reg ( clk, reset, P2_P3_EAX_REG_1_, n11681 );
not U_inv41 ( n73127, P2_P3_EAX_REG_1_ );
dff P2_P3_EAX_REG_2__reg ( clk, reset, P2_P3_EAX_REG_2_, n11686 );
not U_inv42 ( n75284, P2_P3_EAX_REG_2_ );
dff P2_P3_EAX_REG_3__reg ( clk, reset, P2_P3_EAX_REG_3_, n11691 );
not U_inv43 ( n74507, P2_P3_EAX_REG_3_ );
dff P2_P3_EAX_REG_4__reg ( clk, reset, P2_P3_EAX_REG_4_, n11696 );
not U_inv44 ( n75272, P2_P3_EAX_REG_4_ );
dff P2_P3_EAX_REG_5__reg ( clk, reset, P2_P3_EAX_REG_5_, n11701 );
not U_inv45 ( n74539, P2_P3_EAX_REG_5_ );
dff P2_P3_EAX_REG_6__reg ( clk, reset, P2_P3_EAX_REG_6_, n11706 );
not U_inv46 ( n75270, P2_P3_EAX_REG_6_ );
dff P2_P3_EAX_REG_7__reg ( clk, reset, P2_P3_EAX_REG_7_, n11711 );
not U_inv47 ( n74581, P2_P3_EAX_REG_7_ );
dff P2_P3_EAX_REG_8__reg ( clk, reset, P2_P3_EAX_REG_8_, n11716 );
not U_inv48 ( n75271, P2_P3_EAX_REG_8_ );
dff P2_P3_EAX_REG_9__reg ( clk, reset, P2_P3_EAX_REG_9_, n11721 );
not U_inv49 ( n75250, P2_P3_EAX_REG_9_ );
dff P2_P3_EAX_REG_10__reg ( clk, reset, ex_wire5, n11726 );
not U_inv50 ( n74628, ex_wire5 );
dff P2_P3_LWORD_REG_10__reg ( clk, reset, P2_P3_LWORD_REG_10_, n11386 );
not U_inv51 ( n75635, P2_P3_LWORD_REG_10_ );
dff P2_P3_DATAO_REG_10__reg ( clk, reset, P2_P3_DATAO_REG_10_, n11566 );
dff P4_IR_REG_10__reg ( clk, reset, P4_IR_REG_10_, n2076 );
not U_inv52 ( n75410, P4_IR_REG_10_ );
dff P4_REG0_REG_11__reg ( clk, reset, P4_REG0_REG_11_, n2401 );
dff P4_REG0_REG_10__reg ( clk, reset, P4_REG0_REG_10_, n2396 );
dff P4_REG0_REG_12__reg ( clk, reset, P4_REG0_REG_12_, n2406 );
dff P4_B_REG_reg ( clk, reset, P4_B_REG, n3086 );
not U_inv53 ( n74634, P4_B_REG );
dff P4_REG0_REG_29__reg ( clk, reset, P4_REG0_REG_29_, n2491 );
dff P4_REG2_REG_28__reg ( clk, reset, ex_wire6, n2806 );
not U_inv54 ( n74777, ex_wire6 );
dff P4_REG2_REG_27__reg ( clk, reset, ex_wire7, n2801 );
not U_inv55 ( n74775, ex_wire7 );
dff P4_REG0_REG_26__reg ( clk, reset, P4_REG0_REG_26_, n2476 );
dff P4_REG2_REG_25__reg ( clk, reset, ex_wire8, n2791 );
not U_inv56 ( n74703, ex_wire8 );
dff P4_REG0_REG_24__reg ( clk, reset, P4_REG0_REG_24_, n2466 );
dff P4_REG2_REG_23__reg ( clk, reset, ex_wire9, n2781 );
not U_inv57 ( n74598, ex_wire9 );
dff P4_REG2_REG_22__reg ( clk, reset, ex_wire10, n2776 );
not U_inv58 ( n74523, ex_wire10 );
dff P4_REG2_REG_21__reg ( clk, reset, ex_wire11, n2771 );
not U_inv59 ( n74544, ex_wire11 );
dff P4_REG0_REG_20__reg ( clk, reset, P4_REG0_REG_20_, n2446 );
dff P4_REG0_REG_19__reg ( clk, reset, P4_REG0_REG_19_, n2441 );
dff P4_REG0_REG_18__reg ( clk, reset, P4_REG0_REG_18_, n2436 );
dff P4_REG0_REG_17__reg ( clk, reset, P4_REG0_REG_17_, n2431 );
dff P4_REG0_REG_16__reg ( clk, reset, P4_REG0_REG_16_, n2426 );
dff P4_REG2_REG_15__reg ( clk, reset, P4_REG2_REG_15_, n2741 );
not U_inv60 ( n74421, P4_REG2_REG_15_ );
dff P4_REG2_REG_14__reg ( clk, reset, P4_REG2_REG_14_, n2736 );
not U_inv61 ( n74411, P4_REG2_REG_14_ );
dff P4_REG0_REG_13__reg ( clk, reset, P4_REG0_REG_13_, n2411 );
dff P1_P1_INSTQUEUE_REG_15__7__reg ( clk, reset, ex_wire12, n8106 );
not U_inv62 ( n74361, ex_wire12 );
dff P1_P1_STATE2_REG_3__reg ( clk, reset, P1_P1_STATE2_REG_3_, n8086 );
dff P1_P1_INSTQUEUE_REG_14__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__7_, n8146 );
not U_inv63 ( n74376, P1_P1_INSTQUEUE_REG_14__7_ );
dff P1_P1_FLUSH_REG_reg ( clk, reset, P1_P1_FLUSH_REG, n9936 );
not U_inv64 ( n75232, P1_P1_FLUSH_REG );
dff P1_P1_INSTQUEUERD_ADDR_REG_4__reg ( clk, reset, P1_P1_INSTQUEUERD_ADDR_REG_4_, n8746 );
not U_inv65 ( n74646, P1_P1_INSTQUEUERD_ADDR_REG_4_ );
dff P1_P1_INSTADDRPOINTER_REG_1__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_1_, n8801 );
not U_inv66 ( n75059, P1_P1_INSTADDRPOINTER_REG_1_ );
dff P1_P1_INSTADDRPOINTER_REG_3__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_3_, n8811 );
not U_inv67 ( n74429, P1_P1_INSTADDRPOINTER_REG_3_ );
dff P1_P1_PHYADDRPOINTER_REG_3__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_3_, n8971 );
not U_inv68 ( n73072, P1_P1_PHYADDRPOINTER_REG_3_ );
dff P1_P1_PHYADDRPOINTER_REG_4__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_4_, n8976 );
not U_inv69 ( n74484, P1_P1_PHYADDRPOINTER_REG_4_ );
dff P1_P1_PHYADDRPOINTER_REG_5__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_5_, n8981 );
not U_inv70 ( n73087, P1_P1_PHYADDRPOINTER_REG_5_ );
dff P1_P1_REIP_REG_5__reg ( clk, reset, P1_P1_REIP_REG_5_, n9776 );
not U_inv71 ( n74727, P1_P1_REIP_REG_5_ );
dff P1_P1_REIP_REG_6__reg ( clk, reset, ex_wire13, n9781 );
not U_inv72 ( n74729, ex_wire13 );
dff P1_P1_ADDRESS_REG_5__reg ( clk, reset, P1_P1_ADDRESS_REG_5_, n7881 );
not U_inv73 ( n73041, P1_P1_ADDRESS_REG_5_ );
dff P1_P1_LWORD_REG_7__reg ( clk, reset, P1_P1_LWORD_REG_7_, n9156 );
not U_inv74 ( n75683, P1_P1_LWORD_REG_7_ );
dff P1_P1_DATAO_REG_7__reg ( clk, reset, P1_P1_DATAO_REG_7_, n9306 );
dff P1_BUF1_REG_7__reg ( clk, reset, P1_BUF1_REG_7_, n156 );
not U_inv75 ( n75463, P1_BUF1_REG_7_ );
dff P1_P2_INSTQUEUE_REG_15__7__reg ( clk, reset, ex_wire14, n5861 );
not U_inv76 ( n74178, ex_wire14 );
dff P1_P2_STATE2_REG_3__reg ( clk, reset, P1_P2_STATE2_REG_3_, n5841 );
dff P1_P2_INSTQUEUE_REG_15__6__reg ( clk, reset, ex_wire15, n5866 );
not U_inv77 ( n74058, ex_wire15 );
dff P1_P2_FLUSH_REG_reg ( clk, reset, P1_P2_FLUSH_REG, n7691 );
not U_inv78 ( n75231, P1_P2_FLUSH_REG );
dff P1_P2_INSTQUEUERD_ADDR_REG_4__reg ( clk, reset, P1_P2_INSTQUEUERD_ADDR_REG_4_, n6501 );
not U_inv79 ( n74612, P1_P2_INSTQUEUERD_ADDR_REG_4_ );
dff P1_P2_INSTADDRPOINTER_REG_31__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_31_, n6706 );
not U_inv80 ( n75066, P1_P2_INSTADDRPOINTER_REG_31_ );
dff P1_P2_EAX_REG_16__reg ( clk, reset, P1_P2_EAX_REG_16_, n7266 );
not U_inv81 ( n75388, P1_P2_EAX_REG_16_ );
dff P1_P2_EAX_REG_17__reg ( clk, reset, P1_P2_EAX_REG_17_, n7271 );
not U_inv82 ( n74820, P1_P2_EAX_REG_17_ );
dff P1_P2_UWORD_REG_1__reg ( clk, reset, P1_P2_UWORD_REG_1_, n7016 );
not U_inv83 ( n75487, P1_P2_UWORD_REG_1_ );
dff P1_P2_DATAO_REG_17__reg ( clk, reset, P1_P2_DATAO_REG_17_, n7111 );
not U_inv84 ( n75546, P1_P2_DATAO_REG_17_ );
dff P1_BUF2_REG_17__reg ( clk, reset, P1_BUF2_REG_17_, n366 );
not U_inv85 ( n75347, P1_BUF2_REG_17_ );
dff P1_P3_INSTQUEUE_REG_15__1__reg ( clk, reset, ex_wire16, n3646 );
not U_inv86 ( n73969, ex_wire16 );
dff P1_P3_PHYADDRPOINTER_REG_27__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_27_, n4601 );
not U_inv87 ( n74849, P1_P3_PHYADDRPOINTER_REG_27_ );
dff P1_P3_PHYADDRPOINTER_REG_28__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_28_, n4606 );
not U_inv88 ( n75246, P1_P3_PHYADDRPOINTER_REG_28_ );
dff P1_P3_REIP_REG_28__reg ( clk, reset, P1_P3_REIP_REG_28_, n5401 );
not U_inv89 ( n75362, P1_P3_REIP_REG_28_ );
dff P1_P3_REIP_REG_29__reg ( clk, reset, P1_P3_REIP_REG_29_, n5406 );
not U_inv90 ( n73318, P1_P3_REIP_REG_29_ );
dff P1_P3_REIP_REG_30__reg ( clk, reset, P1_P3_REIP_REG_30_, n5411 );
not U_inv91 ( n75069, P1_P3_REIP_REG_30_ );
dff P1_P3_PHYADDRPOINTER_REG_30__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_30_, n4616 );
not U_inv92 ( n75185, P1_P3_PHYADDRPOINTER_REG_30_ );
dff P1_P3_PHYADDRPOINTER_REG_31__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_31_, n4621 );
dff P1_P3_REIP_REG_0__reg ( clk, reset, P1_P3_REIP_REG_0_, n5261 );
not U_inv93 ( n75258, P1_P3_REIP_REG_0_ );
dff P1_P3_BYTEENABLE_REG_3__reg ( clk, reset, P1_P3_BYTEENABLE_REG_3_, n5421 );
dff P1_P3_BE_N_REG_3__reg ( clk, reset, P1_P3_BE_N_REG_3_, n3251 );
dff P1_READY22_REG_reg ( clk, reset, P1_READY22_REG, n451 );
dff P1_P3_STATE_REG_2__reg ( clk, reset, P1_P3_STATE_REG_2_, n3421 );
not U_inv94 ( n72928, P1_P3_STATE_REG_2_ );
dff P1_P3_STATE_REG_1__reg ( clk, reset, P1_P3_STATE_REG_1_, n3426 );
not U_inv95 ( n74654, P1_P3_STATE_REG_1_ );
dff P1_P3_STATE_REG_0__reg ( clk, reset, P1_P3_STATE_REG_0_, n3431 );
not U_inv96 ( n73192, P1_P3_STATE_REG_0_ );
dff P1_P3_DATAWIDTH_REG_0__reg ( clk, reset, P1_P3_DATAWIDTH_REG_0_, n3436 );
dff P1_P3_DATAWIDTH_REG_31__reg ( clk, reset, ex_wire17, n3591 );
not U_inv97 ( n75135, ex_wire17 );
dff P1_P3_DATAWIDTH_REG_30__reg ( clk, reset, ex_wire18, n3586 );
not U_inv98 ( n73335, ex_wire18 );
dff P1_P3_DATAWIDTH_REG_29__reg ( clk, reset, ex_wire19, n3581 );
not U_inv99 ( n73323, ex_wire19 );
dff P1_P3_DATAWIDTH_REG_28__reg ( clk, reset, ex_wire20, n3576 );
not U_inv100 ( n75079, ex_wire20 );
dff P1_P3_DATAWIDTH_REG_27__reg ( clk, reset, ex_wire21, n3571 );
not U_inv101 ( n73349, ex_wire21 );
dff P1_P3_DATAWIDTH_REG_26__reg ( clk, reset, ex_wire22, n3566 );
not U_inv102 ( n75123, ex_wire22 );
dff P1_P3_DATAWIDTH_REG_25__reg ( clk, reset, ex_wire23, n3561 );
not U_inv103 ( n73331, ex_wire23 );
dff P1_P3_DATAWIDTH_REG_24__reg ( clk, reset, ex_wire24, n3556 );
not U_inv104 ( n75089, ex_wire24 );
dff P1_P3_DATAWIDTH_REG_23__reg ( clk, reset, ex_wire25, n3551 );
not U_inv105 ( n73377, ex_wire25 );
dff P1_P3_DATAWIDTH_REG_22__reg ( clk, reset, ex_wire26, n3546 );
not U_inv106 ( n75159, ex_wire26 );
dff P1_P3_DATAWIDTH_REG_21__reg ( clk, reset, ex_wire27, n3541 );
not U_inv107 ( n73355, ex_wire27 );
dff P1_P3_DATAWIDTH_REG_20__reg ( clk, reset, ex_wire28, n3536 );
not U_inv108 ( n75129, ex_wire28 );
dff P1_P3_DATAWIDTH_REG_19__reg ( clk, reset, ex_wire29, n3531 );
not U_inv109 ( n73383, ex_wire29 );
dff P1_P3_DATAWIDTH_REG_18__reg ( clk, reset, ex_wire30, n3526 );
not U_inv110 ( n75165, ex_wire30 );
dff P1_P3_DATAWIDTH_REG_17__reg ( clk, reset, ex_wire31, n3521 );
not U_inv111 ( n73367, ex_wire31 );
dff P1_P3_DATAWIDTH_REG_16__reg ( clk, reset, ex_wire32, n3516 );
not U_inv112 ( n75141, ex_wire32 );
dff P1_P3_DATAWIDTH_REG_15__reg ( clk, reset, ex_wire33, n3511 );
not U_inv113 ( n73347, ex_wire33 );
dff P1_P3_DATAWIDTH_REG_14__reg ( clk, reset, ex_wire34, n3506 );
not U_inv114 ( n75117, ex_wire34 );
dff P1_P3_DATAWIDTH_REG_13__reg ( clk, reset, ex_wire35, n3501 );
not U_inv115 ( n73330, ex_wire35 );
dff P1_P3_DATAWIDTH_REG_12__reg ( clk, reset, ex_wire36, n3496 );
not U_inv116 ( n75088, ex_wire36 );
dff P1_P3_DATAWIDTH_REG_11__reg ( clk, reset, ex_wire37, n3491 );
not U_inv117 ( n73333, ex_wire37 );
dff P1_P3_DATAWIDTH_REG_10__reg ( clk, reset, ex_wire38, n3486 );
not U_inv118 ( n75099, ex_wire38 );
dff P1_P3_DATAWIDTH_REG_9__reg ( clk, reset, ex_wire39, n3481 );
not U_inv119 ( n73369, ex_wire39 );
dff P1_P3_DATAWIDTH_REG_8__reg ( clk, reset, ex_wire40, n3476 );
not U_inv120 ( n75147, ex_wire40 );
dff P1_P3_DATAWIDTH_REG_7__reg ( clk, reset, ex_wire41, n3471 );
not U_inv121 ( n73341, ex_wire41 );
dff P1_P3_DATAWIDTH_REG_6__reg ( clk, reset, ex_wire42, n3466 );
not U_inv122 ( n75111, ex_wire42 );
dff P1_P3_DATAWIDTH_REG_5__reg ( clk, reset, ex_wire43, n3461 );
not U_inv123 ( n73371, ex_wire43 );
dff P1_P3_DATAWIDTH_REG_4__reg ( clk, reset, ex_wire44, n3456 );
not U_inv124 ( n75153, ex_wire44 );
dff P1_P3_DATAWIDTH_REG_3__reg ( clk, reset, ex_wire45, n3451 );
not U_inv125 ( n73361, ex_wire45 );
dff P1_P3_DATAWIDTH_REG_2__reg ( clk, reset, ex_wire46, n3446 );
not U_inv126 ( n75105, ex_wire46 );
dff P1_P3_DATAWIDTH_REG_1__reg ( clk, reset, P1_P3_DATAWIDTH_REG_1_, n3441 );
dff P1_P3_ADS_N_REG_reg ( clk, reset, P1_P3_ADS_N_REG, n5481 );
not U_inv127 ( n75968, P1_P3_ADS_N_REG );
dff P1_P3_STATEBS16_REG_reg ( clk, reset, P1_P3_STATEBS16_REG, n5456 );
not U_inv128 ( n74887, P1_P3_STATEBS16_REG );
dff P1_P3_INSTQUEUE_REG_15__7__reg ( clk, reset, ex_wire47, n3616 );
not U_inv129 ( n74341, ex_wire47 );
dff P1_P3_STATE2_REG_3__reg ( clk, reset, P1_P3_STATE2_REG_3_, n3596 );
dff P1_P3_INSTQUEUERD_ADDR_REG_4__reg ( clk, reset, P1_P3_INSTQUEUERD_ADDR_REG_4_, n4256 );
not U_inv130 ( n74611, P1_P3_INSTQUEUERD_ADDR_REG_4_ );
dff P1_P3_FLUSH_REG_reg ( clk, reset, P1_P3_FLUSH_REG, n5446 );
not U_inv131 ( n75230, P1_P3_FLUSH_REG );
dff P1_P3_INSTQUEUEWR_ADDR_REG_4__reg ( clk, reset, P1_P3_INSTQUEUEWR_ADDR_REG_4_, n4281 );
not U_inv132 ( n75032, P1_P3_INSTQUEUEWR_ADDR_REG_4_ );
dff P1_P3_INSTADDRPOINTER_REG_31__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_31_, n4461 );
not U_inv133 ( n75065, P1_P3_INSTADDRPOINTER_REG_31_ );
dff P1_P3_DATAO_REG_31__reg ( clk, reset, ex_wire48, n4936 );
not U_inv134 ( n73436, ex_wire48 );
dff P1_P3_INSTQUEUEWR_ADDR_REG_1__reg ( clk, reset, P1_P3_INSTQUEUEWR_ADDR_REG_1_, n4296 );
not U_inv135 ( n74561, P1_P3_INSTQUEUEWR_ADDR_REG_1_ );
dff P1_P3_INSTQUEUEWR_ADDR_REG_3__reg ( clk, reset, P1_P3_INSTQUEUEWR_ADDR_REG_3_, n4286 );
not U_inv136 ( n73138, P1_P3_INSTQUEUEWR_ADDR_REG_3_ );
dff P1_P3_EAX_REG_0__reg ( clk, reset, P1_P3_EAX_REG_0_, n4941 );
not U_inv137 ( n74488, P1_P3_EAX_REG_0_ );
dff P1_P3_EAX_REG_1__reg ( clk, reset, P1_P3_EAX_REG_1_, n4946 );
not U_inv138 ( n72957, P1_P3_EAX_REG_1_ );
dff P1_P3_EAX_REG_2__reg ( clk, reset, P1_P3_EAX_REG_2_, n4951 );
not U_inv139 ( n75286, P1_P3_EAX_REG_2_ );
dff P1_P3_EAX_REG_3__reg ( clk, reset, P1_P3_EAX_REG_3_, n4956 );
not U_inv140 ( n73135, P1_P3_EAX_REG_3_ );
dff P1_P3_EAX_REG_4__reg ( clk, reset, P1_P3_EAX_REG_4_, n4961 );
not U_inv141 ( n75279, P1_P3_EAX_REG_4_ );
dff P1_P3_EAX_REG_5__reg ( clk, reset, P1_P3_EAX_REG_5_, n4966 );
not U_inv142 ( n74540, P1_P3_EAX_REG_5_ );
dff P1_P3_EAX_REG_6__reg ( clk, reset, P1_P3_EAX_REG_6_, n4971 );
not U_inv143 ( n75282, P1_P3_EAX_REG_6_ );
dff P1_P3_EAX_REG_7__reg ( clk, reset, P1_P3_EAX_REG_7_, n4976 );
not U_inv144 ( n74582, P1_P3_EAX_REG_7_ );
dff P1_P3_EAX_REG_8__reg ( clk, reset, P1_P3_EAX_REG_8_, n4981 );
not U_inv145 ( n75281, P1_P3_EAX_REG_8_ );
dff P1_P3_EAX_REG_9__reg ( clk, reset, P1_P3_EAX_REG_9_, n4986 );
not U_inv146 ( n75252, P1_P3_EAX_REG_9_ );
dff P1_P3_EAX_REG_10__reg ( clk, reset, ex_wire49, n4991 );
not U_inv147 ( n74629, ex_wire49 );
dff P1_P3_LWORD_REG_10__reg ( clk, reset, P1_P3_LWORD_REG_10_, n4651 );
not U_inv148 ( n75699, P1_P3_LWORD_REG_10_ );
dff P1_P3_DATAO_REG_10__reg ( clk, reset, P1_P3_DATAO_REG_10_, n4831 );
dff P3_REG0_REG_10__reg ( clk, reset, P3_REG0_REG_10_, n1171 );
dff P3_REG0_REG_9__reg ( clk, reset, P3_REG0_REG_9_, n1166 );
dff P3_B_REG_reg ( clk, reset, P3_B_REG, n1861 );
not U_inv149 ( n74537, P3_B_REG );
dff P3_REG0_REG_29__reg ( clk, reset, P3_REG0_REG_29_, n1266 );
dff P3_REG2_REG_28__reg ( clk, reset, ex_wire50, n1581 );
not U_inv150 ( n74809, ex_wire50 );
dff P3_REG2_REG_27__reg ( clk, reset, P3_REG2_REG_27_, n1576 );
not U_inv151 ( n74821, P3_REG2_REG_27_ );
dff P3_REG2_REG_26__reg ( clk, reset, P3_REG2_REG_26_, n1571 );
not U_inv152 ( n74761, P3_REG2_REG_26_ );
dff P3_REG2_REG_25__reg ( clk, reset, ex_wire51, n1566 );
not U_inv153 ( n74714, ex_wire51 );
dff P3_REG2_REG_24__reg ( clk, reset, P3_REG2_REG_24_, n1561 );
not U_inv154 ( n74645, P3_REG2_REG_24_ );
dff P3_REG2_REG_23__reg ( clk, reset, P3_REG2_REG_23_, n1556 );
not U_inv155 ( n74552, P3_REG2_REG_23_ );
dff P3_REG2_REG_22__reg ( clk, reset, ex_wire52, n1551 );
not U_inv156 ( n74549, ex_wire52 );
dff P3_REG2_REG_21__reg ( clk, reset, P3_REG2_REG_21_, n1546 );
not U_inv157 ( n74520, P3_REG2_REG_21_ );
dff P3_REG2_REG_20__reg ( clk, reset, ex_wire53, n1541 );
not U_inv158 ( n74499, ex_wire53 );
dff P3_REG0_REG_19__reg ( clk, reset, P3_REG0_REG_19_, n1216 );
dff P3_REG2_REG_18__reg ( clk, reset, ex_wire54, n1531 );
not U_inv159 ( n74474, ex_wire54 );
dff P3_REG2_REG_17__reg ( clk, reset, P3_REG2_REG_17_, n1526 );
not U_inv160 ( n74448, P3_REG2_REG_17_ );
dff P3_REG0_REG_16__reg ( clk, reset, P3_REG0_REG_16_, n1201 );
dff P3_REG2_REG_15__reg ( clk, reset, P3_REG2_REG_15_, n1516 );
not U_inv161 ( n74407, P3_REG2_REG_15_ );
dff P3_REG2_REG_14__reg ( clk, reset, P3_REG2_REG_14_, n1511 );
not U_inv162 ( n74428, P3_REG2_REG_14_ );
dff P3_REG0_REG_13__reg ( clk, reset, P3_REG0_REG_13_, n1186 );
dff P3_REG2_REG_12__reg ( clk, reset, P3_REG2_REG_12_, n1501 );
not U_inv163 ( n74396, P3_REG2_REG_12_ );
dff P3_REG2_REG_11__reg ( clk, reset, P3_REG2_REG_11_, n1496 );
not U_inv164 ( n74378, P3_REG2_REG_11_ );
dff P2_P1_INSTQUEUE_REG_15__7__reg ( clk, reset, ex_wire55, n14841 );
not U_inv165 ( n74132, ex_wire55 );
dff P2_P1_STATE2_REG_3__reg ( clk, reset, P2_P1_STATE2_REG_3_, n14821 );
dff P2_P1_INSTQUEUE_REG_14__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__7_, n14881 );
not U_inv166 ( n74147, P2_P1_INSTQUEUE_REG_14__7_ );
dff P2_P1_FLUSH_REG_reg ( clk, reset, P2_P1_FLUSH_REG, n16671 );
not U_inv167 ( n75229, P2_P1_FLUSH_REG );
dff P2_P1_INSTQUEUERD_ADDR_REG_4__reg ( clk, reset, P2_P1_INSTQUEUERD_ADDR_REG_4_, n15481 );
not U_inv168 ( n74626, P2_P1_INSTQUEUERD_ADDR_REG_4_ );
dff P2_P1_INSTADDRPOINTER_REG_1__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_1_, n15536 );
not U_inv169 ( n75058, P2_P1_INSTADDRPOINTER_REG_1_ );
dff P2_P1_INSTADDRPOINTER_REG_3__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_3_, n15546 );
not U_inv170 ( n74400, P2_P1_INSTADDRPOINTER_REG_3_ );
dff P2_P1_PHYADDRPOINTER_REG_3__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_3_, n15706 );
not U_inv171 ( n73073, P2_P1_PHYADDRPOINTER_REG_3_ );
dff P2_P1_PHYADDRPOINTER_REG_4__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_4_, n15711 );
not U_inv172 ( n74473, P2_P1_PHYADDRPOINTER_REG_4_ );
dff P2_P1_PHYADDRPOINTER_REG_5__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_5_, n15716 );
not U_inv173 ( n73089, P2_P1_PHYADDRPOINTER_REG_5_ );
dff P2_P1_REIP_REG_5__reg ( clk, reset, P2_P1_REIP_REG_5_, n16511 );
not U_inv174 ( n74726, P2_P1_REIP_REG_5_ );
dff P2_P1_REIP_REG_6__reg ( clk, reset, ex_wire56, n16516 );
not U_inv175 ( n74728, ex_wire56 );
dff P2_P1_ADDRESS_REG_5__reg ( clk, reset, P2_P1_ADDRESS_REG_5_, n14616 );
not U_inv176 ( n73499, P2_P1_ADDRESS_REG_5_ );
dff P2_P1_UWORD_REG_7__reg ( clk, reset, P2_P1_UWORD_REG_7_, n15966 );
not U_inv177 ( n75495, P2_P1_UWORD_REG_7_ );
dff P2_P1_DATAO_REG_23__reg ( clk, reset, P2_P1_DATAO_REG_23_, n16121 );
dff P2_BUF1_REG_23__reg ( clk, reset, P2_BUF1_REG_23_, n576 );
not U_inv178 ( n75376, P2_BUF1_REG_23_ );
dff P2_P2_INSTQUEUE_REG_14__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__7_, n12636 );
not U_inv179 ( n74201, P2_P2_INSTQUEUE_REG_14__7_ );
dff P2_P2_INSTADDRPOINTER_REG_3__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_3_, n13301 );
not U_inv180 ( n74410, P2_P2_INSTADDRPOINTER_REG_3_ );
dff P2_P2_PHYADDRPOINTER_REG_3__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_3_, n13461 );
not U_inv181 ( n73081, P2_P2_PHYADDRPOINTER_REG_3_ );
dff P2_P2_PHYADDRPOINTER_REG_4__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_4_, n13466 );
not U_inv182 ( n74481, P2_P2_PHYADDRPOINTER_REG_4_ );
dff P2_P2_PHYADDRPOINTER_REG_5__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_5_, n13471 );
not U_inv183 ( n73092, P2_P2_PHYADDRPOINTER_REG_5_ );
dff P2_P2_REIP_REG_5__reg ( clk, reset, P2_P2_REIP_REG_5_, n14266 );
not U_inv184 ( n74693, P2_P2_REIP_REG_5_ );
dff P2_P2_REIP_REG_6__reg ( clk, reset, ex_wire57, n14271 );
not U_inv185 ( n74709, ex_wire57 );
dff P2_P2_INSTADDRPOINTER_REG_6__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_6_, n13316 );
not U_inv186 ( n73068, P2_P2_INSTADDRPOINTER_REG_6_ );
dff P2_P2_INSTADDRPOINTER_REG_7__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_7_, n13321 );
not U_inv187 ( n74698, P2_P2_INSTADDRPOINTER_REG_7_ );
dff P2_P2_PHYADDRPOINTER_REG_8__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_8_, n13486 );
not U_inv188 ( n74529, P2_P2_PHYADDRPOINTER_REG_8_ );
dff P2_P2_PHYADDRPOINTER_REG_9__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_9_, n13491 );
not U_inv189 ( n73111, P2_P2_PHYADDRPOINTER_REG_9_ );
dff P2_P2_PHYADDRPOINTER_REG_10__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_10_, n13496 );
not U_inv190 ( n74560, P2_P2_PHYADDRPOINTER_REG_10_ );
dff P2_P2_PHYADDRPOINTER_REG_11__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_11_, n13501 );
not U_inv191 ( n74464, P2_P2_PHYADDRPOINTER_REG_11_ );
dff P2_P2_REIP_REG_11__reg ( clk, reset, P2_P2_REIP_REG_11_, n14296 );
not U_inv192 ( n74788, P2_P2_REIP_REG_11_ );
dff P2_P2_REIP_REG_12__reg ( clk, reset, ex_wire58, n14301 );
not U_inv193 ( n74798, ex_wire58 );
dff P2_P2_INSTADDRPOINTER_REG_12__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_12_, n13346 );
not U_inv194 ( n74440, P2_P2_INSTADDRPOINTER_REG_12_ );
dff P2_P2_INSTADDRPOINTER_REG_15__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_15_, n13361 );
not U_inv195 ( n74854, P2_P2_INSTADDRPOINTER_REG_15_ );
dff P2_P2_PHYADDRPOINTER_REG_15__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_15_, n13521 );
not U_inv196 ( n75199, P2_P2_PHYADDRPOINTER_REG_15_ );
dff P2_P2_REIP_REG_15__reg ( clk, reset, P2_P2_REIP_REG_15_, n14316 );
not U_inv197 ( n74837, P2_P2_REIP_REG_15_ );
dff P2_P2_REIP_REG_16__reg ( clk, reset, P2_P2_REIP_REG_16_, n14321 );
not U_inv198 ( n73247, P2_P2_REIP_REG_16_ );
dff P2_P2_PHYADDRPOINTER_REG_16__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_16_, n13526 );
dff P2_P2_REIP_REG_17__reg ( clk, reset, P2_P2_REIP_REG_17_, n14326 );
not U_inv199 ( n74882, P2_P2_REIP_REG_17_ );
dff P2_P2_REIP_REG_18__reg ( clk, reset, P2_P2_REIP_REG_18_, n14331 );
not U_inv200 ( n74898, P2_P2_REIP_REG_18_ );
dff P2_P2_REIP_REG_19__reg ( clk, reset, P2_P2_REIP_REG_19_, n14336 );
not U_inv201 ( n73261, P2_P2_REIP_REG_19_ );
dff P2_P2_INSTADDRPOINTER_REG_19__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_19_, n13381 );
not U_inv202 ( n74576, P2_P2_INSTADDRPOINTER_REG_19_ );
dff P2_P2_INSTADDRPOINTER_REG_21__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_21_, n13391 );
not U_inv203 ( n73151, P2_P2_INSTADDRPOINTER_REG_21_ );
dff P2_P2_INSTADDRPOINTER_REG_22__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_22_, n13396 );
not U_inv204 ( n74597, P2_P2_INSTADDRPOINTER_REG_22_ );
dff P2_P2_PHYADDRPOINTER_REG_22__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_22_, n13556 );
not U_inv205 ( n75242, P2_P2_PHYADDRPOINTER_REG_22_ );
dff P2_P2_REIP_REG_22__reg ( clk, reset, P2_P2_REIP_REG_22_, n14351 );
not U_inv206 ( n73275, P2_P2_REIP_REG_22_ );
dff P2_P2_REIP_REG_23__reg ( clk, reset, P2_P2_REIP_REG_23_, n14356 );
not U_inv207 ( n74969, P2_P2_REIP_REG_23_ );
dff P2_P2_REIP_REG_24__reg ( clk, reset, P2_P2_REIP_REG_24_, n14361 );
not U_inv208 ( n74990, P2_P2_REIP_REG_24_ );
dff P2_P2_REIP_REG_25__reg ( clk, reset, P2_P2_REIP_REG_25_, n14366 );
not U_inv209 ( n73290, P2_P2_REIP_REG_25_ );
dff P2_P2_INSTADDRPOINTER_REG_28__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_28_, n13426 );
not U_inv210 ( n74977, P2_P2_INSTADDRPOINTER_REG_28_ );
dff P2_P2_PHYADDRPOINTER_REG_30__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_30_, n13596 );
not U_inv211 ( n75187, P2_P2_PHYADDRPOINTER_REG_30_ );
dff P2_P2_PHYADDRPOINTER_REG_31__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_31_, n13601 );
dff P2_P2_REIP_REG_0__reg ( clk, reset, P2_P2_REIP_REG_0_, n14241 );
not U_inv212 ( n75261, P2_P2_REIP_REG_0_ );
dff P2_P2_BYTEENABLE_REG_3__reg ( clk, reset, P2_P2_BYTEENABLE_REG_3_, n14401 );
dff P2_P2_BE_N_REG_3__reg ( clk, reset, P2_P2_BE_N_REG_3_, n12231 );
dff P2_READY12_REG_reg ( clk, reset, P2_READY12_REG, n781 );
dff P2_READY21_REG_reg ( clk, reset, P2_READY21_REG, n76557 );
dff P2_BUF2_REG_0__reg ( clk, reset, P2_BUF2_REG_0_, n621 );
not U_inv213 ( n75287, P2_BUF2_REG_0_ );
dff P2_P3_INSTQUEUE_REG_15__0__reg ( clk, reset, ex_wire59, n10386 );
not U_inv214 ( n73659, ex_wire59 );
dff P2_P3_MEMORYFETCH_REG_reg ( clk, reset, P2_P3_MEMORYFETCH_REG, n12226 );
dff P2_P3_READREQUEST_REG_reg ( clk, reset, P2_P3_READREQUEST_REG, n12221 );
dff P2_P3_CODEFETCH_REG_reg ( clk, reset, P2_P3_CODEFETCH_REG, n12211 );
dff P2_P3_MORE_REG_reg ( clk, reset, P2_P3_MORE_REG, n12186 );
dff P2_P3_LWORD_REG_0__reg ( clk, reset, P2_P3_LWORD_REG_0_, n11436 );
not U_inv215 ( n75634, P2_P3_LWORD_REG_0_ );
dff P2_P3_DATAO_REG_0__reg ( clk, reset, P2_P3_DATAO_REG_0_, n11516 );
dff P2_P3_LWORD_REG_15__reg ( clk, reset, P2_P3_LWORD_REG_15_, n11361 );
not U_inv216 ( n75633, P2_P3_LWORD_REG_15_ );
dff P2_P3_DATAO_REG_15__reg ( clk, reset, P2_P3_DATAO_REG_15_, n11591 );
dff P4_IR_REG_15__reg ( clk, reset, P4_IR_REG_15_, n2101 );
not U_inv217 ( n74391, P4_IR_REG_15_ );
dff P4_IR_REG_16__reg ( clk, reset, P4_IR_REG_16_, n2106 );
not U_inv218 ( n75417, P4_IR_REG_16_ );
dff P4_REG0_REG_30__reg ( clk, reset, P4_REG0_REG_30_, n2496 );
dff P4_DATAO_REG_30__reg ( clk, reset, P4_DATAO_REG_30_, n3076 );
not U_inv219 ( n73396, P4_DATAO_REG_30_ );
dff P1_P1_INSTQUEUE_REG_13__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__7_, n8186 );
not U_inv220 ( n74370, P1_P1_INSTQUEUE_REG_13__7_ );
dff P1_P1_EBX_REG_15__reg ( clk, reset, P1_P1_EBX_REG_15_, n9666 );
not U_inv221 ( n73246, P1_P1_EBX_REG_15_ );
dff P1_P1_EBX_REG_16__reg ( clk, reset, P1_P1_EBX_REG_16_, n9671 );
not U_inv222 ( n74834, P1_P1_EBX_REG_16_ );
dff P1_P1_REIP_REG_16__reg ( clk, reset, P1_P1_REIP_REG_16_, n9831 );
not U_inv223 ( n73254, P1_P1_REIP_REG_16_ );
dff P1_P1_PHYADDRPOINTER_REG_16__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_16_, n9036 );
dff P1_P1_REIP_REG_17__reg ( clk, reset, P1_P1_REIP_REG_17_, n9836 );
not U_inv224 ( n74905, P1_P1_REIP_REG_17_ );
dff P1_P1_REIP_REG_18__reg ( clk, reset, P1_P1_REIP_REG_18_, n9841 );
not U_inv225 ( n74915, P1_P1_REIP_REG_18_ );
dff P1_P1_REIP_REG_19__reg ( clk, reset, P1_P1_REIP_REG_19_, n9846 );
not U_inv226 ( n73268, P1_P1_REIP_REG_19_ );
dff P1_P1_INSTADDRPOINTER_REG_19__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_19_, n8891 );
not U_inv227 ( n74586, P1_P1_INSTADDRPOINTER_REG_19_ );
dff P1_P1_INSTADDRPOINTER_REG_21__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_21_, n8901 );
not U_inv228 ( n73158, P1_P1_INSTADDRPOINTER_REG_21_ );
dff P1_P1_INSTADDRPOINTER_REG_22__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_22_, n8906 );
not U_inv229 ( n74625, P1_P1_INSTADDRPOINTER_REG_22_ );
dff P1_P1_PHYADDRPOINTER_REG_24__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_24_, n9076 );
not U_inv230 ( n74737, P1_P1_PHYADDRPOINTER_REG_24_ );
dff P1_P1_REIP_REG_24__reg ( clk, reset, P1_P1_REIP_REG_24_, n9871 );
not U_inv231 ( n75006, P1_P1_REIP_REG_24_ );
dff P1_P1_REIP_REG_25__reg ( clk, reset, P1_P1_REIP_REG_25_, n9876 );
not U_inv232 ( n73305, P1_P1_REIP_REG_25_ );
dff P1_P1_PHYADDRPOINTER_REG_26__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_26_, n9086 );
not U_inv233 ( n74808, P1_P1_PHYADDRPOINTER_REG_26_ );
dff P1_P1_REIP_REG_26__reg ( clk, reset, P1_P1_REIP_REG_26_, n9881 );
not U_inv234 ( n73309, P1_P1_REIP_REG_26_ );
dff P1_P1_REIP_REG_27__reg ( clk, reset, P1_P1_REIP_REG_27_, n9886 );
not U_inv235 ( n75015, P1_P1_REIP_REG_27_ );
dff P1_P1_INSTADDRPOINTER_REG_27__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_27_, n8931 );
not U_inv236 ( n72970, P1_P1_INSTADDRPOINTER_REG_27_ );
dff P1_P1_PHYADDRPOINTER_REG_27__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_27_, n9091 );
not U_inv237 ( n75207, P1_P1_PHYADDRPOINTER_REG_27_ );
dff P1_P1_REIP_REG_29__reg ( clk, reset, P1_P1_REIP_REG_29_, n9896 );
not U_inv238 ( n73392, P1_P1_REIP_REG_29_ );
dff P1_P1_REIP_REG_30__reg ( clk, reset, P1_P1_REIP_REG_30_, n9901 );
not U_inv239 ( n75238, P1_P1_REIP_REG_30_ );
dff P1_P1_REIP_REG_31__reg ( clk, reset, P1_P1_REIP_REG_31_, n9906 );
not U_inv240 ( n75329, P1_P1_REIP_REG_31_ );
dff P1_P1_INSTADDRPOINTER_REG_31__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_31_, n8951 );
not U_inv241 ( n75051, P1_P1_INSTADDRPOINTER_REG_31_ );
dff P1_P1_PHYADDRPOINTER_REG_31__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_31_, n9111 );
not U_inv242 ( n74964, P1_P1_PHYADDRPOINTER_REG_31_ );
dff P1_P1_REIP_REG_1__reg ( clk, reset, P1_P1_REIP_REG_1_, n9756 );
not U_inv243 ( n72963, P1_P1_REIP_REG_1_ );
dff P1_P1_BYTEENABLE_REG_2__reg ( clk, reset, P1_P1_BYTEENABLE_REG_2_, n9916 );
dff P1_P1_BE_N_REG_2__reg ( clk, reset, P1_P1_BE_N_REG_2_, n7746 );
dff P1_READY11_REG_reg ( clk, reset, P1_READY11_REG, n456 );
dff P1_BUF1_REG_0__reg ( clk, reset, P1_BUF1_REG_0_, n121 );
not U_inv244 ( n75462, P1_BUF1_REG_0_ );
dff P1_P2_INSTQUEUE_REG_15__0__reg ( clk, reset, ex_wire60, n5896 );
not U_inv245 ( n73661, ex_wire60 );
dff P1_P2_PHYADDRPOINTER_REG_27__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_27_, n6846 );
not U_inv246 ( n74850, P1_P2_PHYADDRPOINTER_REG_27_ );
dff P1_P2_PHYADDRPOINTER_REG_28__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_28_, n6851 );
not U_inv247 ( n75243, P1_P2_PHYADDRPOINTER_REG_28_ );
dff P1_P2_REIP_REG_28__reg ( clk, reset, P1_P2_REIP_REG_28_, n7646 );
not U_inv248 ( n75301, P1_P2_REIP_REG_28_ );
dff P1_P2_REIP_REG_29__reg ( clk, reset, P1_P2_REIP_REG_29_, n7651 );
not U_inv249 ( n73317, P1_P2_REIP_REG_29_ );
dff P1_P2_REIP_REG_30__reg ( clk, reset, P1_P2_REIP_REG_30_, n7656 );
not U_inv250 ( n75064, P1_P2_REIP_REG_30_ );
dff P1_P2_ADDRESS_REG_29__reg ( clk, reset, P1_P2_ADDRESS_REG_29_, n5516 );
dff P1_READY12_REG_reg ( clk, reset, P1_READY12_REG, n441 );
dff P1_P2_STATE_REG_2__reg ( clk, reset, P1_P2_STATE_REG_2_, n5666 );
not U_inv251 ( n74651, P1_P2_STATE_REG_2_ );
dff P1_P2_STATE_REG_1__reg ( clk, reset, P1_P2_STATE_REG_1_, n5671 );
not U_inv252 ( n73179, P1_P2_STATE_REG_1_ );
dff P1_P2_BE_N_REG_3__reg ( clk, reset, P1_P2_BE_N_REG_3_, n5496 );
dff P1_READY21_REG_reg ( clk, reset, P1_READY21_REG, n76464 );
dff P1_BUF2_REG_0__reg ( clk, reset, P1_BUF2_REG_0_, n281 );
not U_inv253 ( n75288, P1_BUF2_REG_0_ );
dff P1_P3_INSTQUEUE_REG_15__0__reg ( clk, reset, ex_wire61, n3651 );
not U_inv254 ( n74002, ex_wire61 );
dff P1_P3_MEMORYFETCH_REG_reg ( clk, reset, P1_P3_MEMORYFETCH_REG, n5491 );
dff P1_P3_M_IO_N_REG_reg ( clk, reset, P1_P3_M_IO_N_REG, n5471 );
dff P1_P3_READREQUEST_REG_reg ( clk, reset, P1_P3_READREQUEST_REG, n5486 );
dff P1_P3_W_R_N_REG_reg ( clk, reset, P1_P3_W_R_N_REG, n5441 );
dff P1_P3_CODEFETCH_REG_reg ( clk, reset, P1_P3_CODEFETCH_REG, n5476 );
dff P1_P3_D_C_N_REG_reg ( clk, reset, P1_P3_D_C_N_REG, n5466 );
dff P1_P3_MORE_REG_reg ( clk, reset, P1_P3_MORE_REG, n5451 );
dff P1_P3_LWORD_REG_0__reg ( clk, reset, P1_P3_LWORD_REG_0_, n4701 );
not U_inv255 ( n75698, P1_P3_LWORD_REG_0_ );
dff P1_P3_DATAO_REG_0__reg ( clk, reset, P1_P3_DATAO_REG_0_, n4781 );
dff P1_P3_LWORD_REG_15__reg ( clk, reset, P1_P3_LWORD_REG_15_, n4626 );
not U_inv256 ( n75697, P1_P3_LWORD_REG_15_ );
dff P1_P3_DATAO_REG_15__reg ( clk, reset, P1_P3_DATAO_REG_15_, n4856 );
dff P3_REG0_REG_30__reg ( clk, reset, P3_REG0_REG_30_, n1271 );
dff P3_DATAO_REG_30__reg ( clk, reset, P3_DATAO_REG_30_, n1851 );
dff P2_P1_INSTQUEUE_REG_13__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__7_, n14921 );
not U_inv257 ( n74144, P2_P1_INSTQUEUE_REG_13__7_ );
dff P2_P1_EAX_REG_15__reg ( clk, reset, ex_wire62, n16241 );
not U_inv258 ( n74865, ex_wire62 );
dff P2_P1_LWORD_REG_15__reg ( clk, reset, P2_P1_LWORD_REG_15_, n15851 );
not U_inv259 ( n75667, P2_P1_LWORD_REG_15_ );
dff P2_P1_DATAO_REG_15__reg ( clk, reset, P2_P1_DATAO_REG_15_, n16081 );
dff P2_BUF1_REG_15__reg ( clk, reset, P2_BUF1_REG_15_, n536 );
not U_inv260 ( n75436, P2_BUF1_REG_15_ );
dff P2_P2_LWORD_REG_15__reg ( clk, reset, P2_P2_LWORD_REG_15_, n13606 );
not U_inv261 ( n75632, P2_P2_LWORD_REG_15_ );
dff P2_P2_DATAO_REG_15__reg ( clk, reset, P2_P2_DATAO_REG_15_, n13836 );
not U_inv262 ( n75525, P2_P2_DATAO_REG_15_ );
dff P2_BUF2_REG_15__reg ( clk, reset, P2_BUF2_REG_15_, n696 );
not U_inv263 ( n75364, P2_BUF2_REG_15_ );
dff P2_P3_EAX_REG_15__reg ( clk, reset, P2_P3_EAX_REG_15_, n11751 );
not U_inv264 ( n74776, P2_P3_EAX_REG_15_ );
dff P2_P3_EAX_REG_16__reg ( clk, reset, P2_P3_EAX_REG_16_, n11756 );
not U_inv265 ( n75384, P2_P3_EAX_REG_16_ );
dff P2_P3_UWORD_REG_0__reg ( clk, reset, P2_P3_UWORD_REG_0_, n11511 );
not U_inv266 ( n75478, P2_P3_UWORD_REG_0_ );
dff P2_P3_DATAO_REG_16__reg ( clk, reset, P2_P3_DATAO_REG_16_, n11596 );
dff P2_P3_EAX_REG_17__reg ( clk, reset, P2_P3_EAX_REG_17_, n11761 );
not U_inv267 ( n74814, P2_P3_EAX_REG_17_ );
dff P2_P3_UWORD_REG_1__reg ( clk, reset, P2_P3_UWORD_REG_1_, n11506 );
not U_inv268 ( n75477, P2_P3_UWORD_REG_1_ );
dff P2_P3_DATAO_REG_17__reg ( clk, reset, P2_P3_DATAO_REG_17_, n11601 );
dff P4_IR_REG_17__reg ( clk, reset, P4_IR_REG_17_, n2111 );
not U_inv269 ( n73495, P4_IR_REG_17_ );
dff P4_IR_REG_18__reg ( clk, reset, P4_IR_REG_18_, n2116 );
not U_inv270 ( n73035, P4_IR_REG_18_ );
dff P4_IR_REG_19__reg ( clk, reset, P4_IR_REG_19_, n2121 );
not U_inv271 ( n73479, P4_IR_REG_19_ );
dff P4_IR_REG_20__reg ( clk, reset, P4_IR_REG_20_, n2126 );
not U_inv272 ( n73042, P4_IR_REG_20_ );
dff P4_IR_REG_21__reg ( clk, reset, P4_IR_REG_21_, n2131 );
not U_inv273 ( n73494, P4_IR_REG_21_ );
dff P4_REG0_REG_0__reg ( clk, reset, P4_REG0_REG_0_, n2346 );
dff P4_REG1_REG_0__reg ( clk, reset, P4_REG1_REG_0_, n2506 );
not U_inv274 ( n73798, P4_REG1_REG_0_ );
dff P4_REG3_REG_9__reg ( clk, reset, P4_REG3_REG_9_, n3141 );
not U_inv275 ( n72932, P4_REG3_REG_9_ );
dff P4_REG2_REG_8__reg ( clk, reset, P4_REG2_REG_8_, n2706 );
not U_inv276 ( n74371, P4_REG2_REG_8_ );
dff P4_REG0_REG_7__reg ( clk, reset, P4_REG0_REG_7_, n2381 );
dff P4_REG0_REG_6__reg ( clk, reset, P4_REG0_REG_6_, n2376 );
dff P4_REG0_REG_5__reg ( clk, reset, P4_REG0_REG_5_, n2371 );
dff P4_REG2_REG_4__reg ( clk, reset, P4_REG2_REG_4_, n2686 );
not U_inv277 ( n74218, P4_REG2_REG_4_ );
dff P4_REG0_REG_3__reg ( clk, reset, P4_REG0_REG_3_, n2361 );
dff P4_REG2_REG_2__reg ( clk, reset, P4_REG2_REG_2_, n2676 );
not U_inv278 ( n73897, P4_REG2_REG_2_ );
dff P4_REG0_REG_1__reg ( clk, reset, P4_REG0_REG_1_, n2351 );
dff P1_P1_INSTQUEUE_REG_15__6__reg ( clk, reset, ex_wire63, n8111 );
not U_inv279 ( n74333, ex_wire63 );
dff P1_P1_INSTQUEUEWR_ADDR_REG_4__reg ( clk, reset, P1_P1_INSTQUEUEWR_ADDR_REG_4_, n8771 );
not U_inv280 ( n75031, P1_P1_INSTQUEUEWR_ADDR_REG_4_ );
dff P1_P1_INSTQUEUE_REG_14__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__4_, n8161 );
not U_inv281 ( n74250, P1_P1_INSTQUEUE_REG_14__4_ );
dff P1_P1_EAX_REG_4__reg ( clk, reset, P1_P1_EAX_REG_4_, n9451 );
not U_inv282 ( n74682, P1_P1_EAX_REG_4_ );
dff P1_P1_LWORD_REG_4__reg ( clk, reset, P1_P1_LWORD_REG_4_, n9171 );
not U_inv283 ( n75682, P1_P1_LWORD_REG_4_ );
dff P1_P1_DATAO_REG_4__reg ( clk, reset, P1_P1_DATAO_REG_4_, n9291 );
dff P1_BUF1_REG_4__reg ( clk, reset, P1_BUF1_REG_4_, n141 );
not U_inv284 ( n75461, P1_BUF1_REG_4_ );
dff P1_P2_INSTQUEUE_REG_15__4__reg ( clk, reset, ex_wire64, n5876 );
not U_inv285 ( n73841, ex_wire64 );
dff P1_P2_INSTQUEUEWR_ADDR_REG_4__reg ( clk, reset, P1_P2_INSTQUEUEWR_ADDR_REG_4_, n6526 );
not U_inv286 ( n75033, P1_P2_INSTQUEUEWR_ADDR_REG_4_ );
dff P1_P2_EAX_REG_0__reg ( clk, reset, P1_P2_EAX_REG_0_, n7186 );
not U_inv287 ( n74491, P1_P2_EAX_REG_0_ );
dff P1_P2_EAX_REG_1__reg ( clk, reset, P1_P2_EAX_REG_1_, n7191 );
not U_inv288 ( n73129, P1_P2_EAX_REG_1_ );
dff P1_P2_EAX_REG_2__reg ( clk, reset, P1_P2_EAX_REG_2_, n7196 );
not U_inv289 ( n75285, P1_P2_EAX_REG_2_ );
dff P1_P2_EAX_REG_3__reg ( clk, reset, P1_P2_EAX_REG_3_, n7201 );
not U_inv290 ( n74510, P1_P2_EAX_REG_3_ );
dff P1_P2_EAX_REG_4__reg ( clk, reset, P1_P2_EAX_REG_4_, n7206 );
not U_inv291 ( n75276, P1_P2_EAX_REG_4_ );
dff P1_P2_EAX_REG_5__reg ( clk, reset, P1_P2_EAX_REG_5_, n7211 );
not U_inv292 ( n74543, P1_P2_EAX_REG_5_ );
dff P1_P2_EAX_REG_6__reg ( clk, reset, P1_P2_EAX_REG_6_, n7216 );
not U_inv293 ( n75277, P1_P2_EAX_REG_6_ );
dff P1_P2_EAX_REG_7__reg ( clk, reset, P1_P2_EAX_REG_7_, n7221 );
not U_inv294 ( n74584, P1_P2_EAX_REG_7_ );
dff P1_P2_EAX_REG_8__reg ( clk, reset, P1_P2_EAX_REG_8_, n7226 );
not U_inv295 ( n75275, P1_P2_EAX_REG_8_ );
dff P1_P2_EAX_REG_9__reg ( clk, reset, P1_P2_EAX_REG_9_, n7231 );
not U_inv296 ( n75251, P1_P2_EAX_REG_9_ );
dff P1_P2_EAX_REG_10__reg ( clk, reset, ex_wire65, n7236 );
not U_inv297 ( n74633, ex_wire65 );
dff P1_P2_LWORD_REG_10__reg ( clk, reset, P1_P2_LWORD_REG_10_, n6896 );
not U_inv298 ( n75651, P1_P2_LWORD_REG_10_ );
dff P1_P2_DATAO_REG_10__reg ( clk, reset, P1_P2_DATAO_REG_10_, n7076 );
not U_inv299 ( n75531, P1_P2_DATAO_REG_10_ );
dff P1_BUF2_REG_10__reg ( clk, reset, P1_BUF2_REG_10_, n331 );
not U_inv300 ( n75321, P1_BUF2_REG_10_ );
dff P1_P2_UWORD_REG_10__reg ( clk, reset, P1_P2_UWORD_REG_10_, n6971 );
not U_inv301 ( n75572, P1_P2_UWORD_REG_10_ );
dff P1_P2_DATAO_REG_26__reg ( clk, reset, P1_P2_DATAO_REG_26_, n7156 );
not U_inv302 ( n75595, P1_P2_DATAO_REG_26_ );
dff P1_BUF2_REG_26__reg ( clk, reset, P1_BUF2_REG_26_, n411 );
not U_inv303 ( n75333, P1_BUF2_REG_26_ );
dff P1_P3_INSTQUEUE_REG_14__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__2_, n3681 );
not U_inv304 ( n74044, P1_P3_INSTQUEUE_REG_14__2_ );
dff P1_P3_EAX_REG_18__reg ( clk, reset, P1_P3_EAX_REG_18_, n5031 );
not U_inv305 ( n75422, P1_P3_EAX_REG_18_ );
dff P1_P3_EAX_REG_19__reg ( clk, reset, P1_P3_EAX_REG_19_, n5036 );
not U_inv306 ( n74876, P1_P3_EAX_REG_19_ );
dff P1_P3_UWORD_REG_3__reg ( clk, reset, P1_P3_UWORD_REG_3_, n4761 );
not U_inv307 ( n75600, P1_P3_UWORD_REG_3_ );
dff P1_P3_DATAO_REG_19__reg ( clk, reset, P1_P3_DATAO_REG_19_, n4876 );
dff P3_IR_REG_19__reg ( clk, reset, P3_IR_REG_19_, n896 );
dff P3_IR_REG_27__reg ( clk, reset, P3_IR_REG_27_, n936 );
not U_inv308 ( n73506, P3_IR_REG_27_ );
dff P3_IR_REG_30__reg ( clk, reset, P3_IR_REG_30_, n951 );
dff P3_IR_REG_29__reg ( clk, reset, P3_IR_REG_29_, n946 );
dff P3_IR_REG_28__reg ( clk, reset, P3_IR_REG_28_, n941 );
dff P3_IR_REG_25__reg ( clk, reset, P3_IR_REG_25_, n926 );
dff P3_IR_REG_24__reg ( clk, reset, P3_IR_REG_24_, n921 );
dff P3_IR_REG_23__reg ( clk, reset, P3_IR_REG_23_, n916 );
dff P3_IR_REG_21__reg ( clk, reset, P3_IR_REG_21_, n906 );
dff P3_IR_REG_22__reg ( clk, reset, P3_IR_REG_22_, n911 );
dff P3_IR_REG_20__reg ( clk, reset, P3_IR_REG_20_, n901 );
dff P3_IR_REG_0__reg ( clk, reset, P3_IR_REG_0_, n801 );
not U_inv309 ( n73024, P3_IR_REG_0_ );
dff P3_IR_REG_26__reg ( clk, reset, P3_IR_REG_26_, n931 );
dff P3_D_REG_7__reg ( clk, reset, ex_wire66, n996 );
not U_inv310 ( n74624, ex_wire66 );
dff P3_D_REG_22__reg ( clk, reset, ex_wire67, n1071 );
not U_inv311 ( n74623, ex_wire67 );
dff P3_D_REG_6__reg ( clk, reset, P3_D_REG_6_, n991 );
dff P3_D_REG_5__reg ( clk, reset, P3_D_REG_5_, n986 );
dff P3_D_REG_4__reg ( clk, reset, P3_D_REG_4_, n981 );
dff P3_D_REG_3__reg ( clk, reset, P3_D_REG_3_, n976 );
dff P3_D_REG_2__reg ( clk, reset, P3_D_REG_2_, n971 );
dff P3_D_REG_1__reg ( clk, reset, P3_D_REG_1_, n966 );
dff P3_D_REG_0__reg ( clk, reset, P3_D_REG_0_, n961 );
dff P3_D_REG_31__reg ( clk, reset, P3_D_REG_31_, n1116 );
dff P3_D_REG_30__reg ( clk, reset, P3_D_REG_30_, n1111 );
dff P3_D_REG_29__reg ( clk, reset, P3_D_REG_29_, n1106 );
dff P3_D_REG_28__reg ( clk, reset, P3_D_REG_28_, n1101 );
dff P3_D_REG_27__reg ( clk, reset, P3_D_REG_27_, n1096 );
dff P3_D_REG_26__reg ( clk, reset, P3_D_REG_26_, n1091 );
dff P3_D_REG_25__reg ( clk, reset, P3_D_REG_25_, n1086 );
dff P3_D_REG_24__reg ( clk, reset, P3_D_REG_24_, n1081 );
dff P3_D_REG_23__reg ( clk, reset, P3_D_REG_23_, n1076 );
dff P3_D_REG_21__reg ( clk, reset, P3_D_REG_21_, n1066 );
dff P3_D_REG_20__reg ( clk, reset, P3_D_REG_20_, n1061 );
dff P3_D_REG_19__reg ( clk, reset, P3_D_REG_19_, n1056 );
dff P3_D_REG_18__reg ( clk, reset, P3_D_REG_18_, n1051 );
dff P3_D_REG_17__reg ( clk, reset, P3_D_REG_17_, n1046 );
dff P3_D_REG_16__reg ( clk, reset, P3_D_REG_16_, n1041 );
dff P3_D_REG_15__reg ( clk, reset, P3_D_REG_15_, n1036 );
dff P3_D_REG_14__reg ( clk, reset, P3_D_REG_14_, n1031 );
dff P3_D_REG_13__reg ( clk, reset, P3_D_REG_13_, n1026 );
dff P3_D_REG_12__reg ( clk, reset, P3_D_REG_12_, n1021 );
dff P3_D_REG_11__reg ( clk, reset, P3_D_REG_11_, n1016 );
dff P3_D_REG_10__reg ( clk, reset, P3_D_REG_10_, n1011 );
dff P3_D_REG_9__reg ( clk, reset, P3_D_REG_9_, n1006 );
dff P3_D_REG_8__reg ( clk, reset, P3_D_REG_8_, n1001 );
dff P3_RD_REG_reg ( clk, reset, P3_RD_REG, n2016 );
dff P3_WR_REG_reg ( clk, reset, P3_WR_REG, n76376 );
not U_inv312 ( n73026, P3_WR_REG );
dff P3_DATAO_REG_29__reg ( clk, reset, P3_DATAO_REG_29_, n1846 );
not U_inv313 ( n73402, P3_DATAO_REG_29_ );
dff P3_DATAO_REG_28__reg ( clk, reset, P3_DATAO_REG_28_, n1841 );
not U_inv314 ( n73405, P3_DATAO_REG_28_ );
dff P3_DATAO_REG_27__reg ( clk, reset, P3_DATAO_REG_27_, n1836 );
not U_inv315 ( n73010, P3_DATAO_REG_27_ );
dff P3_DATAO_REG_26__reg ( clk, reset, P3_DATAO_REG_26_, n1831 );
not U_inv316 ( n73014, P3_DATAO_REG_26_ );
dff P3_DATAO_REG_25__reg ( clk, reset, P3_DATAO_REG_25_, n1826 );
not U_inv317 ( n73415, P3_DATAO_REG_25_ );
dff P3_DATAO_REG_24__reg ( clk, reset, P3_DATAO_REG_24_, n1821 );
not U_inv318 ( n73016, P3_DATAO_REG_24_ );
dff P3_DATAO_REG_23__reg ( clk, reset, P3_DATAO_REG_23_, n1816 );
not U_inv319 ( n73416, P3_DATAO_REG_23_ );
dff P3_DATAO_REG_21__reg ( clk, reset, P3_DATAO_REG_21_, n1806 );
not U_inv320 ( n73001, P3_DATAO_REG_21_ );
dff P3_DATAO_REG_20__reg ( clk, reset, P3_DATAO_REG_20_, n1801 );
not U_inv321 ( n73401, P3_DATAO_REG_20_ );
dff P3_DATAO_REG_19__reg ( clk, reset, P3_DATAO_REG_19_, n1796 );
not U_inv322 ( n73005, P3_DATAO_REG_19_ );
dff P3_DATAO_REG_18__reg ( clk, reset, P3_DATAO_REG_18_, n1791 );
not U_inv323 ( n73403, P3_DATAO_REG_18_ );
dff P3_DATAO_REG_17__reg ( clk, reset, P3_DATAO_REG_17_, n1786 );
not U_inv324 ( n73002, P3_DATAO_REG_17_ );
dff P3_DATAO_REG_14__reg ( clk, reset, P3_DATAO_REG_14_, n1771 );
not U_inv325 ( n73400, P3_DATAO_REG_14_ );
dff P3_REG1_REG_30__reg ( clk, reset, P3_REG1_REG_30_, n1431 );
not U_inv326 ( n74866, P3_REG1_REG_30_ );
dff P3_REG1_REG_29__reg ( clk, reset, P3_REG1_REG_29_, n1426 );
not U_inv327 ( n74863, P3_REG1_REG_29_ );
dff P3_REG1_REG_19__reg ( clk, reset, P3_REG1_REG_19_, n1376 );
not U_inv328 ( n74498, P3_REG1_REG_19_ );
dff P3_REG1_REG_16__reg ( clk, reset, P3_REG1_REG_16_, n1361 );
not U_inv329 ( n74416, P3_REG1_REG_16_ );
dff P3_REG1_REG_13__reg ( clk, reset, P3_REG1_REG_13_, n1346 );
not U_inv330 ( n74406, P3_REG1_REG_13_ );
dff P3_REG1_REG_10__reg ( clk, reset, P3_REG1_REG_10_, n1331 );
not U_inv331 ( n74380, P3_REG1_REG_10_ );
dff P3_REG1_REG_9__reg ( clk, reset, P3_REG1_REG_9_, n1326 );
not U_inv332 ( n74386, P3_REG1_REG_9_ );
dff P3_REG2_REG_31__reg ( clk, reset, P3_REG2_REG_31_, n1596 );
not U_inv333 ( n74846, P3_REG2_REG_31_ );
dff P3_REG1_REG_31__reg ( clk, reset, P3_REG1_REG_31_, n1436 );
not U_inv334 ( n74844, P3_REG1_REG_31_ );
dff P3_REG0_REG_31__reg ( clk, reset, P3_REG0_REG_31_, n1276 );
dff P3_DATAO_REG_31__reg ( clk, reset, P3_DATAO_REG_31_, n1856 );
not U_inv335 ( n73431, P3_DATAO_REG_31_ );
dff P3_REG2_REG_30__reg ( clk, reset, P3_REG2_REG_30_, n1591 );
not U_inv336 ( n74867, P3_REG2_REG_30_ );
dff P3_REG1_REG_0__reg ( clk, reset, P3_REG1_REG_0_, n1281 );
not U_inv337 ( n73579, P3_REG1_REG_0_ );
dff P3_REG0_REG_0__reg ( clk, reset, P3_REG0_REG_0_, n1121 );
dff P3_REG1_REG_1__reg ( clk, reset, P3_REG1_REG_1_, n1286 );
not U_inv338 ( n73825, P3_REG1_REG_1_ );
dff P3_REG0_REG_1__reg ( clk, reset, P3_REG0_REG_1_, n1126 );
dff P3_REG3_REG_0__reg ( clk, reset, P3_REG3_REG_0_, n1911 );
not U_inv339 ( n73637, P3_REG3_REG_0_ );
dff P3_REG1_REG_2__reg ( clk, reset, P3_REG1_REG_2_, n1291 );
not U_inv340 ( n73829, P3_REG1_REG_2_ );
dff P3_REG0_REG_2__reg ( clk, reset, P3_REG0_REG_2_, n1131 );
dff P3_REG1_REG_3__reg ( clk, reset, P3_REG1_REG_3_, n1296 );
not U_inv341 ( n73911, P3_REG1_REG_3_ );
dff P3_REG0_REG_3__reg ( clk, reset, P3_REG0_REG_3_, n1136 );
dff P3_REG1_REG_4__reg ( clk, reset, P3_REG1_REG_4_, n1301 );
not U_inv342 ( n74219, P3_REG1_REG_4_ );
dff P3_REG0_REG_4__reg ( clk, reset, P3_REG0_REG_4_, n1141 );
dff P3_REG1_REG_5__reg ( clk, reset, P3_REG1_REG_5_, n1306 );
not U_inv343 ( n74263, P3_REG1_REG_5_ );
dff P3_REG0_REG_5__reg ( clk, reset, P3_REG0_REG_5_, n1146 );
dff P3_REG1_REG_6__reg ( clk, reset, P3_REG1_REG_6_, n1311 );
not U_inv344 ( n74282, P3_REG1_REG_6_ );
dff P3_REG0_REG_6__reg ( clk, reset, P3_REG0_REG_6_, n1151 );
dff P3_REG1_REG_7__reg ( clk, reset, P3_REG1_REG_7_, n1316 );
not U_inv345 ( n74337, P3_REG1_REG_7_ );
dff P3_REG0_REG_7__reg ( clk, reset, P3_REG0_REG_7_, n1156 );
dff P3_REG1_REG_8__reg ( clk, reset, P3_REG1_REG_8_, n1321 );
not U_inv346 ( n74383, P3_REG1_REG_8_ );
dff P3_REG0_REG_8__reg ( clk, reset, P3_REG0_REG_8_, n1161 );
dff P2_P1_INSTQUEUE_REG_15__6__reg ( clk, reset, ex_wire68, n14846 );
not U_inv347 ( n73968, ex_wire68 );
dff P2_P1_INSTQUEUEWR_ADDR_REG_4__reg ( clk, reset, P2_P1_INSTQUEUEWR_ADDR_REG_4_, n15506 );
not U_inv348 ( n75030, P2_P1_INSTQUEUEWR_ADDR_REG_4_ );
dff P2_P1_INSTQUEUE_REG_14__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__4_, n14896 );
not U_inv349 ( n73815, P2_P1_INSTQUEUE_REG_14__4_ );
dff P2_P1_EAX_REG_4__reg ( clk, reset, P2_P1_EAX_REG_4_, n16186 );
not U_inv350 ( n74681, P2_P1_EAX_REG_4_ );
dff P2_P1_LWORD_REG_4__reg ( clk, reset, P2_P1_LWORD_REG_4_, n15906 );
not U_inv351 ( n75666, P2_P1_LWORD_REG_4_ );
dff P2_P1_DATAO_REG_4__reg ( clk, reset, P2_P1_DATAO_REG_4_, n16026 );
dff P2_BUF1_REG_4__reg ( clk, reset, P2_BUF1_REG_4_, n481 );
not U_inv352 ( n75454, P2_BUF1_REG_4_ );
dff P2_P2_INSTQUEUE_REG_15__4__reg ( clk, reset, ex_wire69, n12611 );
not U_inv353 ( n73842, ex_wire69 );
dff P2_P2_INSTQUEUEWR_ADDR_REG_4__reg ( clk, reset, P2_P2_INSTQUEUEWR_ADDR_REG_4_, n13261 );
not U_inv354 ( n75035, P2_P2_INSTQUEUEWR_ADDR_REG_4_ );
dff P2_P2_EAX_REG_0__reg ( clk, reset, P2_P2_EAX_REG_0_, n13921 );
not U_inv355 ( n74490, P2_P2_EAX_REG_0_ );
dff P2_P2_EAX_REG_1__reg ( clk, reset, P2_P2_EAX_REG_1_, n13926 );
not U_inv356 ( n73128, P2_P2_EAX_REG_1_ );
dff P2_P2_EAX_REG_2__reg ( clk, reset, P2_P2_EAX_REG_2_, n13931 );
not U_inv357 ( n75283, P2_P2_EAX_REG_2_ );
dff P2_P2_EAX_REG_3__reg ( clk, reset, P2_P2_EAX_REG_3_, n13936 );
not U_inv358 ( n74509, P2_P2_EAX_REG_3_ );
dff P2_P2_EAX_REG_4__reg ( clk, reset, P2_P2_EAX_REG_4_, n13941 );
not U_inv359 ( n75267, P2_P2_EAX_REG_4_ );
dff P2_P2_EAX_REG_5__reg ( clk, reset, P2_P2_EAX_REG_5_, n13946 );
not U_inv360 ( n74542, P2_P2_EAX_REG_5_ );
dff P2_P2_EAX_REG_6__reg ( clk, reset, P2_P2_EAX_REG_6_, n13951 );
not U_inv361 ( n75263, P2_P2_EAX_REG_6_ );
dff P2_P2_EAX_REG_7__reg ( clk, reset, P2_P2_EAX_REG_7_, n13956 );
not U_inv362 ( n74583, P2_P2_EAX_REG_7_ );
dff P2_P2_EAX_REG_8__reg ( clk, reset, P2_P2_EAX_REG_8_, n13961 );
not U_inv363 ( n75265, P2_P2_EAX_REG_8_ );
dff P2_P2_EAX_REG_9__reg ( clk, reset, P2_P2_EAX_REG_9_, n13966 );
not U_inv364 ( n75249, P2_P2_EAX_REG_9_ );
dff P2_P2_EAX_REG_10__reg ( clk, reset, ex_wire70, n13971 );
not U_inv365 ( n74632, ex_wire70 );
dff P2_P2_LWORD_REG_10__reg ( clk, reset, P2_P2_LWORD_REG_10_, n13631 );
not U_inv366 ( n75631, P2_P2_LWORD_REG_10_ );
dff P2_P2_DATAO_REG_10__reg ( clk, reset, P2_P2_DATAO_REG_10_, n13811 );
not U_inv367 ( n75506, P2_P2_DATAO_REG_10_ );
dff P2_BUF2_REG_10__reg ( clk, reset, P2_BUF2_REG_10_, n671 );
not U_inv368 ( n75310, P2_BUF2_REG_10_ );
dff P2_P2_UWORD_REG_10__reg ( clk, reset, P2_P2_UWORD_REG_10_, n13706 );
not U_inv369 ( n75565, P2_P2_UWORD_REG_10_ );
dff P2_P2_DATAO_REG_26__reg ( clk, reset, P2_P2_DATAO_REG_26_, n13891 );
not U_inv370 ( n75589, P2_P2_DATAO_REG_26_ );
dff P2_BUF2_REG_26__reg ( clk, reset, P2_BUF2_REG_26_, n751 );
not U_inv371 ( n75339, P2_BUF2_REG_26_ );
dff P2_P3_INSTQUEUE_REG_14__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__2_, n10416 );
not U_inv372 ( n73740, P2_P3_INSTQUEUE_REG_14__2_ );
dff P2_P3_EAX_REG_18__reg ( clk, reset, P2_P3_EAX_REG_18_, n11766 );
not U_inv373 ( n75382, P2_P3_EAX_REG_18_ );
dff P2_P3_EAX_REG_19__reg ( clk, reset, P2_P3_EAX_REG_19_, n11771 );
not U_inv374 ( n74875, P2_P3_EAX_REG_19_ );
dff P2_P3_EAX_REG_20__reg ( clk, reset, P2_P3_EAX_REG_20_, n11776 );
not U_inv375 ( n75383, P2_P3_EAX_REG_20_ );
dff P2_P3_EAX_REG_21__reg ( clk, reset, P2_P3_EAX_REG_21_, n11781 );
not U_inv376 ( n74921, P2_P3_EAX_REG_21_ );
dff P2_P3_EAX_REG_22__reg ( clk, reset, P2_P3_EAX_REG_22_, n11786 );
not U_inv377 ( n75381, P2_P3_EAX_REG_22_ );
dff P2_P3_EAX_REG_23__reg ( clk, reset, P2_P3_EAX_REG_23_, n11791 );
not U_inv378 ( n74968, P2_P3_EAX_REG_23_ );
dff P2_P3_UWORD_REG_7__reg ( clk, reset, P2_P3_UWORD_REG_7_, n11476 );
not U_inv379 ( n75476, P2_P3_UWORD_REG_7_ );
dff P2_P3_DATAO_REG_23__reg ( clk, reset, P2_P3_DATAO_REG_23_, n11631 );
dff P4_IR_REG_23__reg ( clk, reset, P4_IR_REG_23_, n2141 );
not U_inv380 ( n73496, P4_IR_REG_23_ );
dff P4_WR_REG_reg ( clk, reset, P4_WR_REG, n76451 );
not U_inv381 ( n73025, P4_WR_REG );
dff P4_DATAO_REG_29__reg ( clk, reset, P4_DATAO_REG_29_, n3071 );
not U_inv382 ( n73399, P4_DATAO_REG_29_ );
dff P4_DATAO_REG_28__reg ( clk, reset, P4_DATAO_REG_28_, n3066 );
not U_inv383 ( n73004, P4_DATAO_REG_28_ );
dff P4_DATAO_REG_27__reg ( clk, reset, P4_DATAO_REG_27_, n3061 );
not U_inv384 ( n73409, P4_DATAO_REG_27_ );
dff P4_DATAO_REG_26__reg ( clk, reset, P4_DATAO_REG_26_, n3056 );
not U_inv385 ( n73013, P4_DATAO_REG_26_ );
dff P4_DATAO_REG_25__reg ( clk, reset, P4_DATAO_REG_25_, n3051 );
not U_inv386 ( n75916, P4_DATAO_REG_25_ );
dff P4_DATAO_REG_24__reg ( clk, reset, P4_DATAO_REG_24_, n3046 );
not U_inv387 ( n73417, P4_DATAO_REG_24_ );
dff P4_DATAO_REG_23__reg ( clk, reset, P4_DATAO_REG_23_, n3041 );
not U_inv388 ( n73000, P4_DATAO_REG_23_ );
dff P4_DATAO_REG_22__reg ( clk, reset, P4_DATAO_REG_22_, n3036 );
not U_inv389 ( n73398, P4_DATAO_REG_22_ );
dff P4_DATAO_REG_21__reg ( clk, reset, P4_DATAO_REG_21_, n3031 );
not U_inv390 ( n73006, P4_DATAO_REG_21_ );
dff P4_DATAO_REG_20__reg ( clk, reset, P4_DATAO_REG_20_, n3026 );
not U_inv391 ( n73407, P4_DATAO_REG_20_ );
dff P4_DATAO_REG_19__reg ( clk, reset, P4_DATAO_REG_19_, n3021 );
not U_inv392 ( n73011, P4_DATAO_REG_19_ );
dff P4_DATAO_REG_17__reg ( clk, reset, P4_DATAO_REG_17_, n3011 );
not U_inv393 ( n73408, P4_DATAO_REG_17_ );
dff P4_DATAO_REG_14__reg ( clk, reset, P4_DATAO_REG_14_, n2996 );
not U_inv394 ( n73404, P4_DATAO_REG_14_ );
dff P1_P1_INSTQUEUE_REG_12__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__6_, n8231 );
not U_inv395 ( n74322, P1_P1_INSTQUEUE_REG_12__6_ );
dff P1_P1_EAX_REG_6__reg ( clk, reset, ex_wire71, n9461 );
not U_inv396 ( n74705, ex_wire71 );
dff P1_P1_LWORD_REG_6__reg ( clk, reset, P1_P1_LWORD_REG_6_, n9161 );
not U_inv397 ( n75681, P1_P1_LWORD_REG_6_ );
dff P1_P1_DATAO_REG_6__reg ( clk, reset, P1_P1_DATAO_REG_6_, n9301 );
dff P1_BUF1_REG_6__reg ( clk, reset, P1_BUF1_REG_6_, n151 );
not U_inv398 ( n75460, P1_BUF1_REG_6_ );
dff P1_P2_INSTQUEUE_REG_14__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__6_, n5906 );
not U_inv399 ( n74092, P1_P2_INSTQUEUE_REG_14__6_ );
dff P1_P2_EAX_REG_14__reg ( clk, reset, P1_P2_EAX_REG_14_, n7256 );
not U_inv400 ( n75273, P1_P2_EAX_REG_14_ );
dff P1_P2_EAX_REG_15__reg ( clk, reset, P1_P2_EAX_REG_15_, n7261 );
not U_inv401 ( n74780, P1_P2_EAX_REG_15_ );
dff P1_P2_LWORD_REG_15__reg ( clk, reset, P1_P2_LWORD_REG_15_, n6871 );
not U_inv402 ( n75650, P1_P2_LWORD_REG_15_ );
dff P1_P2_DATAO_REG_15__reg ( clk, reset, P1_P2_DATAO_REG_15_, n7101 );
not U_inv403 ( n75547, P1_P2_DATAO_REG_15_ );
dff P1_BUF1_REG_15__reg ( clk, reset, P1_BUF1_REG_15_, n196 );
not U_inv404 ( n75444, P1_BUF1_REG_15_ );
dff P1_P1_EAX_REG_15__reg ( clk, reset, ex_wire72, n9506 );
not U_inv405 ( n74864, ex_wire72 );
dff P1_P1_EAX_REG_16__reg ( clk, reset, P1_P1_EAX_REG_16_, n9511 );
not U_inv406 ( n74903, P1_P1_EAX_REG_16_ );
dff P1_P1_EAX_REG_17__reg ( clk, reset, ex_wire73, n9516 );
not U_inv407 ( n74909, ex_wire73 );
dff P1_P1_UWORD_REG_1__reg ( clk, reset, P1_P1_UWORD_REG_1_, n9261 );
not U_inv408 ( n75503, P1_P1_UWORD_REG_1_ );
dff P1_P1_DATAO_REG_17__reg ( clk, reset, P1_P1_DATAO_REG_17_, n9356 );
dff P1_BUF1_REG_17__reg ( clk, reset, P1_BUF1_REG_17_, n206 );
not U_inv409 ( n75401, P1_BUF1_REG_17_ );
dff P1_P2_INSTQUEUE_REG_14__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__1_, n5931 );
not U_inv410 ( n73630, P1_P2_INSTQUEUE_REG_14__1_ );
dff P1_P2_REQUESTPENDING_REG_reg ( clk, reset, P1_P2_REQUESTPENDING_REG, n7706 );
not U_inv411 ( n75254, P1_P2_REQUESTPENDING_REG );
dff P1_P2_STATE_REG_0__reg ( clk, reset, P1_P2_STATE_REG_0_, n5676 );
not U_inv412 ( n74691, P1_P2_STATE_REG_0_ );
dff P1_P2_DATAWIDTH_REG_0__reg ( clk, reset, P1_P2_DATAWIDTH_REG_0_, n5681 );
dff P1_P2_DATAWIDTH_REG_31__reg ( clk, reset, ex_wire74, n5836 );
not U_inv413 ( n75137, ex_wire74 );
dff P1_P2_DATAWIDTH_REG_30__reg ( clk, reset, ex_wire75, n5831 );
not U_inv414 ( n73337, ex_wire75 );
dff P1_P2_DATAWIDTH_REG_29__reg ( clk, reset, ex_wire76, n5826 );
not U_inv415 ( n73325, ex_wire76 );
dff P1_P2_DATAWIDTH_REG_28__reg ( clk, reset, ex_wire77, n5821 );
not U_inv416 ( n75081, ex_wire77 );
dff P1_P2_DATAWIDTH_REG_27__reg ( clk, reset, ex_wire78, n5816 );
not U_inv417 ( n73351, ex_wire78 );
dff P1_P2_DATAWIDTH_REG_26__reg ( clk, reset, ex_wire79, n5811 );
not U_inv418 ( n75125, ex_wire79 );
dff P1_P2_DATAWIDTH_REG_25__reg ( clk, reset, ex_wire80, n5806 );
not U_inv419 ( n72974, ex_wire80 );
dff P1_P2_DATAWIDTH_REG_24__reg ( clk, reset, ex_wire81, n5801 );
not U_inv420 ( n75093, ex_wire81 );
dff P1_P2_DATAWIDTH_REG_23__reg ( clk, reset, ex_wire82, n5796 );
not U_inv421 ( n73379, ex_wire82 );
dff P1_P2_DATAWIDTH_REG_22__reg ( clk, reset, ex_wire83, n5791 );
not U_inv422 ( n75161, ex_wire83 );
dff P1_P2_DATAWIDTH_REG_21__reg ( clk, reset, ex_wire84, n5786 );
not U_inv423 ( n73357, ex_wire84 );
dff P1_P2_DATAWIDTH_REG_20__reg ( clk, reset, ex_wire85, n5781 );
not U_inv424 ( n75131, ex_wire85 );
dff P1_P2_DATAWIDTH_REG_19__reg ( clk, reset, ex_wire86, n5776 );
not U_inv425 ( n72996, ex_wire86 );
dff P1_P2_DATAWIDTH_REG_18__reg ( clk, reset, ex_wire87, n5771 );
not U_inv426 ( n75167, ex_wire87 );
dff P1_P2_DATAWIDTH_REG_17__reg ( clk, reset, ex_wire88, n5766 );
not U_inv427 ( n72988, ex_wire88 );
dff P1_P2_DATAWIDTH_REG_16__reg ( clk, reset, ex_wire89, n5761 );
not U_inv428 ( n75143, ex_wire89 );
dff P1_P2_DATAWIDTH_REG_15__reg ( clk, reset, ex_wire90, n5756 );
not U_inv429 ( n72984, ex_wire90 );
dff P1_P2_DATAWIDTH_REG_14__reg ( clk, reset, ex_wire91, n5751 );
not U_inv430 ( n75119, ex_wire91 );
dff P1_P2_DATAWIDTH_REG_13__reg ( clk, reset, ex_wire92, n5746 );
not U_inv431 ( n72973, ex_wire92 );
dff P1_P2_DATAWIDTH_REG_12__reg ( clk, reset, ex_wire93, n5741 );
not U_inv432 ( n75092, ex_wire93 );
dff P1_P2_DATAWIDTH_REG_11__reg ( clk, reset, ex_wire94, n5736 );
not U_inv433 ( n72981, ex_wire94 );
dff P1_P2_DATAWIDTH_REG_10__reg ( clk, reset, ex_wire95, n5731 );
not U_inv434 ( n75102, ex_wire95 );
dff P1_P2_DATAWIDTH_REG_9__reg ( clk, reset, ex_wire96, n5726 );
not U_inv435 ( n72992, ex_wire96 );
dff P1_P2_DATAWIDTH_REG_8__reg ( clk, reset, ex_wire97, n5721 );
not U_inv436 ( n75149, ex_wire97 );
dff P1_P2_DATAWIDTH_REG_7__reg ( clk, reset, ex_wire98, n5716 );
not U_inv437 ( n73343, ex_wire98 );
dff P1_P2_DATAWIDTH_REG_6__reg ( clk, reset, ex_wire99, n5711 );
not U_inv438 ( n75113, ex_wire99 );
dff P1_P2_DATAWIDTH_REG_5__reg ( clk, reset, ex_wire100, n5706 );
not U_inv439 ( n73373, ex_wire100 );
dff P1_P2_DATAWIDTH_REG_4__reg ( clk, reset, ex_wire101, n5701 );
not U_inv440 ( n75155, ex_wire101 );
dff P1_P2_DATAWIDTH_REG_3__reg ( clk, reset, ex_wire102, n5696 );
not U_inv441 ( n73363, ex_wire102 );
dff P1_P2_DATAWIDTH_REG_2__reg ( clk, reset, ex_wire103, n5691 );
not U_inv442 ( n75107, ex_wire103 );
dff P1_P2_DATAWIDTH_REG_1__reg ( clk, reset, P1_P2_DATAWIDTH_REG_1_, n5686 );
dff P1_P2_ADS_N_REG_reg ( clk, reset, P1_P2_ADS_N_REG, n7726 );
dff P1_P2_STATEBS16_REG_reg ( clk, reset, P1_P2_STATEBS16_REG, n7701 );
not U_inv443 ( n74888, P1_P2_STATEBS16_REG );
dff P1_P2_INSTQUEUEWR_ADDR_REG_1__reg ( clk, reset, P1_P2_INSTQUEUEWR_ADDR_REG_1_, n6541 );
not U_inv444 ( n74555, P1_P2_INSTQUEUEWR_ADDR_REG_1_ );
dff P1_P2_INSTQUEUEWR_ADDR_REG_3__reg ( clk, reset, P1_P2_INSTQUEUEWR_ADDR_REG_3_, n6531 );
not U_inv445 ( n73136, P1_P2_INSTQUEUEWR_ADDR_REG_3_ );
dff P1_P2_MEMORYFETCH_REG_reg ( clk, reset, P1_P2_MEMORYFETCH_REG, n7736 );
dff P1_P2_M_IO_N_REG_reg ( clk, reset, P1_P2_M_IO_N_REG, n7716 );
dff P1_P2_READREQUEST_REG_reg ( clk, reset, P1_P2_READREQUEST_REG, n7731 );
dff P1_P2_W_R_N_REG_reg ( clk, reset, P1_P2_W_R_N_REG, n7686 );
dff P1_P2_UWORD_REG_0__reg ( clk, reset, P1_P2_UWORD_REG_0_, n7021 );
not U_inv446 ( n75486, P1_P2_UWORD_REG_0_ );
dff P1_P2_LWORD_REG_0__reg ( clk, reset, P1_P2_LWORD_REG_0_, n6946 );
not U_inv447 ( n75636, P1_P2_LWORD_REG_0_ );
dff P1_P2_LWORD_REG_4__reg ( clk, reset, P1_P2_LWORD_REG_4_, n6926 );
not U_inv448 ( n75647, P1_P2_LWORD_REG_4_ );
dff P1_P2_LWORD_REG_6__reg ( clk, reset, P1_P2_LWORD_REG_6_, n6916 );
not U_inv449 ( n75648, P1_P2_LWORD_REG_6_ );
dff P1_P2_LWORD_REG_7__reg ( clk, reset, P1_P2_LWORD_REG_7_, n6911 );
not U_inv450 ( n75649, P1_P2_LWORD_REG_7_ );
dff P1_P2_DATAO_REG_31__reg ( clk, reset, P1_P2_DATAO_REG_31_, n7181 );
not U_inv451 ( n75428, P1_P2_DATAO_REG_31_ );
dff P1_BUF2_REG_31__reg ( clk, reset, P1_BUF2_REG_31_, n436 );
dff P1_P2_DATAO_REG_16__reg ( clk, reset, P1_P2_DATAO_REG_16_, n7106 );
not U_inv452 ( n75542, P1_P2_DATAO_REG_16_ );
dff P1_BUF2_REG_16__reg ( clk, reset, P1_BUF2_REG_16_, n361 );
not U_inv453 ( n75411, P1_BUF2_REG_16_ );
dff P1_P2_DATAO_REG_7__reg ( clk, reset, P1_P2_DATAO_REG_7_, n7061 );
not U_inv454 ( n75551, P1_P2_DATAO_REG_7_ );
dff P1_BUF2_REG_7__reg ( clk, reset, P1_BUF2_REG_7_, n316 );
not U_inv455 ( n75315, P1_BUF2_REG_7_ );
dff P1_P3_LWORD_REG_7__reg ( clk, reset, P1_P3_LWORD_REG_7_, n4666 );
not U_inv456 ( n75696, P1_P3_LWORD_REG_7_ );
dff P1_P3_DATAO_REG_7__reg ( clk, reset, P1_P3_DATAO_REG_7_, n4816 );
dff P1_P2_DATAO_REG_6__reg ( clk, reset, P1_P2_DATAO_REG_6_, n7056 );
not U_inv457 ( n75548, P1_P2_DATAO_REG_6_ );
dff P1_BUF2_REG_6__reg ( clk, reset, P1_BUF2_REG_6_, n311 );
not U_inv458 ( n75314, P1_BUF2_REG_6_ );
dff P1_P3_LWORD_REG_6__reg ( clk, reset, P1_P3_LWORD_REG_6_, n4671 );
not U_inv459 ( n75695, P1_P3_LWORD_REG_6_ );
dff P1_P3_DATAO_REG_6__reg ( clk, reset, P1_P3_DATAO_REG_6_, n4811 );
dff P1_P2_DATAO_REG_4__reg ( clk, reset, P1_P2_DATAO_REG_4_, n7046 );
not U_inv460 ( n75549, P1_P2_DATAO_REG_4_ );
dff P1_BUF2_REG_4__reg ( clk, reset, P1_BUF2_REG_4_, n301 );
not U_inv461 ( n75313, P1_BUF2_REG_4_ );
dff P1_P3_LWORD_REG_4__reg ( clk, reset, P1_P3_LWORD_REG_4_, n4681 );
not U_inv462 ( n75694, P1_P3_LWORD_REG_4_ );
dff P1_P3_DATAO_REG_4__reg ( clk, reset, P1_P3_DATAO_REG_4_, n4801 );
dff P1_P2_DATAO_REG_1__reg ( clk, reset, P1_P2_DATAO_REG_1_, n7031 );
not U_inv463 ( n75545, P1_P2_DATAO_REG_1_ );
dff P1_BUF2_REG_1__reg ( clk, reset, P1_BUF2_REG_1_, n286 );
not U_inv464 ( n75297, P1_BUF2_REG_1_ );
dff P1_P3_LWORD_REG_1__reg ( clk, reset, P1_P3_LWORD_REG_1_, n4696 );
not U_inv465 ( n75693, P1_P3_LWORD_REG_1_ );
dff P1_P3_DATAO_REG_1__reg ( clk, reset, P1_P3_DATAO_REG_1_, n4786 );
dff P3_IR_REG_1__reg ( clk, reset, P3_IR_REG_1_, n806 );
not U_inv466 ( n73566, P3_IR_REG_1_ );
dff P3_REG3_REG_1__reg ( clk, reset, P3_REG3_REG_1_, n1961 );
not U_inv467 ( n73823, P3_REG3_REG_1_ );
dff P1_P2_LWORD_REG_1__reg ( clk, reset, P1_P2_LWORD_REG_1_, n6941 );
not U_inv468 ( n75646, P1_P2_LWORD_REG_1_ );
dff P1_P2_INSTQUEUE_REG_15__1__reg ( clk, reset, ex_wire104, n5891 );
not U_inv469 ( n73635, ex_wire104 );
dff P1_P2_EAX_REG_24__reg ( clk, reset, P1_P2_EAX_REG_24_, n7306 );
not U_inv470 ( n75344, P1_P2_EAX_REG_24_ );
dff P1_P2_EAX_REG_25__reg ( clk, reset, P1_P2_EAX_REG_25_, n7311 );
not U_inv471 ( n75037, P1_P2_EAX_REG_25_ );
dff P1_P2_UWORD_REG_9__reg ( clk, reset, P1_P2_UWORD_REG_9_, n6976 );
not U_inv472 ( n75571, P1_P2_UWORD_REG_9_ );
dff P1_P2_DATAO_REG_25__reg ( clk, reset, P1_P2_DATAO_REG_25_, n7151 );
not U_inv473 ( n75598, P1_P2_DATAO_REG_25_ );
dff P1_BUF1_REG_25__reg ( clk, reset, P1_BUF1_REG_25_, n246 );
not U_inv474 ( n75393, P1_BUF1_REG_25_ );
dff P1_P1_INSTQUEUE_REG_15__1__reg ( clk, reset, ex_wire105, n8136 );
not U_inv475 ( n73998, ex_wire105 );
dff P1_P1_REQUESTPENDING_REG_reg ( clk, reset, P1_P1_REQUESTPENDING_REG, n9951 );
not U_inv476 ( n75255, P1_P1_REQUESTPENDING_REG );
dff P1_P1_STATE_REG_2__reg ( clk, reset, P1_P1_STATE_REG_2_, n7911 );
not U_inv477 ( n74670, P1_P1_STATE_REG_2_ );
dff P1_P1_STATE_REG_1__reg ( clk, reset, P1_P1_STATE_REG_1_, n7916 );
not U_inv478 ( n73185, P1_P1_STATE_REG_1_ );
dff P1_P1_STATE_REG_0__reg ( clk, reset, P1_P1_STATE_REG_0_, n7921 );
not U_inv479 ( n74713, P1_P1_STATE_REG_0_ );
dff P1_P1_DATAWIDTH_REG_0__reg ( clk, reset, P1_P1_DATAWIDTH_REG_0_, n7926 );
dff P1_P1_DATAWIDTH_REG_31__reg ( clk, reset, ex_wire106, n8081 );
not U_inv480 ( n75139, ex_wire106 );
dff P1_P1_DATAWIDTH_REG_30__reg ( clk, reset, ex_wire107, n8076 );
not U_inv481 ( n73339, ex_wire107 );
dff P1_P1_DATAWIDTH_REG_29__reg ( clk, reset, ex_wire108, n8071 );
not U_inv482 ( n73327, ex_wire108 );
dff P1_P1_DATAWIDTH_REG_28__reg ( clk, reset, ex_wire109, n8066 );
not U_inv483 ( n75083, ex_wire109 );
dff P1_P1_DATAWIDTH_REG_27__reg ( clk, reset, ex_wire110, n8061 );
not U_inv484 ( n73353, ex_wire110 );
dff P1_P1_DATAWIDTH_REG_26__reg ( clk, reset, ex_wire111, n8056 );
not U_inv485 ( n75127, ex_wire111 );
dff P1_P1_DATAWIDTH_REG_25__reg ( clk, reset, ex_wire112, n8051 );
not U_inv486 ( n72978, ex_wire112 );
dff P1_P1_DATAWIDTH_REG_24__reg ( clk, reset, ex_wire113, n8046 );
not U_inv487 ( n75097, ex_wire113 );
dff P1_P1_DATAWIDTH_REG_23__reg ( clk, reset, ex_wire114, n8041 );
not U_inv488 ( n73381, ex_wire114 );
dff P1_P1_DATAWIDTH_REG_22__reg ( clk, reset, ex_wire115, n8036 );
not U_inv489 ( n75163, ex_wire115 );
dff P1_P1_DATAWIDTH_REG_21__reg ( clk, reset, ex_wire116, n8031 );
not U_inv490 ( n73359, ex_wire116 );
dff P1_P1_DATAWIDTH_REG_20__reg ( clk, reset, ex_wire117, n8026 );
not U_inv491 ( n75133, ex_wire117 );
dff P1_P1_DATAWIDTH_REG_19__reg ( clk, reset, ex_wire118, n8021 );
not U_inv492 ( n72998, ex_wire118 );
dff P1_P1_DATAWIDTH_REG_18__reg ( clk, reset, ex_wire119, n8016 );
not U_inv493 ( n75169, ex_wire119 );
dff P1_P1_DATAWIDTH_REG_17__reg ( clk, reset, ex_wire120, n8011 );
not U_inv494 ( n72990, ex_wire120 );
dff P1_P1_DATAWIDTH_REG_16__reg ( clk, reset, ex_wire121, n8006 );
not U_inv495 ( n75145, ex_wire121 );
dff P1_P1_DATAWIDTH_REG_15__reg ( clk, reset, ex_wire122, n8001 );
not U_inv496 ( n72986, ex_wire122 );
dff P1_P1_DATAWIDTH_REG_14__reg ( clk, reset, ex_wire123, n7996 );
not U_inv497 ( n75121, ex_wire123 );
dff P1_P1_DATAWIDTH_REG_13__reg ( clk, reset, ex_wire124, n7991 );
not U_inv498 ( n72977, ex_wire124 );
dff P1_P1_DATAWIDTH_REG_12__reg ( clk, reset, ex_wire125, n7986 );
not U_inv499 ( n75096, ex_wire125 );
dff P1_P1_DATAWIDTH_REG_11__reg ( clk, reset, ex_wire126, n7981 );
not U_inv500 ( n72982, ex_wire126 );
dff P1_P1_DATAWIDTH_REG_10__reg ( clk, reset, ex_wire127, n7976 );
not U_inv501 ( n75103, ex_wire127 );
dff P1_P1_DATAWIDTH_REG_9__reg ( clk, reset, ex_wire128, n7971 );
not U_inv502 ( n72994, ex_wire128 );
dff P1_P1_DATAWIDTH_REG_8__reg ( clk, reset, ex_wire129, n7966 );
not U_inv503 ( n75151, ex_wire129 );
dff P1_P1_DATAWIDTH_REG_7__reg ( clk, reset, ex_wire130, n7961 );
not U_inv504 ( n73345, ex_wire130 );
dff P1_P1_DATAWIDTH_REG_6__reg ( clk, reset, ex_wire131, n7956 );
not U_inv505 ( n75115, ex_wire131 );
dff P1_P1_DATAWIDTH_REG_5__reg ( clk, reset, ex_wire132, n7951 );
not U_inv506 ( n73375, ex_wire132 );
dff P1_P1_DATAWIDTH_REG_4__reg ( clk, reset, ex_wire133, n7946 );
not U_inv507 ( n75157, ex_wire133 );
dff P1_P1_DATAWIDTH_REG_3__reg ( clk, reset, ex_wire134, n7941 );
not U_inv508 ( n73365, ex_wire134 );
dff P1_P1_DATAWIDTH_REG_2__reg ( clk, reset, ex_wire135, n7936 );
not U_inv509 ( n75109, ex_wire135 );
dff P1_P1_DATAWIDTH_REG_1__reg ( clk, reset, P1_P1_DATAWIDTH_REG_1_, n7931 );
dff P1_P1_ADS_N_REG_reg ( clk, reset, P1_P1_ADS_N_REG, n9971 );
dff P2_P1_STATE_REG_2__reg ( clk, reset, P2_P1_STATE_REG_2_, n14646 );
not U_inv510 ( n74650, P2_P1_STATE_REG_2_ );
dff P2_P1_STATE_REG_1__reg ( clk, reset, P2_P1_STATE_REG_1_, n14651 );
not U_inv511 ( n73177, P2_P1_STATE_REG_1_ );
dff P2_P1_STATE_REG_0__reg ( clk, reset, P2_P1_STATE_REG_0_, n14656 );
not U_inv512 ( n74684, P2_P1_STATE_REG_0_ );
dff P2_P1_DATAWIDTH_REG_0__reg ( clk, reset, P2_P1_DATAWIDTH_REG_0_, n14661 );
dff P2_P1_DATAWIDTH_REG_31__reg ( clk, reset, ex_wire136, n14816 );
not U_inv513 ( n75136, ex_wire136 );
dff P2_P1_DATAWIDTH_REG_30__reg ( clk, reset, ex_wire137, n14811 );
not U_inv514 ( n73336, ex_wire137 );
dff P2_P1_DATAWIDTH_REG_29__reg ( clk, reset, ex_wire138, n14806 );
not U_inv515 ( n73324, ex_wire138 );
dff P2_P1_DATAWIDTH_REG_28__reg ( clk, reset, ex_wire139, n14801 );
not U_inv516 ( n75080, ex_wire139 );
dff P2_P1_DATAWIDTH_REG_27__reg ( clk, reset, ex_wire140, n14796 );
not U_inv517 ( n73350, ex_wire140 );
dff P2_P1_DATAWIDTH_REG_26__reg ( clk, reset, ex_wire141, n14791 );
not U_inv518 ( n75124, ex_wire141 );
dff P2_P1_DATAWIDTH_REG_25__reg ( clk, reset, ex_wire142, n14786 );
not U_inv519 ( n72972, ex_wire142 );
dff P2_P1_DATAWIDTH_REG_24__reg ( clk, reset, ex_wire143, n14781 );
not U_inv520 ( n75091, ex_wire143 );
dff P2_P1_DATAWIDTH_REG_23__reg ( clk, reset, ex_wire144, n14776 );
not U_inv521 ( n73378, ex_wire144 );
dff P2_P1_DATAWIDTH_REG_22__reg ( clk, reset, ex_wire145, n14771 );
not U_inv522 ( n75160, ex_wire145 );
dff P2_P1_DATAWIDTH_REG_21__reg ( clk, reset, ex_wire146, n14766 );
not U_inv523 ( n73356, ex_wire146 );
dff P2_P1_DATAWIDTH_REG_20__reg ( clk, reset, ex_wire147, n14761 );
not U_inv524 ( n75130, ex_wire147 );
dff P2_P1_DATAWIDTH_REG_19__reg ( clk, reset, ex_wire148, n14756 );
not U_inv525 ( n72995, ex_wire148 );
dff P2_P1_DATAWIDTH_REG_18__reg ( clk, reset, ex_wire149, n14751 );
not U_inv526 ( n75166, ex_wire149 );
dff P2_P1_DATAWIDTH_REG_17__reg ( clk, reset, ex_wire150, n14746 );
not U_inv527 ( n72987, ex_wire150 );
dff P2_P1_DATAWIDTH_REG_16__reg ( clk, reset, ex_wire151, n14741 );
not U_inv528 ( n75142, ex_wire151 );
dff P2_P1_DATAWIDTH_REG_15__reg ( clk, reset, ex_wire152, n14736 );
not U_inv529 ( n72983, ex_wire152 );
dff P2_P1_DATAWIDTH_REG_14__reg ( clk, reset, ex_wire153, n14731 );
not U_inv530 ( n75118, ex_wire153 );
dff P2_P1_DATAWIDTH_REG_13__reg ( clk, reset, ex_wire154, n14726 );
not U_inv531 ( n72971, ex_wire154 );
dff P2_P1_DATAWIDTH_REG_12__reg ( clk, reset, ex_wire155, n14721 );
not U_inv532 ( n75090, ex_wire155 );
dff P2_P1_DATAWIDTH_REG_11__reg ( clk, reset, ex_wire156, n14716 );
not U_inv533 ( n72980, ex_wire156 );
dff P2_P1_DATAWIDTH_REG_10__reg ( clk, reset, ex_wire157, n14711 );
not U_inv534 ( n75101, ex_wire157 );
dff P2_P1_DATAWIDTH_REG_9__reg ( clk, reset, ex_wire158, n14706 );
not U_inv535 ( n72991, ex_wire158 );
dff P2_P1_DATAWIDTH_REG_8__reg ( clk, reset, ex_wire159, n14701 );
not U_inv536 ( n75148, ex_wire159 );
dff P2_P1_DATAWIDTH_REG_7__reg ( clk, reset, ex_wire160, n14696 );
not U_inv537 ( n73342, ex_wire160 );
dff P2_P1_DATAWIDTH_REG_6__reg ( clk, reset, ex_wire161, n14691 );
not U_inv538 ( n75112, ex_wire161 );
dff P2_P1_DATAWIDTH_REG_5__reg ( clk, reset, ex_wire162, n14686 );
not U_inv539 ( n73372, ex_wire162 );
dff P2_P1_DATAWIDTH_REG_4__reg ( clk, reset, ex_wire163, n14681 );
not U_inv540 ( n75154, ex_wire163 );
dff P2_P1_DATAWIDTH_REG_3__reg ( clk, reset, ex_wire164, n14676 );
not U_inv541 ( n73362, ex_wire164 );
dff P2_P1_DATAWIDTH_REG_2__reg ( clk, reset, ex_wire165, n14671 );
not U_inv542 ( n75106, ex_wire165 );
dff P2_P1_DATAWIDTH_REG_1__reg ( clk, reset, P2_P1_DATAWIDTH_REG_1_, n14666 );
dff P2_P1_ADS_N_REG_reg ( clk, reset, P2_P1_ADS_N_REG, n16706 );
dff P2_P1_STATEBS16_REG_reg ( clk, reset, P2_P1_STATEBS16_REG, n16681 );
not U_inv543 ( n74907, P2_P1_STATEBS16_REG );
dff P2_P1_INSTQUEUEWR_ADDR_REG_1__reg ( clk, reset, P2_P1_INSTQUEUEWR_ADDR_REG_1_, n15521 );
not U_inv544 ( n73140, P2_P1_INSTQUEUEWR_ADDR_REG_1_ );
dff P2_P1_INSTQUEUEWR_ADDR_REG_3__reg ( clk, reset, P2_P1_INSTQUEUEWR_ADDR_REG_3_, n15511 );
not U_inv545 ( n74525, P2_P1_INSTQUEUEWR_ADDR_REG_3_ );
dff P2_P1_INSTQUEUE_REG_3__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__7_, n15321 );
not U_inv546 ( n74130, P2_P1_INSTQUEUE_REG_3__7_ );
dff P2_P1_INSTQUEUE_REG_9__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__7_, n15081 );
not U_inv547 ( n74158, P2_P1_INSTQUEUE_REG_9__7_ );
dff P2_P1_INSTQUEUE_REG_8__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__7_, n15121 );
not U_inv548 ( n74145, P2_P1_INSTQUEUE_REG_8__7_ );
dff P2_P1_INSTQUEUE_REG_12__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__7_, n14961 );
not U_inv549 ( n74133, P2_P1_INSTQUEUE_REG_12__7_ );
dff P2_P1_INSTQUEUE_REG_10__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__7_, n15041 );
not U_inv550 ( n74160, P2_P1_INSTQUEUE_REG_10__7_ );
dff P2_P1_INSTQUEUE_REG_1__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__7_, n15401 );
not U_inv551 ( n74135, P2_P1_INSTQUEUE_REG_1__7_ );
dff P2_P1_INSTQUEUE_REG_0__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__7_, n15441 );
not U_inv552 ( n74106, P2_P1_INSTQUEUE_REG_0__7_ );
dff P2_P1_INSTQUEUE_REG_4__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__7_, n15281 );
not U_inv553 ( n74138, P2_P1_INSTQUEUE_REG_4__7_ );
dff P2_P1_INSTQUEUE_REG_5__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__7_, n15241 );
not U_inv554 ( n74151, P2_P1_INSTQUEUE_REG_5__7_ );
dff P2_P1_INSTQUEUE_REG_2__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__7_, n15361 );
not U_inv555 ( n74141, P2_P1_INSTQUEUE_REG_2__7_ );
dff P2_P1_INSTQUEUE_REG_6__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__7_, n15201 );
not U_inv556 ( n74159, P2_P1_INSTQUEUE_REG_6__7_ );
dff P2_P1_INSTQUEUE_REG_11__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__7_, n15001 );
not U_inv557 ( n74148, P2_P1_INSTQUEUE_REG_11__7_ );
dff P2_P1_INSTQUEUE_REG_7__7__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__7_, n15161 );
not U_inv558 ( n74146, P2_P1_INSTQUEUE_REG_7__7_ );
dff P2_P1_DATAO_REG_31__reg ( clk, reset, P2_P1_DATAO_REG_31_, n16161 );
dff P2_P1_DATAO_REG_1__reg ( clk, reset, P2_P1_DATAO_REG_1_, n16011 );
dff P2_BUF1_REG_1__reg ( clk, reset, P2_BUF1_REG_1_, n466 );
not U_inv559 ( n75453, P2_BUF1_REG_1_ );
dff P2_P2_INSTQUEUE_REG_15__1__reg ( clk, reset, ex_wire166, n12626 );
not U_inv560 ( n73634, ex_wire166 );
dff P2_P2_REQUESTPENDING_REG_reg ( clk, reset, P2_P2_REQUESTPENDING_REG, n14441 );
not U_inv561 ( n75228, P2_P2_REQUESTPENDING_REG );
dff P2_P2_STATE_REG_2__reg ( clk, reset, P2_P2_STATE_REG_2_, n12401 );
not U_inv562 ( n74636, P2_P2_STATE_REG_2_ );
dff P2_P2_STATE_REG_0__reg ( clk, reset, P2_P2_STATE_REG_0_, n12411 );
not U_inv563 ( n74683, P2_P2_STATE_REG_0_ );
dff P2_P2_STATE_REG_1__reg ( clk, reset, P2_P2_STATE_REG_1_, n12406 );
not U_inv564 ( n73184, P2_P2_STATE_REG_1_ );
dff P2_P2_ADS_N_REG_reg ( clk, reset, P2_P2_ADS_N_REG, n14461 );
dff P2_P2_DATAWIDTH_REG_0__reg ( clk, reset, P2_P2_DATAWIDTH_REG_0_, n12416 );
dff P2_P2_STATEBS16_REG_reg ( clk, reset, P2_P2_STATEBS16_REG, n14436 );
not U_inv565 ( n74890, P2_P2_STATEBS16_REG );
dff P2_P2_INSTQUEUEWR_ADDR_REG_1__reg ( clk, reset, P2_P2_INSTQUEUEWR_ADDR_REG_1_, n13276 );
not U_inv566 ( n74556, P2_P2_INSTQUEUEWR_ADDR_REG_1_ );
dff P2_P2_INSTQUEUEWR_ADDR_REG_3__reg ( clk, reset, P2_P2_INSTQUEUEWR_ADDR_REG_3_, n13266 );
not U_inv567 ( n73137, P2_P2_INSTQUEUEWR_ADDR_REG_3_ );
dff P2_P2_MEMORYFETCH_REG_reg ( clk, reset, P2_P2_MEMORYFETCH_REG, n14471 );
dff P2_P2_READREQUEST_REG_reg ( clk, reset, P2_P2_READREQUEST_REG, n14466 );
dff P2_P2_UWORD_REG_0__reg ( clk, reset, P2_P2_UWORD_REG_0_, n13756 );
not U_inv568 ( n75475, P2_P2_UWORD_REG_0_ );
dff P2_P2_LWORD_REG_0__reg ( clk, reset, P2_P2_LWORD_REG_0_, n13681 );
not U_inv569 ( n75604, P2_P2_LWORD_REG_0_ );
dff P2_P2_LWORD_REG_1__reg ( clk, reset, P2_P2_LWORD_REG_1_, n13676 );
not U_inv570 ( n75606, P2_P2_LWORD_REG_1_ );
dff P2_P2_LWORD_REG_4__reg ( clk, reset, P2_P2_LWORD_REG_4_, n13661 );
not U_inv571 ( n75628, P2_P2_LWORD_REG_4_ );
dff P2_P2_LWORD_REG_7__reg ( clk, reset, P2_P2_LWORD_REG_7_, n13646 );
not U_inv572 ( n75630, P2_P2_LWORD_REG_7_ );
dff P2_P2_DATAO_REG_31__reg ( clk, reset, P2_P2_DATAO_REG_31_, n13916 );
not U_inv573 ( n75427, P2_P2_DATAO_REG_31_ );
dff P2_BUF1_REG_31__reg ( clk, reset, P2_BUF1_REG_31_, n616 );
not U_inv574 ( n75445, P2_BUF1_REG_31_ );
dff P2_BUF2_REG_31__reg ( clk, reset, P2_BUF2_REG_31_, n776 );
dff P2_P2_INSTQUEUE_REG_5__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__7_, n12996 );
not U_inv575 ( n74207, P2_P2_INSTQUEUE_REG_5__7_ );
dff P2_P2_INSTQUEUE_REG_6__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__7_, n12956 );
not U_inv576 ( n74213, P2_P2_INSTQUEUE_REG_6__7_ );
dff P2_P2_INSTQUEUE_REG_7__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__7_, n12916 );
not U_inv577 ( n74197, P2_P2_INSTQUEUE_REG_7__7_ );
dff P2_P2_INSTQUEUE_REG_8__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__7_, n12876 );
not U_inv578 ( n74194, P2_P2_INSTQUEUE_REG_8__7_ );
dff P2_P2_INSTQUEUE_REG_9__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__7_, n12836 );
not U_inv579 ( n74210, P2_P2_INSTQUEUE_REG_9__7_ );
dff P2_P2_INSTQUEUE_REG_10__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__7_, n12796 );
not U_inv580 ( n74216, P2_P2_INSTQUEUE_REG_10__7_ );
dff P2_P2_INSTQUEUE_REG_11__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__7_, n12756 );
not U_inv581 ( n74204, P2_P2_INSTQUEUE_REG_11__7_ );
dff P2_P2_INSTQUEUE_REG_12__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__7_, n12716 );
not U_inv582 ( n74176, P2_P2_INSTQUEUE_REG_12__7_ );
dff P2_P2_INSTQUEUE_REG_13__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__7_, n12676 );
not U_inv583 ( n74191, P2_P2_INSTQUEUE_REG_13__7_ );
dff P2_P2_INSTQUEUE_REG_0__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__7_, n13196 );
not U_inv584 ( n74169, P2_P2_INSTQUEUE_REG_0__7_ );
dff P2_P2_INSTQUEUE_REG_1__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__7_, n13156 );
not U_inv585 ( n74183, P2_P2_INSTQUEUE_REG_1__7_ );
dff P2_P2_INSTQUEUE_REG_2__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__7_, n13116 );
not U_inv586 ( n74188, P2_P2_INSTQUEUE_REG_2__7_ );
dff P2_P2_INSTQUEUE_REG_3__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__7_, n13076 );
not U_inv587 ( n74173, P2_P2_INSTQUEUE_REG_3__7_ );
dff P2_P2_INSTQUEUE_REG_4__7__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__7_, n13036 );
not U_inv588 ( n74185, P2_P2_INSTQUEUE_REG_4__7_ );
dff P2_P2_DATAO_REG_16__reg ( clk, reset, P2_P2_DATAO_REG_16_, n13841 );
not U_inv589 ( n75516, P2_P2_DATAO_REG_16_ );
dff P2_BUF2_REG_16__reg ( clk, reset, P2_BUF2_REG_16_, n701 );
not U_inv590 ( n75412, P2_BUF2_REG_16_ );
dff P2_P2_DATAO_REG_7__reg ( clk, reset, P2_P2_DATAO_REG_7_, n13796 );
not U_inv591 ( n75504, P2_P2_DATAO_REG_7_ );
dff P2_BUF2_REG_7__reg ( clk, reset, P2_BUF2_REG_7_, n656 );
not U_inv592 ( n75294, P2_BUF2_REG_7_ );
dff P2_P3_LWORD_REG_7__reg ( clk, reset, P2_P3_LWORD_REG_7_, n11401 );
not U_inv593 ( n75629, P2_P3_LWORD_REG_7_ );
dff P2_P3_DATAO_REG_7__reg ( clk, reset, P2_P3_DATAO_REG_7_, n11551 );
dff P2_P2_DATAO_REG_4__reg ( clk, reset, P2_P2_DATAO_REG_4_, n13781 );
not U_inv594 ( n75524, P2_P2_DATAO_REG_4_ );
dff P2_BUF2_REG_4__reg ( clk, reset, P2_BUF2_REG_4_, n641 );
not U_inv595 ( n75293, P2_BUF2_REG_4_ );
dff P2_P3_UWORD_REG_4__reg ( clk, reset, P2_P3_UWORD_REG_4_, n11491 );
not U_inv596 ( n75474, P2_P3_UWORD_REG_4_ );
dff P2_P3_DATAO_REG_20__reg ( clk, reset, P2_P3_DATAO_REG_20_, n11616 );
dff P2_P3_LWORD_REG_4__reg ( clk, reset, P2_P3_LWORD_REG_4_, n11416 );
not U_inv597 ( n75627, P2_P3_LWORD_REG_4_ );
dff P2_P3_DATAO_REG_4__reg ( clk, reset, P2_P3_DATAO_REG_4_, n11536 );
dff P2_P2_DATAO_REG_2__reg ( clk, reset, P2_P2_DATAO_REG_2_, n13771 );
not U_inv598 ( n75515, P2_P2_DATAO_REG_2_ );
dff P2_BUF2_REG_2__reg ( clk, reset, P2_BUF2_REG_2_, n631 );
not U_inv599 ( n75292, P2_BUF2_REG_2_ );
dff P2_P3_UWORD_REG_2__reg ( clk, reset, P2_P3_UWORD_REG_2_, n11501 );
not U_inv600 ( n75473, P2_P3_UWORD_REG_2_ );
dff P2_P3_DATAO_REG_18__reg ( clk, reset, P2_P3_DATAO_REG_18_, n11606 );
dff P2_P3_LWORD_REG_2__reg ( clk, reset, P2_P3_LWORD_REG_2_, n11426 );
not U_inv601 ( n75625, P2_P3_LWORD_REG_2_ );
dff P2_P3_DATAO_REG_2__reg ( clk, reset, P2_P3_DATAO_REG_2_, n11526 );
dff P2_P2_LWORD_REG_2__reg ( clk, reset, P2_P2_LWORD_REG_2_, n13671 );
not U_inv602 ( n75626, P2_P2_LWORD_REG_2_ );
dff P2_P2_INSTQUEUE_REG_15__2__reg ( clk, reset, ex_wire167, n12621 );
not U_inv603 ( n73747, ex_wire167 );
dff P2_P2_EAX_REG_18__reg ( clk, reset, P2_P2_EAX_REG_18_, n14011 );
not U_inv604 ( n75379, P2_P2_EAX_REG_18_ );
dff P2_P2_UWORD_REG_2__reg ( clk, reset, P2_P2_UWORD_REG_2_, n13746 );
not U_inv605 ( n75472, P2_P2_UWORD_REG_2_ );
dff P2_P2_DATAO_REG_18__reg ( clk, reset, P2_P2_DATAO_REG_18_, n13851 );
not U_inv606 ( n75511, P2_P2_DATAO_REG_18_ );
dff P2_BUF2_REG_18__reg ( clk, reset, P2_BUF2_REG_18_, n711 );
not U_inv607 ( n75359, P2_BUF2_REG_18_ );
dff P2_P2_EAX_REG_19__reg ( clk, reset, P2_P2_EAX_REG_19_, n14016 );
not U_inv608 ( n74877, P2_P2_EAX_REG_19_ );
dff P2_P2_UWORD_REG_3__reg ( clk, reset, P2_P2_UWORD_REG_3_, n13741 );
not U_inv609 ( n75471, P2_P2_UWORD_REG_3_ );
dff P2_P2_DATAO_REG_19__reg ( clk, reset, P2_P2_DATAO_REG_19_, n13856 );
not U_inv610 ( n75507, P2_P2_DATAO_REG_19_ );
dff P2_BUF2_REG_19__reg ( clk, reset, P2_BUF2_REG_19_, n716 );
not U_inv611 ( n75358, P2_BUF2_REG_19_ );
dff P2_P2_INSTQUEUE_REG_14__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__3_, n12656 );
not U_inv612 ( n73781, P2_P2_INSTQUEUE_REG_14__3_ );
dff P2_P2_EAX_REG_11__reg ( clk, reset, P2_P2_EAX_REG_11_, n13976 );
not U_inv613 ( n74678, P2_P2_EAX_REG_11_ );
dff P2_P2_EAX_REG_12__reg ( clk, reset, P2_P2_EAX_REG_12_, n13981 );
not U_inv614 ( n75264, P2_P2_EAX_REG_12_ );
dff P2_P2_EAX_REG_13__reg ( clk, reset, P2_P2_EAX_REG_13_, n13986 );
not U_inv615 ( n74732, P2_P2_EAX_REG_13_ );
dff P2_P2_EAX_REG_14__reg ( clk, reset, P2_P2_EAX_REG_14_, n13991 );
not U_inv616 ( n75266, P2_P2_EAX_REG_14_ );
dff P2_P2_LWORD_REG_14__reg ( clk, reset, P2_P2_LWORD_REG_14_, n13611 );
not U_inv617 ( n75624, P2_P2_LWORD_REG_14_ );
dff P2_P2_DATAO_REG_14__reg ( clk, reset, P2_P2_DATAO_REG_14_, n13831 );
not U_inv618 ( n75505, P2_P2_DATAO_REG_14_ );
dff P2_BUF2_REG_14__reg ( clk, reset, P2_BUF2_REG_14_, n691 );
not U_inv619 ( n75304, P2_BUF2_REG_14_ );
dff P2_P2_UWORD_REG_14__reg ( clk, reset, P2_P2_UWORD_REG_14_, n13686 );
not U_inv620 ( n75564, P2_P2_UWORD_REG_14_ );
dff P2_P2_DATAO_REG_30__reg ( clk, reset, P2_P2_DATAO_REG_30_, n13911 );
not U_inv621 ( n73427, P2_P2_DATAO_REG_30_ );
dff P2_BUF2_REG_30__reg ( clk, reset, P2_BUF2_REG_30_, n771 );
not U_inv622 ( n75336, P2_BUF2_REG_30_ );
dff P2_P2_INSTQUEUE_REG_4__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__6_, n13041 );
not U_inv623 ( n74069, P2_P2_INSTQUEUE_REG_4__6_ );
dff P2_P2_EAX_REG_22__reg ( clk, reset, P2_P2_EAX_REG_22_, n14031 );
not U_inv624 ( n75377, P2_P2_EAX_REG_22_ );
dff P2_P2_EAX_REG_23__reg ( clk, reset, P2_P2_EAX_REG_23_, n14036 );
not U_inv625 ( n74971, P2_P2_EAX_REG_23_ );
dff P2_P2_EAX_REG_24__reg ( clk, reset, P2_P2_EAX_REG_24_, n14041 );
not U_inv626 ( n75342, P2_P2_EAX_REG_24_ );
dff P2_P2_EAX_REG_25__reg ( clk, reset, P2_P2_EAX_REG_25_, n14046 );
not U_inv627 ( n75036, P2_P2_EAX_REG_25_ );
dff P2_P2_UWORD_REG_9__reg ( clk, reset, P2_P2_UWORD_REG_9_, n13711 );
not U_inv628 ( n75563, P2_P2_UWORD_REG_9_ );
dff P2_P2_DATAO_REG_25__reg ( clk, reset, P2_P2_DATAO_REG_25_, n13886 );
not U_inv629 ( n75592, P2_P2_DATAO_REG_25_ );
dff P2_BUF2_REG_25__reg ( clk, reset, P2_BUF2_REG_25_, n746 );
not U_inv630 ( n75340, P2_BUF2_REG_25_ );
dff P2_P2_INSTQUEUE_REG_4__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__1_, n13066 );
not U_inv631 ( n73597, P2_P2_INSTQUEUE_REG_4__1_ );
dff P2_P2_EAX_REG_26__reg ( clk, reset, P2_P2_EAX_REG_26_, n14051 );
not U_inv632 ( n75343, P2_P2_EAX_REG_26_ );
dff P2_P2_EAX_REG_27__reg ( clk, reset, P2_P2_EAX_REG_27_, n14056 );
not U_inv633 ( n75322, P2_P2_EAX_REG_27_ );
dff P2_P2_EAX_REG_28__reg ( clk, reset, P2_P2_EAX_REG_28_, n14061 );
not U_inv634 ( n73393, P2_P2_EAX_REG_28_ );
dff P2_P2_EAX_REG_29__reg ( clk, reset, P2_P2_EAX_REG_29_, n14066 );
not U_inv635 ( n75203, P2_P2_EAX_REG_29_ );
dff P2_P2_UWORD_REG_13__reg ( clk, reset, P2_P2_UWORD_REG_13_, n13691 );
not U_inv636 ( n75562, P2_P2_UWORD_REG_13_ );
dff P2_P2_DATAO_REG_29__reg ( clk, reset, P2_P2_DATAO_REG_29_, n13906 );
not U_inv637 ( n75590, P2_P2_DATAO_REG_29_ );
dff P2_BUF2_REG_29__reg ( clk, reset, P2_BUF2_REG_29_, n766 );
not U_inv638 ( n75337, P2_BUF2_REG_29_ );
dff P2_P2_INSTQUEUE_REG_15__5__reg ( clk, reset, ex_wire168, n12606 );
not U_inv639 ( n73909, ex_wire168 );
dff P2_P2_EAX_REG_20__reg ( clk, reset, P2_P2_EAX_REG_20_, n14021 );
not U_inv640 ( n75378, P2_P2_EAX_REG_20_ );
dff P2_P2_UWORD_REG_4__reg ( clk, reset, P2_P2_UWORD_REG_4_, n13736 );
not U_inv641 ( n75470, P2_P2_UWORD_REG_4_ );
dff P2_P2_DATAO_REG_20__reg ( clk, reset, P2_P2_DATAO_REG_20_, n13861 );
not U_inv642 ( n75508, P2_P2_DATAO_REG_20_ );
dff P2_BUF2_REG_20__reg ( clk, reset, P2_BUF2_REG_20_, n721 );
not U_inv643 ( n75357, P2_BUF2_REG_20_ );
dff P2_P2_EAX_REG_21__reg ( clk, reset, P2_P2_EAX_REG_21_, n14026 );
not U_inv644 ( n74922, P2_P2_EAX_REG_21_ );
dff P2_P2_UWORD_REG_5__reg ( clk, reset, P2_P2_UWORD_REG_5_, n13731 );
not U_inv645 ( n75469, P2_P2_UWORD_REG_5_ );
dff P2_P2_DATAO_REG_21__reg ( clk, reset, P2_P2_DATAO_REG_21_, n13866 );
not U_inv646 ( n75522, P2_P2_DATAO_REG_21_ );
dff P2_BUF1_REG_21__reg ( clk, reset, P2_BUF1_REG_21_, n566 );
not U_inv647 ( n75375, P2_BUF1_REG_21_ );
dff P2_P1_INSTQUEUE_REG_15__5__reg ( clk, reset, ex_wire169, n14851 );
not U_inv648 ( n73882, ex_wire169 );
dff P2_P1_EAX_REG_0__reg ( clk, reset, P2_P1_EAX_REG_0_, n16166 );
not U_inv649 ( n73161, P2_P1_EAX_REG_0_ );
dff P2_P1_EAX_REG_1__reg ( clk, reset, ex_wire170, n16171 );
not U_inv650 ( n74609, ex_wire170 );
dff P2_P1_EAX_REG_2__reg ( clk, reset, P2_P1_EAX_REG_2_, n16176 );
not U_inv651 ( n73165, P2_P1_EAX_REG_2_ );
dff P2_P1_EAX_REG_3__reg ( clk, reset, ex_wire171, n16181 );
not U_inv652 ( n74631, ex_wire171 );
dff P2_P1_LWORD_REG_3__reg ( clk, reset, P2_P1_LWORD_REG_3_, n15911 );
not U_inv653 ( n75664, P2_P1_LWORD_REG_3_ );
dff P2_P1_DATAO_REG_3__reg ( clk, reset, P2_P1_DATAO_REG_3_, n16021 );
dff P2_BUF1_REG_3__reg ( clk, reset, P2_BUF1_REG_3_, n476 );
not U_inv654 ( n75452, P2_BUF1_REG_3_ );
dff P2_P1_INSTQUEUE_REG_12__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__3_, n14981 );
not U_inv655 ( n73638, P2_P1_INSTQUEUE_REG_12__3_ );
dff P2_P1_EAX_REG_6__reg ( clk, reset, ex_wire172, n16196 );
not U_inv656 ( n74704, ex_wire172 );
dff P2_P1_LWORD_REG_6__reg ( clk, reset, P2_P1_LWORD_REG_6_, n15896 );
not U_inv657 ( n75663, P2_P1_LWORD_REG_6_ );
dff P2_P1_DATAO_REG_6__reg ( clk, reset, P2_P1_DATAO_REG_6_, n16036 );
dff P2_BUF1_REG_6__reg ( clk, reset, P2_BUF1_REG_6_, n491 );
not U_inv658 ( n75451, P2_BUF1_REG_6_ );
dff P2_P2_UWORD_REG_6__reg ( clk, reset, P2_P2_UWORD_REG_6_, n13726 );
not U_inv659 ( n75468, P2_P2_UWORD_REG_6_ );
dff P2_P2_DATAO_REG_22__reg ( clk, reset, P2_P2_DATAO_REG_22_, n13871 );
not U_inv660 ( n75519, P2_P2_DATAO_REG_22_ );
dff P2_BUF1_REG_22__reg ( clk, reset, P2_BUF1_REG_22_, n571 );
not U_inv661 ( n75374, P2_BUF1_REG_22_ );
dff P2_P1_INSTQUEUE_REG_0__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__6_, n15446 );
not U_inv662 ( n73950, P2_P1_INSTQUEUE_REG_0__6_ );
dff P2_P1_INSTQUEUE_REG_1__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__6_, n15406 );
not U_inv663 ( n73970, P2_P1_INSTQUEUE_REG_1__6_ );
dff P2_P1_INSTQUEUE_REG_2__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__6_, n15366 );
not U_inv664 ( n73974, P2_P1_INSTQUEUE_REG_2__6_ );
dff P2_P1_INSTQUEUE_REG_3__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__6_, n15326 );
not U_inv665 ( n73967, P2_P1_INSTQUEUE_REG_3__6_ );
dff P2_P1_INSTQUEUE_REG_4__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__6_, n15286 );
not U_inv666 ( n73971, P2_P1_INSTQUEUE_REG_4__6_ );
dff P2_P1_INSTQUEUE_REG_5__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__6_, n15246 );
not U_inv667 ( n73990, P2_P1_INSTQUEUE_REG_5__6_ );
dff P2_P1_INSTQUEUE_REG_6__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__6_, n15206 );
not U_inv668 ( n73994, P2_P1_INSTQUEUE_REG_6__6_ );
dff P2_P1_INSTQUEUE_REG_7__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__6_, n15166 );
not U_inv669 ( n73975, P2_P1_INSTQUEUE_REG_7__6_ );
dff P2_P1_INSTQUEUE_REG_8__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__6_, n15126 );
not U_inv670 ( n73973, P2_P1_INSTQUEUE_REG_8__6_ );
dff P2_P1_INSTQUEUE_REG_9__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__6_, n15086 );
not U_inv671 ( n73993, P2_P1_INSTQUEUE_REG_9__6_ );
dff P2_P1_INSTQUEUE_REG_10__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__6_, n15046 );
not U_inv672 ( n73996, P2_P1_INSTQUEUE_REG_10__6_ );
dff P2_P1_INSTQUEUE_REG_11__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__6_, n15006 );
not U_inv673 ( n73977, P2_P1_INSTQUEUE_REG_11__6_ );
dff P2_P1_INSTQUEUE_REG_12__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__6_, n14966 );
not U_inv674 ( n73966, P2_P1_INSTQUEUE_REG_12__6_ );
dff P2_P1_INSTQUEUE_REG_13__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__6_, n14926 );
not U_inv675 ( n73972, P2_P1_INSTQUEUE_REG_13__6_ );
dff P2_P1_INSTQUEUE_REG_14__6__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__6_, n14886 );
not U_inv676 ( n73976, P2_P1_INSTQUEUE_REG_14__6_ );
dff P2_P1_EAX_REG_14__reg ( clk, reset, P2_P1_EAX_REG_14_, n16236 );
not U_inv677 ( n73251, P2_P1_EAX_REG_14_ );
dff P2_P1_EAX_REG_16__reg ( clk, reset, P2_P1_EAX_REG_16_, n16246 );
not U_inv678 ( n74902, P2_P1_EAX_REG_16_ );
dff P2_P1_EAX_REG_17__reg ( clk, reset, ex_wire173, n16251 );
not U_inv679 ( n74908, ex_wire173 );
dff P2_P1_UWORD_REG_1__reg ( clk, reset, P2_P1_UWORD_REG_1_, n15996 );
not U_inv680 ( n75494, P2_P1_UWORD_REG_1_ );
dff P2_P1_DATAO_REG_17__reg ( clk, reset, P2_P1_DATAO_REG_17_, n16091 );
dff P2_BUF1_REG_17__reg ( clk, reset, P2_BUF1_REG_17_, n546 );
not U_inv681 ( n75373, P2_BUF1_REG_17_ );
dff P2_P1_INSTQUEUE_REG_15__1__reg ( clk, reset, ex_wire174, n14871 );
not U_inv682 ( n73552, ex_wire174 );
dff P2_P1_INSTQUEUE_REG_14__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__1_, n14911 );
not U_inv683 ( n73549, P2_P1_INSTQUEUE_REG_14__1_ );
dff P2_P1_EAX_REG_9__reg ( clk, reset, ex_wire175, n16211 );
not U_inv684 ( n74757, ex_wire175 );
dff P2_P1_LWORD_REG_9__reg ( clk, reset, P2_P1_LWORD_REG_9_, n15881 );
not U_inv685 ( n75662, P2_P1_LWORD_REG_9_ );
dff P2_P1_DATAO_REG_9__reg ( clk, reset, P2_P1_DATAO_REG_9_, n16051 );
dff P2_BUF1_REG_9__reg ( clk, reset, P2_BUF1_REG_9_, n506 );
not U_inv686 ( n75435, P2_BUF1_REG_9_ );
dff P2_P1_UWORD_REG_9__reg ( clk, reset, P2_P1_UWORD_REG_9_, n15956 );
not U_inv687 ( n75579, P2_P1_UWORD_REG_9_ );
dff P2_P1_DATAO_REG_25__reg ( clk, reset, P2_P1_DATAO_REG_25_, n16131 );
dff P2_BUF1_REG_25__reg ( clk, reset, P2_BUF1_REG_25_, n586 );
not U_inv688 ( n75368, P2_BUF1_REG_25_ );
dff P2_P1_INSTQUEUE_REG_0__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__1_, n15471 );
not U_inv689 ( n73534, P2_P1_INSTQUEUE_REG_0__1_ );
dff P2_P1_INSTQUEUE_REG_1__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__1_, n15431 );
not U_inv690 ( n73537, P2_P1_INSTQUEUE_REG_1__1_ );
dff P2_P1_INSTQUEUE_REG_2__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__1_, n15391 );
not U_inv691 ( n73545, P2_P1_INSTQUEUE_REG_2__1_ );
dff P2_P1_INSTQUEUE_REG_3__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__1_, n15351 );
not U_inv692 ( n73539, P2_P1_INSTQUEUE_REG_3__1_ );
dff P2_P1_INSTQUEUE_REG_4__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__1_, n15311 );
not U_inv693 ( n73536, P2_P1_INSTQUEUE_REG_4__1_ );
dff P2_P1_INSTQUEUE_REG_5__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__1_, n15271 );
not U_inv694 ( n73540, P2_P1_INSTQUEUE_REG_5__1_ );
dff P2_P1_INSTQUEUE_REG_6__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__1_, n15231 );
not U_inv695 ( n73547, P2_P1_INSTQUEUE_REG_6__1_ );
dff P2_P1_INSTQUEUE_REG_7__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__1_, n15191 );
not U_inv696 ( n73542, P2_P1_INSTQUEUE_REG_7__1_ );
dff P2_P1_INSTQUEUE_REG_8__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__1_, n15151 );
not U_inv697 ( n73541, P2_P1_INSTQUEUE_REG_8__1_ );
dff P2_P1_INSTQUEUE_REG_9__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__1_, n15111 );
not U_inv698 ( n73546, P2_P1_INSTQUEUE_REG_9__1_ );
dff P2_P1_INSTQUEUE_REG_10__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__1_, n15071 );
not U_inv699 ( n73550, P2_P1_INSTQUEUE_REG_10__1_ );
dff P2_P1_INSTQUEUE_REG_11__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__1_, n15031 );
not U_inv700 ( n73548, P2_P1_INSTQUEUE_REG_11__1_ );
dff P2_P1_INSTQUEUE_REG_12__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__1_, n14991 );
not U_inv701 ( n73538, P2_P1_INSTQUEUE_REG_12__1_ );
dff P2_P1_INSTQUEUE_REG_13__1__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__1_, n14951 );
not U_inv702 ( n73543, P2_P1_INSTQUEUE_REG_13__1_ );
dff P2_P1_EAX_REG_24__reg ( clk, reset, P2_P1_EAX_REG_24_, n16286 );
not U_inv703 ( n73306, P2_P1_EAX_REG_24_ );
dff P2_P1_UWORD_REG_8__reg ( clk, reset, P2_P1_UWORD_REG_8_, n15961 );
not U_inv704 ( n75578, P2_P1_UWORD_REG_8_ );
dff P2_P1_DATAO_REG_24__reg ( clk, reset, P2_P1_DATAO_REG_24_, n16126 );
dff P2_BUF1_REG_24__reg ( clk, reset, P2_BUF1_REG_24_, n581 );
not U_inv705 ( n75409, P2_BUF1_REG_24_ );
dff P2_P1_INSTQUEUE_REG_15__0__reg ( clk, reset, ex_wire176, n14876 );
not U_inv706 ( n73556, ex_wire176 );
dff P2_P1_UWORD_REG_0__reg ( clk, reset, P2_P1_UWORD_REG_0_, n16001 );
not U_inv707 ( n75493, P2_P1_UWORD_REG_0_ );
dff P2_P1_DATAO_REG_16__reg ( clk, reset, P2_P1_DATAO_REG_16_, n16086 );
dff P2_BUF1_REG_16__reg ( clk, reset, P2_BUF1_REG_16_, n541 );
not U_inv708 ( n75372, P2_BUF1_REG_16_ );
dff P2_P1_INSTQUEUE_REG_0__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__0_, n15476 );
not U_inv709 ( n73553, P2_P1_INSTQUEUE_REG_0__0_ );
dff P2_P1_INSTQUEUE_REG_1__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__0_, n15436 );
not U_inv710 ( n73557, P2_P1_INSTQUEUE_REG_1__0_ );
dff P2_P1_INSTQUEUE_REG_2__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__0_, n15396 );
not U_inv711 ( n73562, P2_P1_INSTQUEUE_REG_2__0_ );
dff P2_P1_INSTQUEUE_REG_3__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__0_, n15356 );
not U_inv712 ( n73555, P2_P1_INSTQUEUE_REG_3__0_ );
dff P2_P1_INSTQUEUE_REG_4__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__0_, n15316 );
not U_inv713 ( n73559, P2_P1_INSTQUEUE_REG_4__0_ );
dff P2_P1_INSTQUEUE_REG_5__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__0_, n15276 );
not U_inv714 ( n73570, P2_P1_INSTQUEUE_REG_5__0_ );
dff P2_P1_INSTQUEUE_REG_6__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__0_, n15236 );
not U_inv715 ( n73572, P2_P1_INSTQUEUE_REG_6__0_ );
dff P2_P1_INSTQUEUE_REG_7__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__0_, n15196 );
not U_inv716 ( n73563, P2_P1_INSTQUEUE_REG_7__0_ );
dff P2_P1_INSTQUEUE_REG_8__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__0_, n15156 );
not U_inv717 ( n73561, P2_P1_INSTQUEUE_REG_8__0_ );
dff P2_P1_INSTQUEUE_REG_9__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__0_, n15116 );
not U_inv718 ( n73571, P2_P1_INSTQUEUE_REG_9__0_ );
dff P2_P1_INSTQUEUE_REG_10__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__0_, n15076 );
not U_inv719 ( n73574, P2_P1_INSTQUEUE_REG_10__0_ );
dff P2_P1_INSTQUEUE_REG_11__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__0_, n15036 );
not U_inv720 ( n73567, P2_P1_INSTQUEUE_REG_11__0_ );
dff P2_P1_INSTQUEUE_REG_12__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__0_, n14996 );
not U_inv721 ( n73554, P2_P1_INSTQUEUE_REG_12__0_ );
dff P2_P1_INSTQUEUE_REG_13__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__0_, n14956 );
not U_inv722 ( n73560, P2_P1_INSTQUEUE_REG_13__0_ );
dff P2_P1_INSTQUEUE_REG_14__0__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__0_, n14916 );
not U_inv723 ( n73565, P2_P1_INSTQUEUE_REG_14__0_ );
dff P2_P1_LWORD_REG_0__reg ( clk, reset, P2_P1_LWORD_REG_0_, n15926 );
not U_inv724 ( n75653, P2_P1_LWORD_REG_0_ );
dff P2_P1_LWORD_REG_2__reg ( clk, reset, P2_P1_LWORD_REG_2_, n15916 );
not U_inv725 ( n75661, P2_P1_LWORD_REG_2_ );
dff P2_P1_DATAO_REG_2__reg ( clk, reset, P2_P1_DATAO_REG_2_, n16016 );
dff P2_BUF1_REG_2__reg ( clk, reset, P2_BUF1_REG_2_, n471 );
not U_inv726 ( n75450, P2_BUF1_REG_2_ );
dff P2_P1_LWORD_REG_13__reg ( clk, reset, P2_P1_LWORD_REG_13_, n15861 );
not U_inv727 ( n75660, P2_P1_LWORD_REG_13_ );
dff P2_P1_DATAO_REG_13__reg ( clk, reset, P2_P1_DATAO_REG_13_, n16071 );
dff P2_BUF1_REG_13__reg ( clk, reset, P2_BUF1_REG_13_, n526 );
not U_inv728 ( n75434, P2_BUF1_REG_13_ );
dff P2_P1_UWORD_REG_13__reg ( clk, reset, P2_P1_UWORD_REG_13_, n15936 );
not U_inv729 ( n75577, P2_P1_UWORD_REG_13_ );
dff P2_P1_DATAO_REG_29__reg ( clk, reset, P2_P1_DATAO_REG_29_, n16151 );
dff P2_BUF1_REG_29__reg ( clk, reset, P2_BUF1_REG_29_, n606 );
not U_inv730 ( n75367, P2_BUF1_REG_29_ );
dff P2_P1_INSTQUEUE_REG_14__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__5_, n14891 );
not U_inv731 ( n73889, P2_P1_INSTQUEUE_REG_14__5_ );
dff P2_P1_EAX_REG_5__reg ( clk, reset, P2_P1_EAX_REG_5_, n16191 );
not U_inv732 ( n73195, P2_P1_EAX_REG_5_ );
dff P2_P1_EAX_REG_7__reg ( clk, reset, P2_P1_EAX_REG_7_, n16201 );
not U_inv733 ( n74738, P2_P1_EAX_REG_7_ );
dff P2_P1_EAX_REG_8__reg ( clk, reset, P2_P1_EAX_REG_8_, n16206 );
not U_inv734 ( n73218, P2_P1_EAX_REG_8_ );
dff P2_P1_LWORD_REG_8__reg ( clk, reset, P2_P1_LWORD_REG_8_, n15886 );
not U_inv735 ( n75659, P2_P1_LWORD_REG_8_ );
dff P2_P1_DATAO_REG_8__reg ( clk, reset, P2_P1_DATAO_REG_8_, n16046 );
dff P2_BUF1_REG_8__reg ( clk, reset, P2_BUF1_REG_8_, n501 );
not U_inv736 ( n75433, P2_BUF1_REG_8_ );
dff P2_P2_UWORD_REG_8__reg ( clk, reset, P2_P2_UWORD_REG_8_, n13716 );
not U_inv737 ( n75561, P2_P2_UWORD_REG_8_ );
dff P2_P2_DATAO_REG_24__reg ( clk, reset, P2_P2_DATAO_REG_24_, n13881 );
not U_inv738 ( n75591, P2_P2_DATAO_REG_24_ );
dff P2_BUF2_REG_24__reg ( clk, reset, P2_BUF2_REG_24_, n741 );
not U_inv739 ( n75341, P2_BUF2_REG_24_ );
dff P2_P3_INSTQUEUE_REG_0__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__0_, n10986 );
not U_inv740 ( n73643, P2_P3_INSTQUEUE_REG_0__0_ );
dff P2_P3_EBX_REG_0__reg ( clk, reset, P2_P3_EBX_REG_0_, n11836 );
not U_inv741 ( n73121, P2_P3_EBX_REG_0_ );
dff P2_P3_INSTQUEUE_REG_1__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__0_, n10946 );
not U_inv742 ( n73665, P2_P3_INSTQUEUE_REG_1__0_ );
dff P2_P3_INSTQUEUE_REG_2__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__0_, n10906 );
not U_inv743 ( n73676, P2_P3_INSTQUEUE_REG_2__0_ );
dff P2_P3_INSTQUEUE_REG_3__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__0_, n10866 );
not U_inv744 ( n73655, P2_P3_INSTQUEUE_REG_3__0_ );
dff P2_P3_INSTQUEUE_REG_4__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__0_, n10826 );
not U_inv745 ( n73667, P2_P3_INSTQUEUE_REG_4__0_ );
dff P2_P3_INSTQUEUE_REG_5__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__0_, n10786 );
not U_inv746 ( n73692, P2_P3_INSTQUEUE_REG_5__0_ );
dff P2_P3_INSTQUEUE_REG_6__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__0_, n10746 );
not U_inv747 ( n73698, P2_P3_INSTQUEUE_REG_6__0_ );
dff P2_P3_INSTQUEUE_REG_7__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__0_, n10706 );
not U_inv748 ( n73681, P2_P3_INSTQUEUE_REG_7__0_ );
dff P2_P3_INSTQUEUE_REG_8__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__0_, n10666 );
not U_inv749 ( n73675, P2_P3_INSTQUEUE_REG_8__0_ );
dff P2_P3_INSTQUEUE_REG_9__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__0_, n10626 );
not U_inv750 ( n73695, P2_P3_INSTQUEUE_REG_9__0_ );
dff P2_P3_INSTQUEUE_REG_10__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__0_, n10586 );
not U_inv751 ( n73702, P2_P3_INSTQUEUE_REG_10__0_ );
dff P2_P3_INSTQUEUE_REG_11__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__0_, n10546 );
not U_inv752 ( n73687, P2_P3_INSTQUEUE_REG_11__0_ );
dff P2_P3_INSTQUEUE_REG_12__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__0_, n10506 );
not U_inv753 ( n73652, P2_P3_INSTQUEUE_REG_12__0_ );
dff P2_P3_INSTQUEUE_REG_13__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__0_, n10466 );
not U_inv754 ( n73674, P2_P3_INSTQUEUE_REG_13__0_ );
dff P2_P3_INSTQUEUE_REG_14__0__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__0_, n10426 );
not U_inv755 ( n73686, P2_P3_INSTQUEUE_REG_14__0_ );
dff P2_P2_LWORD_REG_8__reg ( clk, reset, P2_P2_LWORD_REG_8_, n13641 );
not U_inv756 ( n75623, P2_P2_LWORD_REG_8_ );
dff P2_P2_DATAO_REG_8__reg ( clk, reset, P2_P2_DATAO_REG_8_, n13801 );
not U_inv757 ( n75513, P2_P2_DATAO_REG_8_ );
dff P2_BUF2_REG_8__reg ( clk, reset, P2_BUF2_REG_8_, n661 );
not U_inv758 ( n75309, P2_BUF2_REG_8_ );
dff P2_P3_LWORD_REG_8__reg ( clk, reset, P2_P3_LWORD_REG_8_, n11396 );
not U_inv759 ( n75622, P2_P3_LWORD_REG_8_ );
dff P2_P3_DATAO_REG_8__reg ( clk, reset, P2_P3_DATAO_REG_8_, n11556 );
dff P2_P1_LWORD_REG_5__reg ( clk, reset, P2_P1_LWORD_REG_5_, n15901 );
not U_inv760 ( n75658, P2_P1_LWORD_REG_5_ );
dff P2_P1_DATAO_REG_5__reg ( clk, reset, P2_P1_DATAO_REG_5_, n16031 );
dff P2_BUF1_REG_5__reg ( clk, reset, P2_BUF1_REG_5_, n486 );
not U_inv761 ( n75449, P2_BUF1_REG_5_ );
dff P2_P1_INSTQUEUE_REG_5__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__5_, n15251 );
not U_inv762 ( n73891, P2_P1_INSTQUEUE_REG_5__5_ );
dff P2_P1_INSTQUEUE_REG_6__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__5_, n15211 );
not U_inv763 ( n73893, P2_P1_INSTQUEUE_REG_6__5_ );
dff P2_P1_INSTQUEUE_REG_7__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__5_, n15171 );
not U_inv764 ( n73888, P2_P1_INSTQUEUE_REG_7__5_ );
dff P2_P1_INSTQUEUE_REG_9__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__5_, n15091 );
not U_inv765 ( n73892, P2_P1_INSTQUEUE_REG_9__5_ );
dff P2_P1_INSTQUEUE_REG_10__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__5_, n15051 );
not U_inv766 ( n73894, P2_P1_INSTQUEUE_REG_10__5_ );
dff P2_P1_INSTQUEUE_REG_11__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__5_, n15011 );
not U_inv767 ( n73890, P2_P1_INSTQUEUE_REG_11__5_ );
dff P2_P1_INSTQUEUE_REG_13__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__5_, n14931 );
not U_inv768 ( n73885, P2_P1_INSTQUEUE_REG_13__5_ );
dff P2_P1_INSTQUEUE_REG_0__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__5_, n15451 );
not U_inv769 ( n73867, P2_P1_INSTQUEUE_REG_0__5_ );
dff P2_P1_INSTQUEUE_REG_1__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__5_, n15411 );
not U_inv770 ( n73883, P2_P1_INSTQUEUE_REG_1__5_ );
dff P2_P1_INSTQUEUE_REG_2__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__5_, n15371 );
not U_inv771 ( n73887, P2_P1_INSTQUEUE_REG_2__5_ );
dff P2_P1_INSTQUEUE_REG_3__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__5_, n15331 );
not U_inv772 ( n73881, P2_P1_INSTQUEUE_REG_3__5_ );
dff P2_P1_INSTQUEUE_REG_4__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__5_, n15291 );
not U_inv773 ( n73884, P2_P1_INSTQUEUE_REG_4__5_ );
dff P2_P1_INSTQUEUE_REG_8__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__5_, n15131 );
not U_inv774 ( n73886, P2_P1_INSTQUEUE_REG_8__5_ );
dff P2_P1_INSTQUEUE_REG_12__5__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__5_, n14971 );
not U_inv775 ( n73880, P2_P1_INSTQUEUE_REG_12__5_ );
dff P2_P1_EAX_REG_21__reg ( clk, reset, P2_P1_EAX_REG_21_, n16271 );
not U_inv776 ( n73288, P2_P1_EAX_REG_21_ );
dff P2_P1_EAX_REG_22__reg ( clk, reset, P2_P1_EAX_REG_22_, n16276 );
not U_inv777 ( n75001, P2_P1_EAX_REG_22_ );
dff P2_P1_UWORD_REG_6__reg ( clk, reset, P2_P1_UWORD_REG_6_, n15971 );
not U_inv778 ( n75492, P2_P1_UWORD_REG_6_ );
dff P2_P1_DATAO_REG_22__reg ( clk, reset, P2_P1_DATAO_REG_22_, n16116 );
dff P2_P1_EAX_REG_23__reg ( clk, reset, ex_wire177, n16281 );
not U_inv779 ( n75012, ex_wire177 );
dff P2_P1_EAX_REG_25__reg ( clk, reset, P2_P1_EAX_REG_25_, n16291 );
not U_inv780 ( n75061, P2_P1_EAX_REG_25_ );
dff P2_P1_EAX_REG_26__reg ( clk, reset, ex_wire178, n16296 );
not U_inv781 ( n75084, ex_wire178 );
dff P2_P1_UWORD_REG_10__reg ( clk, reset, P2_P1_UWORD_REG_10_, n15951 );
not U_inv782 ( n75576, P2_P1_UWORD_REG_10_ );
dff P2_P1_DATAO_REG_26__reg ( clk, reset, P2_P1_DATAO_REG_26_, n16136 );
dff P2_BUF1_REG_26__reg ( clk, reset, P2_BUF1_REG_26_, n591 );
not U_inv783 ( n75366, P2_BUF1_REG_26_ );
dff P2_P1_INSTQUEUE_REG_15__2__reg ( clk, reset, ex_wire179, n14866 );
not U_inv784 ( n73611, ex_wire179 );
dff P2_P1_EAX_REG_18__reg ( clk, reset, P2_P1_EAX_REG_18_, n16256 );
not U_inv785 ( n73265, P2_P1_EAX_REG_18_ );
dff P2_P1_UWORD_REG_2__reg ( clk, reset, P2_P1_UWORD_REG_2_, n15991 );
not U_inv786 ( n75491, P2_P1_UWORD_REG_2_ );
dff P2_P1_DATAO_REG_18__reg ( clk, reset, P2_P1_DATAO_REG_18_, n16096 );
dff P2_BUF1_REG_18__reg ( clk, reset, P2_BUF1_REG_18_, n551 );
not U_inv787 ( n75371, P2_BUF1_REG_18_ );
dff P2_P1_INSTQUEUE_REG_0__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__2_, n15466 );
not U_inv788 ( n73558, P2_P1_INSTQUEUE_REG_0__2_ );
dff P2_P1_INSTQUEUE_REG_1__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__2_, n15426 );
not U_inv789 ( n73575, P2_P1_INSTQUEUE_REG_1__2_ );
dff P2_P1_INSTQUEUE_REG_2__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__2_, n15386 );
not U_inv790 ( n73584, P2_P1_INSTQUEUE_REG_2__2_ );
dff P2_P1_INSTQUEUE_REG_3__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__2_, n15346 );
not U_inv791 ( n73577, P2_P1_INSTQUEUE_REG_3__2_ );
dff P2_P1_INSTQUEUE_REG_4__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__2_, n15306 );
not U_inv792 ( n73573, P2_P1_INSTQUEUE_REG_4__2_ );
dff P2_P1_INSTQUEUE_REG_5__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__2_, n15266 );
not U_inv793 ( n73578, P2_P1_INSTQUEUE_REG_5__2_ );
dff P2_P1_INSTQUEUE_REG_6__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__2_, n15226 );
not U_inv794 ( n73587, P2_P1_INSTQUEUE_REG_6__2_ );
dff P2_P1_INSTQUEUE_REG_7__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__2_, n15186 );
not U_inv795 ( n73581, P2_P1_INSTQUEUE_REG_7__2_ );
dff P2_P1_INSTQUEUE_REG_8__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__2_, n15146 );
not U_inv796 ( n73580, P2_P1_INSTQUEUE_REG_8__2_ );
dff P2_P1_INSTQUEUE_REG_9__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__2_, n15106 );
not U_inv797 ( n73586, P2_P1_INSTQUEUE_REG_9__2_ );
dff P2_P1_INSTQUEUE_REG_10__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__2_, n15066 );
not U_inv798 ( n73599, P2_P1_INSTQUEUE_REG_10__2_ );
dff P2_P1_INSTQUEUE_REG_11__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__2_, n15026 );
not U_inv799 ( n73591, P2_P1_INSTQUEUE_REG_11__2_ );
dff P2_P1_INSTQUEUE_REG_12__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__2_, n14986 );
not U_inv800 ( n73576, P2_P1_INSTQUEUE_REG_12__2_ );
dff P2_P1_INSTQUEUE_REG_13__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__2_, n14946 );
not U_inv801 ( n73582, P2_P1_INSTQUEUE_REG_13__2_ );
dff P2_P1_INSTQUEUE_REG_14__2__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__2_, n14906 );
not U_inv802 ( n73593, P2_P1_INSTQUEUE_REG_14__2_ );
dff P2_P1_EAX_REG_10__reg ( clk, reset, P2_P1_EAX_REG_10_, n16216 );
not U_inv803 ( n74786, P2_P1_EAX_REG_10_ );
dff P2_P1_EAX_REG_11__reg ( clk, reset, P2_P1_EAX_REG_11_, n16221 );
not U_inv804 ( n73237, P2_P1_EAX_REG_11_ );
dff P2_P1_LWORD_REG_11__reg ( clk, reset, P2_P1_LWORD_REG_11_, n15871 );
not U_inv805 ( n75657, P2_P1_LWORD_REG_11_ );
dff P2_P1_DATAO_REG_11__reg ( clk, reset, P2_P1_DATAO_REG_11_, n16061 );
dff P2_BUF1_REG_11__reg ( clk, reset, P2_BUF1_REG_11_, n516 );
not U_inv806 ( n75432, P2_BUF1_REG_11_ );
dff P2_P2_UWORD_REG_11__reg ( clk, reset, P2_P2_UWORD_REG_11_, n13701 );
not U_inv807 ( n75560, P2_P2_UWORD_REG_11_ );
dff P2_P2_DATAO_REG_27__reg ( clk, reset, P2_P2_DATAO_REG_27_, n13896 );
not U_inv808 ( n75587, P2_P2_DATAO_REG_27_ );
dff P2_BUF2_REG_27__reg ( clk, reset, P2_BUF2_REG_27_, n756 );
not U_inv809 ( n75338, P2_BUF2_REG_27_ );
dff P2_P2_LWORD_REG_11__reg ( clk, reset, P2_P2_LWORD_REG_11_, n13626 );
not U_inv810 ( n75621, P2_P2_LWORD_REG_11_ );
dff P2_P2_DATAO_REG_11__reg ( clk, reset, P2_P2_DATAO_REG_11_, n13816 );
not U_inv811 ( n75510, P2_P2_DATAO_REG_11_ );
dff P2_BUF2_REG_11__reg ( clk, reset, P2_BUF2_REG_11_, n676 );
not U_inv812 ( n75307, P2_BUF2_REG_11_ );
dff P2_P1_EAX_REG_12__reg ( clk, reset, ex_wire180, n16226 );
not U_inv813 ( n74803, ex_wire180 );
dff P2_P1_LWORD_REG_12__reg ( clk, reset, P2_P1_LWORD_REG_12_, n15866 );
not U_inv814 ( n75656, P2_P1_LWORD_REG_12_ );
dff P2_P1_DATAO_REG_12__reg ( clk, reset, P2_P1_DATAO_REG_12_, n16066 );
dff P2_BUF1_REG_12__reg ( clk, reset, P2_BUF1_REG_12_, n521 );
not U_inv815 ( n75431, P2_BUF1_REG_12_ );
dff P2_P2_UWORD_REG_12__reg ( clk, reset, P2_P2_UWORD_REG_12_, n13696 );
not U_inv816 ( n75559, P2_P2_UWORD_REG_12_ );
dff P2_P2_DATAO_REG_28__reg ( clk, reset, P2_P2_DATAO_REG_28_, n13901 );
not U_inv817 ( n75588, P2_P2_DATAO_REG_28_ );
dff P2_BUF1_REG_28__reg ( clk, reset, P2_BUF1_REG_28_, n601 );
not U_inv818 ( n75408, P2_BUF1_REG_28_ );
dff P2_P1_INSTQUEUE_REG_15__4__reg ( clk, reset, ex_wire181, n14856 );
not U_inv819 ( n73808, ex_wire181 );
dff P2_P1_EAX_REG_20__reg ( clk, reset, ex_wire182, n16266 );
not U_inv820 ( n74965, ex_wire182 );
dff P2_P1_UWORD_REG_4__reg ( clk, reset, P2_P1_UWORD_REG_4_, n15981 );
not U_inv821 ( n75490, P2_P1_UWORD_REG_4_ );
dff P2_P1_DATAO_REG_20__reg ( clk, reset, P2_P1_DATAO_REG_20_, n16106 );
dff P2_BUF1_REG_20__reg ( clk, reset, P2_BUF1_REG_20_, n561 );
not U_inv822 ( n75370, P2_BUF1_REG_20_ );
dff P2_P1_INSTQUEUE_REG_0__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__4_, n15456 );
not U_inv823 ( n73805, P2_P1_INSTQUEUE_REG_0__4_ );
dff P2_P1_INSTQUEUE_REG_1__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__4_, n15416 );
not U_inv824 ( n73809, P2_P1_INSTQUEUE_REG_1__4_ );
dff P2_P1_INSTQUEUE_REG_2__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__4_, n15376 );
not U_inv825 ( n73813, P2_P1_INSTQUEUE_REG_2__4_ );
dff P2_P1_INSTQUEUE_REG_3__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__4_, n15336 );
not U_inv826 ( n73807, P2_P1_INSTQUEUE_REG_3__4_ );
dff P2_P1_INSTQUEUE_REG_4__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__4_, n15296 );
not U_inv827 ( n73810, P2_P1_INSTQUEUE_REG_4__4_ );
dff P2_P1_INSTQUEUE_REG_5__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__4_, n15256 );
not U_inv828 ( n73817, P2_P1_INSTQUEUE_REG_5__4_ );
dff P2_P1_INSTQUEUE_REG_6__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__4_, n15216 );
not U_inv829 ( n73819, P2_P1_INSTQUEUE_REG_6__4_ );
dff P2_P1_INSTQUEUE_REG_7__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__4_, n15176 );
not U_inv830 ( n73814, P2_P1_INSTQUEUE_REG_7__4_ );
dff P2_P1_INSTQUEUE_REG_8__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__4_, n15136 );
not U_inv831 ( n73812, P2_P1_INSTQUEUE_REG_8__4_ );
dff P2_P1_INSTQUEUE_REG_9__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__4_, n15096 );
not U_inv832 ( n73818, P2_P1_INSTQUEUE_REG_9__4_ );
dff P2_P1_INSTQUEUE_REG_10__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__4_, n15056 );
not U_inv833 ( n73820, P2_P1_INSTQUEUE_REG_10__4_ );
dff P2_P1_INSTQUEUE_REG_11__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__4_, n15016 );
not U_inv834 ( n73816, P2_P1_INSTQUEUE_REG_11__4_ );
dff P2_P1_INSTQUEUE_REG_12__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_12__4_, n14976 );
not U_inv835 ( n73806, P2_P1_INSTQUEUE_REG_12__4_ );
dff P2_P1_INSTQUEUE_REG_13__4__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__4_, n14936 );
not U_inv836 ( n73811, P2_P1_INSTQUEUE_REG_13__4_ );
dff P2_P1_EAX_REG_27__reg ( clk, reset, P2_P1_EAX_REG_27_, n16301 );
not U_inv837 ( n73320, P2_P1_EAX_REG_27_ );
dff P2_P1_UWORD_REG_11__reg ( clk, reset, P2_P1_UWORD_REG_11_, n15946 );
not U_inv838 ( n75575, P2_P1_UWORD_REG_11_ );
dff P2_P1_DATAO_REG_27__reg ( clk, reset, P2_P1_DATAO_REG_27_, n16141 );
dff P2_BUF1_REG_27__reg ( clk, reset, P2_BUF1_REG_27_, n596 );
not U_inv839 ( n75407, P2_BUF1_REG_27_ );
dff P2_P1_INSTQUEUE_REG_15__3__reg ( clk, reset, ex_wire183, n14861 );
not U_inv840 ( n73640, ex_wire183 );
dff P2_P1_EAX_REG_19__reg ( clk, reset, P2_P1_EAX_REG_19_, n16261 );
not U_inv841 ( n74953, P2_P1_EAX_REG_19_ );
dff P2_P1_UWORD_REG_3__reg ( clk, reset, P2_P1_UWORD_REG_3_, n15986 );
not U_inv842 ( n75489, P2_P1_UWORD_REG_3_ );
dff P2_P1_DATAO_REG_19__reg ( clk, reset, P2_P1_DATAO_REG_19_, n16101 );
dff P2_BUF1_REG_19__reg ( clk, reset, P2_BUF1_REG_19_, n556 );
not U_inv843 ( n75369, P2_BUF1_REG_19_ );
dff P2_P1_INSTQUEUE_REG_0__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_0__3_, n15461 );
not U_inv844 ( n73636, P2_P1_INSTQUEUE_REG_0__3_ );
dff P2_P1_INSTQUEUE_REG_1__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_1__3_, n15421 );
not U_inv845 ( n73644, P2_P1_INSTQUEUE_REG_1__3_ );
dff P2_P1_INSTQUEUE_REG_2__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_2__3_, n15381 );
not U_inv846 ( n73648, P2_P1_INSTQUEUE_REG_2__3_ );
dff P2_P1_INSTQUEUE_REG_3__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_3__3_, n15341 );
not U_inv847 ( n73639, P2_P1_INSTQUEUE_REG_3__3_ );
dff P2_P1_INSTQUEUE_REG_4__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_4__3_, n15301 );
not U_inv848 ( n73645, P2_P1_INSTQUEUE_REG_4__3_ );
dff P2_P1_INSTQUEUE_REG_5__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_5__3_, n15261 );
not U_inv849 ( n73656, P2_P1_INSTQUEUE_REG_5__3_ );
dff P2_P1_INSTQUEUE_REG_6__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_6__3_, n15221 );
not U_inv850 ( n73663, P2_P1_INSTQUEUE_REG_6__3_ );
dff P2_P1_INSTQUEUE_REG_7__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_7__3_, n15181 );
not U_inv851 ( n73649, P2_P1_INSTQUEUE_REG_7__3_ );
dff P2_P1_INSTQUEUE_REG_8__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_8__3_, n15141 );
not U_inv852 ( n73647, P2_P1_INSTQUEUE_REG_8__3_ );
dff P2_P1_INSTQUEUE_REG_9__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_9__3_, n15101 );
not U_inv853 ( n73662, P2_P1_INSTQUEUE_REG_9__3_ );
dff P2_P1_INSTQUEUE_REG_10__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_10__3_, n15061 );
not U_inv854 ( n73664, P2_P1_INSTQUEUE_REG_10__3_ );
dff P2_P1_INSTQUEUE_REG_11__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_11__3_, n15021 );
not U_inv855 ( n73651, P2_P1_INSTQUEUE_REG_11__3_ );
dff P2_P1_INSTQUEUE_REG_13__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_13__3_, n14941 );
not U_inv856 ( n73646, P2_P1_INSTQUEUE_REG_13__3_ );
dff P2_P1_INSTQUEUE_REG_14__3__reg ( clk, reset, P2_P1_INSTQUEUE_REG_14__3_, n14901 );
not U_inv857 ( n73650, P2_P1_INSTQUEUE_REG_14__3_ );
dff P2_P1_EAX_REG_28__reg ( clk, reset, P2_P1_EAX_REG_28_, n16306 );
not U_inv858 ( n75324, P2_P1_EAX_REG_28_ );
dff P2_P1_UWORD_REG_12__reg ( clk, reset, P2_P1_UWORD_REG_12_, n15941 );
not U_inv859 ( n75574, P2_P1_UWORD_REG_12_ );
dff P2_P1_DATAO_REG_28__reg ( clk, reset, P2_P1_DATAO_REG_28_, n16146 );
dff P2_P1_EAX_REG_29__reg ( clk, reset, P2_P1_EAX_REG_29_, n16311 );
not U_inv860 ( n75218, P2_P1_EAX_REG_29_ );
dff P2_BUF2_REG_28__reg ( clk, reset, P2_BUF2_REG_28_, n761 );
not U_inv861 ( n75326, P2_BUF2_REG_28_ );
dff P2_P2_INSTQUEUE_REG_5__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__4_, n13011 );
not U_inv862 ( n73870, P2_P2_INSTQUEUE_REG_5__4_ );
dff P2_P2_INSTQUEUE_REG_6__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__4_, n12971 );
not U_inv863 ( n73876, P2_P2_INSTQUEUE_REG_6__4_ );
dff P2_P2_INSTQUEUE_REG_7__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__4_, n12931 );
not U_inv864 ( n73860, P2_P2_INSTQUEUE_REG_7__4_ );
dff P2_P2_INSTQUEUE_REG_8__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__4_, n12891 );
not U_inv865 ( n73854, P2_P2_INSTQUEUE_REG_8__4_ );
dff P2_P2_INSTQUEUE_REG_9__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__4_, n12851 );
not U_inv866 ( n73873, P2_P2_INSTQUEUE_REG_9__4_ );
dff P2_P2_INSTQUEUE_REG_10__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__4_, n12811 );
not U_inv867 ( n73879, P2_P2_INSTQUEUE_REG_10__4_ );
dff P2_P2_INSTQUEUE_REG_11__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__4_, n12771 );
not U_inv868 ( n73866, P2_P2_INSTQUEUE_REG_11__4_ );
dff P2_P2_INSTQUEUE_REG_12__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__4_, n12731 );
not U_inv869 ( n73836, P2_P2_INSTQUEUE_REG_12__4_ );
dff P2_P2_INSTQUEUE_REG_13__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__4_, n12691 );
not U_inv870 ( n73852, P2_P2_INSTQUEUE_REG_13__4_ );
dff P2_P2_INSTQUEUE_REG_14__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__4_, n12651 );
not U_inv871 ( n73863, P2_P2_INSTQUEUE_REG_14__4_ );
dff P2_P2_INSTQUEUE_REG_0__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__4_, n13211 );
not U_inv872 ( n73832, P2_P2_INSTQUEUE_REG_0__4_ );
dff P2_P2_INSTQUEUE_REG_1__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__4_, n13171 );
not U_inv873 ( n73846, P2_P2_INSTQUEUE_REG_1__4_ );
dff P2_P2_INSTQUEUE_REG_2__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__4_, n13131 );
not U_inv874 ( n73857, P2_P2_INSTQUEUE_REG_2__4_ );
dff P2_P2_INSTQUEUE_REG_3__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__4_, n13091 );
not U_inv875 ( n73839, P2_P2_INSTQUEUE_REG_3__4_ );
dff P2_P2_INSTQUEUE_REG_4__4__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__4_, n13051 );
not U_inv876 ( n73848, P2_P2_INSTQUEUE_REG_4__4_ );
dff P2_P3_INSTQUEUE_REG_0__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__4_, n10966 );
not U_inv877 ( n73830, P2_P3_INSTQUEUE_REG_0__4_ );
dff P2_P3_INSTQUEUE_REG_1__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__4_, n10926 );
not U_inv878 ( n73843, P2_P3_INSTQUEUE_REG_1__4_ );
dff P2_P3_INSTQUEUE_REG_2__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__4_, n10886 );
not U_inv879 ( n73855, P2_P3_INSTQUEUE_REG_2__4_ );
dff P2_P3_INSTQUEUE_REG_3__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__4_, n10846 );
not U_inv880 ( n73837, P2_P3_INSTQUEUE_REG_3__4_ );
dff P2_P3_INSTQUEUE_REG_4__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__4_, n10806 );
not U_inv881 ( n73844, P2_P3_INSTQUEUE_REG_4__4_ );
dff P2_P3_INSTQUEUE_REG_15__4__reg ( clk, reset, ex_wire184, n10366 );
not U_inv882 ( n73840, ex_wire184 );
dff P2_P3_INSTQUEUE_REG_5__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__4_, n10766 );
not U_inv883 ( n73868, P2_P3_INSTQUEUE_REG_5__4_ );
dff P2_P3_INSTQUEUE_REG_6__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__4_, n10726 );
not U_inv884 ( n73874, P2_P3_INSTQUEUE_REG_6__4_ );
dff P2_P3_INSTQUEUE_REG_7__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__4_, n10686 );
not U_inv885 ( n73858, P2_P3_INSTQUEUE_REG_7__4_ );
dff P2_P3_INSTQUEUE_REG_8__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__4_, n10646 );
not U_inv886 ( n73850, P2_P3_INSTQUEUE_REG_8__4_ );
dff P2_P3_INSTQUEUE_REG_9__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__4_, n10606 );
not U_inv887 ( n73871, P2_P3_INSTQUEUE_REG_9__4_ );
dff P2_P3_INSTQUEUE_REG_10__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__4_, n10566 );
not U_inv888 ( n73877, P2_P3_INSTQUEUE_REG_10__4_ );
dff P2_P3_INSTQUEUE_REG_11__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__4_, n10526 );
not U_inv889 ( n73864, P2_P3_INSTQUEUE_REG_11__4_ );
dff P2_P3_INSTQUEUE_REG_12__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__4_, n10486 );
not U_inv890 ( n73834, P2_P3_INSTQUEUE_REG_12__4_ );
dff P2_P3_INSTQUEUE_REG_13__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__4_, n10446 );
not U_inv891 ( n73849, P2_P3_INSTQUEUE_REG_13__4_ );
dff P2_P3_INSTQUEUE_REG_14__4__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__4_, n10406 );
not U_inv892 ( n73861, P2_P3_INSTQUEUE_REG_14__4_ );
dff P2_P2_LWORD_REG_12__reg ( clk, reset, P2_P2_LWORD_REG_12_, n13621 );
not U_inv893 ( n75620, P2_P2_LWORD_REG_12_ );
dff P2_P2_DATAO_REG_12__reg ( clk, reset, P2_P2_DATAO_REG_12_, n13821 );
not U_inv894 ( n75509, P2_P2_DATAO_REG_12_ );
dff P2_BUF2_REG_12__reg ( clk, reset, P2_BUF2_REG_12_, n681 );
not U_inv895 ( n75306, P2_BUF2_REG_12_ );
dff P2_P1_LWORD_REG_10__reg ( clk, reset, P2_P1_LWORD_REG_10_, n15876 );
not U_inv896 ( n75655, P2_P1_LWORD_REG_10_ );
dff P2_P1_DATAO_REG_10__reg ( clk, reset, P2_P1_DATAO_REG_10_, n16056 );
dff P2_BUF1_REG_10__reg ( clk, reset, P2_BUF1_REG_10_, n511 );
not U_inv897 ( n75430, P2_BUF1_REG_10_ );
dff P2_P2_INSTQUEUE_REG_5__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__2_, n13021 );
not U_inv898 ( n73717, P2_P2_INSTQUEUE_REG_5__2_ );
dff P2_P2_INSTQUEUE_REG_6__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__2_, n12981 );
not U_inv899 ( n73735, P2_P2_INSTQUEUE_REG_6__2_ );
dff P2_P2_INSTQUEUE_REG_7__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__2_, n12941 );
not U_inv900 ( n73723, P2_P2_INSTQUEUE_REG_7__2_ );
dff P2_P2_INSTQUEUE_REG_8__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__2_, n12901 );
not U_inv901 ( n73720, P2_P2_INSTQUEUE_REG_8__2_ );
dff P2_P2_INSTQUEUE_REG_9__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__2_, n12861 );
not U_inv902 ( n73732, P2_P2_INSTQUEUE_REG_9__2_ );
dff P2_P2_INSTQUEUE_REG_10__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__2_, n12821 );
not U_inv903 ( n73744, P2_P2_INSTQUEUE_REG_10__2_ );
dff P2_P2_INSTQUEUE_REG_11__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__2_, n12781 );
not U_inv904 ( n73738, P2_P2_INSTQUEUE_REG_11__2_ );
dff P2_P2_INSTQUEUE_REG_12__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__2_, n12741 );
not U_inv905 ( n73712, P2_P2_INSTQUEUE_REG_12__2_ );
dff P2_P2_INSTQUEUE_REG_13__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__2_, n12701 );
not U_inv906 ( n73726, P2_P2_INSTQUEUE_REG_13__2_ );
dff P2_P2_INSTQUEUE_REG_14__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__2_, n12661 );
not U_inv907 ( n73741, P2_P2_INSTQUEUE_REG_14__2_ );
dff P2_P2_INSTQUEUE_REG_0__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__2_, n13221 );
not U_inv908 ( n73670, P2_P2_INSTQUEUE_REG_0__2_ );
dff P2_P2_INSTQUEUE_REG_1__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__2_, n13181 );
not U_inv909 ( n73708, P2_P2_INSTQUEUE_REG_1__2_ );
dff P2_P2_INSTQUEUE_REG_2__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__2_, n13141 );
not U_inv910 ( n73729, P2_P2_INSTQUEUE_REG_2__2_ );
dff P2_P2_INSTQUEUE_REG_3__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__2_, n13101 );
not U_inv911 ( n73715, P2_P2_INSTQUEUE_REG_3__2_ );
dff P2_P2_INSTQUEUE_REG_4__2__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__2_, n13061 );
not U_inv912 ( n73705, P2_P2_INSTQUEUE_REG_4__2_ );
dff P2_P1_UWORD_REG_5__reg ( clk, reset, P2_P1_UWORD_REG_5_, n15976 );
not U_inv913 ( n75488, P2_P1_UWORD_REG_5_ );
dff P2_P1_DATAO_REG_21__reg ( clk, reset, P2_P1_DATAO_REG_21_, n16111 );
dff P2_P1_EAX_REG_13__reg ( clk, reset, P2_P1_EAX_REG_13_, n16231 );
not U_inv914 ( n74842, P2_P1_EAX_REG_13_ );
dff P2_P2_LWORD_REG_5__reg ( clk, reset, P2_P2_LWORD_REG_5_, n13656 );
not U_inv915 ( n75619, P2_P2_LWORD_REG_5_ );
dff P2_P2_DATAO_REG_5__reg ( clk, reset, P2_P2_DATAO_REG_5_, n13786 );
not U_inv916 ( n75512, P2_P2_DATAO_REG_5_ );
dff P2_BUF2_REG_5__reg ( clk, reset, P2_BUF2_REG_5_, n646 );
not U_inv917 ( n75291, P2_BUF2_REG_5_ );
dff P2_P3_LWORD_REG_5__reg ( clk, reset, P2_P3_LWORD_REG_5_, n11411 );
not U_inv918 ( n75618, P2_P3_LWORD_REG_5_ );
dff P2_P3_DATAO_REG_5__reg ( clk, reset, P2_P3_DATAO_REG_5_, n11541 );
dff P2_P2_LWORD_REG_13__reg ( clk, reset, P2_P2_LWORD_REG_13_, n13616 );
not U_inv919 ( n75617, P2_P2_LWORD_REG_13_ );
dff P2_P2_DATAO_REG_13__reg ( clk, reset, P2_P2_DATAO_REG_13_, n13826 );
not U_inv920 ( n75514, P2_P2_DATAO_REG_13_ );
dff P2_BUF2_REG_13__reg ( clk, reset, P2_BUF2_REG_13_, n686 );
not U_inv921 ( n75305, P2_BUF2_REG_13_ );
dff P2_P2_INSTQUEUE_REG_5__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__0_, n13031 );
not U_inv922 ( n73693, P2_P2_INSTQUEUE_REG_5__0_ );
dff P2_P2_INSTQUEUE_REG_6__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__0_, n12991 );
not U_inv923 ( n73699, P2_P2_INSTQUEUE_REG_6__0_ );
dff P2_P2_INSTQUEUE_REG_7__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__0_, n12951 );
not U_inv924 ( n73684, P2_P2_INSTQUEUE_REG_7__0_ );
dff P2_P2_INSTQUEUE_REG_8__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__0_, n12911 );
not U_inv925 ( n73679, P2_P2_INSTQUEUE_REG_8__0_ );
dff P2_P2_INSTQUEUE_REG_9__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__0_, n12871 );
not U_inv926 ( n73696, P2_P2_INSTQUEUE_REG_9__0_ );
dff P2_P2_INSTQUEUE_REG_10__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__0_, n12831 );
not U_inv927 ( n73703, P2_P2_INSTQUEUE_REG_10__0_ );
dff P2_P2_INSTQUEUE_REG_11__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__0_, n12791 );
not U_inv928 ( n73690, P2_P2_INSTQUEUE_REG_11__0_ );
dff P2_P2_INSTQUEUE_REG_12__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__0_, n12751 );
not U_inv929 ( n73653, P2_P2_INSTQUEUE_REG_12__0_ );
dff P2_P2_INSTQUEUE_REG_13__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__0_, n12711 );
not U_inv930 ( n73677, P2_P2_INSTQUEUE_REG_13__0_ );
dff P2_P2_INSTQUEUE_REG_14__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__0_, n12671 );
not U_inv931 ( n73688, P2_P2_INSTQUEUE_REG_14__0_ );
dff P2_P2_INSTQUEUE_REG_0__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__0_, n13231 );
not U_inv932 ( n73642, P2_P2_INSTQUEUE_REG_0__0_ );
dff P2_P2_EBX_REG_0__reg ( clk, reset, P2_P2_EBX_REG_0_, n14081 );
not U_inv933 ( n73122, P2_P2_EBX_REG_0_ );
dff P2_P2_INSTQUEUE_REG_1__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__0_, n13191 );
not U_inv934 ( n73668, P2_P2_INSTQUEUE_REG_1__0_ );
dff P2_P2_INSTQUEUE_REG_2__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__0_, n13151 );
not U_inv935 ( n73682, P2_P2_INSTQUEUE_REG_2__0_ );
dff P2_P2_INSTQUEUE_REG_3__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__0_, n13111 );
not U_inv936 ( n73657, P2_P2_INSTQUEUE_REG_3__0_ );
dff P2_P2_INSTQUEUE_REG_4__0__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__0_, n13071 );
not U_inv937 ( n73672, P2_P2_INSTQUEUE_REG_4__0_ );
dff P2_P2_PHYADDRPOINTER_REG_0__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_0_, n13446 );
not U_inv938 ( n75224, P2_P2_PHYADDRPOINTER_REG_0_ );
dff P2_P2_LWORD_REG_9__reg ( clk, reset, P2_P2_LWORD_REG_9_, n13636 );
not U_inv939 ( n75616, P2_P2_LWORD_REG_9_ );
dff P2_P2_DATAO_REG_9__reg ( clk, reset, P2_P2_DATAO_REG_9_, n13806 );
not U_inv940 ( n75517, P2_P2_DATAO_REG_9_ );
dff P2_BUF2_REG_9__reg ( clk, reset, P2_BUF2_REG_9_, n666 );
not U_inv941 ( n75308, P2_BUF2_REG_9_ );
dff P2_P3_LWORD_REG_9__reg ( clk, reset, P2_P3_LWORD_REG_9_, n11391 );
not U_inv942 ( n75615, P2_P3_LWORD_REG_9_ );
dff P2_P3_DATAO_REG_9__reg ( clk, reset, P2_P3_DATAO_REG_9_, n11561 );
dff P2_P1_REQUESTPENDING_REG_reg ( clk, reset, P2_P1_REQUESTPENDING_REG, n16686 );
not U_inv943 ( n75253, P2_P1_REQUESTPENDING_REG );
dff P2_P1_CODEFETCH_REG_reg ( clk, reset, P2_P1_CODEFETCH_REG, n16701 );
dff P2_P1_D_C_N_REG_reg ( clk, reset, P2_P1_D_C_N_REG, n16691 );
dff P2_P1_MORE_REG_reg ( clk, reset, P2_P1_MORE_REG, n16676 );
dff P2_P1_READREQUEST_REG_reg ( clk, reset, P2_P1_READREQUEST_REG, n16711 );
dff P2_P1_W_R_N_REG_reg ( clk, reset, P2_P1_W_R_N_REG, n16666 );
dff P2_P1_EBX_REG_0__reg ( clk, reset, P2_P1_EBX_REG_0_, n16326 );
not U_inv944 ( n73123, P2_P1_EBX_REG_0_ );
dff P2_P1_EBX_REG_2__reg ( clk, reset, P2_P1_EBX_REG_2_, n16336 );
not U_inv945 ( n74536, P2_P1_EBX_REG_2_ );
dff P2_P1_EBX_REG_3__reg ( clk, reset, P2_P1_EBX_REG_3_, n16341 );
not U_inv946 ( n73142, P2_P1_EBX_REG_3_ );
dff P2_P1_EBX_REG_4__reg ( clk, reset, P2_P1_EBX_REG_4_, n16346 );
not U_inv947 ( n74571, P2_P1_EBX_REG_4_ );
dff P2_P1_EBX_REG_5__reg ( clk, reset, P2_P1_EBX_REG_5_, n16351 );
not U_inv948 ( n73156, P2_P1_EBX_REG_5_ );
dff P2_P1_EBX_REG_6__reg ( clk, reset, P2_P1_EBX_REG_6_, n16356 );
not U_inv949 ( n74604, P2_P1_EBX_REG_6_ );
dff P2_P1_EBX_REG_7__reg ( clk, reset, P2_P1_EBX_REG_7_, n16361 );
not U_inv950 ( n73174, P2_P1_EBX_REG_7_ );
dff P2_P1_EBX_REG_8__reg ( clk, reset, P2_P1_EBX_REG_8_, n16366 );
not U_inv951 ( n74667, P2_P1_EBX_REG_8_ );
dff P2_P1_EBX_REG_9__reg ( clk, reset, P2_P1_EBX_REG_9_, n16371 );
not U_inv952 ( n73204, P2_P1_EBX_REG_9_ );
dff P2_P1_EBX_REG_10__reg ( clk, reset, P2_P1_EBX_REG_10_, n16376 );
not U_inv953 ( n74722, P2_P1_EBX_REG_10_ );
dff P2_P1_EBX_REG_11__reg ( clk, reset, P2_P1_EBX_REG_11_, n16381 );
not U_inv954 ( n73212, P2_P1_EBX_REG_11_ );
dff P2_P1_EBX_REG_12__reg ( clk, reset, P2_P1_EBX_REG_12_, n16386 );
not U_inv955 ( n74765, P2_P1_EBX_REG_12_ );
dff P2_P1_EBX_REG_13__reg ( clk, reset, P2_P1_EBX_REG_13_, n16391 );
not U_inv956 ( n73226, P2_P1_EBX_REG_13_ );
dff P2_P2_INSTQUEUE_REG_0__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__1_, n13226 );
not U_inv957 ( n73568, P2_P2_INSTQUEUE_REG_0__1_ );
dff P2_P2_EBX_REG_2__reg ( clk, reset, P2_P2_EBX_REG_2_, n14091 );
not U_inv958 ( n74535, P2_P2_EBX_REG_2_ );
dff P2_P2_INSTQUEUE_REG_1__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__1_, n13186 );
not U_inv959 ( n73600, P2_P2_INSTQUEUE_REG_1__1_ );
dff P2_P2_INSTQUEUE_REG_2__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__1_, n13146 );
not U_inv960 ( n73619, P2_P2_INSTQUEUE_REG_2__1_ );
dff P2_P2_INSTQUEUE_REG_3__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__1_, n13106 );
not U_inv961 ( n73606, P2_P2_INSTQUEUE_REG_3__1_ );
dff P2_P2_INSTQUEUE_REG_7__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__1_, n12946 );
not U_inv962 ( n73615, P2_P2_INSTQUEUE_REG_7__1_ );
dff P2_P2_INSTQUEUE_REG_5__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__1_, n13026 );
not U_inv963 ( n73608, P2_P2_INSTQUEUE_REG_5__1_ );
dff P2_P2_INSTQUEUE_REG_6__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__1_, n12986 );
not U_inv964 ( n73624, P2_P2_INSTQUEUE_REG_6__1_ );
dff P2_P2_INSTQUEUE_REG_8__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__1_, n12906 );
not U_inv965 ( n73613, P2_P2_INSTQUEUE_REG_8__1_ );
dff P2_P2_INSTQUEUE_REG_9__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__1_, n12866 );
not U_inv966 ( n73622, P2_P2_INSTQUEUE_REG_9__1_ );
dff P2_P2_INSTQUEUE_REG_10__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__1_, n12826 );
not U_inv967 ( n73631, P2_P2_INSTQUEUE_REG_10__1_ );
dff P2_P2_INSTQUEUE_REG_11__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__1_, n12786 );
not U_inv968 ( n73626, P2_P2_INSTQUEUE_REG_11__1_ );
dff P2_P2_INSTQUEUE_REG_12__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__1_, n12746 );
not U_inv969 ( n73604, P2_P2_INSTQUEUE_REG_12__1_ );
dff P2_P2_INSTQUEUE_REG_13__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__1_, n12706 );
not U_inv970 ( n73617, P2_P2_INSTQUEUE_REG_13__1_ );
dff P2_P2_INSTQUEUE_REG_14__1__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__1_, n12666 );
not U_inv971 ( n73629, P2_P2_INSTQUEUE_REG_14__1_ );
dff P2_P1_LWORD_REG_14__reg ( clk, reset, P2_P1_LWORD_REG_14_, n15856 );
not U_inv972 ( n75654, P2_P1_LWORD_REG_14_ );
dff P2_P1_DATAO_REG_14__reg ( clk, reset, P2_P1_DATAO_REG_14_, n16076 );
dff P2_BUF1_REG_14__reg ( clk, reset, P2_BUF1_REG_14_, n531 );
not U_inv973 ( n75429, P2_BUF1_REG_14_ );
dff P2_P1_EAX_REG_30__reg ( clk, reset, P2_P1_EAX_REG_30_, n16316 );
not U_inv974 ( n75404, P2_P1_EAX_REG_30_ );
dff P2_P1_UWORD_REG_14__reg ( clk, reset, P2_P1_UWORD_REG_14_, n15931 );
not U_inv975 ( n75573, P2_P1_UWORD_REG_14_ );
dff P2_P1_DATAO_REG_30__reg ( clk, reset, P2_P1_DATAO_REG_30_, n16156 );
not U_inv976 ( n73428, P2_P1_DATAO_REG_30_ );
dff P2_BUF1_REG_30__reg ( clk, reset, P2_BUF1_REG_30_, n611 );
not U_inv977 ( n75406, P2_BUF1_REG_30_ );
dff P2_P1_EBX_REG_14__reg ( clk, reset, P2_P1_EBX_REG_14_, n16396 );
not U_inv978 ( n74795, P2_P1_EBX_REG_14_ );
dff P2_BUF2_REG_22__reg ( clk, reset, P2_BUF2_REG_22_, n731 );
not U_inv979 ( n75355, P2_BUF2_REG_22_ );
dff P2_P2_LWORD_REG_6__reg ( clk, reset, P2_P2_LWORD_REG_6_, n13651 );
not U_inv980 ( n75614, P2_P2_LWORD_REG_6_ );
dff P2_P2_DATAO_REG_6__reg ( clk, reset, P2_P2_DATAO_REG_6_, n13791 );
not U_inv981 ( n75520, P2_P2_DATAO_REG_6_ );
dff P2_BUF2_REG_6__reg ( clk, reset, P2_BUF2_REG_6_, n651 );
not U_inv982 ( n75290, P2_BUF2_REG_6_ );
dff P2_P3_UWORD_REG_6__reg ( clk, reset, P2_P3_UWORD_REG_6_, n11481 );
not U_inv983 ( n75467, P2_P3_UWORD_REG_6_ );
dff P2_P3_DATAO_REG_22__reg ( clk, reset, P2_P3_DATAO_REG_22_, n11626 );
dff P2_P3_LWORD_REG_6__reg ( clk, reset, P2_P3_LWORD_REG_6_, n11406 );
not U_inv984 ( n75613, P2_P3_LWORD_REG_6_ );
dff P2_P3_DATAO_REG_6__reg ( clk, reset, P2_P3_DATAO_REG_6_, n11546 );
dff P2_P2_INSTQUEUE_REG_7__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__6_, n12921 );
not U_inv985 ( n74086, P2_P2_INSTQUEUE_REG_7__6_ );
dff P2_P2_INSTQUEUE_REG_0__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__6_, n13201 );
not U_inv986 ( n74028, P2_P2_INSTQUEUE_REG_0__6_ );
dff P2_P2_INSTQUEUE_REG_1__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__6_, n13161 );
not U_inv987 ( n74067, P2_P2_INSTQUEUE_REG_1__6_ );
dff P2_P2_INSTQUEUE_REG_2__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__6_, n13121 );
not U_inv988 ( n74080, P2_P2_INSTQUEUE_REG_2__6_ );
dff P2_P2_INSTQUEUE_REG_3__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__6_, n13081 );
not U_inv989 ( n74054, P2_P2_INSTQUEUE_REG_3__6_ );
dff P2_P2_INSTQUEUE_REG_5__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__6_, n13001 );
not U_inv990 ( n74109, P2_P2_INSTQUEUE_REG_5__6_ );
dff P2_P2_INSTQUEUE_REG_6__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__6_, n12961 );
not U_inv991 ( n74116, P2_P2_INSTQUEUE_REG_6__6_ );
dff P2_P2_INSTQUEUE_REG_8__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__6_, n12881 );
not U_inv992 ( n74077, P2_P2_INSTQUEUE_REG_8__6_ );
dff P2_P2_INSTQUEUE_REG_9__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__6_, n12841 );
not U_inv993 ( n74113, P2_P2_INSTQUEUE_REG_9__6_ );
dff P2_P2_INSTQUEUE_REG_10__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__6_, n12801 );
not U_inv994 ( n74119, P2_P2_INSTQUEUE_REG_10__6_ );
dff P2_P2_INSTQUEUE_REG_11__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__6_, n12761 );
not U_inv995 ( n74095, P2_P2_INSTQUEUE_REG_11__6_ );
dff P2_P2_INSTQUEUE_REG_12__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__6_, n12721 );
not U_inv996 ( n74050, P2_P2_INSTQUEUE_REG_12__6_ );
dff P2_P2_INSTQUEUE_REG_13__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__6_, n12681 );
not U_inv997 ( n74075, P2_P2_INSTQUEUE_REG_13__6_ );
dff P2_P2_INSTQUEUE_REG_14__6__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__6_, n12641 );
not U_inv998 ( n74091, P2_P2_INSTQUEUE_REG_14__6_ );
dff P2_P2_LWORD_REG_3__reg ( clk, reset, P2_P2_LWORD_REG_3_, n13666 );
not U_inv999 ( n75612, P2_P2_LWORD_REG_3_ );
dff P2_P2_DATAO_REG_3__reg ( clk, reset, P2_P2_DATAO_REG_3_, n13776 );
not U_inv1000 ( n75521, P2_P2_DATAO_REG_3_ );
dff P2_BUF2_REG_3__reg ( clk, reset, P2_BUF2_REG_3_, n636 );
not U_inv1001 ( n75289, P2_BUF2_REG_3_ );
dff P2_P3_LWORD_REG_3__reg ( clk, reset, P2_P3_LWORD_REG_3_, n11421 );
not U_inv1002 ( n75611, P2_P3_LWORD_REG_3_ );
dff P2_P3_DATAO_REG_3__reg ( clk, reset, P2_P3_DATAO_REG_3_, n11531 );
dff P2_P2_INSTQUEUE_REG_7__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__3_, n12936 );
not U_inv1003 ( n73778, P2_P2_INSTQUEUE_REG_7__3_ );
dff P2_P2_INSTQUEUE_REG_0__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__3_, n13216 );
not U_inv1004 ( n73751, P2_P2_INSTQUEUE_REG_0__3_ );
dff P2_P2_EBX_REG_3__reg ( clk, reset, P2_P2_EBX_REG_3_, n14096 );
not U_inv1005 ( n73147, P2_P2_EBX_REG_3_ );
dff P2_P2_EBX_REG_4__reg ( clk, reset, P2_P2_EBX_REG_4_, n14101 );
not U_inv1006 ( n74573, P2_P2_EBX_REG_4_ );
dff P2_P2_INSTQUEUE_REG_1__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__3_, n13176 );
not U_inv1007 ( n73764, P2_P2_INSTQUEUE_REG_1__3_ );
dff P2_P2_INSTQUEUE_REG_2__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__3_, n13136 );
not U_inv1008 ( n73775, P2_P2_INSTQUEUE_REG_2__3_ );
dff P2_P2_INSTQUEUE_REG_3__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__3_, n13096 );
not U_inv1009 ( n73757, P2_P2_INSTQUEUE_REG_3__3_ );
dff P2_P2_INSTQUEUE_REG_4__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__3_, n13056 );
not U_inv1010 ( n73766, P2_P2_INSTQUEUE_REG_4__3_ );
dff P2_P2_INSTQUEUE_REG_5__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__3_, n13016 );
not U_inv1011 ( n73787, P2_P2_INSTQUEUE_REG_5__3_ );
dff P2_P2_INSTQUEUE_REG_6__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__3_, n12976 );
not U_inv1012 ( n73793, P2_P2_INSTQUEUE_REG_6__3_ );
dff P2_P2_INSTQUEUE_REG_8__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__3_, n12896 );
not U_inv1013 ( n73772, P2_P2_INSTQUEUE_REG_8__3_ );
dff P2_P2_INSTQUEUE_REG_9__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__3_, n12856 );
not U_inv1014 ( n73790, P2_P2_INSTQUEUE_REG_9__3_ );
dff P2_P2_INSTQUEUE_REG_10__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__3_, n12816 );
not U_inv1015 ( n73796, P2_P2_INSTQUEUE_REG_10__3_ );
dff P2_P2_INSTQUEUE_REG_11__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__3_, n12776 );
not U_inv1016 ( n73784, P2_P2_INSTQUEUE_REG_11__3_ );
dff P2_P2_INSTQUEUE_REG_12__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__3_, n12736 );
not U_inv1017 ( n73754, P2_P2_INSTQUEUE_REG_12__3_ );
dff P2_P2_INSTQUEUE_REG_13__3__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__3_, n12696 );
not U_inv1018 ( n73770, P2_P2_INSTQUEUE_REG_13__3_ );
dff P2_P2_INSTQUEUE_REG_15__3__reg ( clk, reset, ex_wire185, n12616 );
not U_inv1019 ( n73760, ex_wire185 );
dff P2_P1_LWORD_REG_1__reg ( clk, reset, P2_P1_LWORD_REG_1_, n15921 );
not U_inv1020 ( n75665, P2_P1_LWORD_REG_1_ );
dff P2_BUF2_REG_21__reg ( clk, reset, P2_BUF2_REG_21_, n726 );
not U_inv1021 ( n75356, P2_BUF2_REG_21_ );
dff P2_P2_INSTQUEUE_REG_0__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_0__5_, n13206 );
not U_inv1022 ( n73900, P2_P2_INSTQUEUE_REG_0__5_ );
dff P2_P2_EBX_REG_5__reg ( clk, reset, P2_P2_EBX_REG_5_, n14106 );
not U_inv1023 ( n73155, P2_P2_EBX_REG_5_ );
dff P2_P2_EBX_REG_6__reg ( clk, reset, P2_P2_EBX_REG_6_, n14111 );
not U_inv1024 ( n74606, P2_P2_EBX_REG_6_ );
dff P2_P2_EBX_REG_7__reg ( clk, reset, P2_P2_EBX_REG_7_, n14116 );
not U_inv1025 ( n73173, P2_P2_EBX_REG_7_ );
dff P2_P2_EBX_REG_8__reg ( clk, reset, P2_P2_EBX_REG_8_, n14121 );
not U_inv1026 ( n74669, P2_P2_EBX_REG_8_ );
dff P2_P2_INSTQUEUE_REG_1__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_1__5_, n13166 );
not U_inv1027 ( n73915, P2_P2_INSTQUEUE_REG_1__5_ );
dff P2_P2_INSTQUEUE_REG_2__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_2__5_, n13126 );
not U_inv1028 ( n73926, P2_P2_INSTQUEUE_REG_2__5_ );
dff P2_P2_INSTQUEUE_REG_3__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_3__5_, n13086 );
not U_inv1029 ( n73906, P2_P2_INSTQUEUE_REG_3__5_ );
dff P2_P2_INSTQUEUE_REG_4__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_4__5_, n13046 );
not U_inv1030 ( n73917, P2_P2_INSTQUEUE_REG_4__5_ );
dff P2_P2_INSTQUEUE_REG_7__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_7__5_, n12926 );
not U_inv1031 ( n73929, P2_P2_INSTQUEUE_REG_7__5_ );
dff P2_P2_INSTQUEUE_REG_5__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_5__5_, n13006 );
not U_inv1032 ( n73938, P2_P2_INSTQUEUE_REG_5__5_ );
dff P2_P2_INSTQUEUE_REG_6__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_6__5_, n12966 );
not U_inv1033 ( n73944, P2_P2_INSTQUEUE_REG_6__5_ );
dff P2_P2_INSTQUEUE_REG_8__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_8__5_, n12886 );
not U_inv1034 ( n73923, P2_P2_INSTQUEUE_REG_8__5_ );
dff P2_P2_INSTQUEUE_REG_9__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_9__5_, n12846 );
not U_inv1035 ( n73941, P2_P2_INSTQUEUE_REG_9__5_ );
dff P2_P2_INSTQUEUE_REG_10__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_10__5_, n12806 );
not U_inv1036 ( n73947, P2_P2_INSTQUEUE_REG_10__5_ );
dff P2_P2_INSTQUEUE_REG_11__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_11__5_, n12766 );
not U_inv1037 ( n73935, P2_P2_INSTQUEUE_REG_11__5_ );
dff P2_P2_INSTQUEUE_REG_12__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_12__5_, n12726 );
not U_inv1038 ( n73903, P2_P2_INSTQUEUE_REG_12__5_ );
dff P2_P2_INSTQUEUE_REG_13__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_13__5_, n12686 );
not U_inv1039 ( n73921, P2_P2_INSTQUEUE_REG_13__5_ );
dff P2_P2_INSTQUEUE_REG_14__5__reg ( clk, reset, P2_P2_INSTQUEUE_REG_14__5_, n12646 );
not U_inv1040 ( n73932, P2_P2_INSTQUEUE_REG_14__5_ );
dff P2_P2_EAX_REG_30__reg ( clk, reset, P2_P2_EAX_REG_30_, n14071 );
not U_inv1041 ( n75402, P2_P2_EAX_REG_30_ );
dff P2_P3_INSTQUEUE_REG_14__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__5_, n10401 );
not U_inv1042 ( n73930, P2_P3_INSTQUEUE_REG_14__5_ );
dff P2_P3_INSTQUEUE_REG_0__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__5_, n10961 );
not U_inv1043 ( n73898, P2_P3_INSTQUEUE_REG_0__5_ );
dff P2_P3_INSTQUEUE_REG_1__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__5_, n10921 );
not U_inv1044 ( n73912, P2_P3_INSTQUEUE_REG_1__5_ );
dff P2_P3_INSTQUEUE_REG_2__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__5_, n10881 );
not U_inv1045 ( n73924, P2_P3_INSTQUEUE_REG_2__5_ );
dff P2_P3_INSTQUEUE_REG_3__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__5_, n10841 );
not U_inv1046 ( n73904, P2_P3_INSTQUEUE_REG_3__5_ );
dff P2_P3_INSTQUEUE_REG_4__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__5_, n10801 );
not U_inv1047 ( n73913, P2_P3_INSTQUEUE_REG_4__5_ );
dff P2_P3_INSTQUEUE_REG_5__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__5_, n10761 );
not U_inv1048 ( n73936, P2_P3_INSTQUEUE_REG_5__5_ );
dff P2_P3_INSTQUEUE_REG_6__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__5_, n10721 );
not U_inv1049 ( n73942, P2_P3_INSTQUEUE_REG_6__5_ );
dff P2_P3_INSTQUEUE_REG_7__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__5_, n10681 );
not U_inv1050 ( n73927, P2_P3_INSTQUEUE_REG_7__5_ );
dff P2_P3_INSTQUEUE_REG_8__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__5_, n10641 );
not U_inv1051 ( n73919, P2_P3_INSTQUEUE_REG_8__5_ );
dff P2_P3_INSTQUEUE_REG_9__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__5_, n10601 );
not U_inv1052 ( n73939, P2_P3_INSTQUEUE_REG_9__5_ );
dff P2_P3_INSTQUEUE_REG_10__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__5_, n10561 );
not U_inv1053 ( n73945, P2_P3_INSTQUEUE_REG_10__5_ );
dff P2_P3_INSTQUEUE_REG_11__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__5_, n10521 );
not U_inv1054 ( n73933, P2_P3_INSTQUEUE_REG_11__5_ );
dff P2_P3_INSTQUEUE_REG_12__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__5_, n10481 );
not U_inv1055 ( n73901, P2_P3_INSTQUEUE_REG_12__5_ );
dff P2_P3_INSTQUEUE_REG_13__5__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__5_, n10441 );
not U_inv1056 ( n73918, P2_P3_INSTQUEUE_REG_13__5_ );
dff P2_P3_INSTQUEUE_REG_15__5__reg ( clk, reset, ex_wire186, n10361 );
not U_inv1057 ( n73907, ex_wire186 );
dff P2_P2_EBX_REG_9__reg ( clk, reset, P2_P2_EBX_REG_9_, n14126 );
not U_inv1058 ( n73203, P2_P2_EBX_REG_9_ );
dff P2_P2_UWORD_REG_7__reg ( clk, reset, P2_P2_UWORD_REG_7_, n13721 );
not U_inv1059 ( n75466, P2_P2_UWORD_REG_7_ );
dff P2_P2_DATAO_REG_23__reg ( clk, reset, P2_P2_DATAO_REG_23_, n13876 );
not U_inv1060 ( n75526, P2_P2_DATAO_REG_23_ );
dff P2_BUF2_REG_23__reg ( clk, reset, P2_BUF2_REG_23_, n736 );
not U_inv1061 ( n75354, P2_BUF2_REG_23_ );
dff P2_P3_INSTQUEUE_REG_5__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__7_, n10751 );
not U_inv1062 ( n74205, P2_P3_INSTQUEUE_REG_5__7_ );
dff P2_P3_INSTQUEUE_REG_6__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__7_, n10711 );
not U_inv1063 ( n74211, P2_P3_INSTQUEUE_REG_6__7_ );
dff P2_P3_INSTQUEUE_REG_8__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__7_, n10631 );
not U_inv1064 ( n74192, P2_P3_INSTQUEUE_REG_8__7_ );
dff P2_P3_INSTQUEUE_REG_9__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__7_, n10591 );
not U_inv1065 ( n74208, P2_P3_INSTQUEUE_REG_9__7_ );
dff P2_P3_INSTQUEUE_REG_10__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__7_, n10551 );
not U_inv1066 ( n74214, P2_P3_INSTQUEUE_REG_10__7_ );
dff P2_P3_INSTQUEUE_REG_11__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__7_, n10511 );
not U_inv1067 ( n74202, P2_P3_INSTQUEUE_REG_11__7_ );
dff P2_P3_INSTQUEUE_REG_12__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__7_, n10471 );
not U_inv1068 ( n74174, P2_P3_INSTQUEUE_REG_12__7_ );
dff P2_P3_INSTQUEUE_REG_13__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__7_, n10431 );
not U_inv1069 ( n74189, P2_P3_INSTQUEUE_REG_13__7_ );
dff P2_P3_INSTQUEUE_REG_14__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__7_, n10391 );
not U_inv1070 ( n74199, P2_P3_INSTQUEUE_REG_14__7_ );
dff P2_P3_INSTQUEUE_REG_0__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__7_, n10951 );
not U_inv1071 ( n74167, P2_P3_INSTQUEUE_REG_0__7_ );
dff P2_P3_INSTQUEUE_REG_1__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__7_, n10911 );
not U_inv1072 ( n74180, P2_P3_INSTQUEUE_REG_1__7_ );
dff P2_P3_INSTQUEUE_REG_2__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__7_, n10871 );
not U_inv1073 ( n74186, P2_P3_INSTQUEUE_REG_2__7_ );
dff P2_P3_INSTQUEUE_REG_3__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__7_, n10831 );
not U_inv1074 ( n74171, P2_P3_INSTQUEUE_REG_3__7_ );
dff P2_P3_INSTQUEUE_REG_4__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__7_, n10791 );
not U_inv1075 ( n74181, P2_P3_INSTQUEUE_REG_4__7_ );
dff P2_P3_INSTQUEUE_REG_7__7__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__7_, n10671 );
not U_inv1076 ( n74195, P2_P3_INSTQUEUE_REG_7__7_ );
dff P2_P3_INSTQUEUE_REG_14__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__6_, n10396 );
not U_inv1077 ( n74090, P2_P3_INSTQUEUE_REG_14__6_ );
dff P2_P3_INSTQUEUE_REG_0__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__6_, n10956 );
not U_inv1078 ( n74027, P2_P3_INSTQUEUE_REG_0__6_ );
dff P2_P3_INSTQUEUE_REG_1__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__6_, n10916 );
not U_inv1079 ( n74065, P2_P3_INSTQUEUE_REG_1__6_ );
dff P2_P3_INSTQUEUE_REG_2__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__6_, n10876 );
not U_inv1080 ( n74079, P2_P3_INSTQUEUE_REG_2__6_ );
dff P2_P3_INSTQUEUE_REG_3__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__6_, n10836 );
not U_inv1081 ( n74053, P2_P3_INSTQUEUE_REG_3__6_ );
dff P2_P3_INSTQUEUE_REG_4__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__6_, n10796 );
not U_inv1082 ( n74066, P2_P3_INSTQUEUE_REG_4__6_ );
dff P2_P3_INSTQUEUE_REG_5__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__6_, n10756 );
not U_inv1083 ( n74108, P2_P3_INSTQUEUE_REG_5__6_ );
dff P2_P3_INSTQUEUE_REG_6__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__6_, n10716 );
not U_inv1084 ( n74115, P2_P3_INSTQUEUE_REG_6__6_ );
dff P2_P3_INSTQUEUE_REG_7__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__6_, n10676 );
not U_inv1085 ( n74083, P2_P3_INSTQUEUE_REG_7__6_ );
dff P2_P3_INSTQUEUE_REG_8__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__6_, n10636 );
not U_inv1086 ( n74074, P2_P3_INSTQUEUE_REG_8__6_ );
dff P2_P3_INSTQUEUE_REG_9__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__6_, n10596 );
not U_inv1087 ( n74112, P2_P3_INSTQUEUE_REG_9__6_ );
dff P2_P3_INSTQUEUE_REG_10__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__6_, n10556 );
not U_inv1088 ( n74118, P2_P3_INSTQUEUE_REG_10__6_ );
dff P2_P3_INSTQUEUE_REG_11__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__6_, n10516 );
not U_inv1089 ( n74094, P2_P3_INSTQUEUE_REG_11__6_ );
dff P2_P3_INSTQUEUE_REG_12__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__6_, n10476 );
not U_inv1090 ( n74049, P2_P3_INSTQUEUE_REG_12__6_ );
dff P2_P3_INSTQUEUE_REG_13__6__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__6_, n10436 );
not U_inv1091 ( n74073, P2_P3_INSTQUEUE_REG_13__6_ );
dff P2_P3_INSTQUEUE_REG_15__6__reg ( clk, reset, ex_wire187, n10356 );
not U_inv1092 ( n74056, ex_wire187 );
dff P2_P3_PHYADDRPOINTER_REG_0__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_0_, n11201 );
not U_inv1093 ( n75223, P2_P3_PHYADDRPOINTER_REG_0_ );
dff P2_P2_EAX_REG_15__reg ( clk, reset, P2_P2_EAX_REG_15_, n13996 );
not U_inv1094 ( n74779, P2_P2_EAX_REG_15_ );
dff P2_P3_INSTQUEUE_REG_5__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__3_, n10771 );
not U_inv1095 ( n73785, P2_P3_INSTQUEUE_REG_5__3_ );
dff P2_P3_INSTQUEUE_REG_6__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__3_, n10731 );
not U_inv1096 ( n73791, P2_P3_INSTQUEUE_REG_6__3_ );
dff P2_P3_INSTQUEUE_REG_8__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__3_, n10651 );
not U_inv1097 ( n73768, P2_P3_INSTQUEUE_REG_8__3_ );
dff P2_P3_INSTQUEUE_REG_9__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__3_, n10611 );
not U_inv1098 ( n73788, P2_P3_INSTQUEUE_REG_9__3_ );
dff P2_P3_INSTQUEUE_REG_10__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__3_, n10571 );
not U_inv1099 ( n73794, P2_P3_INSTQUEUE_REG_10__3_ );
dff P2_P3_INSTQUEUE_REG_11__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__3_, n10531 );
not U_inv1100 ( n73782, P2_P3_INSTQUEUE_REG_11__3_ );
dff P2_P3_INSTQUEUE_REG_12__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__3_, n10491 );
not U_inv1101 ( n73752, P2_P3_INSTQUEUE_REG_12__3_ );
dff P2_P3_INSTQUEUE_REG_13__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__3_, n10451 );
not U_inv1102 ( n73767, P2_P3_INSTQUEUE_REG_13__3_ );
dff P2_P3_INSTQUEUE_REG_14__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__3_, n10411 );
not U_inv1103 ( n73779, P2_P3_INSTQUEUE_REG_14__3_ );
dff P2_P3_INSTQUEUE_REG_0__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__3_, n10971 );
not U_inv1104 ( n73749, P2_P3_INSTQUEUE_REG_0__3_ );
dff P2_P3_INSTQUEUE_REG_1__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__3_, n10931 );
not U_inv1105 ( n73761, P2_P3_INSTQUEUE_REG_1__3_ );
dff P2_P3_INSTQUEUE_REG_2__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__3_, n10891 );
not U_inv1106 ( n73773, P2_P3_INSTQUEUE_REG_2__3_ );
dff P2_P3_INSTQUEUE_REG_3__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__3_, n10851 );
not U_inv1107 ( n73755, P2_P3_INSTQUEUE_REG_3__3_ );
dff P2_P3_INSTQUEUE_REG_4__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__3_, n10811 );
not U_inv1108 ( n73762, P2_P3_INSTQUEUE_REG_4__3_ );
dff P2_P3_INSTQUEUE_REG_7__3__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__3_, n10691 );
not U_inv1109 ( n73776, P2_P3_INSTQUEUE_REG_7__3_ );
dff P2_P3_INSTQUEUE_REG_15__3__reg ( clk, reset, ex_wire188, n10371 );
not U_inv1110 ( n73758, ex_wire188 );
dff P2_P3_EAX_REG_11__reg ( clk, reset, P2_P3_EAX_REG_11_, n11731 );
not U_inv1111 ( n74675, P2_P3_EAX_REG_11_ );
dff P2_P3_LWORD_REG_11__reg ( clk, reset, P2_P3_LWORD_REG_11_, n11381 );
not U_inv1112 ( n75610, P2_P3_LWORD_REG_11_ );
dff P2_P3_DATAO_REG_11__reg ( clk, reset, P2_P3_DATAO_REG_11_, n11571 );
dff P2_P3_EAX_REG_12__reg ( clk, reset, P2_P3_EAX_REG_12_, n11736 );
not U_inv1113 ( n75269, P2_P3_EAX_REG_12_ );
dff P2_P3_LWORD_REG_12__reg ( clk, reset, P2_P3_LWORD_REG_12_, n11376 );
not U_inv1114 ( n75609, P2_P3_LWORD_REG_12_ );
dff P2_P3_DATAO_REG_12__reg ( clk, reset, P2_P3_DATAO_REG_12_, n11576 );
dff P2_P3_EAX_REG_13__reg ( clk, reset, P2_P3_EAX_REG_13_, n11741 );
not U_inv1115 ( n74730, P2_P3_EAX_REG_13_ );
dff P2_P3_LWORD_REG_13__reg ( clk, reset, P2_P3_LWORD_REG_13_, n11371 );
not U_inv1116 ( n75608, P2_P3_LWORD_REG_13_ );
dff P2_P3_DATAO_REG_13__reg ( clk, reset, P2_P3_DATAO_REG_13_, n11581 );
dff P2_P3_EAX_REG_14__reg ( clk, reset, P2_P3_EAX_REG_14_, n11746 );
not U_inv1117 ( n75268, P2_P3_EAX_REG_14_ );
dff P2_P3_LWORD_REG_14__reg ( clk, reset, P2_P3_LWORD_REG_14_, n11366 );
not U_inv1118 ( n75607, P2_P3_LWORD_REG_14_ );
dff P2_P3_DATAO_REG_14__reg ( clk, reset, P2_P3_DATAO_REG_14_, n11586 );
dff P2_P2_EBX_REG_10__reg ( clk, reset, P2_P2_EBX_REG_10_, n14131 );
not U_inv1119 ( n74724, P2_P2_EBX_REG_10_ );
dff P2_P2_EBX_REG_11__reg ( clk, reset, P2_P2_EBX_REG_11_, n14136 );
not U_inv1120 ( n73211, P2_P2_EBX_REG_11_ );
dff P2_P2_EBX_REG_12__reg ( clk, reset, P2_P2_EBX_REG_12_, n14141 );
not U_inv1121 ( n74767, P2_P2_EBX_REG_12_ );
dff P2_P2_EBX_REG_13__reg ( clk, reset, P2_P2_EBX_REG_13_, n14146 );
not U_inv1122 ( n73230, P2_P2_EBX_REG_13_ );
dff P2_P2_EBX_REG_14__reg ( clk, reset, P2_P2_EBX_REG_14_, n14151 );
not U_inv1123 ( n74797, P2_P2_EBX_REG_14_ );
dff P2_P2_EBX_REG_15__reg ( clk, reset, P2_P2_EBX_REG_15_, n14156 );
not U_inv1124 ( n73245, P2_P2_EBX_REG_15_ );
dff P2_P2_EBX_REG_16__reg ( clk, reset, P2_P2_EBX_REG_16_, n14161 );
not U_inv1125 ( n74836, P2_P2_EBX_REG_16_ );
dff P2_P2_EBX_REG_17__reg ( clk, reset, P2_P2_EBX_REG_17_, n14166 );
not U_inv1126 ( n73259, P2_P2_EBX_REG_17_ );
dff P2_P2_EBX_REG_18__reg ( clk, reset, P2_P2_EBX_REG_18_, n14171 );
not U_inv1127 ( n74897, P2_P2_EBX_REG_18_ );
dff P2_P2_EBX_REG_19__reg ( clk, reset, P2_P2_EBX_REG_19_, n14176 );
not U_inv1128 ( n73273, P2_P2_EBX_REG_19_ );
dff P2_P2_EBX_REG_20__reg ( clk, reset, P2_P2_EBX_REG_20_, n14181 );
not U_inv1129 ( n74937, P2_P2_EBX_REG_20_ );
dff P2_P2_EBX_REG_21__reg ( clk, reset, P2_P2_EBX_REG_21_, n14186 );
not U_inv1130 ( n73286, P2_P2_EBX_REG_21_ );
dff P2_P2_EBX_REG_22__reg ( clk, reset, P2_P2_EBX_REG_22_, n14191 );
not U_inv1131 ( n74983, P2_P2_EBX_REG_22_ );
dff P2_P2_EBX_REG_23__reg ( clk, reset, P2_P2_EBX_REG_23_, n14196 );
not U_inv1132 ( n73302, P2_P2_EBX_REG_23_ );
dff P2_P2_EBX_REG_24__reg ( clk, reset, P2_P2_EBX_REG_24_, n14201 );
not U_inv1133 ( n75026, P2_P2_EBX_REG_24_ );
dff P2_P2_EBX_REG_25__reg ( clk, reset, P2_P2_EBX_REG_25_, n14206 );
not U_inv1134 ( n73314, P2_P2_EBX_REG_25_ );
dff P2_P2_EBX_REG_26__reg ( clk, reset, P2_P2_EBX_REG_26_, n14211 );
not U_inv1135 ( n75076, P2_P2_EBX_REG_26_ );
dff P2_P2_EBX_REG_27__reg ( clk, reset, P2_P2_EBX_REG_27_, n14216 );
not U_inv1136 ( n75174, P2_P2_EBX_REG_27_ );
dff P2_P2_EBX_REG_28__reg ( clk, reset, P2_P2_EBX_REG_28_, n14221 );
not U_inv1137 ( n73389, P2_P2_EBX_REG_28_ );
dff P2_P2_EBX_REG_29__reg ( clk, reset, P2_P2_EBX_REG_29_, n14226 );
not U_inv1138 ( n75184, P2_P2_EBX_REG_29_ );
dff P2_P2_EBX_REG_30__reg ( clk, reset, P2_P2_EBX_REG_30_, n14231 );
not U_inv1139 ( n75216, P2_P2_EBX_REG_30_ );
dff P2_P2_EBX_REG_31__reg ( clk, reset, P2_P2_EBX_REG_31_, n14236 );
dff P2_P3_INSTQUEUE_REG_7__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__2_, n10696 );
not U_inv1140 ( n73722, P2_P3_INSTQUEUE_REG_7__2_ );
dff P2_P3_INSTQUEUE_REG_0__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__2_, n10976 );
not U_inv1141 ( n73666, P2_P3_INSTQUEUE_REG_0__2_ );
dff P2_P3_INSTQUEUE_REG_1__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__2_, n10936 );
not U_inv1142 ( n73707, P2_P3_INSTQUEUE_REG_1__2_ );
dff P2_P3_INSTQUEUE_REG_2__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__2_, n10896 );
not U_inv1143 ( n73728, P2_P3_INSTQUEUE_REG_2__2_ );
dff P2_P3_INSTQUEUE_REG_3__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__2_, n10856 );
not U_inv1144 ( n73714, P2_P3_INSTQUEUE_REG_3__2_ );
dff P2_P3_INSTQUEUE_REG_4__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__2_, n10816 );
not U_inv1145 ( n73701, P2_P3_INSTQUEUE_REG_4__2_ );
dff P2_P3_INSTQUEUE_REG_5__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__2_, n10776 );
not U_inv1146 ( n73711, P2_P3_INSTQUEUE_REG_5__2_ );
dff P2_P3_INSTQUEUE_REG_6__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__2_, n10736 );
not U_inv1147 ( n73734, P2_P3_INSTQUEUE_REG_6__2_ );
dff P2_P3_INSTQUEUE_REG_8__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__2_, n10656 );
not U_inv1148 ( n73719, P2_P3_INSTQUEUE_REG_8__2_ );
dff P2_P3_INSTQUEUE_REG_9__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__2_, n10616 );
not U_inv1149 ( n73731, P2_P3_INSTQUEUE_REG_9__2_ );
dff P2_P3_INSTQUEUE_REG_10__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__2_, n10576 );
not U_inv1150 ( n73743, P2_P3_INSTQUEUE_REG_10__2_ );
dff P2_P3_INSTQUEUE_REG_11__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__2_, n10536 );
not U_inv1151 ( n73737, P2_P3_INSTQUEUE_REG_11__2_ );
dff P2_P3_INSTQUEUE_REG_12__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__2_, n10496 );
not U_inv1152 ( n73710, P2_P3_INSTQUEUE_REG_12__2_ );
dff P2_P3_INSTQUEUE_REG_13__2__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__2_, n10456 );
not U_inv1153 ( n73725, P2_P3_INSTQUEUE_REG_13__2_ );
dff P2_P3_INSTQUEUE_REG_15__2__reg ( clk, reset, ex_wire189, n10376 );
not U_inv1154 ( n73746, ex_wire189 );
dff P2_P2_DATAO_REG_1__reg ( clk, reset, P2_P2_DATAO_REG_1_, n13766 );
not U_inv1155 ( n75523, P2_P2_DATAO_REG_1_ );
dff P2_BUF2_REG_1__reg ( clk, reset, P2_BUF2_REG_1_, n626 );
not U_inv1156 ( n75295, P2_BUF2_REG_1_ );
dff P2_P3_LWORD_REG_1__reg ( clk, reset, P2_P3_LWORD_REG_1_, n11431 );
not U_inv1157 ( n75605, P2_P3_LWORD_REG_1_ );
dff P2_P3_DATAO_REG_1__reg ( clk, reset, P2_P3_DATAO_REG_1_, n11521 );
dff P2_P3_INSTQUEUE_REG_7__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_7__1_, n10701 );
not U_inv1158 ( n73594, P2_P3_INSTQUEUE_REG_7__1_ );
dff P2_P3_INSTQUEUE_REG_0__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_0__1_, n10981 );
not U_inv1159 ( n73564, P2_P3_INSTQUEUE_REG_0__1_ );
dff P2_P3_EBX_REG_2__reg ( clk, reset, P2_P3_EBX_REG_2_, n11846 );
not U_inv1160 ( n74534, P2_P3_EBX_REG_2_ );
dff P2_P3_EBX_REG_3__reg ( clk, reset, P2_P3_EBX_REG_3_, n11851 );
not U_inv1161 ( n73146, P2_P3_EBX_REG_3_ );
dff P2_P3_EBX_REG_4__reg ( clk, reset, P2_P3_EBX_REG_4_, n11856 );
not U_inv1162 ( n74570, P2_P3_EBX_REG_4_ );
dff P2_P3_EBX_REG_5__reg ( clk, reset, P2_P3_EBX_REG_5_, n11861 );
not U_inv1163 ( n73154, P2_P3_EBX_REG_5_ );
dff P2_P3_EBX_REG_6__reg ( clk, reset, P2_P3_EBX_REG_6_, n11866 );
not U_inv1164 ( n74603, P2_P3_EBX_REG_6_ );
dff P2_P3_EBX_REG_7__reg ( clk, reset, P2_P3_EBX_REG_7_, n11871 );
not U_inv1165 ( n73172, P2_P3_EBX_REG_7_ );
dff P2_P3_EBX_REG_8__reg ( clk, reset, P2_P3_EBX_REG_8_, n11876 );
not U_inv1166 ( n74666, P2_P3_EBX_REG_8_ );
dff P2_P3_INSTQUEUE_REG_1__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_1__1_, n10941 );
not U_inv1167 ( n73585, P2_P3_INSTQUEUE_REG_1__1_ );
dff P2_P3_INSTQUEUE_REG_2__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_2__1_, n10901 );
not U_inv1168 ( n73596, P2_P3_INSTQUEUE_REG_2__1_ );
dff P2_P3_INSTQUEUE_REG_3__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_3__1_, n10861 );
not U_inv1169 ( n73589, P2_P3_INSTQUEUE_REG_3__1_ );
dff P2_P3_INSTQUEUE_REG_4__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_4__1_, n10821 );
not U_inv1170 ( n73583, P2_P3_INSTQUEUE_REG_4__1_ );
dff P2_P3_INSTQUEUE_REG_5__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_5__1_, n10781 );
not U_inv1171 ( n73590, P2_P3_INSTQUEUE_REG_5__1_ );
dff P2_P3_INSTQUEUE_REG_6__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_6__1_, n10741 );
not U_inv1172 ( n73603, P2_P3_INSTQUEUE_REG_6__1_ );
dff P2_P3_INSTQUEUE_REG_8__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_8__1_, n10661 );
not U_inv1173 ( n73592, P2_P3_INSTQUEUE_REG_8__1_ );
dff P2_P3_INSTQUEUE_REG_9__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_9__1_, n10621 );
not U_inv1174 ( n73602, P2_P3_INSTQUEUE_REG_9__1_ );
dff P2_P3_INSTQUEUE_REG_10__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_10__1_, n10581 );
not U_inv1175 ( n73621, P2_P3_INSTQUEUE_REG_10__1_ );
dff P2_P3_INSTQUEUE_REG_11__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_11__1_, n10541 );
not U_inv1176 ( n73610, P2_P3_INSTQUEUE_REG_11__1_ );
dff P2_P3_INSTQUEUE_REG_12__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_12__1_, n10501 );
not U_inv1177 ( n73588, P2_P3_INSTQUEUE_REG_12__1_ );
dff P2_P3_INSTQUEUE_REG_13__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_13__1_, n10461 );
not U_inv1178 ( n73595, P2_P3_INSTQUEUE_REG_13__1_ );
dff P2_P3_INSTQUEUE_REG_14__1__reg ( clk, reset, P2_P3_INSTQUEUE_REG_14__1_, n10421 );
not U_inv1179 ( n73612, P2_P3_INSTQUEUE_REG_14__1_ );
dff P2_P3_EAX_REG_24__reg ( clk, reset, P2_P3_EAX_REG_24_, n11796 );
not U_inv1180 ( n75390, P2_P3_EAX_REG_24_ );
dff P2_P3_UWORD_REG_8__reg ( clk, reset, P2_P3_UWORD_REG_8_, n11471 );
not U_inv1181 ( n75558, P2_P3_UWORD_REG_8_ );
dff P2_P3_DATAO_REG_24__reg ( clk, reset, P2_P3_DATAO_REG_24_, n11636 );
dff P2_P3_EAX_REG_25__reg ( clk, reset, P2_P3_EAX_REG_25_, n11801 );
not U_inv1182 ( n75028, P2_P3_EAX_REG_25_ );
dff P2_P3_EAX_REG_26__reg ( clk, reset, P2_P3_EAX_REG_26_, n11806 );
not U_inv1183 ( n75389, P2_P3_EAX_REG_26_ );
dff P2_P3_UWORD_REG_10__reg ( clk, reset, P2_P3_UWORD_REG_10_, n11461 );
not U_inv1184 ( n75557, P2_P3_UWORD_REG_10_ );
dff P2_P3_DATAO_REG_26__reg ( clk, reset, P2_P3_DATAO_REG_26_, n11646 );
dff P2_P3_EAX_REG_27__reg ( clk, reset, P2_P3_EAX_REG_27_, n11811 );
not U_inv1185 ( n75346, P2_P3_EAX_REG_27_ );
dff P2_P3_UWORD_REG_11__reg ( clk, reset, P2_P3_UWORD_REG_11_, n11456 );
not U_inv1186 ( n75556, P2_P3_UWORD_REG_11_ );
dff P2_P3_DATAO_REG_27__reg ( clk, reset, P2_P3_DATAO_REG_27_, n11651 );
dff P2_P3_EAX_REG_28__reg ( clk, reset, P2_P3_EAX_REG_28_, n11816 );
not U_inv1187 ( n73390, P2_P3_EAX_REG_28_ );
dff P2_P3_UWORD_REG_12__reg ( clk, reset, P2_P3_UWORD_REG_12_, n11451 );
not U_inv1188 ( n75555, P2_P3_UWORD_REG_12_ );
dff P2_P3_DATAO_REG_28__reg ( clk, reset, P2_P3_DATAO_REG_28_, n11656 );
dff P2_P3_EAX_REG_29__reg ( clk, reset, P2_P3_EAX_REG_29_, n11821 );
not U_inv1189 ( n75204, P2_P3_EAX_REG_29_ );
dff P2_P3_EAX_REG_30__reg ( clk, reset, P2_P3_EAX_REG_30_, n11826 );
not U_inv1190 ( n75426, P2_P3_EAX_REG_30_ );
dff P2_P3_UWORD_REG_14__reg ( clk, reset, P2_P3_UWORD_REG_14_, n11441 );
not U_inv1191 ( n75554, P2_P3_UWORD_REG_14_ );
dff P2_P3_DATAO_REG_30__reg ( clk, reset, P2_P3_DATAO_REG_30_, n11666 );
dff P2_P3_UWORD_REG_13__reg ( clk, reset, P2_P3_UWORD_REG_13_, n11446 );
not U_inv1192 ( n75553, P2_P3_UWORD_REG_13_ );
dff P2_P3_DATAO_REG_29__reg ( clk, reset, P2_P3_DATAO_REG_29_, n11661 );
dff P2_P3_UWORD_REG_9__reg ( clk, reset, P2_P3_UWORD_REG_9_, n11466 );
not U_inv1193 ( n75552, P2_P3_UWORD_REG_9_ );
dff P2_P3_DATAO_REG_25__reg ( clk, reset, P2_P3_DATAO_REG_25_, n11641 );
dff P4_IR_REG_25__reg ( clk, reset, P4_IR_REG_25_, n2151 );
not U_inv1194 ( n75365, P4_IR_REG_25_ );
dff P4_IR_REG_26__reg ( clk, reset, P4_IR_REG_26_, n2156 );
not U_inv1195 ( n73505, P4_IR_REG_26_ );
dff P4_IR_REG_28__reg ( clk, reset, P4_IR_REG_28_, n2166 );
not U_inv1196 ( n73519, P4_IR_REG_28_ );
dff P4_IR_REG_29__reg ( clk, reset, P4_IR_REG_29_, n2171 );
not U_inv1197 ( n73058, P4_IR_REG_29_ );
dff P4_IR_REG_30__reg ( clk, reset, P4_IR_REG_30_, n2176 );
not U_inv1198 ( n75299, P4_IR_REG_30_ );
dff P4_IR_REG_27__reg ( clk, reset, P4_IR_REG_27_, n2161 );
not U_inv1199 ( n73051, P4_IR_REG_27_ );
dff P4_IR_REG_22__reg ( clk, reset, P4_IR_REG_22_, n2136 );
not U_inv1200 ( n73047, P4_IR_REG_22_ );
dff P4_IR_REG_24__reg ( clk, reset, P4_IR_REG_24_, n2146 );
not U_inv1201 ( n73050, P4_IR_REG_24_ );
dff P4_IR_REG_0__reg ( clk, reset, P4_IR_REG_0_, n2026 );
not U_inv1202 ( n73023, P4_IR_REG_0_ );
dff P4_IR_REG_1__reg ( clk, reset, P4_IR_REG_1_, n2031 );
not U_inv1203 ( n73535, P4_IR_REG_1_ );
dff P4_IR_REG_3__reg ( clk, reset, P4_IR_REG_3_, n2041 );
not U_inv1204 ( n73803, P4_IR_REG_3_ );
dff P4_IR_REG_5__reg ( clk, reset, P4_IR_REG_5_, n2051 );
not U_inv1205 ( n73948, P4_IR_REG_5_ );
dff P4_IR_REG_7__reg ( clk, reset, P4_IR_REG_7_, n2061 );
not U_inv1206 ( n74257, P4_IR_REG_7_ );
dff P4_IR_REG_9__reg ( clk, reset, P4_IR_REG_9_, n2071 );
not U_inv1207 ( n74298, P4_IR_REG_9_ );
dff P4_IR_REG_11__reg ( clk, reset, P4_IR_REG_11_, n2081 );
not U_inv1208 ( n74335, P4_IR_REG_11_ );
dff P4_IR_REG_13__reg ( clk, reset, P4_IR_REG_13_, n2091 );
not U_inv1209 ( n74390, P4_IR_REG_13_ );
dff P4_IR_REG_14__reg ( clk, reset, P4_IR_REG_14_, n2096 );
not U_inv1210 ( n75420, P4_IR_REG_14_ );
dff P4_IR_REG_12__reg ( clk, reset, P4_IR_REG_12_, n2086 );
not U_inv1211 ( n75419, P4_IR_REG_12_ );
dff P4_IR_REG_8__reg ( clk, reset, P4_IR_REG_8_, n2066 );
not U_inv1212 ( n75418, P4_IR_REG_8_ );
dff P4_IR_REG_6__reg ( clk, reset, P4_IR_REG_6_, n2056 );
not U_inv1213 ( n75425, P4_IR_REG_6_ );
dff P4_IR_REG_4__reg ( clk, reset, P4_IR_REG_4_, n2046 );
not U_inv1214 ( n75424, P4_IR_REG_4_ );
dff P4_IR_REG_2__reg ( clk, reset, P4_IR_REG_2_, n2036 );
not U_inv1215 ( n75423, P4_IR_REG_2_ );
dff P4_RD_REG_reg ( clk, reset, P4_RD_REG, n3241 );
dff P2_P3_EBX_REG_9__reg ( clk, reset, P2_P3_EBX_REG_9_, n11881 );
not U_inv1216 ( n73201, P2_P3_EBX_REG_9_ );
dff P2_P2_DATAO_REG_0__reg ( clk, reset, P2_P2_DATAO_REG_0_, n13761 );
not U_inv1217 ( n75527, P2_P2_DATAO_REG_0_ );
dff P2_P2_DATAWIDTH_REG_31__reg ( clk, reset, ex_wire190, n12571 );
not U_inv1218 ( n75138, ex_wire190 );
dff P2_P2_DATAWIDTH_REG_30__reg ( clk, reset, ex_wire191, n12566 );
not U_inv1219 ( n73338, ex_wire191 );
dff P2_P2_DATAWIDTH_REG_29__reg ( clk, reset, ex_wire192, n12561 );
not U_inv1220 ( n73326, ex_wire192 );
dff P2_P2_DATAWIDTH_REG_28__reg ( clk, reset, ex_wire193, n12556 );
not U_inv1221 ( n75082, ex_wire193 );
dff P2_P2_DATAWIDTH_REG_27__reg ( clk, reset, ex_wire194, n12551 );
not U_inv1222 ( n73352, ex_wire194 );
dff P2_P2_DATAWIDTH_REG_26__reg ( clk, reset, ex_wire195, n12546 );
not U_inv1223 ( n75126, ex_wire195 );
dff P2_P2_DATAWIDTH_REG_25__reg ( clk, reset, ex_wire196, n12541 );
not U_inv1224 ( n72976, ex_wire196 );
dff P2_P2_DATAWIDTH_REG_24__reg ( clk, reset, ex_wire197, n12536 );
not U_inv1225 ( n75095, ex_wire197 );
dff P2_P2_DATAWIDTH_REG_23__reg ( clk, reset, ex_wire198, n12531 );
not U_inv1226 ( n73380, ex_wire198 );
dff P2_P2_DATAWIDTH_REG_22__reg ( clk, reset, ex_wire199, n12526 );
not U_inv1227 ( n75162, ex_wire199 );
dff P2_P2_DATAWIDTH_REG_21__reg ( clk, reset, ex_wire200, n12521 );
not U_inv1228 ( n73358, ex_wire200 );
dff P2_P2_DATAWIDTH_REG_20__reg ( clk, reset, ex_wire201, n12516 );
not U_inv1229 ( n75132, ex_wire201 );
dff P2_P2_DATAWIDTH_REG_19__reg ( clk, reset, ex_wire202, n12511 );
not U_inv1230 ( n72997, ex_wire202 );
dff P2_P2_DATAWIDTH_REG_18__reg ( clk, reset, ex_wire203, n12506 );
not U_inv1231 ( n75168, ex_wire203 );
dff P2_P2_DATAWIDTH_REG_17__reg ( clk, reset, ex_wire204, n12501 );
not U_inv1232 ( n72989, ex_wire204 );
dff P2_P2_DATAWIDTH_REG_16__reg ( clk, reset, ex_wire205, n12496 );
not U_inv1233 ( n75144, ex_wire205 );
dff P2_P2_DATAWIDTH_REG_15__reg ( clk, reset, ex_wire206, n12491 );
not U_inv1234 ( n72985, ex_wire206 );
dff P2_P2_DATAWIDTH_REG_14__reg ( clk, reset, ex_wire207, n12486 );
not U_inv1235 ( n75120, ex_wire207 );
dff P2_P2_DATAWIDTH_REG_13__reg ( clk, reset, ex_wire208, n12481 );
not U_inv1236 ( n72975, ex_wire208 );
dff P2_P2_DATAWIDTH_REG_12__reg ( clk, reset, ex_wire209, n12476 );
not U_inv1237 ( n75094, ex_wire209 );
dff P2_P2_DATAWIDTH_REG_11__reg ( clk, reset, ex_wire210, n12471 );
not U_inv1238 ( n72979, ex_wire210 );
dff P2_P2_DATAWIDTH_REG_10__reg ( clk, reset, ex_wire211, n12466 );
not U_inv1239 ( n75100, ex_wire211 );
dff P2_P2_DATAWIDTH_REG_9__reg ( clk, reset, ex_wire212, n12461 );
not U_inv1240 ( n72993, ex_wire212 );
dff P2_P2_DATAWIDTH_REG_8__reg ( clk, reset, ex_wire213, n12456 );
not U_inv1241 ( n75150, ex_wire213 );
dff P2_P2_DATAWIDTH_REG_7__reg ( clk, reset, ex_wire214, n12451 );
not U_inv1242 ( n73344, ex_wire214 );
dff P2_P2_DATAWIDTH_REG_6__reg ( clk, reset, ex_wire215, n12446 );
not U_inv1243 ( n75114, ex_wire215 );
dff P2_P2_DATAWIDTH_REG_5__reg ( clk, reset, ex_wire216, n12441 );
not U_inv1244 ( n73374, ex_wire216 );
dff P2_P2_DATAWIDTH_REG_4__reg ( clk, reset, ex_wire217, n12436 );
not U_inv1245 ( n75156, ex_wire217 );
dff P2_P2_DATAWIDTH_REG_3__reg ( clk, reset, ex_wire218, n12431 );
not U_inv1246 ( n73364, ex_wire218 );
dff P2_P2_DATAWIDTH_REG_2__reg ( clk, reset, ex_wire219, n12426 );
not U_inv1247 ( n75108, ex_wire219 );
dff P2_P2_DATAWIDTH_REG_1__reg ( clk, reset, P2_P2_DATAWIDTH_REG_1_, n12421 );
dff P2_P2_M_IO_N_REG_reg ( clk, reset, P2_P2_M_IO_N_REG, n14451 );
dff P2_P2_W_R_N_REG_reg ( clk, reset, P2_P2_W_R_N_REG, n14421 );
dff P2_P2_ADDRESS_REG_16__reg ( clk, reset, P2_P2_ADDRESS_REG_16_, n12316 );
not U_inv1248 ( n74444, P2_P2_ADDRESS_REG_16_ );
dff P2_P2_ADDRESS_REG_22__reg ( clk, reset, P2_P2_ADDRESS_REG_22_, n12286 );
dff P2_P2_ADDRESS_REG_27__reg ( clk, reset, P2_P2_ADDRESS_REG_27_, n12261 );
dff P2_P2_ADDRESS_REG_28__reg ( clk, reset, P2_P2_ADDRESS_REG_28_, n12256 );
dff P2_P2_CODEFETCH_REG_reg ( clk, reset, P2_P2_CODEFETCH_REG, n14456 );
dff P2_P2_D_C_N_REG_reg ( clk, reset, P2_P2_D_C_N_REG, n14446 );
dff P2_P2_MORE_REG_reg ( clk, reset, P2_P2_MORE_REG, n14431 );
dff P2_P1_DATAO_REG_0__reg ( clk, reset, P2_P1_DATAO_REG_0_, n16006 );
dff P2_P1_ADDRESS_REG_4__reg ( clk, reset, P2_P1_ADDRESS_REG_4_, n14621 );
not U_inv1249 ( n73046, P2_P1_ADDRESS_REG_4_ );
dff P1_P1_STATEBS16_REG_reg ( clk, reset, P1_P1_STATEBS16_REG, n9946 );
not U_inv1250 ( n74906, P1_P1_STATEBS16_REG );
dff P1_P1_INSTQUEUEWR_ADDR_REG_1__reg ( clk, reset, P1_P1_INSTQUEUEWR_ADDR_REG_1_, n8786 );
not U_inv1251 ( n73141, P1_P1_INSTQUEUEWR_ADDR_REG_1_ );
dff P1_P1_INSTQUEUEWR_ADDR_REG_3__reg ( clk, reset, P1_P1_INSTQUEUEWR_ADDR_REG_3_, n8776 );
not U_inv1252 ( n74538, P1_P1_INSTQUEUEWR_ADDR_REG_3_ );
dff P1_P1_INSTQUEUE_REG_5__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__7_, n8506 );
not U_inv1253 ( n74365, P1_P1_INSTQUEUE_REG_5__7_ );
dff P1_P1_INSTQUEUE_REG_6__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__7_, n8466 );
not U_inv1254 ( n74374, P1_P1_INSTQUEUE_REG_6__7_ );
dff P1_P1_INSTQUEUE_REG_4__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__7_, n8546 );
not U_inv1255 ( n74363, P1_P1_INSTQUEUE_REG_4__7_ );
dff P1_P1_INSTQUEUE_REG_12__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__7_, n8226 );
not U_inv1256 ( n74362, P1_P1_INSTQUEUE_REG_12__7_ );
dff P1_P1_INSTQUEUE_REG_8__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__7_, n8386 );
not U_inv1257 ( n74368, P1_P1_INSTQUEUE_REG_8__7_ );
dff P1_P1_INSTQUEUE_REG_9__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__7_, n8346 );
not U_inv1258 ( n74373, P1_P1_INSTQUEUE_REG_9__7_ );
dff P1_P1_INSTQUEUE_REG_10__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__7_, n8306 );
not U_inv1259 ( n74377, P1_P1_INSTQUEUE_REG_10__7_ );
dff P1_P1_INSTQUEUE_REG_11__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__7_, n8266 );
not U_inv1260 ( n74375, P1_P1_INSTQUEUE_REG_11__7_ );
dff P1_P1_INSTQUEUE_REG_0__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__7_, n8706 );
not U_inv1261 ( n74357, P1_P1_INSTQUEUE_REG_0__7_ );
dff P1_P1_INSTQUEUE_REG_1__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__7_, n8666 );
not U_inv1262 ( n74364, P1_P1_INSTQUEUE_REG_1__7_ );
dff P1_P1_INSTQUEUE_REG_2__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__7_, n8626 );
not U_inv1263 ( n74367, P1_P1_INSTQUEUE_REG_2__7_ );
dff P1_P1_INSTQUEUE_REG_3__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__7_, n8586 );
not U_inv1264 ( n74359, P1_P1_INSTQUEUE_REG_3__7_ );
dff P1_P1_INSTQUEUE_REG_7__7__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__7_, n8426 );
not U_inv1265 ( n74369, P1_P1_INSTQUEUE_REG_7__7_ );
dff P1_P1_DATAO_REG_31__reg ( clk, reset, P1_P1_DATAO_REG_31_, n9426 );
dff P1_BUF1_REG_31__reg ( clk, reset, P1_BUF1_REG_31_, n276 );
not U_inv1266 ( n75446, P1_BUF1_REG_31_ );
dff P1_P1_DATAO_REG_1__reg ( clk, reset, P1_P1_DATAO_REG_1_, n9276 );
dff P1_BUF1_REG_1__reg ( clk, reset, P1_BUF1_REG_1_, n126 );
not U_inv1267 ( n75459, P1_BUF1_REG_1_ );
dff P1_P1_INSTQUEUE_REG_5__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__1_, n8536 );
not U_inv1268 ( n73982, P1_P1_INSTQUEUE_REG_5__1_ );
dff P1_P1_INSTQUEUE_REG_6__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__1_, n8496 );
not U_inv1269 ( n73989, P1_P1_INSTQUEUE_REG_6__1_ );
dff P1_P1_INSTQUEUE_REG_7__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__1_, n8456 );
not U_inv1270 ( n73984, P1_P1_INSTQUEUE_REG_7__1_ );
dff P1_P1_INSTQUEUE_REG_9__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__1_, n8376 );
not U_inv1271 ( n73988, P1_P1_INSTQUEUE_REG_9__1_ );
dff P1_P1_INSTQUEUE_REG_10__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__1_, n8336 );
not U_inv1272 ( n73995, P1_P1_INSTQUEUE_REG_10__1_ );
dff P1_P1_INSTQUEUE_REG_11__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__1_, n8296 );
not U_inv1273 ( n73991, P1_P1_INSTQUEUE_REG_11__1_ );
dff P1_P1_INSTQUEUE_REG_13__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__1_, n8216 );
not U_inv1274 ( n73985, P1_P1_INSTQUEUE_REG_13__1_ );
dff P1_P1_INSTQUEUE_REG_14__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__1_, n8176 );
not U_inv1275 ( n73992, P1_P1_INSTQUEUE_REG_14__1_ );
dff P1_P1_INSTQUEUE_REG_0__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__1_, n8736 );
not U_inv1276 ( n73964, P1_P1_INSTQUEUE_REG_0__1_ );
dff P1_P1_INSTQUEUE_REG_1__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__1_, n8696 );
not U_inv1277 ( n73979, P1_P1_INSTQUEUE_REG_1__1_ );
dff P1_P1_INSTQUEUE_REG_2__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__1_, n8656 );
not U_inv1278 ( n73986, P1_P1_INSTQUEUE_REG_2__1_ );
dff P1_P1_INSTQUEUE_REG_3__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__1_, n8616 );
not U_inv1279 ( n73981, P1_P1_INSTQUEUE_REG_3__1_ );
dff P1_P1_INSTQUEUE_REG_4__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__1_, n8576 );
not U_inv1280 ( n73978, P1_P1_INSTQUEUE_REG_4__1_ );
dff P1_P1_INSTQUEUE_REG_8__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__1_, n8416 );
not U_inv1281 ( n73983, P1_P1_INSTQUEUE_REG_8__1_ );
dff P1_P1_INSTQUEUE_REG_12__1__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__1_, n8256 );
not U_inv1282 ( n73980, P1_P1_INSTQUEUE_REG_12__1_ );
dff P1_P1_EAX_REG_1__reg ( clk, reset, ex_wire220, n9436 );
not U_inv1283 ( n74608, ex_wire220 );
dff P1_P1_EAX_REG_2__reg ( clk, reset, P1_P1_EAX_REG_2_, n9441 );
not U_inv1284 ( n73166, P1_P1_EAX_REG_2_ );
dff P1_P1_EAX_REG_3__reg ( clk, reset, ex_wire221, n9446 );
not U_inv1285 ( n74630, ex_wire221 );
dff P1_P1_LWORD_REG_3__reg ( clk, reset, P1_P1_LWORD_REG_3_, n9176 );
not U_inv1286 ( n75679, P1_P1_LWORD_REG_3_ );
dff P1_P1_DATAO_REG_3__reg ( clk, reset, P1_P1_DATAO_REG_3_, n9286 );
dff P1_BUF1_REG_3__reg ( clk, reset, P1_BUF1_REG_3_, n136 );
not U_inv1287 ( n75458, P1_BUF1_REG_3_ );
dff P1_P2_LWORD_REG_3__reg ( clk, reset, P1_P2_LWORD_REG_3_, n6931 );
not U_inv1288 ( n75645, P1_P2_LWORD_REG_3_ );
dff P1_P2_DATAO_REG_3__reg ( clk, reset, P1_P2_DATAO_REG_3_, n7041 );
not U_inv1289 ( n75544, P1_P2_DATAO_REG_3_ );
dff P1_BUF2_REG_3__reg ( clk, reset, P1_BUF2_REG_3_, n296 );
not U_inv1290 ( n75298, P1_BUF2_REG_3_ );
dff P1_P3_LWORD_REG_3__reg ( clk, reset, P1_P3_LWORD_REG_3_, n4686 );
not U_inv1291 ( n75692, P1_P3_LWORD_REG_3_ );
dff P1_P3_DATAO_REG_3__reg ( clk, reset, P1_P3_DATAO_REG_3_, n4796 );
dff P1_P2_INSTQUEUE_REG_15__3__reg ( clk, reset, ex_wire222, n5881 );
not U_inv1292 ( n73759, ex_wire222 );
dff P1_P2_EAX_REG_11__reg ( clk, reset, P1_P2_EAX_REG_11_, n7241 );
not U_inv1293 ( n74679, P1_P2_EAX_REG_11_ );
dff P1_P2_EAX_REG_12__reg ( clk, reset, P1_P2_EAX_REG_12_, n7246 );
not U_inv1294 ( n75274, P1_P2_EAX_REG_12_ );
dff P1_P2_EAX_REG_13__reg ( clk, reset, P1_P2_EAX_REG_13_, n7251 );
not U_inv1295 ( n74733, P1_P2_EAX_REG_13_ );
dff P1_P2_LWORD_REG_13__reg ( clk, reset, P1_P2_LWORD_REG_13_, n6881 );
not U_inv1296 ( n75644, P1_P2_LWORD_REG_13_ );
dff P1_P2_DATAO_REG_13__reg ( clk, reset, P1_P2_DATAO_REG_13_, n7091 );
not U_inv1297 ( n75540, P1_P2_DATAO_REG_13_ );
dff P1_BUF2_REG_13__reg ( clk, reset, P1_BUF2_REG_13_, n346 );
not U_inv1298 ( n75316, P1_BUF2_REG_13_ );
dff P1_P2_UWORD_REG_13__reg ( clk, reset, P1_P2_UWORD_REG_13_, n6956 );
not U_inv1299 ( n75570, P1_P2_UWORD_REG_13_ );
dff P1_P2_DATAO_REG_29__reg ( clk, reset, P1_P2_DATAO_REG_29_, n7171 );
not U_inv1300 ( n75596, P1_P2_DATAO_REG_29_ );
dff P1_BUF2_REG_29__reg ( clk, reset, P1_BUF2_REG_29_, n426 );
not U_inv1301 ( n75331, P1_BUF2_REG_29_ );
dff P1_P2_INSTQUEUE_REG_15__5__reg ( clk, reset, ex_wire223, n5871 );
not U_inv1302 ( n73908, ex_wire223 );
dff P1_P2_EAX_REG_27__reg ( clk, reset, P1_P2_EAX_REG_27_, n7321 );
not U_inv1303 ( n75323, P1_P2_EAX_REG_27_ );
dff P1_P2_EAX_REG_28__reg ( clk, reset, P1_P2_EAX_REG_28_, n7326 );
not U_inv1304 ( n73394, P1_P2_EAX_REG_28_ );
dff P1_P2_EAX_REG_29__reg ( clk, reset, P1_P2_EAX_REG_29_, n7331 );
not U_inv1305 ( n75205, P1_P2_EAX_REG_29_ );
dff P1_P2_EAX_REG_30__reg ( clk, reset, P1_P2_EAX_REG_30_, n7336 );
not U_inv1306 ( n75403, P1_P2_EAX_REG_30_ );
dff P1_P2_UWORD_REG_14__reg ( clk, reset, P1_P2_UWORD_REG_14_, n6951 );
not U_inv1307 ( n75569, P1_P2_UWORD_REG_14_ );
dff P1_P2_DATAO_REG_30__reg ( clk, reset, P1_P2_DATAO_REG_30_, n7176 );
not U_inv1308 ( n73432, P1_P2_DATAO_REG_30_ );
dff P1_BUF2_REG_30__reg ( clk, reset, P1_BUF2_REG_30_, n431 );
not U_inv1309 ( n75330, P1_BUF2_REG_30_ );
dff P1_P2_INSTQUEUE_REG_4__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__6_, n6306 );
not U_inv1310 ( n74070, P1_P2_INSTQUEUE_REG_4__6_ );
dff P1_P2_EAX_REG_22__reg ( clk, reset, P1_P2_EAX_REG_22_, n7296 );
not U_inv1311 ( n75387, P1_P2_EAX_REG_22_ );
dff P1_P2_UWORD_REG_6__reg ( clk, reset, P1_P2_UWORD_REG_6_, n6991 );
not U_inv1312 ( n75485, P1_P2_UWORD_REG_6_ );
dff P1_P2_DATAO_REG_22__reg ( clk, reset, P1_P2_DATAO_REG_22_, n7136 );
not U_inv1313 ( n75543, P1_P2_DATAO_REG_22_ );
dff P1_BUF1_REG_22__reg ( clk, reset, P1_BUF1_REG_22_, n231 );
not U_inv1314 ( n75400, P1_BUF1_REG_22_ );
dff P1_P1_INSTQUEUE_REG_0__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__6_, n8711 );
not U_inv1315 ( n74319, P1_P1_INSTQUEUE_REG_0__6_ );
dff P1_P1_INSTQUEUE_REG_1__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__6_, n8671 );
not U_inv1316 ( n74321, P1_P1_INSTQUEUE_REG_1__6_ );
dff P1_P1_INSTQUEUE_REG_2__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__6_, n8631 );
not U_inv1317 ( n74328, P1_P1_INSTQUEUE_REG_2__6_ );
dff P1_P1_INSTQUEUE_REG_3__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__6_, n8591 );
not U_inv1318 ( n74323, P1_P1_INSTQUEUE_REG_3__6_ );
dff P1_P1_INSTQUEUE_REG_4__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__6_, n8551 );
not U_inv1319 ( n74320, P1_P1_INSTQUEUE_REG_4__6_ );
dff P1_P1_INSTQUEUE_REG_5__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__6_, n8511 );
not U_inv1320 ( n74324, P1_P1_INSTQUEUE_REG_5__6_ );
dff P1_P1_INSTQUEUE_REG_6__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__6_, n8471 );
not U_inv1321 ( n74330, P1_P1_INSTQUEUE_REG_6__6_ );
dff P1_P1_INSTQUEUE_REG_7__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__6_, n8431 );
not U_inv1322 ( n74326, P1_P1_INSTQUEUE_REG_7__6_ );
dff P1_P1_INSTQUEUE_REG_8__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__6_, n8391 );
not U_inv1323 ( n74325, P1_P1_INSTQUEUE_REG_8__6_ );
dff P1_P1_INSTQUEUE_REG_9__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__6_, n8351 );
not U_inv1324 ( n74329, P1_P1_INSTQUEUE_REG_9__6_ );
dff P1_P1_INSTQUEUE_REG_10__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__6_, n8311 );
not U_inv1325 ( n74334, P1_P1_INSTQUEUE_REG_10__6_ );
dff P1_P1_INSTQUEUE_REG_11__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__6_, n8271 );
not U_inv1326 ( n74331, P1_P1_INSTQUEUE_REG_11__6_ );
dff P1_P1_INSTQUEUE_REG_13__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__6_, n8191 );
not U_inv1327 ( n74327, P1_P1_INSTQUEUE_REG_13__6_ );
dff P1_P1_INSTQUEUE_REG_14__6__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__6_, n8151 );
not U_inv1328 ( n74332, P1_P1_INSTQUEUE_REG_14__6_ );
dff P1_P1_EAX_REG_22__reg ( clk, reset, P1_P1_EAX_REG_22_, n9541 );
not U_inv1329 ( n75002, P1_P1_EAX_REG_22_ );
dff P1_P1_EAX_REG_23__reg ( clk, reset, ex_wire224, n9546 );
not U_inv1330 ( n75013, ex_wire224 );
dff P1_P1_EAX_REG_24__reg ( clk, reset, P1_P1_EAX_REG_24_, n9551 );
not U_inv1331 ( n73307, P1_P1_EAX_REG_24_ );
dff P1_P1_UWORD_REG_8__reg ( clk, reset, P1_P1_UWORD_REG_8_, n9226 );
not U_inv1332 ( n75586, P1_P1_UWORD_REG_8_ );
dff P1_P1_DATAO_REG_24__reg ( clk, reset, P1_P1_DATAO_REG_24_, n9391 );
dff P1_BUF1_REG_24__reg ( clk, reset, P1_BUF1_REG_24_, n241 );
not U_inv1333 ( n75416, P1_BUF1_REG_24_ );
dff P1_P1_INSTQUEUE_REG_15__0__reg ( clk, reset, ex_wire225, n8141 );
not U_inv1334 ( n74019, ex_wire225 );
dff P1_P1_MEMORYFETCH_REG_reg ( clk, reset, P1_P1_MEMORYFETCH_REG, n9981 );
dff P1_P1_M_IO_N_REG_reg ( clk, reset, P1_P1_M_IO_N_REG, n9961 );
not U_inv1335 ( n75988, P1_P1_M_IO_N_REG );
dff P1_P1_UWORD_REG_0__reg ( clk, reset, P1_P1_UWORD_REG_0_, n9266 );
not U_inv1336 ( n75502, P1_P1_UWORD_REG_0_ );
dff P1_P1_DATAO_REG_16__reg ( clk, reset, P1_P1_DATAO_REG_16_, n9351 );
dff P1_BUF1_REG_16__reg ( clk, reset, P1_BUF1_REG_16_, n201 );
not U_inv1337 ( n75399, P1_BUF1_REG_16_ );
dff P1_P1_INSTQUEUE_REG_0__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__0_, n8741 );
not U_inv1338 ( n74005, P1_P1_INSTQUEUE_REG_0__0_ );
dff P1_P1_INSTQUEUE_REG_1__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__0_, n8701 );
not U_inv1339 ( n74026, P1_P1_INSTQUEUE_REG_1__0_ );
dff P1_P1_INSTQUEUE_REG_2__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__0_, n8661 );
not U_inv1340 ( n74038, P1_P1_INSTQUEUE_REG_2__0_ );
dff P1_P1_INSTQUEUE_REG_3__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__0_, n8621 );
not U_inv1341 ( n74017, P1_P1_INSTQUEUE_REG_3__0_ );
dff P1_P1_INSTQUEUE_REG_4__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__0_, n8581 );
not U_inv1342 ( n74031, P1_P1_INSTQUEUE_REG_4__0_ );
dff P1_P1_INSTQUEUE_REG_5__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__0_, n8541 );
not U_inv1343 ( n74052, P1_P1_INSTQUEUE_REG_5__0_ );
dff P1_P1_INSTQUEUE_REG_6__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__0_, n8501 );
not U_inv1344 ( n74060, P1_P1_INSTQUEUE_REG_6__0_ );
dff P1_P1_INSTQUEUE_REG_7__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__0_, n8461 );
not U_inv1345 ( n74039, P1_P1_INSTQUEUE_REG_7__0_ );
dff P1_P1_INSTQUEUE_REG_8__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__0_, n8421 );
not U_inv1346 ( n74037, P1_P1_INSTQUEUE_REG_8__0_ );
dff P1_P1_INSTQUEUE_REG_9__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__0_, n8381 );
not U_inv1347 ( n74059, P1_P1_INSTQUEUE_REG_9__0_ );
dff P1_P1_INSTQUEUE_REG_10__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__0_, n8341 );
not U_inv1348 ( n74061, P1_P1_INSTQUEUE_REG_10__0_ );
dff P1_P1_INSTQUEUE_REG_11__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__0_, n8301 );
not U_inv1349 ( n74045, P1_P1_INSTQUEUE_REG_11__0_ );
dff P1_P1_INSTQUEUE_REG_12__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__0_, n8261 );
not U_inv1350 ( n74016, P1_P1_INSTQUEUE_REG_12__0_ );
dff P1_P1_INSTQUEUE_REG_13__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__0_, n8221 );
not U_inv1351 ( n74035, P1_P1_INSTQUEUE_REG_13__0_ );
dff P1_P1_INSTQUEUE_REG_14__0__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__0_, n8181 );
not U_inv1352 ( n74043, P1_P1_INSTQUEUE_REG_14__0_ );
dff P1_P1_UWORD_REG_6__reg ( clk, reset, P1_P1_UWORD_REG_6_, n9236 );
not U_inv1353 ( n75501, P1_P1_UWORD_REG_6_ );
dff P1_P1_DATAO_REG_22__reg ( clk, reset, P1_P1_DATAO_REG_22_, n9381 );
dff P1_P1_LWORD_REG_2__reg ( clk, reset, P1_P1_LWORD_REG_2_, n9181 );
not U_inv1354 ( n75678, P1_P1_LWORD_REG_2_ );
dff P1_P1_DATAO_REG_2__reg ( clk, reset, P1_P1_DATAO_REG_2_, n9281 );
dff P1_BUF1_REG_2__reg ( clk, reset, P1_BUF1_REG_2_, n131 );
not U_inv1355 ( n75457, P1_BUF1_REG_2_ );
dff P1_P2_LWORD_REG_2__reg ( clk, reset, P1_P2_LWORD_REG_2_, n6936 );
not U_inv1356 ( n75643, P1_P2_LWORD_REG_2_ );
dff P1_P2_DATAO_REG_2__reg ( clk, reset, P1_P2_DATAO_REG_2_, n7036 );
not U_inv1357 ( n75541, P1_P2_DATAO_REG_2_ );
dff P1_BUF2_REG_2__reg ( clk, reset, P1_BUF2_REG_2_, n291 );
not U_inv1358 ( n75296, P1_BUF2_REG_2_ );
dff P1_P3_UWORD_REG_2__reg ( clk, reset, P1_P3_UWORD_REG_2_, n4766 );
not U_inv1359 ( n75603, P1_P3_UWORD_REG_2_ );
dff P1_P3_DATAO_REG_18__reg ( clk, reset, P1_P3_DATAO_REG_18_, n4871 );
dff P1_P3_LWORD_REG_2__reg ( clk, reset, P1_P3_LWORD_REG_2_, n4691 );
not U_inv1360 ( n75691, P1_P3_LWORD_REG_2_ );
dff P1_P3_DATAO_REG_2__reg ( clk, reset, P1_P3_DATAO_REG_2_, n4791 );
dff P3_IR_REG_2__reg ( clk, reset, P3_IR_REG_2_, n811 );
dff P3_IR_REG_3__reg ( clk, reset, P3_IR_REG_3_, n816 );
not U_inv1361 ( n73797, P3_IR_REG_3_ );
dff P3_IR_REG_4__reg ( clk, reset, P3_IR_REG_4_, n821 );
dff P3_REG3_REG_2__reg ( clk, reset, P3_REG3_REG_2_, n1886 );
not U_inv1362 ( n73833, P3_REG3_REG_2_ );
dff P3_REG3_REG_3__reg ( clk, reset, P3_REG3_REG_3_, n1981 );
not U_inv1363 ( n75248, P3_REG3_REG_3_ );
dff P3_REG3_REG_4__reg ( clk, reset, P3_REG3_REG_4_, n1921 );
not U_inv1364 ( n74064, P3_REG3_REG_4_ );
dff P3_REG2_REG_4__reg ( clk, reset, P3_REG2_REG_4_, n1461 );
not U_inv1365 ( n74217, P3_REG2_REG_4_ );
dff P3_REG2_REG_3__reg ( clk, reset, P3_REG2_REG_3_, n1456 );
not U_inv1366 ( n73910, P3_REG2_REG_3_ );
dff P3_REG2_REG_2__reg ( clk, reset, P3_REG2_REG_2_, n1451 );
not U_inv1367 ( n73826, P3_REG2_REG_2_ );
dff P1_P1_LWORD_REG_13__reg ( clk, reset, P1_P1_LWORD_REG_13_, n9126 );
not U_inv1368 ( n75677, P1_P1_LWORD_REG_13_ );
dff P1_P1_DATAO_REG_13__reg ( clk, reset, P1_P1_DATAO_REG_13_, n9336 );
dff P1_BUF1_REG_13__reg ( clk, reset, P1_BUF1_REG_13_, n186 );
not U_inv1369 ( n75443, P1_BUF1_REG_13_ );
dff P1_P1_UWORD_REG_13__reg ( clk, reset, P1_P1_UWORD_REG_13_, n9201 );
not U_inv1370 ( n75585, P1_P1_UWORD_REG_13_ );
dff P1_P1_DATAO_REG_29__reg ( clk, reset, P1_P1_DATAO_REG_29_, n9416 );
dff P1_BUF1_REG_29__reg ( clk, reset, P1_BUF1_REG_29_, n266 );
not U_inv1371 ( n75392, P1_BUF1_REG_29_ );
dff P1_P1_INSTQUEUE_REG_15__5__reg ( clk, reset, ex_wire226, n8116 );
not U_inv1372 ( n74297, ex_wire226 );
dff P1_P1_EAX_REG_5__reg ( clk, reset, P1_P1_EAX_REG_5_, n9456 );
not U_inv1373 ( n73196, P1_P1_EAX_REG_5_ );
dff P1_P1_LWORD_REG_5__reg ( clk, reset, P1_P1_LWORD_REG_5_, n9166 );
not U_inv1374 ( n75676, P1_P1_LWORD_REG_5_ );
dff P1_P1_DATAO_REG_5__reg ( clk, reset, P1_P1_DATAO_REG_5_, n9296 );
dff P1_BUF1_REG_5__reg ( clk, reset, P1_BUF1_REG_5_, n146 );
not U_inv1375 ( n75456, P1_BUF1_REG_5_ );
dff P1_P2_LWORD_REG_5__reg ( clk, reset, P1_P2_LWORD_REG_5_, n6921 );
not U_inv1376 ( n75642, P1_P2_LWORD_REG_5_ );
dff P1_P2_DATAO_REG_5__reg ( clk, reset, P1_P2_DATAO_REG_5_, n7051 );
not U_inv1377 ( n75539, P1_P2_DATAO_REG_5_ );
dff P1_BUF2_REG_5__reg ( clk, reset, P1_BUF2_REG_5_, n306 );
not U_inv1378 ( n75312, P1_BUF2_REG_5_ );
dff P1_P3_LWORD_REG_5__reg ( clk, reset, P1_P3_LWORD_REG_5_, n4676 );
not U_inv1379 ( n75690, P1_P3_LWORD_REG_5_ );
dff P1_P3_DATAO_REG_5__reg ( clk, reset, P1_P3_DATAO_REG_5_, n4806 );
dff P3_IR_REG_5__reg ( clk, reset, P3_IR_REG_5_, n826 );
not U_inv1380 ( n74105, P3_IR_REG_5_ );
dff P3_IR_REG_6__reg ( clk, reset, P3_IR_REG_6_, n831 );
dff P3_IR_REG_7__reg ( clk, reset, P3_IR_REG_7_, n836 );
not U_inv1381 ( n74225, P3_IR_REG_7_ );
dff P3_REG3_REG_5__reg ( clk, reset, P3_REG3_REG_5_, n1936 );
not U_inv1382 ( n74170, P3_REG3_REG_5_ );
dff P3_REG3_REG_6__reg ( clk, reset, P3_REG3_REG_6_, n1876 );
not U_inv1383 ( n74256, P3_REG3_REG_6_ );
dff P3_REG3_REG_7__reg ( clk, reset, P3_REG3_REG_7_, n2006 );
not U_inv1384 ( n72929, P3_REG3_REG_7_ );
dff P3_REG2_REG_5__reg ( clk, reset, P3_REG2_REG_5_, n1466 );
not U_inv1385 ( n74259, P3_REG2_REG_5_ );
dff P1_P2_INSTQUEUE_REG_14__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__5_, n5911 );
not U_inv1386 ( n73931, P1_P2_INSTQUEUE_REG_14__5_ );
dff P1_P2_EAX_REG_21__reg ( clk, reset, P1_P2_EAX_REG_21_, n7291 );
not U_inv1387 ( n74923, P1_P2_EAX_REG_21_ );
dff P1_P2_UWORD_REG_5__reg ( clk, reset, P1_P2_UWORD_REG_5_, n6996 );
not U_inv1388 ( n75484, P1_P2_UWORD_REG_5_ );
dff P1_P2_DATAO_REG_21__reg ( clk, reset, P1_P2_DATAO_REG_21_, n7131 );
not U_inv1389 ( n75538, P1_P2_DATAO_REG_21_ );
dff P1_BUF1_REG_21__reg ( clk, reset, P1_BUF1_REG_21_, n226 );
not U_inv1390 ( n75398, P1_BUF1_REG_21_ );
dff P1_P1_INSTQUEUE_REG_0__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__5_, n8716 );
not U_inv1391 ( n74280, P1_P1_INSTQUEUE_REG_0__5_ );
dff P1_P1_INSTQUEUE_REG_1__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__5_, n8676 );
not U_inv1392 ( n74284, P1_P1_INSTQUEUE_REG_1__5_ );
dff P1_P1_INSTQUEUE_REG_2__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__5_, n8636 );
not U_inv1393 ( n74291, P1_P1_INSTQUEUE_REG_2__5_ );
dff P1_P1_INSTQUEUE_REG_3__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__5_, n8596 );
not U_inv1394 ( n74286, P1_P1_INSTQUEUE_REG_3__5_ );
dff P1_P1_INSTQUEUE_REG_4__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__5_, n8556 );
not U_inv1395 ( n74283, P1_P1_INSTQUEUE_REG_4__5_ );
dff P1_P1_INSTQUEUE_REG_5__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__5_, n8516 );
not U_inv1396 ( n74287, P1_P1_INSTQUEUE_REG_5__5_ );
dff P1_P1_INSTQUEUE_REG_6__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__5_, n8476 );
not U_inv1397 ( n74293, P1_P1_INSTQUEUE_REG_6__5_ );
dff P1_P1_INSTQUEUE_REG_7__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__5_, n8436 );
not U_inv1398 ( n74289, P1_P1_INSTQUEUE_REG_7__5_ );
dff P1_P1_INSTQUEUE_REG_8__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__5_, n8396 );
not U_inv1399 ( n74288, P1_P1_INSTQUEUE_REG_8__5_ );
dff P1_P1_INSTQUEUE_REG_9__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__5_, n8356 );
not U_inv1400 ( n74292, P1_P1_INSTQUEUE_REG_9__5_ );
dff P1_P1_INSTQUEUE_REG_10__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__5_, n8316 );
not U_inv1401 ( n74296, P1_P1_INSTQUEUE_REG_10__5_ );
dff P1_P1_INSTQUEUE_REG_11__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__5_, n8276 );
not U_inv1402 ( n74294, P1_P1_INSTQUEUE_REG_11__5_ );
dff P1_P1_INSTQUEUE_REG_12__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__5_, n8236 );
not U_inv1403 ( n74285, P1_P1_INSTQUEUE_REG_12__5_ );
dff P1_P1_INSTQUEUE_REG_13__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__5_, n8196 );
not U_inv1404 ( n74290, P1_P1_INSTQUEUE_REG_13__5_ );
dff P1_P1_INSTQUEUE_REG_14__5__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__5_, n8156 );
not U_inv1405 ( n74295, P1_P1_INSTQUEUE_REG_14__5_ );
dff P1_P1_EAX_REG_21__reg ( clk, reset, P1_P1_EAX_REG_21_, n9536 );
not U_inv1406 ( n73289, P1_P1_EAX_REG_21_ );
dff P1_P1_EAX_REG_25__reg ( clk, reset, P1_P1_EAX_REG_25_, n9556 );
not U_inv1407 ( n75062, P1_P1_EAX_REG_25_ );
dff P1_P1_EAX_REG_26__reg ( clk, reset, ex_wire227, n9561 );
not U_inv1408 ( n75085, ex_wire227 );
dff P1_P1_UWORD_REG_10__reg ( clk, reset, P1_P1_UWORD_REG_10_, n9216 );
not U_inv1409 ( n75584, P1_P1_UWORD_REG_10_ );
dff P1_P1_DATAO_REG_26__reg ( clk, reset, P1_P1_DATAO_REG_26_, n9401 );
dff P1_BUF1_REG_26__reg ( clk, reset, P1_BUF1_REG_26_, n251 );
not U_inv1410 ( n75391, P1_BUF1_REG_26_ );
dff P1_P2_INSTQUEUE_REG_15__2__reg ( clk, reset, ex_wire228, n5886 );
not U_inv1411 ( n73748, ex_wire228 );
dff P1_P2_EAX_REG_18__reg ( clk, reset, P1_P2_EAX_REG_18_, n7276 );
not U_inv1412 ( n75386, P1_P2_EAX_REG_18_ );
dff P1_P2_UWORD_REG_2__reg ( clk, reset, P1_P2_UWORD_REG_2_, n7011 );
not U_inv1413 ( n75483, P1_P2_UWORD_REG_2_ );
dff P1_P2_DATAO_REG_18__reg ( clk, reset, P1_P2_DATAO_REG_18_, n7116 );
not U_inv1414 ( n75536, P1_P2_DATAO_REG_18_ );
dff P1_BUF2_REG_18__reg ( clk, reset, P1_BUF2_REG_18_, n371 );
not U_inv1415 ( n75353, P1_BUF2_REG_18_ );
dff P1_P3_INSTQUEUE_REG_5__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__2_, n4041 );
not U_inv1416 ( n74025, P1_P3_INSTQUEUE_REG_5__2_ );
dff P1_P3_INSTQUEUE_REG_6__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__2_, n4001 );
not U_inv1417 ( n74040, P1_P3_INSTQUEUE_REG_6__2_ );
dff P1_P3_INSTQUEUE_REG_8__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__2_, n3921 );
not U_inv1418 ( n74030, P1_P3_INSTQUEUE_REG_8__2_ );
dff P1_P3_INSTQUEUE_REG_9__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__2_, n3881 );
not U_inv1419 ( n74036, P1_P3_INSTQUEUE_REG_9__2_ );
dff P1_P3_INSTQUEUE_REG_10__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__2_, n3841 );
not U_inv1420 ( n74047, P1_P3_INSTQUEUE_REG_10__2_ );
dff P1_P3_INSTQUEUE_REG_11__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__2_, n3801 );
not U_inv1421 ( n74042, P1_P3_INSTQUEUE_REG_11__2_ );
dff P1_P3_INSTQUEUE_REG_12__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__2_, n3761 );
not U_inv1422 ( n74023, P1_P3_INSTQUEUE_REG_12__2_ );
dff P1_P3_INSTQUEUE_REG_13__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__2_, n3721 );
not U_inv1423 ( n74033, P1_P3_INSTQUEUE_REG_13__2_ );
dff P1_P3_INSTQUEUE_REG_0__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__2_, n4241 );
not U_inv1424 ( n74012, P1_P3_INSTQUEUE_REG_0__2_ );
dff P1_P3_INSTQUEUE_REG_1__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__2_, n4201 );
not U_inv1425 ( n74022, P1_P3_INSTQUEUE_REG_1__2_ );
dff P1_P3_INSTQUEUE_REG_2__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__2_, n4161 );
not U_inv1426 ( n74034, P1_P3_INSTQUEUE_REG_2__2_ );
dff P1_P3_INSTQUEUE_REG_3__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__2_, n4121 );
not U_inv1427 ( n74024, P1_P3_INSTQUEUE_REG_3__2_ );
dff P1_P3_INSTQUEUE_REG_4__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__2_, n4081 );
not U_inv1428 ( n74021, P1_P3_INSTQUEUE_REG_4__2_ );
dff P1_P3_INSTQUEUE_REG_7__2__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__2_, n3961 );
not U_inv1429 ( n74032, P1_P3_INSTQUEUE_REG_7__2_ );
dff P1_P3_INSTQUEUE_REG_15__2__reg ( clk, reset, ex_wire229, n3641 );
not U_inv1430 ( n74048, ex_wire229 );
dff P1_P2_EAX_REG_19__reg ( clk, reset, P1_P2_EAX_REG_19_, n7281 );
not U_inv1431 ( n74878, P1_P2_EAX_REG_19_ );
dff P1_P2_UWORD_REG_3__reg ( clk, reset, P1_P2_UWORD_REG_3_, n7006 );
not U_inv1432 ( n75482, P1_P2_UWORD_REG_3_ );
dff P1_P2_DATAO_REG_19__reg ( clk, reset, P1_P2_DATAO_REG_19_, n7121 );
not U_inv1433 ( n75537, P1_P2_DATAO_REG_19_ );
dff P1_BUF1_REG_19__reg ( clk, reset, P1_BUF1_REG_19_, n216 );
not U_inv1434 ( n75397, P1_BUF1_REG_19_ );
dff P1_P1_INSTQUEUE_REG_15__3__reg ( clk, reset, ex_wire230, n8126 );
not U_inv1435 ( n74143, ex_wire230 );
dff P1_P1_EAX_REG_18__reg ( clk, reset, P1_P1_EAX_REG_18_, n9521 );
not U_inv1436 ( n73266, P1_P1_EAX_REG_18_ );
dff P1_P1_UWORD_REG_2__reg ( clk, reset, P1_P1_UWORD_REG_2_, n9256 );
not U_inv1437 ( n75500, P1_P1_UWORD_REG_2_ );
dff P1_P1_DATAO_REG_18__reg ( clk, reset, P1_P1_DATAO_REG_18_, n9361 );
dff P1_BUF1_REG_18__reg ( clk, reset, P1_BUF1_REG_18_, n211 );
not U_inv1438 ( n75396, P1_BUF1_REG_18_ );
dff P1_P1_INSTQUEUE_REG_0__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__2_, n8731 );
not U_inv1439 ( n74046, P1_P1_INSTQUEUE_REG_0__2_ );
dff P1_P1_INSTQUEUE_REG_1__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__2_, n8691 );
not U_inv1440 ( n74072, P1_P1_INSTQUEUE_REG_1__2_ );
dff P1_P1_INSTQUEUE_REG_2__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__2_, n8651 );
not U_inv1441 ( n74097, P1_P1_INSTQUEUE_REG_2__2_ );
dff P1_P1_INSTQUEUE_REG_3__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__2_, n8611 );
not U_inv1442 ( n74084, P1_P1_INSTQUEUE_REG_3__2_ );
dff P1_P1_INSTQUEUE_REG_4__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__2_, n8571 );
not U_inv1443 ( n74071, P1_P1_INSTQUEUE_REG_4__2_ );
dff P1_P1_INSTQUEUE_REG_5__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__2_, n8531 );
not U_inv1444 ( n74085, P1_P1_INSTQUEUE_REG_5__2_ );
dff P1_P1_INSTQUEUE_REG_6__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__2_, n8491 );
not U_inv1445 ( n74099, P1_P1_INSTQUEUE_REG_6__2_ );
dff P1_P1_INSTQUEUE_REG_7__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__2_, n8451 );
not U_inv1446 ( n74089, P1_P1_INSTQUEUE_REG_7__2_ );
dff P1_P1_INSTQUEUE_REG_8__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__2_, n8411 );
not U_inv1447 ( n74088, P1_P1_INSTQUEUE_REG_8__2_ );
dff P1_P1_INSTQUEUE_REG_9__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__2_, n8371 );
not U_inv1448 ( n74098, P1_P1_INSTQUEUE_REG_9__2_ );
dff P1_P1_INSTQUEUE_REG_10__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__2_, n8331 );
not U_inv1449 ( n74103, P1_P1_INSTQUEUE_REG_10__2_ );
dff P1_P1_INSTQUEUE_REG_11__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__2_, n8291 );
not U_inv1450 ( n74100, P1_P1_INSTQUEUE_REG_11__2_ );
dff P1_P1_INSTQUEUE_REG_12__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__2_, n8251 );
not U_inv1451 ( n74082, P1_P1_INSTQUEUE_REG_12__2_ );
dff P1_P1_INSTQUEUE_REG_13__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__2_, n8211 );
not U_inv1452 ( n74093, P1_P1_INSTQUEUE_REG_13__2_ );
dff P1_P1_INSTQUEUE_REG_14__2__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__2_, n8171 );
not U_inv1453 ( n74101, P1_P1_INSTQUEUE_REG_14__2_ );
dff P1_P1_INSTQUEUE_REG_15__2__reg ( clk, reset, ex_wire231, n8131 );
not U_inv1454 ( n74111, ex_wire231 );
dff P1_P2_INSTQUEUE_REG_0__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__2_, n6486 );
not U_inv1455 ( n73671, P1_P2_INSTQUEUE_REG_0__2_ );
dff P1_P2_INSTQUEUE_REG_1__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__2_, n6446 );
not U_inv1456 ( n73709, P1_P2_INSTQUEUE_REG_1__2_ );
dff P1_P2_INSTQUEUE_REG_2__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__2_, n6406 );
not U_inv1457 ( n73730, P1_P2_INSTQUEUE_REG_2__2_ );
dff P1_P2_INSTQUEUE_REG_3__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__2_, n6366 );
not U_inv1458 ( n73716, P1_P2_INSTQUEUE_REG_3__2_ );
dff P1_P2_INSTQUEUE_REG_4__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__2_, n6326 );
not U_inv1459 ( n73706, P1_P2_INSTQUEUE_REG_4__2_ );
dff P1_P2_INSTQUEUE_REG_7__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__2_, n6206 );
not U_inv1460 ( n73724, P1_P2_INSTQUEUE_REG_7__2_ );
dff P1_P2_INSTQUEUE_REG_5__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__2_, n6286 );
not U_inv1461 ( n73718, P1_P2_INSTQUEUE_REG_5__2_ );
dff P1_P2_INSTQUEUE_REG_6__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__2_, n6246 );
not U_inv1462 ( n73736, P1_P2_INSTQUEUE_REG_6__2_ );
dff P1_P2_INSTQUEUE_REG_8__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__2_, n6166 );
not U_inv1463 ( n73721, P1_P2_INSTQUEUE_REG_8__2_ );
dff P1_P2_INSTQUEUE_REG_9__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__2_, n6126 );
not U_inv1464 ( n73733, P1_P2_INSTQUEUE_REG_9__2_ );
dff P1_P2_INSTQUEUE_REG_10__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__2_, n6086 );
not U_inv1465 ( n73745, P1_P2_INSTQUEUE_REG_10__2_ );
dff P1_P2_INSTQUEUE_REG_11__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__2_, n6046 );
not U_inv1466 ( n73739, P1_P2_INSTQUEUE_REG_11__2_ );
dff P1_P2_INSTQUEUE_REG_12__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__2_, n6006 );
not U_inv1467 ( n73713, P1_P2_INSTQUEUE_REG_12__2_ );
dff P1_P2_INSTQUEUE_REG_13__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__2_, n5966 );
not U_inv1468 ( n73727, P1_P2_INSTQUEUE_REG_13__2_ );
dff P1_P2_INSTQUEUE_REG_14__2__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__2_, n5926 );
not U_inv1469 ( n73742, P1_P2_INSTQUEUE_REG_14__2_ );
dff P1_P1_EAX_REG_7__reg ( clk, reset, P1_P1_EAX_REG_7_, n9466 );
not U_inv1470 ( n74739, P1_P1_EAX_REG_7_ );
dff P1_P1_EAX_REG_8__reg ( clk, reset, P1_P1_EAX_REG_8_, n9471 );
not U_inv1471 ( n73219, P1_P1_EAX_REG_8_ );
dff P1_P1_LWORD_REG_8__reg ( clk, reset, P1_P1_LWORD_REG_8_, n9151 );
not U_inv1472 ( n75675, P1_P1_LWORD_REG_8_ );
dff P1_P1_DATAO_REG_8__reg ( clk, reset, P1_P1_DATAO_REG_8_, n9311 );
dff P1_BUF1_REG_8__reg ( clk, reset, P1_BUF1_REG_8_, n161 );
not U_inv1473 ( n75442, P1_BUF1_REG_8_ );
dff P1_P2_UWORD_REG_8__reg ( clk, reset, P1_P2_UWORD_REG_8_, n6981 );
not U_inv1474 ( n75568, P1_P2_UWORD_REG_8_ );
dff P1_P2_DATAO_REG_24__reg ( clk, reset, P1_P2_DATAO_REG_24_, n7146 );
not U_inv1475 ( n75597, P1_P2_DATAO_REG_24_ );
dff P1_BUF2_REG_24__reg ( clk, reset, P1_BUF2_REG_24_, n401 );
not U_inv1476 ( n75335, P1_BUF2_REG_24_ );
dff P1_P3_INSTQUEUE_REG_0__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__0_, n4251 );
not U_inv1477 ( n73987, P1_P3_INSTQUEUE_REG_0__0_ );
dff P1_P3_EBX_REG_0__reg ( clk, reset, P1_P3_EBX_REG_0_, n5101 );
not U_inv1478 ( n73119, P1_P3_EBX_REG_0_ );
dff P1_P3_INSTQUEUE_REG_1__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__0_, n4211 );
not U_inv1479 ( n74003, P1_P3_INSTQUEUE_REG_1__0_ );
dff P1_P3_INSTQUEUE_REG_2__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__0_, n4171 );
not U_inv1480 ( n74008, P1_P3_INSTQUEUE_REG_2__0_ );
dff P1_P3_INSTQUEUE_REG_3__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__0_, n4131 );
not U_inv1481 ( n74001, P1_P3_INSTQUEUE_REG_3__0_ );
dff P1_P3_INSTQUEUE_REG_4__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__0_, n4091 );
not U_inv1482 ( n74004, P1_P3_INSTQUEUE_REG_4__0_ );
dff P1_P3_INSTQUEUE_REG_5__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__0_, n4051 );
not U_inv1483 ( n74013, P1_P3_INSTQUEUE_REG_5__0_ );
dff P1_P3_INSTQUEUE_REG_6__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__0_, n4011 );
not U_inv1484 ( n74015, P1_P3_INSTQUEUE_REG_6__0_ );
dff P1_P3_INSTQUEUE_REG_7__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__0_, n3971 );
not U_inv1485 ( n74009, P1_P3_INSTQUEUE_REG_7__0_ );
dff P1_P3_INSTQUEUE_REG_8__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__0_, n3931 );
not U_inv1486 ( n74007, P1_P3_INSTQUEUE_REG_8__0_ );
dff P1_P3_INSTQUEUE_REG_9__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__0_, n3891 );
not U_inv1487 ( n74014, P1_P3_INSTQUEUE_REG_9__0_ );
dff P1_P3_INSTQUEUE_REG_10__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__0_, n3851 );
not U_inv1488 ( n74018, P1_P3_INSTQUEUE_REG_10__0_ );
dff P1_P3_INSTQUEUE_REG_11__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__0_, n3811 );
not U_inv1489 ( n74011, P1_P3_INSTQUEUE_REG_11__0_ );
dff P1_P3_INSTQUEUE_REG_12__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__0_, n3771 );
not U_inv1490 ( n74000, P1_P3_INSTQUEUE_REG_12__0_ );
dff P1_P3_INSTQUEUE_REG_13__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__0_, n3731 );
not U_inv1491 ( n74006, P1_P3_INSTQUEUE_REG_13__0_ );
dff P1_P3_INSTQUEUE_REG_14__0__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__0_, n3691 );
not U_inv1492 ( n74010, P1_P3_INSTQUEUE_REG_14__0_ );
dff P1_P2_LWORD_REG_8__reg ( clk, reset, P1_P2_LWORD_REG_8_, n6906 );
not U_inv1493 ( n75641, P1_P2_LWORD_REG_8_ );
dff P1_P2_DATAO_REG_8__reg ( clk, reset, P1_P2_DATAO_REG_8_, n7066 );
not U_inv1494 ( n75535, P1_P2_DATAO_REG_8_ );
dff P1_BUF2_REG_8__reg ( clk, reset, P1_BUF2_REG_8_, n321 );
not U_inv1495 ( n75320, P1_BUF2_REG_8_ );
dff P1_P3_LWORD_REG_8__reg ( clk, reset, P1_P3_LWORD_REG_8_, n4661 );
not U_inv1496 ( n75689, P1_P3_LWORD_REG_8_ );
dff P1_P3_DATAO_REG_8__reg ( clk, reset, P1_P3_DATAO_REG_8_, n4821 );
dff P3_IR_REG_8__reg ( clk, reset, P3_IR_REG_8_, n841 );
dff P3_REG3_REG_8__reg ( clk, reset, P3_REG3_REG_8_, n1966 );
not U_inv1497 ( n72936, P3_REG3_REG_8_ );
dff P3_REG2_REG_8__reg ( clk, reset, P3_REG2_REG_8_, n1481 );
not U_inv1498 ( n74382, P3_REG2_REG_8_ );
dff P1_P1_EAX_REG_9__reg ( clk, reset, ex_wire232, n9476 );
not U_inv1499 ( n74756, ex_wire232 );
dff P1_P1_EAX_REG_10__reg ( clk, reset, P1_P1_EAX_REG_10_, n9481 );
not U_inv1500 ( n74787, P1_P1_EAX_REG_10_ );
dff P1_P1_EAX_REG_11__reg ( clk, reset, P1_P1_EAX_REG_11_, n9486 );
not U_inv1501 ( n73238, P1_P1_EAX_REG_11_ );
dff P1_P1_LWORD_REG_11__reg ( clk, reset, P1_P1_LWORD_REG_11_, n9136 );
not U_inv1502 ( n75674, P1_P1_LWORD_REG_11_ );
dff P1_P1_DATAO_REG_11__reg ( clk, reset, P1_P1_DATAO_REG_11_, n9326 );
dff P1_BUF1_REG_11__reg ( clk, reset, P1_BUF1_REG_11_, n176 );
not U_inv1503 ( n75441, P1_BUF1_REG_11_ );
dff P1_P2_UWORD_REG_11__reg ( clk, reset, P1_P2_UWORD_REG_11_, n6966 );
not U_inv1504 ( n75567, P1_P2_UWORD_REG_11_ );
dff P1_P2_DATAO_REG_27__reg ( clk, reset, P1_P2_DATAO_REG_27_, n7161 );
not U_inv1505 ( n75594, P1_P2_DATAO_REG_27_ );
dff P1_BUF2_REG_27__reg ( clk, reset, P1_BUF2_REG_27_, n416 );
not U_inv1506 ( n75332, P1_BUF2_REG_27_ );
dff P1_P2_LWORD_REG_11__reg ( clk, reset, P1_P2_LWORD_REG_11_, n6891 );
not U_inv1507 ( n75640, P1_P2_LWORD_REG_11_ );
dff P1_P2_DATAO_REG_11__reg ( clk, reset, P1_P2_DATAO_REG_11_, n7081 );
not U_inv1508 ( n75534, P1_P2_DATAO_REG_11_ );
dff P1_BUF2_REG_11__reg ( clk, reset, P1_BUF2_REG_11_, n336 );
not U_inv1509 ( n75318, P1_BUF2_REG_11_ );
dff P1_P1_EAX_REG_12__reg ( clk, reset, ex_wire233, n9491 );
not U_inv1510 ( n74802, ex_wire233 );
dff P1_P1_LWORD_REG_12__reg ( clk, reset, P1_P1_LWORD_REG_12_, n9131 );
not U_inv1511 ( n75673, P1_P1_LWORD_REG_12_ );
dff P1_P1_DATAO_REG_12__reg ( clk, reset, P1_P1_DATAO_REG_12_, n9331 );
dff P1_BUF1_REG_12__reg ( clk, reset, P1_BUF1_REG_12_, n181 );
not U_inv1512 ( n75440, P1_BUF1_REG_12_ );
dff P1_P2_UWORD_REG_12__reg ( clk, reset, P1_P2_UWORD_REG_12_, n6961 );
not U_inv1513 ( n75566, P1_P2_UWORD_REG_12_ );
dff P1_P2_DATAO_REG_28__reg ( clk, reset, P1_P2_DATAO_REG_28_, n7166 );
not U_inv1514 ( n75593, P1_P2_DATAO_REG_28_ );
dff P1_BUF2_REG_28__reg ( clk, reset, P1_BUF2_REG_28_, n421 );
not U_inv1515 ( n75327, P1_BUF2_REG_28_ );
dff P1_P2_INSTQUEUE_REG_4__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__4_, n6316 );
not U_inv1516 ( n73847, P1_P2_INSTQUEUE_REG_4__4_ );
dff P1_P2_EAX_REG_20__reg ( clk, reset, P1_P2_EAX_REG_20_, n7286 );
not U_inv1517 ( n75385, P1_P2_EAX_REG_20_ );
dff P1_P2_UWORD_REG_4__reg ( clk, reset, P1_P2_UWORD_REG_4_, n7001 );
not U_inv1518 ( n75481, P1_P2_UWORD_REG_4_ );
dff P1_P2_DATAO_REG_20__reg ( clk, reset, P1_P2_DATAO_REG_20_, n7126 );
not U_inv1519 ( n75532, P1_P2_DATAO_REG_20_ );
dff P1_BUF1_REG_20__reg ( clk, reset, P1_BUF1_REG_20_, n221 );
not U_inv1520 ( n75395, P1_BUF1_REG_20_ );
dff P1_P1_INSTQUEUE_REG_15__4__reg ( clk, reset, ex_wire234, n8121 );
not U_inv1521 ( n74243, ex_wire234 );
dff P1_P1_EAX_REG_27__reg ( clk, reset, P1_P1_EAX_REG_27_, n9566 );
not U_inv1522 ( n73321, P1_P1_EAX_REG_27_ );
dff P1_P1_UWORD_REG_11__reg ( clk, reset, P1_P1_UWORD_REG_11_, n9211 );
not U_inv1523 ( n75583, P1_P1_UWORD_REG_11_ );
dff P1_P1_DATAO_REG_27__reg ( clk, reset, P1_P1_DATAO_REG_27_, n9406 );
dff P1_BUF1_REG_27__reg ( clk, reset, P1_BUF1_REG_27_, n256 );
not U_inv1524 ( n75415, P1_BUF1_REG_27_ );
dff P1_P1_INSTQUEUE_REG_0__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__3_, n8726 );
not U_inv1525 ( n74128, P1_P1_INSTQUEUE_REG_0__3_ );
dff P1_P1_INSTQUEUE_REG_1__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__3_, n8686 );
not U_inv1526 ( n74149, P1_P1_INSTQUEUE_REG_1__3_ );
dff P1_P1_INSTQUEUE_REG_2__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__3_, n8646 );
not U_inv1527 ( n74154, P1_P1_INSTQUEUE_REG_2__3_ );
dff P1_P1_INSTQUEUE_REG_3__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__3_, n8606 );
not U_inv1528 ( n74140, P1_P1_INSTQUEUE_REG_3__3_ );
dff P1_P1_INSTQUEUE_REG_4__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__3_, n8566 );
not U_inv1529 ( n74150, P1_P1_INSTQUEUE_REG_4__3_ );
dff P1_P1_INSTQUEUE_REG_5__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__3_, n8526 );
not U_inv1530 ( n74161, P1_P1_INSTQUEUE_REG_5__3_ );
dff P1_P1_INSTQUEUE_REG_6__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__3_, n8486 );
not U_inv1531 ( n74163, P1_P1_INSTQUEUE_REG_6__3_ );
dff P1_P1_INSTQUEUE_REG_7__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__3_, n8446 );
not U_inv1532 ( n74155, P1_P1_INSTQUEUE_REG_7__3_ );
dff P1_P1_INSTQUEUE_REG_8__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__3_, n8406 );
not U_inv1533 ( n74153, P1_P1_INSTQUEUE_REG_8__3_ );
dff P1_P1_INSTQUEUE_REG_9__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__3_, n8366 );
not U_inv1534 ( n74162, P1_P1_INSTQUEUE_REG_9__3_ );
dff P1_P1_INSTQUEUE_REG_10__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__3_, n8326 );
not U_inv1535 ( n74164, P1_P1_INSTQUEUE_REG_10__3_ );
dff P1_P1_INSTQUEUE_REG_11__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__3_, n8286 );
not U_inv1536 ( n74157, P1_P1_INSTQUEUE_REG_11__3_ );
dff P1_P1_INSTQUEUE_REG_12__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__3_, n8246 );
not U_inv1537 ( n74139, P1_P1_INSTQUEUE_REG_12__3_ );
dff P1_P1_INSTQUEUE_REG_13__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__3_, n8206 );
not U_inv1538 ( n74152, P1_P1_INSTQUEUE_REG_13__3_ );
dff P1_P1_INSTQUEUE_REG_14__3__reg ( clk, reset, P1_P1_INSTQUEUE_REG_14__3_, n8166 );
not U_inv1539 ( n74156, P1_P1_INSTQUEUE_REG_14__3_ );
dff P1_P1_EAX_REG_28__reg ( clk, reset, P1_P1_EAX_REG_28_, n9571 );
not U_inv1540 ( n75325, P1_P1_EAX_REG_28_ );
dff P1_P1_UWORD_REG_12__reg ( clk, reset, P1_P1_UWORD_REG_12_, n9206 );
not U_inv1541 ( n75582, P1_P1_UWORD_REG_12_ );
dff P1_P1_DATAO_REG_28__reg ( clk, reset, P1_P1_DATAO_REG_28_, n9411 );
dff P1_BUF1_REG_28__reg ( clk, reset, P1_BUF1_REG_28_, n261 );
not U_inv1542 ( n75414, P1_BUF1_REG_28_ );
dff P1_P1_INSTQUEUE_REG_0__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_0__4_, n8721 );
not U_inv1543 ( n74232, P1_P1_INSTQUEUE_REG_0__4_ );
dff P1_P1_INSTQUEUE_REG_1__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_1__4_, n8681 );
not U_inv1544 ( n74244, P1_P1_INSTQUEUE_REG_1__4_ );
dff P1_P1_INSTQUEUE_REG_2__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_2__4_, n8641 );
not U_inv1545 ( n74248, P1_P1_INSTQUEUE_REG_2__4_ );
dff P1_P1_INSTQUEUE_REG_3__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_3__4_, n8601 );
not U_inv1546 ( n74241, P1_P1_INSTQUEUE_REG_3__4_ );
dff P1_P1_INSTQUEUE_REG_4__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_4__4_, n8561 );
not U_inv1547 ( n74245, P1_P1_INSTQUEUE_REG_4__4_ );
dff P1_P1_INSTQUEUE_REG_5__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_5__4_, n8521 );
not U_inv1548 ( n74252, P1_P1_INSTQUEUE_REG_5__4_ );
dff P1_P1_INSTQUEUE_REG_6__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_6__4_, n8481 );
not U_inv1549 ( n74254, P1_P1_INSTQUEUE_REG_6__4_ );
dff P1_P1_INSTQUEUE_REG_7__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_7__4_, n8441 );
not U_inv1550 ( n74249, P1_P1_INSTQUEUE_REG_7__4_ );
dff P1_P1_INSTQUEUE_REG_8__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_8__4_, n8401 );
not U_inv1551 ( n74247, P1_P1_INSTQUEUE_REG_8__4_ );
dff P1_P1_INSTQUEUE_REG_9__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_9__4_, n8361 );
not U_inv1552 ( n74253, P1_P1_INSTQUEUE_REG_9__4_ );
dff P1_P1_INSTQUEUE_REG_10__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_10__4_, n8321 );
not U_inv1553 ( n74255, P1_P1_INSTQUEUE_REG_10__4_ );
dff P1_P1_INSTQUEUE_REG_11__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_11__4_, n8281 );
not U_inv1554 ( n74251, P1_P1_INSTQUEUE_REG_11__4_ );
dff P1_P1_INSTQUEUE_REG_12__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_12__4_, n8241 );
not U_inv1555 ( n74240, P1_P1_INSTQUEUE_REG_12__4_ );
dff P1_P1_INSTQUEUE_REG_13__4__reg ( clk, reset, P1_P1_INSTQUEUE_REG_13__4_, n8201 );
not U_inv1556 ( n74246, P1_P1_INSTQUEUE_REG_13__4_ );
dff P1_P1_EAX_REG_29__reg ( clk, reset, P1_P1_EAX_REG_29_, n9576 );
not U_inv1557 ( n75219, P1_P1_EAX_REG_29_ );
dff P1_P1_EAX_REG_19__reg ( clk, reset, P1_P1_EAX_REG_19_, n9526 );
not U_inv1558 ( n74954, P1_P1_EAX_REG_19_ );
dff P1_P1_UWORD_REG_3__reg ( clk, reset, P1_P1_UWORD_REG_3_, n9251 );
not U_inv1559 ( n75499, P1_P1_UWORD_REG_3_ );
dff P1_P1_DATAO_REG_19__reg ( clk, reset, P1_P1_DATAO_REG_19_, n9366 );
dff P1_P1_EAX_REG_20__reg ( clk, reset, ex_wire235, n9531 );
not U_inv1560 ( n74966, ex_wire235 );
dff P1_P1_UWORD_REG_4__reg ( clk, reset, P1_P1_UWORD_REG_4_, n9246 );
not U_inv1561 ( n75498, P1_P1_UWORD_REG_4_ );
dff P1_P1_DATAO_REG_20__reg ( clk, reset, P1_P1_DATAO_REG_20_, n9371 );
dff P1_BUF2_REG_20__reg ( clk, reset, P1_BUF2_REG_20_, n381 );
not U_inv1562 ( n75351, P1_BUF2_REG_20_ );
dff P1_P2_INSTQUEUE_REG_0__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__4_, n6476 );
not U_inv1563 ( n73831, P1_P2_INSTQUEUE_REG_0__4_ );
dff P1_P2_INSTQUEUE_REG_1__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__4_, n6436 );
not U_inv1564 ( n73845, P1_P2_INSTQUEUE_REG_1__4_ );
dff P1_P2_INSTQUEUE_REG_2__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__4_, n6396 );
not U_inv1565 ( n73856, P1_P2_INSTQUEUE_REG_2__4_ );
dff P1_P2_INSTQUEUE_REG_3__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__4_, n6356 );
not U_inv1566 ( n73838, P1_P2_INSTQUEUE_REG_3__4_ );
dff P1_P2_INSTQUEUE_REG_7__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__4_, n6196 );
not U_inv1567 ( n73859, P1_P2_INSTQUEUE_REG_7__4_ );
dff P1_P2_INSTQUEUE_REG_5__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__4_, n6276 );
not U_inv1568 ( n73869, P1_P2_INSTQUEUE_REG_5__4_ );
dff P1_P2_INSTQUEUE_REG_6__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__4_, n6236 );
not U_inv1569 ( n73875, P1_P2_INSTQUEUE_REG_6__4_ );
dff P1_P2_INSTQUEUE_REG_8__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__4_, n6156 );
not U_inv1570 ( n73853, P1_P2_INSTQUEUE_REG_8__4_ );
dff P1_P2_INSTQUEUE_REG_9__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__4_, n6116 );
not U_inv1571 ( n73872, P1_P2_INSTQUEUE_REG_9__4_ );
dff P1_P2_INSTQUEUE_REG_10__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__4_, n6076 );
not U_inv1572 ( n73878, P1_P2_INSTQUEUE_REG_10__4_ );
dff P1_P2_INSTQUEUE_REG_11__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__4_, n6036 );
not U_inv1573 ( n73865, P1_P2_INSTQUEUE_REG_11__4_ );
dff P1_P2_INSTQUEUE_REG_12__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__4_, n5996 );
not U_inv1574 ( n73835, P1_P2_INSTQUEUE_REG_12__4_ );
dff P1_P2_INSTQUEUE_REG_13__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__4_, n5956 );
not U_inv1575 ( n73851, P1_P2_INSTQUEUE_REG_13__4_ );
dff P1_P2_INSTQUEUE_REG_14__4__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__4_, n5916 );
not U_inv1576 ( n73862, P1_P2_INSTQUEUE_REG_14__4_ );
dff P1_P3_INSTQUEUE_REG_0__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__4_, n4231 );
not U_inv1577 ( n74221, P1_P3_INSTQUEUE_REG_0__4_ );
dff P1_P3_INSTQUEUE_REG_1__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__4_, n4191 );
not U_inv1578 ( n74226, P1_P3_INSTQUEUE_REG_1__4_ );
dff P1_P3_INSTQUEUE_REG_2__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__4_, n4151 );
not U_inv1579 ( n74230, P1_P3_INSTQUEUE_REG_2__4_ );
dff P1_P3_INSTQUEUE_REG_3__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__4_, n4111 );
not U_inv1580 ( n74223, P1_P3_INSTQUEUE_REG_3__4_ );
dff P1_P3_INSTQUEUE_REG_4__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__4_, n4071 );
not U_inv1581 ( n74227, P1_P3_INSTQUEUE_REG_4__4_ );
dff P1_P3_INSTQUEUE_REG_15__4__reg ( clk, reset, ex_wire236, n3631 );
not U_inv1582 ( n74224, ex_wire236 );
dff P1_P3_INSTQUEUE_REG_5__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__4_, n4031 );
not U_inv1583 ( n74237, P1_P3_INSTQUEUE_REG_5__4_ );
dff P1_P3_INSTQUEUE_REG_6__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__4_, n3991 );
not U_inv1584 ( n74239, P1_P3_INSTQUEUE_REG_6__4_ );
dff P1_P3_INSTQUEUE_REG_7__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__4_, n3951 );
not U_inv1585 ( n74231, P1_P3_INSTQUEUE_REG_7__4_ );
dff P1_P3_INSTQUEUE_REG_8__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__4_, n3911 );
not U_inv1586 ( n74229, P1_P3_INSTQUEUE_REG_8__4_ );
dff P1_P3_INSTQUEUE_REG_9__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__4_, n3871 );
not U_inv1587 ( n74238, P1_P3_INSTQUEUE_REG_9__4_ );
dff P1_P3_INSTQUEUE_REG_10__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__4_, n3831 );
not U_inv1588 ( n74242, P1_P3_INSTQUEUE_REG_10__4_ );
dff P1_P3_INSTQUEUE_REG_11__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__4_, n3791 );
not U_inv1589 ( n74235, P1_P3_INSTQUEUE_REG_11__4_ );
dff P1_P3_INSTQUEUE_REG_12__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__4_, n3751 );
not U_inv1590 ( n74222, P1_P3_INSTQUEUE_REG_12__4_ );
dff P1_P3_INSTQUEUE_REG_13__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__4_, n3711 );
not U_inv1591 ( n74228, P1_P3_INSTQUEUE_REG_13__4_ );
dff P1_P3_INSTQUEUE_REG_14__4__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__4_, n3671 );
not U_inv1592 ( n74233, P1_P3_INSTQUEUE_REG_14__4_ );
dff P1_P2_LWORD_REG_12__reg ( clk, reset, P1_P2_LWORD_REG_12_, n6886 );
not U_inv1593 ( n75639, P1_P2_LWORD_REG_12_ );
dff P1_P2_DATAO_REG_12__reg ( clk, reset, P1_P2_DATAO_REG_12_, n7086 );
not U_inv1594 ( n75533, P1_P2_DATAO_REG_12_ );
dff P1_BUF2_REG_12__reg ( clk, reset, P1_BUF2_REG_12_, n341 );
not U_inv1595 ( n75317, P1_BUF2_REG_12_ );
dff P1_P1_LWORD_REG_10__reg ( clk, reset, P1_P1_LWORD_REG_10_, n9141 );
not U_inv1596 ( n75672, P1_P1_LWORD_REG_10_ );
dff P1_P1_DATAO_REG_10__reg ( clk, reset, P1_P1_DATAO_REG_10_, n9321 );
dff P1_BUF1_REG_10__reg ( clk, reset, P1_BUF1_REG_10_, n171 );
not U_inv1597 ( n75439, P1_BUF1_REG_10_ );
dff P1_P1_LWORD_REG_9__reg ( clk, reset, P1_P1_LWORD_REG_9_, n9146 );
not U_inv1598 ( n75671, P1_P1_LWORD_REG_9_ );
dff P1_P1_DATAO_REG_9__reg ( clk, reset, P1_P1_DATAO_REG_9_, n9316 );
dff P1_BUF1_REG_9__reg ( clk, reset, P1_BUF1_REG_9_, n166 );
not U_inv1599 ( n75438, P1_BUF1_REG_9_ );
dff P1_P1_UWORD_REG_9__reg ( clk, reset, P1_P1_UWORD_REG_9_, n9221 );
not U_inv1600 ( n75581, P1_P1_UWORD_REG_9_ );
dff P1_P1_DATAO_REG_25__reg ( clk, reset, P1_P1_DATAO_REG_25_, n9396 );
dff P1_P2_LWORD_REG_9__reg ( clk, reset, P1_P2_LWORD_REG_9_, n6901 );
not U_inv1601 ( n75638, P1_P2_LWORD_REG_9_ );
dff P1_P2_DATAO_REG_9__reg ( clk, reset, P1_P2_DATAO_REG_9_, n7071 );
not U_inv1602 ( n75530, P1_P2_DATAO_REG_9_ );
dff P1_BUF2_REG_9__reg ( clk, reset, P1_BUF2_REG_9_, n326 );
not U_inv1603 ( n75319, P1_BUF2_REG_9_ );
dff P1_P3_LWORD_REG_9__reg ( clk, reset, P1_P3_LWORD_REG_9_, n4656 );
not U_inv1604 ( n75688, P1_P3_LWORD_REG_9_ );
dff P1_P3_DATAO_REG_9__reg ( clk, reset, P1_P3_DATAO_REG_9_, n4826 );
dff P3_IR_REG_9__reg ( clk, reset, P3_IR_REG_9_, n846 );
not U_inv1605 ( n74300, P3_IR_REG_9_ );
dff P3_IR_REG_10__reg ( clk, reset, P3_IR_REG_10_, n851 );
dff P3_REG3_REG_9__reg ( clk, reset, P3_REG3_REG_9_, n1916 );
not U_inv1606 ( n72931, P3_REG3_REG_9_ );
dff P3_REG3_REG_10__reg ( clk, reset, P3_REG3_REG_10_, n1986 );
not U_inv1607 ( n72935, P3_REG3_REG_10_ );
dff P1_BUF2_REG_19__reg ( clk, reset, P1_BUF2_REG_19_, n376 );
not U_inv1608 ( n75352, P1_BUF2_REG_19_ );
dff P1_P2_INSTQUEUE_REG_0__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__3_, n6481 );
not U_inv1609 ( n73750, P1_P2_INSTQUEUE_REG_0__3_ );
dff P1_P2_INSTQUEUE_REG_1__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__3_, n6441 );
not U_inv1610 ( n73763, P1_P2_INSTQUEUE_REG_1__3_ );
dff P1_P2_INSTQUEUE_REG_2__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__3_, n6401 );
not U_inv1611 ( n73774, P1_P2_INSTQUEUE_REG_2__3_ );
dff P1_P2_INSTQUEUE_REG_3__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__3_, n6361 );
not U_inv1612 ( n73756, P1_P2_INSTQUEUE_REG_3__3_ );
dff P1_P2_INSTQUEUE_REG_4__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__3_, n6321 );
not U_inv1613 ( n73765, P1_P2_INSTQUEUE_REG_4__3_ );
dff P1_P2_INSTQUEUE_REG_7__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__3_, n6201 );
not U_inv1614 ( n73777, P1_P2_INSTQUEUE_REG_7__3_ );
dff P1_P2_INSTQUEUE_REG_5__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__3_, n6281 );
not U_inv1615 ( n73786, P1_P2_INSTQUEUE_REG_5__3_ );
dff P1_P2_INSTQUEUE_REG_6__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__3_, n6241 );
not U_inv1616 ( n73792, P1_P2_INSTQUEUE_REG_6__3_ );
dff P1_P2_INSTQUEUE_REG_8__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__3_, n6161 );
not U_inv1617 ( n73771, P1_P2_INSTQUEUE_REG_8__3_ );
dff P1_P2_INSTQUEUE_REG_9__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__3_, n6121 );
not U_inv1618 ( n73789, P1_P2_INSTQUEUE_REG_9__3_ );
dff P1_P2_INSTQUEUE_REG_10__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__3_, n6081 );
not U_inv1619 ( n73795, P1_P2_INSTQUEUE_REG_10__3_ );
dff P1_P2_INSTQUEUE_REG_11__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__3_, n6041 );
not U_inv1620 ( n73783, P1_P2_INSTQUEUE_REG_11__3_ );
dff P1_P2_INSTQUEUE_REG_12__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__3_, n6001 );
not U_inv1621 ( n73753, P1_P2_INSTQUEUE_REG_12__3_ );
dff P1_P2_INSTQUEUE_REG_13__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__3_, n5961 );
not U_inv1622 ( n73769, P1_P2_INSTQUEUE_REG_13__3_ );
dff P1_P2_INSTQUEUE_REG_14__3__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__3_, n5921 );
not U_inv1623 ( n73780, P1_P2_INSTQUEUE_REG_14__3_ );
dff P1_P3_INSTQUEUE_REG_5__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__3_, n4036 );
not U_inv1624 ( n74134, P1_P3_INSTQUEUE_REG_5__3_ );
dff P1_P3_INSTQUEUE_REG_6__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__3_, n3996 );
not U_inv1625 ( n74137, P1_P3_INSTQUEUE_REG_6__3_ );
dff P1_P3_INSTQUEUE_REG_8__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__3_, n3916 );
not U_inv1626 ( n74125, P1_P3_INSTQUEUE_REG_8__3_ );
dff P1_P3_INSTQUEUE_REG_9__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__3_, n3876 );
not U_inv1627 ( n74136, P1_P3_INSTQUEUE_REG_9__3_ );
dff P1_P3_INSTQUEUE_REG_10__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__3_, n3836 );
not U_inv1628 ( n74142, P1_P3_INSTQUEUE_REG_10__3_ );
dff P1_P3_INSTQUEUE_REG_11__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__3_, n3796 );
not U_inv1629 ( n74131, P1_P3_INSTQUEUE_REG_11__3_ );
dff P1_P3_INSTQUEUE_REG_12__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__3_, n3756 );
not U_inv1630 ( n74102, P1_P3_INSTQUEUE_REG_12__3_ );
dff P1_P3_INSTQUEUE_REG_13__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__3_, n3716 );
not U_inv1631 ( n74124, P1_P3_INSTQUEUE_REG_13__3_ );
dff P1_P3_INSTQUEUE_REG_14__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__3_, n3676 );
not U_inv1632 ( n74129, P1_P3_INSTQUEUE_REG_14__3_ );
dff P1_P3_INSTQUEUE_REG_0__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__3_, n4236 );
not U_inv1633 ( n74063, P1_P3_INSTQUEUE_REG_0__3_ );
dff P1_P3_INSTQUEUE_REG_1__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__3_, n4196 );
not U_inv1634 ( n74121, P1_P3_INSTQUEUE_REG_1__3_ );
dff P1_P3_INSTQUEUE_REG_2__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__3_, n4156 );
not U_inv1635 ( n74126, P1_P3_INSTQUEUE_REG_2__3_ );
dff P1_P3_INSTQUEUE_REG_3__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__3_, n4116 );
not U_inv1636 ( n74104, P1_P3_INSTQUEUE_REG_3__3_ );
dff P1_P3_INSTQUEUE_REG_4__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__3_, n4076 );
not U_inv1637 ( n74122, P1_P3_INSTQUEUE_REG_4__3_ );
dff P1_P3_INSTQUEUE_REG_7__3__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__3_, n3956 );
not U_inv1638 ( n74127, P1_P3_INSTQUEUE_REG_7__3_ );
dff P1_P3_INSTQUEUE_REG_15__3__reg ( clk, reset, ex_wire237, n3636 );
not U_inv1639 ( n74107, ex_wire237 );
dff P1_P1_UWORD_REG_5__reg ( clk, reset, P1_P1_UWORD_REG_5_, n9241 );
not U_inv1640 ( n75497, P1_P1_UWORD_REG_5_ );
dff P1_P1_DATAO_REG_21__reg ( clk, reset, P1_P1_DATAO_REG_21_, n9376 );
dff P1_P1_EAX_REG_13__reg ( clk, reset, P1_P1_EAX_REG_13_, n9496 );
not U_inv1641 ( n74843, P1_P1_EAX_REG_13_ );
dff P1_BUF2_REG_21__reg ( clk, reset, P1_BUF2_REG_21_, n386 );
not U_inv1642 ( n75350, P1_BUF2_REG_21_ );
dff P1_P2_INSTQUEUE_REG_0__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__5_, n6471 );
not U_inv1643 ( n73899, P1_P2_INSTQUEUE_REG_0__5_ );
dff P1_P2_INSTQUEUE_REG_1__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__5_, n6431 );
not U_inv1644 ( n73914, P1_P2_INSTQUEUE_REG_1__5_ );
dff P1_P2_INSTQUEUE_REG_2__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__5_, n6391 );
not U_inv1645 ( n73925, P1_P2_INSTQUEUE_REG_2__5_ );
dff P1_P2_INSTQUEUE_REG_3__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__5_, n6351 );
not U_inv1646 ( n73905, P1_P2_INSTQUEUE_REG_3__5_ );
dff P1_P2_INSTQUEUE_REG_4__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__5_, n6311 );
not U_inv1647 ( n73916, P1_P2_INSTQUEUE_REG_4__5_ );
dff P1_P2_INSTQUEUE_REG_7__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__5_, n6191 );
not U_inv1648 ( n73928, P1_P2_INSTQUEUE_REG_7__5_ );
dff P1_P2_INSTQUEUE_REG_5__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__5_, n6271 );
not U_inv1649 ( n73937, P1_P2_INSTQUEUE_REG_5__5_ );
dff P1_P2_INSTQUEUE_REG_6__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__5_, n6231 );
not U_inv1650 ( n73943, P1_P2_INSTQUEUE_REG_6__5_ );
dff P1_P2_INSTQUEUE_REG_8__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__5_, n6151 );
not U_inv1651 ( n73922, P1_P2_INSTQUEUE_REG_8__5_ );
dff P1_P2_INSTQUEUE_REG_9__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__5_, n6111 );
not U_inv1652 ( n73940, P1_P2_INSTQUEUE_REG_9__5_ );
dff P1_P2_INSTQUEUE_REG_10__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__5_, n6071 );
not U_inv1653 ( n73946, P1_P2_INSTQUEUE_REG_10__5_ );
dff P1_P2_INSTQUEUE_REG_11__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__5_, n6031 );
not U_inv1654 ( n73934, P1_P2_INSTQUEUE_REG_11__5_ );
dff P1_P2_INSTQUEUE_REG_12__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__5_, n5991 );
not U_inv1655 ( n73902, P1_P2_INSTQUEUE_REG_12__5_ );
dff P1_P2_INSTQUEUE_REG_13__5__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__5_, n5951 );
not U_inv1656 ( n73920, P1_P2_INSTQUEUE_REG_13__5_ );
dff P1_P1_EAX_REG_0__reg ( clk, reset, P1_P1_EAX_REG_0_, n9431 );
not U_inv1657 ( n73162, P1_P1_EAX_REG_0_ );
dff P1_P1_LWORD_REG_0__reg ( clk, reset, P1_P1_LWORD_REG_0_, n9191 );
not U_inv1658 ( n75669, P1_P1_LWORD_REG_0_ );
dff P1_P2_INSTQUEUE_REG_5__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__0_, n6296 );
not U_inv1659 ( n73694, P1_P2_INSTQUEUE_REG_5__0_ );
dff P1_P2_INSTQUEUE_REG_6__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__0_, n6256 );
not U_inv1660 ( n73700, P1_P2_INSTQUEUE_REG_6__0_ );
dff P1_P2_INSTQUEUE_REG_7__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__0_, n6216 );
not U_inv1661 ( n73685, P1_P2_INSTQUEUE_REG_7__0_ );
dff P1_P2_INSTQUEUE_REG_8__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__0_, n6176 );
not U_inv1662 ( n73680, P1_P2_INSTQUEUE_REG_8__0_ );
dff P1_P2_INSTQUEUE_REG_9__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__0_, n6136 );
not U_inv1663 ( n73697, P1_P2_INSTQUEUE_REG_9__0_ );
dff P1_P2_INSTQUEUE_REG_10__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__0_, n6096 );
not U_inv1664 ( n73704, P1_P2_INSTQUEUE_REG_10__0_ );
dff P1_P2_INSTQUEUE_REG_11__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__0_, n6056 );
not U_inv1665 ( n73691, P1_P2_INSTQUEUE_REG_11__0_ );
dff P1_P2_INSTQUEUE_REG_12__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__0_, n6016 );
not U_inv1666 ( n73654, P1_P2_INSTQUEUE_REG_12__0_ );
dff P1_P2_INSTQUEUE_REG_13__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__0_, n5976 );
not U_inv1667 ( n73678, P1_P2_INSTQUEUE_REG_13__0_ );
dff P1_P2_INSTQUEUE_REG_14__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__0_, n5936 );
not U_inv1668 ( n73689, P1_P2_INSTQUEUE_REG_14__0_ );
dff P1_P2_INSTQUEUE_REG_0__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__0_, n6496 );
not U_inv1669 ( n73641, P1_P2_INSTQUEUE_REG_0__0_ );
dff P1_P2_EBX_REG_0__reg ( clk, reset, P1_P2_EBX_REG_0_, n7346 );
not U_inv1670 ( n73120, P1_P2_EBX_REG_0_ );
dff P1_P2_INSTQUEUE_REG_1__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__0_, n6456 );
not U_inv1671 ( n73669, P1_P2_INSTQUEUE_REG_1__0_ );
dff P1_P2_INSTQUEUE_REG_2__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__0_, n6416 );
not U_inv1672 ( n73683, P1_P2_INSTQUEUE_REG_2__0_ );
dff P1_P2_INSTQUEUE_REG_3__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__0_, n6376 );
not U_inv1673 ( n73658, P1_P2_INSTQUEUE_REG_3__0_ );
dff P1_P2_INSTQUEUE_REG_4__0__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__0_, n6336 );
not U_inv1674 ( n73673, P1_P2_INSTQUEUE_REG_4__0_ );
dff P1_P1_UWORD_REG_7__reg ( clk, reset, P1_P1_UWORD_REG_7_, n9231 );
not U_inv1675 ( n75496, P1_P1_UWORD_REG_7_ );
dff P1_P1_DATAO_REG_23__reg ( clk, reset, P1_P1_DATAO_REG_23_, n9386 );
dff P1_P1_EAX_REG_14__reg ( clk, reset, P1_P1_EAX_REG_14_, n9501 );
not U_inv1676 ( n73252, P1_P1_EAX_REG_14_ );
dff P1_P1_LWORD_REG_14__reg ( clk, reset, P1_P1_LWORD_REG_14_, n9121 );
not U_inv1677 ( n75670, P1_P1_LWORD_REG_14_ );
dff P1_P1_DATAO_REG_14__reg ( clk, reset, P1_P1_DATAO_REG_14_, n9341 );
dff P1_BUF1_REG_14__reg ( clk, reset, P1_BUF1_REG_14_, n191 );
not U_inv1678 ( n75437, P1_BUF1_REG_14_ );
dff P1_P1_EAX_REG_30__reg ( clk, reset, P1_P1_EAX_REG_30_, n9581 );
not U_inv1679 ( n75405, P1_P1_EAX_REG_30_ );
dff P1_P1_UWORD_REG_14__reg ( clk, reset, P1_P1_UWORD_REG_14_, n9196 );
not U_inv1680 ( n75580, P1_P1_UWORD_REG_14_ );
dff P1_P1_DATAO_REG_30__reg ( clk, reset, P1_P1_DATAO_REG_30_, n9421 );
not U_inv1681 ( n73433, P1_P1_DATAO_REG_30_ );
dff P1_BUF1_REG_30__reg ( clk, reset, P1_BUF1_REG_30_, n271 );
not U_inv1682 ( n75413, P1_BUF1_REG_30_ );
dff P1_P2_LWORD_REG_14__reg ( clk, reset, P1_P2_LWORD_REG_14_, n6876 );
not U_inv1683 ( n75637, P1_P2_LWORD_REG_14_ );
dff P1_P2_DATAO_REG_14__reg ( clk, reset, P1_P2_DATAO_REG_14_, n7096 );
not U_inv1684 ( n75529, P1_P2_DATAO_REG_14_ );
dff P1_BUF2_REG_14__reg ( clk, reset, P1_BUF2_REG_14_, n351 );
not U_inv1685 ( n75311, P1_BUF2_REG_14_ );
dff P1_BUF2_REG_22__reg ( clk, reset, P1_BUF2_REG_22_, n391 );
not U_inv1686 ( n75349, P1_BUF2_REG_22_ );
dff P1_P2_INSTQUEUE_REG_0__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__6_, n6466 );
not U_inv1687 ( n74029, P1_P2_INSTQUEUE_REG_0__6_ );
dff P1_P2_INSTQUEUE_REG_1__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__6_, n6426 );
not U_inv1688 ( n74068, P1_P2_INSTQUEUE_REG_1__6_ );
dff P1_P2_INSTQUEUE_REG_2__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__6_, n6386 );
not U_inv1689 ( n74081, P1_P2_INSTQUEUE_REG_2__6_ );
dff P1_P2_INSTQUEUE_REG_3__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__6_, n6346 );
not U_inv1690 ( n74055, P1_P2_INSTQUEUE_REG_3__6_ );
dff P1_P2_INSTQUEUE_REG_7__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__6_, n6186 );
not U_inv1691 ( n74087, P1_P2_INSTQUEUE_REG_7__6_ );
dff P1_P2_INSTQUEUE_REG_5__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__6_, n6266 );
not U_inv1692 ( n74110, P1_P2_INSTQUEUE_REG_5__6_ );
dff P1_P2_INSTQUEUE_REG_6__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__6_, n6226 );
not U_inv1693 ( n74117, P1_P2_INSTQUEUE_REG_6__6_ );
dff P1_P2_INSTQUEUE_REG_8__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__6_, n6146 );
not U_inv1694 ( n74078, P1_P2_INSTQUEUE_REG_8__6_ );
dff P1_P2_INSTQUEUE_REG_9__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__6_, n6106 );
not U_inv1695 ( n74114, P1_P2_INSTQUEUE_REG_9__6_ );
dff P1_P2_INSTQUEUE_REG_10__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__6_, n6066 );
not U_inv1696 ( n74120, P1_P2_INSTQUEUE_REG_10__6_ );
dff P1_P2_INSTQUEUE_REG_11__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__6_, n6026 );
not U_inv1697 ( n74096, P1_P2_INSTQUEUE_REG_11__6_ );
dff P1_P2_INSTQUEUE_REG_12__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__6_, n5986 );
not U_inv1698 ( n74051, P1_P2_INSTQUEUE_REG_12__6_ );
dff P1_P2_INSTQUEUE_REG_13__6__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__6_, n5946 );
not U_inv1699 ( n74076, P1_P2_INSTQUEUE_REG_13__6_ );
dff P1_P2_EAX_REG_23__reg ( clk, reset, P1_P2_EAX_REG_23_, n7301 );
not U_inv1700 ( n74972, P1_P2_EAX_REG_23_ );
dff P1_P2_UWORD_REG_7__reg ( clk, reset, P1_P2_UWORD_REG_7_, n6986 );
not U_inv1701 ( n75480, P1_P2_UWORD_REG_7_ );
dff P1_P2_DATAO_REG_23__reg ( clk, reset, P1_P2_DATAO_REG_23_, n7141 );
not U_inv1702 ( n75528, P1_P2_DATAO_REG_23_ );
dff P1_BUF1_REG_23__reg ( clk, reset, P1_BUF1_REG_23_, n236 );
not U_inv1703 ( n75394, P1_BUF1_REG_23_ );
dff P1_BUF2_REG_23__reg ( clk, reset, P1_BUF2_REG_23_, n396 );
not U_inv1704 ( n75348, P1_BUF2_REG_23_ );
dff P1_P2_INSTQUEUE_REG_0__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__7_, n6461 );
not U_inv1705 ( n74168, P1_P2_INSTQUEUE_REG_0__7_ );
dff P1_P2_INSTQUEUE_REG_1__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__7_, n6421 );
not U_inv1706 ( n74182, P1_P2_INSTQUEUE_REG_1__7_ );
dff P1_P2_INSTQUEUE_REG_2__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__7_, n6381 );
not U_inv1707 ( n74187, P1_P2_INSTQUEUE_REG_2__7_ );
dff P1_P2_INSTQUEUE_REG_3__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__7_, n6341 );
not U_inv1708 ( n74172, P1_P2_INSTQUEUE_REG_3__7_ );
dff P1_P2_INSTQUEUE_REG_4__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__7_, n6301 );
not U_inv1709 ( n74184, P1_P2_INSTQUEUE_REG_4__7_ );
dff P1_P2_INSTQUEUE_REG_7__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__7_, n6181 );
not U_inv1710 ( n74196, P1_P2_INSTQUEUE_REG_7__7_ );
dff P1_P2_INSTQUEUE_REG_5__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__7_, n6261 );
not U_inv1711 ( n74206, P1_P2_INSTQUEUE_REG_5__7_ );
dff P1_P2_INSTQUEUE_REG_6__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__7_, n6221 );
not U_inv1712 ( n74212, P1_P2_INSTQUEUE_REG_6__7_ );
dff P1_P2_INSTQUEUE_REG_8__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__7_, n6141 );
not U_inv1713 ( n74193, P1_P2_INSTQUEUE_REG_8__7_ );
dff P1_P2_INSTQUEUE_REG_9__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__7_, n6101 );
not U_inv1714 ( n74209, P1_P2_INSTQUEUE_REG_9__7_ );
dff P1_P2_INSTQUEUE_REG_10__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__7_, n6061 );
not U_inv1715 ( n74215, P1_P2_INSTQUEUE_REG_10__7_ );
dff P1_P2_INSTQUEUE_REG_11__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__7_, n6021 );
not U_inv1716 ( n74203, P1_P2_INSTQUEUE_REG_11__7_ );
dff P1_P2_INSTQUEUE_REG_12__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__7_, n5981 );
not U_inv1717 ( n74175, P1_P2_INSTQUEUE_REG_12__7_ );
dff P1_P2_INSTQUEUE_REG_13__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__7_, n5941 );
not U_inv1718 ( n74190, P1_P2_INSTQUEUE_REG_13__7_ );
dff P1_P2_INSTQUEUE_REG_14__7__reg ( clk, reset, P1_P2_INSTQUEUE_REG_14__7_, n5901 );
not U_inv1719 ( n74200, P1_P2_INSTQUEUE_REG_14__7_ );
dff P1_P2_EAX_REG_26__reg ( clk, reset, P1_P2_EAX_REG_26_, n7316 );
not U_inv1720 ( n75345, P1_P2_EAX_REG_26_ );
dff P1_P3_INSTQUEUE_REG_5__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__7_, n4016 );
not U_inv1721 ( n74352, P1_P3_INSTQUEUE_REG_5__7_ );
dff P1_P3_INSTQUEUE_REG_6__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__7_, n3976 );
not U_inv1722 ( n74354, P1_P3_INSTQUEUE_REG_6__7_ );
dff P1_P3_INSTQUEUE_REG_8__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__7_, n3896 );
not U_inv1723 ( n74348, P1_P3_INSTQUEUE_REG_8__7_ );
dff P1_P3_INSTQUEUE_REG_9__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__7_, n3856 );
not U_inv1724 ( n74353, P1_P3_INSTQUEUE_REG_9__7_ );
dff P1_P3_INSTQUEUE_REG_10__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__7_, n3816 );
not U_inv1725 ( n74355, P1_P3_INSTQUEUE_REG_10__7_ );
dff P1_P3_INSTQUEUE_REG_11__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__7_, n3776 );
not U_inv1726 ( n74351, P1_P3_INSTQUEUE_REG_11__7_ );
dff P1_P3_INSTQUEUE_REG_12__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__7_, n3736 );
not U_inv1727 ( n74340, P1_P3_INSTQUEUE_REG_12__7_ );
dff P1_P3_INSTQUEUE_REG_13__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__7_, n3696 );
not U_inv1728 ( n74347, P1_P3_INSTQUEUE_REG_13__7_ );
dff P1_P3_INSTQUEUE_REG_14__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__7_, n3656 );
not U_inv1729 ( n74350, P1_P3_INSTQUEUE_REG_14__7_ );
dff P1_P3_INSTQUEUE_REG_0__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__7_, n4216 );
not U_inv1730 ( n74338, P1_P3_INSTQUEUE_REG_0__7_ );
dff P1_P3_INSTQUEUE_REG_1__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__7_, n4176 );
not U_inv1731 ( n74343, P1_P3_INSTQUEUE_REG_1__7_ );
dff P1_P3_INSTQUEUE_REG_2__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__7_, n4136 );
not U_inv1732 ( n74345, P1_P3_INSTQUEUE_REG_2__7_ );
dff P1_P3_INSTQUEUE_REG_3__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__7_, n4096 );
not U_inv1733 ( n74339, P1_P3_INSTQUEUE_REG_3__7_ );
dff P1_P3_INSTQUEUE_REG_4__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__7_, n4056 );
not U_inv1734 ( n74344, P1_P3_INSTQUEUE_REG_4__7_ );
dff P1_P3_INSTQUEUE_REG_7__7__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__7_, n3936 );
not U_inv1735 ( n74349, P1_P3_INSTQUEUE_REG_7__7_ );
dff P1_P3_INSTQUEUE_REG_14__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__6_, n3661 );
not U_inv1736 ( n74311, P1_P3_INSTQUEUE_REG_14__6_ );
dff P1_P3_INSTQUEUE_REG_0__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__6_, n4221 );
not U_inv1737 ( n74299, P1_P3_INSTQUEUE_REG_0__6_ );
dff P1_P3_INSTQUEUE_REG_1__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__6_, n4181 );
not U_inv1738 ( n74305, P1_P3_INSTQUEUE_REG_1__6_ );
dff P1_P3_INSTQUEUE_REG_2__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__6_, n4141 );
not U_inv1739 ( n74309, P1_P3_INSTQUEUE_REG_2__6_ );
dff P1_P3_INSTQUEUE_REG_3__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__6_, n4101 );
not U_inv1740 ( n74303, P1_P3_INSTQUEUE_REG_3__6_ );
dff P1_P3_INSTQUEUE_REG_4__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__6_, n4061 );
not U_inv1741 ( n74306, P1_P3_INSTQUEUE_REG_4__6_ );
dff P1_P3_INSTQUEUE_REG_5__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__6_, n4021 );
not U_inv1742 ( n74313, P1_P3_INSTQUEUE_REG_5__6_ );
dff P1_P3_INSTQUEUE_REG_6__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__6_, n3981 );
not U_inv1743 ( n74316, P1_P3_INSTQUEUE_REG_6__6_ );
dff P1_P3_INSTQUEUE_REG_7__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__6_, n3941 );
not U_inv1744 ( n74310, P1_P3_INSTQUEUE_REG_7__6_ );
dff P1_P3_INSTQUEUE_REG_8__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__6_, n3901 );
not U_inv1745 ( n74308, P1_P3_INSTQUEUE_REG_8__6_ );
dff P1_P3_INSTQUEUE_REG_9__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__6_, n3861 );
not U_inv1746 ( n74315, P1_P3_INSTQUEUE_REG_9__6_ );
dff P1_P3_INSTQUEUE_REG_10__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__6_, n3821 );
not U_inv1747 ( n74317, P1_P3_INSTQUEUE_REG_10__6_ );
dff P1_P3_INSTQUEUE_REG_11__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__6_, n3781 );
not U_inv1748 ( n74312, P1_P3_INSTQUEUE_REG_11__6_ );
dff P1_P3_INSTQUEUE_REG_12__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__6_, n3741 );
not U_inv1749 ( n74302, P1_P3_INSTQUEUE_REG_12__6_ );
dff P1_P3_INSTQUEUE_REG_13__6__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__6_, n3701 );
not U_inv1750 ( n74307, P1_P3_INSTQUEUE_REG_13__6_ );
dff P1_P3_INSTQUEUE_REG_15__6__reg ( clk, reset, ex_wire238, n3621 );
not U_inv1751 ( n74304, ex_wire238 );
dff P1_P3_INSTQUEUE_REG_14__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__5_, n3666 );
not U_inv1752 ( n74271, P1_P3_INSTQUEUE_REG_14__5_ );
dff P1_P3_INSTQUEUE_REG_0__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__5_, n4226 );
not U_inv1753 ( n74258, P1_P3_INSTQUEUE_REG_0__5_ );
dff P1_P3_INSTQUEUE_REG_1__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__5_, n4186 );
not U_inv1754 ( n74264, P1_P3_INSTQUEUE_REG_1__5_ );
dff P1_P3_INSTQUEUE_REG_2__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__5_, n4146 );
not U_inv1755 ( n74269, P1_P3_INSTQUEUE_REG_2__5_ );
dff P1_P3_INSTQUEUE_REG_3__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__5_, n4106 );
not U_inv1756 ( n74261, P1_P3_INSTQUEUE_REG_3__5_ );
dff P1_P3_INSTQUEUE_REG_4__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__5_, n4066 );
not U_inv1757 ( n74265, P1_P3_INSTQUEUE_REG_4__5_ );
dff P1_P3_INSTQUEUE_REG_5__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__5_, n4026 );
not U_inv1758 ( n74275, P1_P3_INSTQUEUE_REG_5__5_ );
dff P1_P3_INSTQUEUE_REG_6__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__5_, n3986 );
not U_inv1759 ( n74277, P1_P3_INSTQUEUE_REG_6__5_ );
dff P1_P3_INSTQUEUE_REG_7__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__5_, n3946 );
not U_inv1760 ( n74270, P1_P3_INSTQUEUE_REG_7__5_ );
dff P1_P3_INSTQUEUE_REG_8__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__5_, n3906 );
not U_inv1761 ( n74268, P1_P3_INSTQUEUE_REG_8__5_ );
dff P1_P3_INSTQUEUE_REG_9__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__5_, n3866 );
not U_inv1762 ( n74276, P1_P3_INSTQUEUE_REG_9__5_ );
dff P1_P3_INSTQUEUE_REG_10__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__5_, n3826 );
not U_inv1763 ( n74278, P1_P3_INSTQUEUE_REG_10__5_ );
dff P1_P3_INSTQUEUE_REG_11__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__5_, n3786 );
not U_inv1764 ( n74272, P1_P3_INSTQUEUE_REG_11__5_ );
dff P1_P3_INSTQUEUE_REG_12__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__5_, n3746 );
not U_inv1765 ( n74260, P1_P3_INSTQUEUE_REG_12__5_ );
dff P1_P3_INSTQUEUE_REG_13__5__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__5_, n3706 );
not U_inv1766 ( n74267, P1_P3_INSTQUEUE_REG_13__5_ );
dff P1_P3_INSTQUEUE_REG_15__5__reg ( clk, reset, ex_wire239, n3626 );
not U_inv1767 ( n74262, ex_wire239 );
dff P1_P3_EAX_REG_20__reg ( clk, reset, P1_P3_EAX_REG_20_, n5041 );
dff P1_P3_EAX_REG_21__reg ( clk, reset, P1_P3_EAX_REG_21_, n5046 );
not U_inv1768 ( n74927, P1_P3_EAX_REG_21_ );
dff P1_P3_EAX_REG_22__reg ( clk, reset, P1_P3_EAX_REG_22_, n5051 );
dff P1_P3_EAX_REG_23__reg ( clk, reset, P1_P3_EAX_REG_23_, n5056 );
not U_inv1769 ( n74984, P1_P3_EAX_REG_23_ );
dff P1_P3_EAX_REG_11__reg ( clk, reset, P1_P3_EAX_REG_11_, n4996 );
not U_inv1770 ( n74676, P1_P3_EAX_REG_11_ );
dff P1_P3_LWORD_REG_11__reg ( clk, reset, P1_P3_LWORD_REG_11_, n4646 );
not U_inv1771 ( n75687, P1_P3_LWORD_REG_11_ );
dff P1_P3_DATAO_REG_11__reg ( clk, reset, P1_P3_DATAO_REG_11_, n4836 );
dff P3_IR_REG_11__reg ( clk, reset, P3_IR_REG_11_, n856 );
not U_inv1772 ( n74301, P3_IR_REG_11_ );
dff P3_REG3_REG_11__reg ( clk, reset, P3_REG3_REG_11_, n1891 );
not U_inv1773 ( n72937, P3_REG3_REG_11_ );
dff P1_P3_EAX_REG_12__reg ( clk, reset, P1_P3_EAX_REG_12_, n5001 );
not U_inv1774 ( n75280, P1_P3_EAX_REG_12_ );
dff P1_P3_LWORD_REG_12__reg ( clk, reset, P1_P3_LWORD_REG_12_, n4641 );
not U_inv1775 ( n75686, P1_P3_LWORD_REG_12_ );
dff P1_P3_DATAO_REG_12__reg ( clk, reset, P1_P3_DATAO_REG_12_, n4841 );
dff P3_IR_REG_12__reg ( clk, reset, P3_IR_REG_12_, n861 );
dff P3_REG3_REG_12__reg ( clk, reset, P3_REG3_REG_12_, n1951 );
not U_inv1776 ( n72942, P3_REG3_REG_12_ );
dff P1_P3_EAX_REG_13__reg ( clk, reset, P1_P3_EAX_REG_13_, n5006 );
not U_inv1777 ( n74731, P1_P3_EAX_REG_13_ );
dff P1_P3_LWORD_REG_13__reg ( clk, reset, P1_P3_LWORD_REG_13_, n4636 );
not U_inv1778 ( n75685, P1_P3_LWORD_REG_13_ );
dff P1_P3_DATAO_REG_13__reg ( clk, reset, P1_P3_DATAO_REG_13_, n4846 );
dff P3_IR_REG_13__reg ( clk, reset, P3_IR_REG_13_, n866 );
not U_inv1779 ( n74392, P3_IR_REG_13_ );
dff P3_REG3_REG_13__reg ( clk, reset, P3_REG3_REG_13_, n1901 );
not U_inv1780 ( n72939, P3_REG3_REG_13_ );
dff P1_P3_EAX_REG_14__reg ( clk, reset, P1_P3_EAX_REG_14_, n5011 );
not U_inv1781 ( n75278, P1_P3_EAX_REG_14_ );
dff P1_P3_LWORD_REG_14__reg ( clk, reset, P1_P3_LWORD_REG_14_, n4631 );
not U_inv1782 ( n75684, P1_P3_LWORD_REG_14_ );
dff P1_P3_DATAO_REG_14__reg ( clk, reset, P1_P3_DATAO_REG_14_, n4851 );
dff P3_IR_REG_14__reg ( clk, reset, P3_IR_REG_14_, n871 );
dff P3_IR_REG_15__reg ( clk, reset, P3_IR_REG_15_, n876 );
not U_inv1783 ( n74395, P3_IR_REG_15_ );
dff P3_REG3_REG_14__reg ( clk, reset, P3_REG3_REG_14_, n1996 );
not U_inv1784 ( n72949, P3_REG3_REG_14_ );
dff P3_REG3_REG_15__reg ( clk, reset, P3_REG3_REG_15_, n1866 );
not U_inv1785 ( n72943, P3_REG3_REG_15_ );
dff P1_P3_PHYADDRPOINTER_REG_0__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_0_, n4466 );
not U_inv1786 ( n75221, P1_P3_PHYADDRPOINTER_REG_0_ );
dff P1_P1_LWORD_REG_1__reg ( clk, reset, P1_P1_LWORD_REG_1_, n9186 );
not U_inv1787 ( n75680, P1_P1_LWORD_REG_1_ );
dff P1_P1_DATAO_REG_0__reg ( clk, reset, P1_P1_DATAO_REG_0_, n9271 );
dff P1_P1_ADDRESS_REG_4__reg ( clk, reset, P1_P1_ADDRESS_REG_4_, n7886 );
not U_inv1788 ( n73477, P1_P1_ADDRESS_REG_4_ );
dff P1_P1_ADDRESS_REG_16__reg ( clk, reset, P1_P1_ADDRESS_REG_16_, n7826 );
not U_inv1789 ( n73483, P1_P1_ADDRESS_REG_16_ );
dff P1_P1_ADDRESS_REG_28__reg ( clk, reset, P1_P1_ADDRESS_REG_28_, n7766 );
dff P1_P1_CODEFETCH_REG_reg ( clk, reset, P1_P1_CODEFETCH_REG, n9966 );
dff P1_P1_D_C_N_REG_reg ( clk, reset, P1_P1_D_C_N_REG, n9956 );
dff P1_P1_MORE_REG_reg ( clk, reset, P1_P1_MORE_REG, n9941 );
dff P1_P1_READREQUEST_REG_reg ( clk, reset, P1_P1_READREQUEST_REG, n9976 );
dff P1_P1_W_R_N_REG_reg ( clk, reset, P1_P1_W_R_N_REG, n9931 );
dff P1_P1_PHYADDRPOINTER_REG_1__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_1_, n8961 );
not U_inv1790 ( n74477, P1_P1_PHYADDRPOINTER_REG_1_ );
dff P1_P1_EBX_REG_0__reg ( clk, reset, P1_P1_EBX_REG_0_, n9591 );
not U_inv1791 ( n73126, P1_P1_EBX_REG_0_ );
dff P1_P1_EBX_REG_2__reg ( clk, reset, P1_P1_EBX_REG_2_, n9601 );
not U_inv1792 ( n74533, P1_P1_EBX_REG_2_ );
dff P1_P1_EBX_REG_3__reg ( clk, reset, P1_P1_EBX_REG_3_, n9606 );
not U_inv1793 ( n73143, P1_P1_EBX_REG_3_ );
dff P1_P1_EBX_REG_4__reg ( clk, reset, P1_P1_EBX_REG_4_, n9611 );
not U_inv1794 ( n74569, P1_P1_EBX_REG_4_ );
dff P1_P1_EBX_REG_5__reg ( clk, reset, P1_P1_EBX_REG_5_, n9616 );
not U_inv1795 ( n73157, P1_P1_EBX_REG_5_ );
dff P1_P1_EBX_REG_6__reg ( clk, reset, P1_P1_EBX_REG_6_, n9621 );
not U_inv1796 ( n74602, P1_P1_EBX_REG_6_ );
dff P1_P1_EBX_REG_7__reg ( clk, reset, P1_P1_EBX_REG_7_, n9626 );
not U_inv1797 ( n73175, P1_P1_EBX_REG_7_ );
dff P1_P1_EBX_REG_8__reg ( clk, reset, P1_P1_EBX_REG_8_, n9631 );
not U_inv1798 ( n74665, P1_P1_EBX_REG_8_ );
dff P1_P1_EBX_REG_9__reg ( clk, reset, P1_P1_EBX_REG_9_, n9636 );
not U_inv1799 ( n73205, P1_P1_EBX_REG_9_ );
dff P1_P1_EBX_REG_10__reg ( clk, reset, P1_P1_EBX_REG_10_, n9641 );
not U_inv1800 ( n74721, P1_P1_EBX_REG_10_ );
dff P1_P1_EBX_REG_11__reg ( clk, reset, P1_P1_EBX_REG_11_, n9646 );
not U_inv1801 ( n73213, P1_P1_EBX_REG_11_ );
dff P1_P1_EBX_REG_12__reg ( clk, reset, P1_P1_EBX_REG_12_, n9651 );
not U_inv1802 ( n74764, P1_P1_EBX_REG_12_ );
dff P1_P1_EBX_REG_13__reg ( clk, reset, P1_P1_EBX_REG_13_, n9656 );
not U_inv1803 ( n73231, P1_P1_EBX_REG_13_ );
dff P1_P1_EBX_REG_14__reg ( clk, reset, P1_P1_EBX_REG_14_, n9661 );
not U_inv1804 ( n74794, P1_P1_EBX_REG_14_ );
dff P1_P1_EBX_REG_17__reg ( clk, reset, P1_P1_EBX_REG_17_, n9676 );
not U_inv1805 ( n73260, P1_P1_EBX_REG_17_ );
dff P1_P1_EBX_REG_18__reg ( clk, reset, P1_P1_EBX_REG_18_, n9681 );
not U_inv1806 ( n74895, P1_P1_EBX_REG_18_ );
dff P1_P1_EBX_REG_19__reg ( clk, reset, P1_P1_EBX_REG_19_, n9686 );
not U_inv1807 ( n73274, P1_P1_EBX_REG_19_ );
dff P1_P1_EBX_REG_20__reg ( clk, reset, P1_P1_EBX_REG_20_, n9691 );
not U_inv1808 ( n74935, P1_P1_EBX_REG_20_ );
dff P1_P1_EBX_REG_21__reg ( clk, reset, P1_P1_EBX_REG_21_, n9696 );
not U_inv1809 ( n73287, P1_P1_EBX_REG_21_ );
dff P1_P1_EBX_REG_22__reg ( clk, reset, P1_P1_EBX_REG_22_, n9701 );
not U_inv1810 ( n74981, P1_P1_EBX_REG_22_ );
dff P1_P1_EBX_REG_23__reg ( clk, reset, P1_P1_EBX_REG_23_, n9706 );
not U_inv1811 ( n73303, P1_P1_EBX_REG_23_ );
dff P1_P1_EBX_REG_24__reg ( clk, reset, P1_P1_EBX_REG_24_, n9711 );
not U_inv1812 ( n75025, P1_P1_EBX_REG_24_ );
dff P1_P1_EBX_REG_25__reg ( clk, reset, P1_P1_EBX_REG_25_, n9716 );
not U_inv1813 ( n73315, P1_P1_EBX_REG_25_ );
dff P1_P1_EBX_REG_26__reg ( clk, reset, P1_P1_EBX_REG_26_, n9721 );
not U_inv1814 ( n75075, P1_P1_EBX_REG_26_ );
dff P1_P1_EBX_REG_27__reg ( clk, reset, P1_P1_EBX_REG_27_, n9726 );
not U_inv1815 ( n75176, P1_P1_EBX_REG_27_ );
dff P1_P1_EBX_REG_28__reg ( clk, reset, P1_P1_EBX_REG_28_, n9731 );
not U_inv1816 ( n73384, P1_P1_EBX_REG_28_ );
dff P1_P1_EBX_REG_29__reg ( clk, reset, P1_P1_EBX_REG_29_, n9736 );
not U_inv1817 ( n75189, P1_P1_EBX_REG_29_ );
dff P1_P1_EBX_REG_30__reg ( clk, reset, P1_P1_EBX_REG_30_, n9741 );
not U_inv1818 ( n75217, P1_P1_EBX_REG_30_ );
dff P1_P1_EBX_REG_31__reg ( clk, reset, P1_P1_EBX_REG_31_, n9746 );
not U_inv1819 ( n74985, P1_P1_EBX_REG_31_ );
dff P1_P1_REIP_REG_0__reg ( clk, reset, P1_P1_REIP_REG_0_, n9751 );
not U_inv1820 ( n75262, P1_P1_REIP_REG_0_ );
dff P1_P1_BYTEENABLE_REG_0__reg ( clk, reset, P1_P1_BYTEENABLE_REG_0_, n9926 );
dff P1_P1_BE_N_REG_0__reg ( clk, reset, P1_P1_BE_N_REG_0_, n7756 );
dff P1_P1_PHYADDRPOINTER_REG_0__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_0_, n8956 );
not U_inv1821 ( n75226, P1_P1_PHYADDRPOINTER_REG_0_ );
dff P1_P1_BYTEENABLE_REG_1__reg ( clk, reset, P1_P1_BYTEENABLE_REG_1_, n9921 );
dff P1_P1_BE_N_REG_1__reg ( clk, reset, P1_P1_BE_N_REG_1_, n7751 );
dff P1_P1_BYTEENABLE_REG_3__reg ( clk, reset, P1_P1_BYTEENABLE_REG_3_, n9911 );
dff P1_P1_BE_N_REG_3__reg ( clk, reset, P1_P1_BE_N_REG_3_, n7741 );
dff P1_BUF2_REG_25__reg ( clk, reset, P1_BUF2_REG_25_, n406 );
not U_inv1822 ( n75334, P1_BUF2_REG_25_ );
dff P1_P2_INSTQUEUE_REG_5__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_5__1_, n6291 );
not U_inv1823 ( n73609, P1_P2_INSTQUEUE_REG_5__1_ );
dff P1_P2_INSTQUEUE_REG_6__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_6__1_, n6251 );
not U_inv1824 ( n73625, P1_P2_INSTQUEUE_REG_6__1_ );
dff P1_P2_INSTQUEUE_REG_7__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_7__1_, n6211 );
not U_inv1825 ( n73616, P1_P2_INSTQUEUE_REG_7__1_ );
dff P1_P2_INSTQUEUE_REG_8__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_8__1_, n6171 );
not U_inv1826 ( n73614, P1_P2_INSTQUEUE_REG_8__1_ );
dff P1_P2_INSTQUEUE_REG_9__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_9__1_, n6131 );
not U_inv1827 ( n73623, P1_P2_INSTQUEUE_REG_9__1_ );
dff P1_P2_INSTQUEUE_REG_10__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_10__1_, n6091 );
not U_inv1828 ( n73632, P1_P2_INSTQUEUE_REG_10__1_ );
dff P1_P2_INSTQUEUE_REG_11__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_11__1_, n6051 );
not U_inv1829 ( n73627, P1_P2_INSTQUEUE_REG_11__1_ );
dff P1_P2_INSTQUEUE_REG_12__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_12__1_, n6011 );
not U_inv1830 ( n73605, P1_P2_INSTQUEUE_REG_12__1_ );
dff P1_P2_INSTQUEUE_REG_13__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_13__1_, n5971 );
not U_inv1831 ( n73618, P1_P2_INSTQUEUE_REG_13__1_ );
dff P1_P2_INSTQUEUE_REG_0__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_0__1_, n6491 );
not U_inv1832 ( n73569, P1_P2_INSTQUEUE_REG_0__1_ );
dff P1_P2_EBX_REG_2__reg ( clk, reset, P1_P2_EBX_REG_2_, n7356 );
not U_inv1833 ( n74532, P1_P2_EBX_REG_2_ );
dff P1_P2_EBX_REG_3__reg ( clk, reset, P1_P2_EBX_REG_3_, n7361 );
not U_inv1834 ( n73145, P1_P2_EBX_REG_3_ );
dff P1_P2_EBX_REG_4__reg ( clk, reset, P1_P2_EBX_REG_4_, n7366 );
not U_inv1835 ( n74572, P1_P2_EBX_REG_4_ );
dff P1_P2_EBX_REG_5__reg ( clk, reset, P1_P2_EBX_REG_5_, n7371 );
not U_inv1836 ( n73153, P1_P2_EBX_REG_5_ );
dff P1_P2_EBX_REG_6__reg ( clk, reset, P1_P2_EBX_REG_6_, n7376 );
not U_inv1837 ( n74605, P1_P2_EBX_REG_6_ );
dff P1_P2_EBX_REG_7__reg ( clk, reset, P1_P2_EBX_REG_7_, n7381 );
not U_inv1838 ( n73171, P1_P2_EBX_REG_7_ );
dff P1_P2_EBX_REG_8__reg ( clk, reset, P1_P2_EBX_REG_8_, n7386 );
not U_inv1839 ( n74668, P1_P2_EBX_REG_8_ );
dff P1_P2_INSTQUEUE_REG_1__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_1__1_, n6451 );
not U_inv1840 ( n73601, P1_P2_INSTQUEUE_REG_1__1_ );
dff P1_P2_INSTQUEUE_REG_2__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_2__1_, n6411 );
not U_inv1841 ( n73620, P1_P2_INSTQUEUE_REG_2__1_ );
dff P1_P2_INSTQUEUE_REG_3__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_3__1_, n6371 );
not U_inv1842 ( n73607, P1_P2_INSTQUEUE_REG_3__1_ );
dff P1_P2_INSTQUEUE_REG_4__1__reg ( clk, reset, P1_P2_INSTQUEUE_REG_4__1_, n6331 );
not U_inv1843 ( n73598, P1_P2_INSTQUEUE_REG_4__1_ );
dff P1_P2_EBX_REG_9__reg ( clk, reset, P1_P2_EBX_REG_9_, n7391 );
not U_inv1844 ( n73202, P1_P2_EBX_REG_9_ );
dff P1_P2_EBX_REG_10__reg ( clk, reset, P1_P2_EBX_REG_10_, n7396 );
not U_inv1845 ( n74723, P1_P2_EBX_REG_10_ );
dff P1_P2_EBX_REG_11__reg ( clk, reset, P1_P2_EBX_REG_11_, n7401 );
not U_inv1846 ( n73210, P1_P2_EBX_REG_11_ );
dff P1_P2_EBX_REG_12__reg ( clk, reset, P1_P2_EBX_REG_12_, n7406 );
not U_inv1847 ( n74766, P1_P2_EBX_REG_12_ );
dff P1_P2_EBX_REG_13__reg ( clk, reset, P1_P2_EBX_REG_13_, n7411 );
not U_inv1848 ( n73229, P1_P2_EBX_REG_13_ );
dff P1_P2_EBX_REG_14__reg ( clk, reset, P1_P2_EBX_REG_14_, n7416 );
not U_inv1849 ( n74796, P1_P2_EBX_REG_14_ );
dff P1_P2_EBX_REG_15__reg ( clk, reset, P1_P2_EBX_REG_15_, n7421 );
not U_inv1850 ( n73244, P1_P2_EBX_REG_15_ );
dff P1_P2_EBX_REG_16__reg ( clk, reset, P1_P2_EBX_REG_16_, n7426 );
not U_inv1851 ( n74835, P1_P2_EBX_REG_16_ );
dff P1_P2_EBX_REG_17__reg ( clk, reset, P1_P2_EBX_REG_17_, n7431 );
not U_inv1852 ( n73258, P1_P2_EBX_REG_17_ );
dff P1_P2_EBX_REG_18__reg ( clk, reset, P1_P2_EBX_REG_18_, n7436 );
not U_inv1853 ( n74896, P1_P2_EBX_REG_18_ );
dff P1_P2_EBX_REG_19__reg ( clk, reset, P1_P2_EBX_REG_19_, n7441 );
not U_inv1854 ( n73272, P1_P2_EBX_REG_19_ );
dff P1_P2_EBX_REG_20__reg ( clk, reset, P1_P2_EBX_REG_20_, n7446 );
not U_inv1855 ( n74936, P1_P2_EBX_REG_20_ );
dff P1_P2_EBX_REG_21__reg ( clk, reset, P1_P2_EBX_REG_21_, n7451 );
not U_inv1856 ( n73285, P1_P2_EBX_REG_21_ );
dff P1_P2_EBX_REG_22__reg ( clk, reset, P1_P2_EBX_REG_22_, n7456 );
not U_inv1857 ( n74982, P1_P2_EBX_REG_22_ );
dff P1_P2_EBX_REG_23__reg ( clk, reset, P1_P2_EBX_REG_23_, n7461 );
not U_inv1858 ( n73301, P1_P2_EBX_REG_23_ );
dff P1_P2_EBX_REG_24__reg ( clk, reset, P1_P2_EBX_REG_24_, n7466 );
not U_inv1859 ( n75024, P1_P2_EBX_REG_24_ );
dff P1_P2_EBX_REG_25__reg ( clk, reset, P1_P2_EBX_REG_25_, n7471 );
not U_inv1860 ( n73313, P1_P2_EBX_REG_25_ );
dff P1_P2_EBX_REG_26__reg ( clk, reset, P1_P2_EBX_REG_26_, n7476 );
not U_inv1861 ( n75074, P1_P2_EBX_REG_26_ );
dff P1_P2_EBX_REG_27__reg ( clk, reset, P1_P2_EBX_REG_27_, n7481 );
not U_inv1862 ( n75173, P1_P2_EBX_REG_27_ );
dff P1_P2_EBX_REG_28__reg ( clk, reset, P1_P2_EBX_REG_28_, n7486 );
not U_inv1863 ( n73386, P1_P2_EBX_REG_28_ );
dff P1_P2_EBX_REG_29__reg ( clk, reset, P1_P2_EBX_REG_29_, n7491 );
not U_inv1864 ( n75183, P1_P2_EBX_REG_29_ );
dff P1_P2_EBX_REG_30__reg ( clk, reset, P1_P2_EBX_REG_30_, n7496 );
not U_inv1865 ( n75215, P1_P2_EBX_REG_30_ );
dff P1_P2_EBX_REG_31__reg ( clk, reset, P1_P2_EBX_REG_31_, n7501 );
dff P1_P3_INSTQUEUE_REG_7__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_7__1_, n3966 );
not U_inv1866 ( n73957, P1_P3_INSTQUEUE_REG_7__1_ );
dff P1_P3_INSTQUEUE_REG_0__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_0__1_, n4246 );
not U_inv1867 ( n73949, P1_P3_INSTQUEUE_REG_0__1_ );
dff P1_P3_EBX_REG_2__reg ( clk, reset, P1_P3_EBX_REG_2_, n5111 );
not U_inv1868 ( n74531, P1_P3_EBX_REG_2_ );
dff P1_P3_EBX_REG_3__reg ( clk, reset, P1_P3_EBX_REG_3_, n5116 );
not U_inv1869 ( n73144, P1_P3_EBX_REG_3_ );
dff P1_P3_EBX_REG_4__reg ( clk, reset, P1_P3_EBX_REG_4_, n5121 );
not U_inv1870 ( n74568, P1_P3_EBX_REG_4_ );
dff P1_P3_EBX_REG_5__reg ( clk, reset, P1_P3_EBX_REG_5_, n5126 );
not U_inv1871 ( n73152, P1_P3_EBX_REG_5_ );
dff P1_P3_EBX_REG_6__reg ( clk, reset, P1_P3_EBX_REG_6_, n5131 );
not U_inv1872 ( n74601, P1_P3_EBX_REG_6_ );
dff P1_P3_EBX_REG_7__reg ( clk, reset, P1_P3_EBX_REG_7_, n5136 );
not U_inv1873 ( n73170, P1_P3_EBX_REG_7_ );
dff P1_P3_EBX_REG_8__reg ( clk, reset, P1_P3_EBX_REG_8_, n5141 );
not U_inv1874 ( n74664, P1_P3_EBX_REG_8_ );
dff P1_P3_INSTQUEUE_REG_1__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_1__1_, n4206 );
not U_inv1875 ( n73952, P1_P3_INSTQUEUE_REG_1__1_ );
dff P1_P3_INSTQUEUE_REG_2__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_2__1_, n4166 );
not U_inv1876 ( n73959, P1_P3_INSTQUEUE_REG_2__1_ );
dff P1_P3_INSTQUEUE_REG_3__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_3__1_, n4126 );
not U_inv1877 ( n73954, P1_P3_INSTQUEUE_REG_3__1_ );
dff P1_P3_INSTQUEUE_REG_4__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_4__1_, n4086 );
not U_inv1878 ( n73951, P1_P3_INSTQUEUE_REG_4__1_ );
dff P1_P3_INSTQUEUE_REG_5__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_5__1_, n4046 );
not U_inv1879 ( n73955, P1_P3_INSTQUEUE_REG_5__1_ );
dff P1_P3_INSTQUEUE_REG_6__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_6__1_, n4006 );
not U_inv1880 ( n73961, P1_P3_INSTQUEUE_REG_6__1_ );
dff P1_P3_INSTQUEUE_REG_8__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_8__1_, n3926 );
not U_inv1881 ( n73956, P1_P3_INSTQUEUE_REG_8__1_ );
dff P1_P3_INSTQUEUE_REG_9__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_9__1_, n3886 );
not U_inv1882 ( n73960, P1_P3_INSTQUEUE_REG_9__1_ );
dff P1_P3_INSTQUEUE_REG_10__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_10__1_, n3846 );
not U_inv1883 ( n73965, P1_P3_INSTQUEUE_REG_10__1_ );
dff P1_P3_INSTQUEUE_REG_11__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_11__1_, n3806 );
not U_inv1884 ( n73962, P1_P3_INSTQUEUE_REG_11__1_ );
dff P1_P3_INSTQUEUE_REG_12__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_12__1_, n3766 );
not U_inv1885 ( n73953, P1_P3_INSTQUEUE_REG_12__1_ );
dff P1_P3_INSTQUEUE_REG_13__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_13__1_, n3726 );
not U_inv1886 ( n73958, P1_P3_INSTQUEUE_REG_13__1_ );
dff P1_P3_INSTQUEUE_REG_14__1__reg ( clk, reset, P1_P3_INSTQUEUE_REG_14__1_, n3686 );
not U_inv1887 ( n73963, P1_P3_INSTQUEUE_REG_14__1_ );
dff P1_P3_EAX_REG_24__reg ( clk, reset, P1_P3_EAX_REG_24_, n5061 );
dff P1_P3_EAX_REG_25__reg ( clk, reset, P1_P3_EAX_REG_25_, n5066 );
not U_inv1888 ( n75041, P1_P3_EAX_REG_25_ );
dff P1_P3_EAX_REG_26__reg ( clk, reset, P1_P3_EAX_REG_26_, n5071 );
dff P1_P3_EAX_REG_27__reg ( clk, reset, P1_P3_EAX_REG_27_, n5076 );
dff P1_P3_EAX_REG_28__reg ( clk, reset, P1_P3_EAX_REG_28_, n5081 );
not U_inv1889 ( n73395, P1_P3_EAX_REG_28_ );
dff P1_P3_EAX_REG_29__reg ( clk, reset, P1_P3_EAX_REG_29_, n5086 );
not U_inv1890 ( n75206, P1_P3_EAX_REG_29_ );
dff P1_P3_EAX_REG_30__reg ( clk, reset, P1_P3_EAX_REG_30_, n5091 );
not U_inv1891 ( n75447, P1_P3_EAX_REG_30_ );
dff P1_P3_UWORD_REG_14__reg ( clk, reset, P1_P3_UWORD_REG_14_, n4706 );
not U_inv1892 ( n75601, P1_P3_UWORD_REG_14_ );
dff P1_P3_DATAO_REG_30__reg ( clk, reset, P1_P3_DATAO_REG_30_, n4931 );
dff P1_P3_EBX_REG_9__reg ( clk, reset, P1_P3_EBX_REG_9_, n5146 );
not U_inv1893 ( n73200, P1_P3_EBX_REG_9_ );
dff P1_P2_DATAO_REG_0__reg ( clk, reset, P1_P2_DATAO_REG_0_, n7026 );
not U_inv1894 ( n75550, P1_P2_DATAO_REG_0_ );
dff P1_P2_CODEFETCH_REG_reg ( clk, reset, P1_P2_CODEFETCH_REG, n7721 );
dff P1_P2_D_C_N_REG_reg ( clk, reset, P1_P2_D_C_N_REG, n7711 );
dff P1_P2_MORE_REG_reg ( clk, reset, P1_P2_MORE_REG, n7696 );
dff P1_P1_LWORD_REG_15__reg ( clk, reset, P1_P1_LWORD_REG_15_, n9116 );
not U_inv1895 ( n75668, P1_P1_LWORD_REG_15_ );
dff P1_P1_DATAO_REG_15__reg ( clk, reset, P1_P1_DATAO_REG_15_, n9346 );
dff P1_BUF2_REG_15__reg ( clk, reset, P1_BUF2_REG_15_, n356 );
not U_inv1896 ( n75363, P1_BUF2_REG_15_ );
dff P1_P3_EAX_REG_15__reg ( clk, reset, P1_P3_EAX_REG_15_, n5016 );
not U_inv1897 ( n74778, P1_P3_EAX_REG_15_ );
dff P1_P3_EAX_REG_16__reg ( clk, reset, P1_P3_EAX_REG_16_, n5021 );
not U_inv1898 ( n75421, P1_P3_EAX_REG_16_ );
dff P1_P3_UWORD_REG_0__reg ( clk, reset, P1_P3_UWORD_REG_0_, n4776 );
not U_inv1899 ( n75602, P1_P3_UWORD_REG_0_ );
dff P1_P3_DATAO_REG_16__reg ( clk, reset, P1_P3_DATAO_REG_16_, n4861 );
dff P3_IR_REG_16__reg ( clk, reset, P3_IR_REG_16_, n881 );
dff P3_REG3_REG_16__reg ( clk, reset, P3_REG3_REG_16_, n1941 );
not U_inv1900 ( n72946, P3_REG3_REG_16_ );
dff P1_P3_EAX_REG_17__reg ( clk, reset, P1_P3_EAX_REG_17_, n5026 );
not U_inv1901 ( n74817, P1_P3_EAX_REG_17_ );
dff P1_P3_UWORD_REG_1__reg ( clk, reset, P1_P3_UWORD_REG_1_, n4771 );
not U_inv1902 ( n75599, P1_P3_UWORD_REG_1_ );
dff P1_P3_DATAO_REG_17__reg ( clk, reset, P1_P3_DATAO_REG_17_, n4866 );
dff P3_IR_REG_17__reg ( clk, reset, P3_IR_REG_17_, n886 );
not U_inv1903 ( n74418, P3_IR_REG_17_ );
dff P3_IR_REG_18__reg ( clk, reset, P3_IR_REG_18_, n891 );
dff P3_REG3_REG_17__reg ( clk, reset, P3_REG3_REG_17_, n1931 );
not U_inv1904 ( n72954, P3_REG3_REG_17_ );
dff P3_REG3_REG_18__reg ( clk, reset, P3_REG3_REG_18_, n1881 );
not U_inv1905 ( n72955, P3_REG3_REG_18_ );
dff P4_D_REG_22__reg ( clk, reset, ex_wire240, n2296 );
not U_inv1906 ( n74741, ex_wire240 );
dff P4_D_REG_7__reg ( clk, reset, ex_wire241, n2221 );
not U_inv1907 ( n74742, ex_wire241 );
dff P4_D_REG_31__reg ( clk, reset, P4_D_REG_31_, n2341 );
dff P4_D_REG_30__reg ( clk, reset, P4_D_REG_30_, n2336 );
dff P4_D_REG_29__reg ( clk, reset, P4_D_REG_29_, n2331 );
dff P4_D_REG_28__reg ( clk, reset, P4_D_REG_28_, n2326 );
dff P4_D_REG_27__reg ( clk, reset, P4_D_REG_27_, n2321 );
dff P4_D_REG_26__reg ( clk, reset, P4_D_REG_26_, n2316 );
dff P4_D_REG_25__reg ( clk, reset, P4_D_REG_25_, n2311 );
dff P4_D_REG_24__reg ( clk, reset, P4_D_REG_24_, n2306 );
dff P4_D_REG_23__reg ( clk, reset, P4_D_REG_23_, n2301 );
dff P4_D_REG_21__reg ( clk, reset, P4_D_REG_21_, n2291 );
dff P4_D_REG_20__reg ( clk, reset, P4_D_REG_20_, n2286 );
dff P4_D_REG_19__reg ( clk, reset, P4_D_REG_19_, n2281 );
dff P4_D_REG_18__reg ( clk, reset, P4_D_REG_18_, n2276 );
dff P4_D_REG_17__reg ( clk, reset, P4_D_REG_17_, n2271 );
dff P4_D_REG_16__reg ( clk, reset, P4_D_REG_16_, n2266 );
dff P4_D_REG_15__reg ( clk, reset, P4_D_REG_15_, n2261 );
dff P4_D_REG_14__reg ( clk, reset, P4_D_REG_14_, n2256 );
dff P4_D_REG_13__reg ( clk, reset, P4_D_REG_13_, n2251 );
dff P4_D_REG_12__reg ( clk, reset, P4_D_REG_12_, n2246 );
dff P4_D_REG_11__reg ( clk, reset, P4_D_REG_11_, n2241 );
dff P4_D_REG_10__reg ( clk, reset, P4_D_REG_10_, n2236 );
dff P4_D_REG_9__reg ( clk, reset, P4_D_REG_9_, n2231 );
dff P4_D_REG_8__reg ( clk, reset, P4_D_REG_8_, n2226 );
dff P4_D_REG_6__reg ( clk, reset, P4_D_REG_6_, n2216 );
dff P4_D_REG_5__reg ( clk, reset, P4_D_REG_5_, n2211 );
dff P4_D_REG_4__reg ( clk, reset, P4_D_REG_4_, n2206 );
dff P4_D_REG_3__reg ( clk, reset, P4_D_REG_3_, n2201 );
dff P4_D_REG_2__reg ( clk, reset, P4_D_REG_2_, n2196 );
dff P4_D_REG_1__reg ( clk, reset, P4_D_REG_1_, n2191 );
dff P4_D_REG_0__reg ( clk, reset, P4_D_REG_0_, n2186 );
dff P4_REG1_REG_30__reg ( clk, reset, P4_REG1_REG_30_, n2656 );
not U_inv1908 ( n74825, P4_REG1_REG_30_ );
dff P4_REG1_REG_29__reg ( clk, reset, P4_REG1_REG_29_, n2651 );
not U_inv1909 ( n74784, P4_REG1_REG_29_ );
dff P4_REG1_REG_26__reg ( clk, reset, P4_REG1_REG_26_, n2636 );
not U_inv1910 ( n74716, P4_REG1_REG_26_ );
dff P4_REG1_REG_24__reg ( clk, reset, P4_REG1_REG_24_, n2626 );
not U_inv1911 ( n74707, P4_REG1_REG_24_ );
dff P4_REG1_REG_20__reg ( clk, reset, P4_REG1_REG_20_, n2606 );
not U_inv1912 ( n74519, P4_REG1_REG_20_ );
dff P4_REG1_REG_19__reg ( clk, reset, P4_REG1_REG_19_, n2601 );
not U_inv1913 ( n74511, P4_REG1_REG_19_ );
dff P4_REG1_REG_18__reg ( clk, reset, P4_REG1_REG_18_, n2596 );
not U_inv1914 ( n74483, P4_REG1_REG_18_ );
dff P4_REG1_REG_17__reg ( clk, reset, P4_REG1_REG_17_, n2591 );
not U_inv1915 ( n74457, P4_REG1_REG_17_ );
dff P4_REG1_REG_16__reg ( clk, reset, P4_REG1_REG_16_, n2586 );
not U_inv1916 ( n74420, P4_REG1_REG_16_ );
dff P4_REG1_REG_13__reg ( clk, reset, P4_REG1_REG_13_, n2571 );
not U_inv1917 ( n74404, P4_REG1_REG_13_ );
dff P4_REG1_REG_12__reg ( clk, reset, P4_REG1_REG_12_, n2566 );
not U_inv1918 ( n74399, P4_REG1_REG_12_ );
dff P4_REG1_REG_11__reg ( clk, reset, P4_REG1_REG_11_, n2561 );
not U_inv1919 ( n74394, P4_REG1_REG_11_ );
dff P4_REG1_REG_10__reg ( clk, reset, P4_REG1_REG_10_, n2556 );
not U_inv1920 ( n74358, P4_REG1_REG_10_ );
dff P4_REG1_REG_7__reg ( clk, reset, P4_REG1_REG_7_, n2541 );
not U_inv1921 ( n74318, P4_REG1_REG_7_ );
dff P4_REG1_REG_6__reg ( clk, reset, P4_REG1_REG_6_, n2536 );
not U_inv1922 ( n74236, P4_REG1_REG_6_ );
dff P4_REG1_REG_5__reg ( clk, reset, P4_REG1_REG_5_, n2531 );
not U_inv1923 ( n74166, P4_REG1_REG_5_ );
dff P4_REG1_REG_3__reg ( clk, reset, P4_REG1_REG_3_, n2521 );
not U_inv1924 ( n73999, P4_REG1_REG_3_ );
dff P4_REG1_REG_1__reg ( clk, reset, P4_REG1_REG_1_, n2511 );
not U_inv1925 ( n73804, P4_REG1_REG_1_ );
dff P4_REG2_REG_31__reg ( clk, reset, ex_wire242, n2821 );
not U_inv1926 ( n74773, ex_wire242 );
dff P4_REG1_REG_31__reg ( clk, reset, P4_REG1_REG_31_, n2661 );
not U_inv1927 ( n74771, P4_REG1_REG_31_ );
dff P4_REG0_REG_31__reg ( clk, reset, P4_REG0_REG_31_, n2501 );
dff P4_DATAO_REG_31__reg ( clk, reset, P4_DATAO_REG_31_, n3081 );
not U_inv1928 ( n73430, P4_DATAO_REG_31_ );
dff P4_REG2_REG_30__reg ( clk, reset, ex_wire243, n2816 );
not U_inv1929 ( n74826, ex_wire243 );
dff P4_REG3_REG_3__reg ( clk, reset, P4_REG3_REG_3_, n3206 );
not U_inv1930 ( n75247, P4_REG3_REG_3_ );
dff P4_REG3_REG_4__reg ( clk, reset, P4_REG3_REG_4_, n3146 );
not U_inv1931 ( n74062, P4_REG3_REG_4_ );
dff P4_REG3_REG_5__reg ( clk, reset, P4_REG3_REG_5_, n3161 );
not U_inv1932 ( n74123, P4_REG3_REG_5_ );
dff P4_REG3_REG_1__reg ( clk, reset, P4_REG3_REG_1_, n3186 );
not U_inv1933 ( n73801, P4_REG3_REG_1_ );
dff P4_REG3_REG_2__reg ( clk, reset, P4_REG3_REG_2_, n3111 );
not U_inv1934 ( n73895, P4_REG3_REG_2_ );
dff P4_REG3_REG_6__reg ( clk, reset, P4_REG3_REG_6_, n3101 );
not U_inv1935 ( n74198, P4_REG3_REG_6_ );
dff P4_REG3_REG_7__reg ( clk, reset, P4_REG3_REG_7_, n3231 );
not U_inv1936 ( n72930, P4_REG3_REG_7_ );
dff P4_REG3_REG_8__reg ( clk, reset, P4_REG3_REG_8_, n3191 );
not U_inv1937 ( n72934, P4_REG3_REG_8_ );
dff P2_P3_UWORD_REG_5__reg ( clk, reset, P2_P3_UWORD_REG_5_, n11486 );
not U_inv1938 ( n75465, P2_P3_UWORD_REG_5_ );
dff P2_P3_DATAO_REG_21__reg ( clk, reset, P2_P3_DATAO_REG_21_, n11621 );
dff P2_P3_UWORD_REG_3__reg ( clk, reset, P2_P3_UWORD_REG_3_, n11496 );
not U_inv1939 ( n75464, P2_P3_UWORD_REG_3_ );
dff P2_P3_DATAO_REG_19__reg ( clk, reset, P2_P3_DATAO_REG_19_, n11611 );
dff P2_P3_EBX_REG_10__reg ( clk, reset, P2_P3_EBX_REG_10_, n11886 );
not U_inv1940 ( n74720, P2_P3_EBX_REG_10_ );
dff P2_P3_EBX_REG_11__reg ( clk, reset, P2_P3_EBX_REG_11_, n11891 );
not U_inv1941 ( n73209, P2_P3_EBX_REG_11_ );
dff P2_P3_EBX_REG_12__reg ( clk, reset, P2_P3_EBX_REG_12_, n11896 );
not U_inv1942 ( n74763, P2_P3_EBX_REG_12_ );
dff P2_P3_EBX_REG_13__reg ( clk, reset, P2_P3_EBX_REG_13_, n11901 );
not U_inv1943 ( n73228, P2_P3_EBX_REG_13_ );
dff P2_P3_EBX_REG_14__reg ( clk, reset, P2_P3_EBX_REG_14_, n11906 );
not U_inv1944 ( n74793, P2_P3_EBX_REG_14_ );
dff P2_P3_EBX_REG_15__reg ( clk, reset, P2_P3_EBX_REG_15_, n11911 );
not U_inv1945 ( n73243, P2_P3_EBX_REG_15_ );
dff P2_P3_EBX_REG_16__reg ( clk, reset, P2_P3_EBX_REG_16_, n11916 );
not U_inv1946 ( n74833, P2_P3_EBX_REG_16_ );
dff P2_P3_EBX_REG_17__reg ( clk, reset, P2_P3_EBX_REG_17_, n11921 );
not U_inv1947 ( n73257, P2_P3_EBX_REG_17_ );
dff P2_P3_EBX_REG_18__reg ( clk, reset, P2_P3_EBX_REG_18_, n11926 );
not U_inv1948 ( n74894, P2_P3_EBX_REG_18_ );
dff P2_P3_EBX_REG_19__reg ( clk, reset, P2_P3_EBX_REG_19_, n11931 );
not U_inv1949 ( n73271, P2_P3_EBX_REG_19_ );
dff P2_P3_EBX_REG_20__reg ( clk, reset, P2_P3_EBX_REG_20_, n11936 );
not U_inv1950 ( n74934, P2_P3_EBX_REG_20_ );
dff P2_P3_EBX_REG_21__reg ( clk, reset, P2_P3_EBX_REG_21_, n11941 );
not U_inv1951 ( n73284, P2_P3_EBX_REG_21_ );
dff P2_P3_EBX_REG_22__reg ( clk, reset, P2_P3_EBX_REG_22_, n11946 );
not U_inv1952 ( n74980, P2_P3_EBX_REG_22_ );
dff P2_P3_EBX_REG_23__reg ( clk, reset, P2_P3_EBX_REG_23_, n11951 );
not U_inv1953 ( n73300, P2_P3_EBX_REG_23_ );
dff P2_P3_EBX_REG_24__reg ( clk, reset, P2_P3_EBX_REG_24_, n11956 );
not U_inv1954 ( n75023, P2_P3_EBX_REG_24_ );
dff P2_P3_EBX_REG_25__reg ( clk, reset, P2_P3_EBX_REG_25_, n11961 );
not U_inv1955 ( n73312, P2_P3_EBX_REG_25_ );
dff P2_P3_EBX_REG_26__reg ( clk, reset, P2_P3_EBX_REG_26_, n11966 );
not U_inv1956 ( n75073, P2_P3_EBX_REG_26_ );
dff P2_P3_EBX_REG_27__reg ( clk, reset, P2_P3_EBX_REG_27_, n11971 );
not U_inv1957 ( n75172, P2_P3_EBX_REG_27_ );
dff P2_P3_EBX_REG_28__reg ( clk, reset, P2_P3_EBX_REG_28_, n11976 );
not U_inv1958 ( n73388, P2_P3_EBX_REG_28_ );
dff P2_P3_EBX_REG_29__reg ( clk, reset, P2_P3_EBX_REG_29_, n11981 );
not U_inv1959 ( n75182, P2_P3_EBX_REG_29_ );
dff P2_P3_EBX_REG_30__reg ( clk, reset, P2_P3_EBX_REG_30_, n11986 );
not U_inv1960 ( n75214, P2_P3_EBX_REG_30_ );
dff P2_P3_EBX_REG_31__reg ( clk, reset, P2_P3_EBX_REG_31_, n11991 );
dff P2_P2_INSTADDRPOINTER_REG_1__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_1_, n13291 );
not U_inv1961 ( n75057, P2_P2_INSTADDRPOINTER_REG_1_ );
dff P2_P2_PHYADDRPOINTER_REG_1__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_1_, n13451 );
not U_inv1962 ( n74472, P2_P2_PHYADDRPOINTER_REG_1_ );
dff P2_P2_REIP_REG_1__reg ( clk, reset, P2_P2_REIP_REG_1_, n14246 );
not U_inv1963 ( n72959, P2_P2_REIP_REG_1_ );
dff P2_P2_BYTEENABLE_REG_0__reg ( clk, reset, P2_P2_BYTEENABLE_REG_0_, n14416 );
dff P2_P2_BE_N_REG_0__reg ( clk, reset, P2_P2_BE_N_REG_0_, n12246 );
dff P2_P2_BYTEENABLE_REG_1__reg ( clk, reset, P2_P2_BYTEENABLE_REG_1_, n14411 );
dff P2_P2_BE_N_REG_1__reg ( clk, reset, P2_P2_BE_N_REG_1_, n12241 );
dff P2_P2_BYTEENABLE_REG_2__reg ( clk, reset, P2_P2_BYTEENABLE_REG_2_, n14406 );
dff P2_P2_BE_N_REG_2__reg ( clk, reset, P2_P2_BE_N_REG_2_, n12236 );
dff P2_P2_PHYADDRPOINTER_REG_2__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_2_, n13456 );
not U_inv1964 ( n74702, P2_P2_PHYADDRPOINTER_REG_2_ );
dff P2_P2_REIP_REG_2__reg ( clk, reset, P2_P2_REIP_REG_2_, n14251 );
not U_inv1965 ( n74619, P2_P2_REIP_REG_2_ );
dff P2_P2_ADDRESS_REG_0__reg ( clk, reset, P2_P2_ADDRESS_REG_0_, n12396 );
not U_inv1966 ( n73435, P2_P2_ADDRESS_REG_0_ );
dff P2_P2_REIP_REG_3__reg ( clk, reset, P2_P2_REIP_REG_3_, n14256 );
not U_inv1967 ( n72960, P2_P2_REIP_REG_3_ );
dff P2_P2_ADDRESS_REG_1__reg ( clk, reset, P2_P2_ADDRESS_REG_1_, n12391 );
not U_inv1968 ( n73437, P2_P2_ADDRESS_REG_1_ );
dff P2_P2_REIP_REG_4__reg ( clk, reset, P2_P2_REIP_REG_4_, n14261 );
not U_inv1969 ( n74640, P2_P2_REIP_REG_4_ );
dff P2_P2_ADDRESS_REG_2__reg ( clk, reset, P2_P2_ADDRESS_REG_2_, n12386 );
not U_inv1970 ( n73027, P2_P2_ADDRESS_REG_2_ );
dff P2_P2_ADDRESS_REG_3__reg ( clk, reset, P2_P2_ADDRESS_REG_3_, n12381 );
not U_inv1971 ( n73472, P2_P2_ADDRESS_REG_3_ );
dff P2_P2_INSTADDRPOINTER_REG_4__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_4_, n13306 );
not U_inv1972 ( n75939, P2_P2_INSTADDRPOINTER_REG_4_ );
dff P2_P2_INSTADDRPOINTER_REG_5__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_5_, n13311 );
not U_inv1973 ( n74454, P2_P2_INSTADDRPOINTER_REG_5_ );
dff P2_P2_PHYADDRPOINTER_REG_6__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_6_, n13476 );
not U_inv1974 ( n74505, P2_P2_PHYADDRPOINTER_REG_6_ );
dff P2_P2_PHYADDRPOINTER_REG_7__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_7_, n13481 );
not U_inv1975 ( n73101, P2_P2_PHYADDRPOINTER_REG_7_ );
dff P2_P2_REIP_REG_7__reg ( clk, reset, P2_P2_REIP_REG_7_, n14276 );
not U_inv1976 ( n73198, P2_P2_REIP_REG_7_ );
dff P2_P2_REIP_REG_8__reg ( clk, reset, P2_P2_REIP_REG_8_, n14281 );
not U_inv1977 ( n74747, P2_P2_REIP_REG_8_ );
dff P2_P2_REIP_REG_9__reg ( clk, reset, ex_wire244, n14286 );
not U_inv1978 ( n73214, ex_wire244 );
dff P2_P2_REIP_REG_10__reg ( clk, reset, P2_P2_REIP_REG_10_, n14291 );
not U_inv1979 ( n74743, P2_P2_REIP_REG_10_ );
dff P2_P2_ADDRESS_REG_9__reg ( clk, reset, P2_P2_ADDRESS_REG_9_, n12351 );
not U_inv1980 ( n73821, P2_P2_ADDRESS_REG_9_ );
dff P2_P2_INSTADDRPOINTER_REG_10__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_10_, n13336 );
not U_inv1981 ( n74760, P2_P2_INSTADDRPOINTER_REG_10_ );
dff P2_P2_PHYADDRPOINTER_REG_12__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_12_, n13506 );
not U_inv1982 ( n74618, P2_P2_PHYADDRPOINTER_REG_12_ );
dff P2_P2_PHYADDRPOINTER_REG_13__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_13_, n13511 );
dff P2_P2_REIP_REG_13__reg ( clk, reset, P2_P2_REIP_REG_13_, n14306 );
not U_inv1983 ( n73233, P2_P2_REIP_REG_13_ );
dff P2_P2_REIP_REG_14__reg ( clk, reset, P2_P2_REIP_REG_14_, n14311 );
not U_inv1984 ( n74827, P2_P2_REIP_REG_14_ );
dff P2_P2_INSTADDRPOINTER_REG_14__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_14_, n13356 );
not U_inv1985 ( n74433, P2_P2_INSTADDRPOINTER_REG_14_ );
dff P2_P2_INSTADDRPOINTER_REG_17__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_17_, n13371 );
not U_inv1986 ( n74874, P2_P2_INSTADDRPOINTER_REG_17_ );
dff P2_P2_INSTADDRPOINTER_REG_18__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_18_, n13376 );
not U_inv1987 ( n74548, P2_P2_INSTADDRPOINTER_REG_18_ );
dff P2_P2_INSTADDRPOINTER_REG_23__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_23_, n13401 );
not U_inv1988 ( n74639, P2_P2_INSTADDRPOINTER_REG_23_ );
dff P2_P2_PHYADDRPOINTER_REG_14__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_14_, n13516 );
not U_inv1989 ( n74858, P2_P2_PHYADDRPOINTER_REG_14_ );
dff P2_P2_PHYADDRPOINTER_REG_17__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_17_, n13531 );
not U_inv1990 ( n74566, P2_P2_PHYADDRPOINTER_REG_17_ );
dff P2_P2_PHYADDRPOINTER_REG_18__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_18_, n13536 );
not U_inv1991 ( n75194, P2_P2_PHYADDRPOINTER_REG_18_ );
dff P2_P2_PHYADDRPOINTER_REG_19__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_19_, n13541 );
dff P2_P2_REIP_REG_20__reg ( clk, reset, P2_P2_REIP_REG_20_, n14341 );
not U_inv1992 ( n74925, P2_P2_REIP_REG_20_ );
dff P2_P2_PHYADDRPOINTER_REG_20__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_20_, n13546 );
not U_inv1993 ( n74943, P2_P2_PHYADDRPOINTER_REG_20_ );
dff P2_P2_REIP_REG_21__reg ( clk, reset, P2_P2_REIP_REG_21_, n14346 );
not U_inv1994 ( n74938, P2_P2_REIP_REG_21_ );
dff P2_P2_PHYADDRPOINTER_REG_21__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_21_, n13551 );
not U_inv1995 ( n74690, P2_P2_PHYADDRPOINTER_REG_21_ );
dff P2_P2_PHYADDRPOINTER_REG_23__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_23_, n13561 );
not U_inv1996 ( n74754, P2_P2_PHYADDRPOINTER_REG_23_ );
dff P2_P2_PHYADDRPOINTER_REG_24__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_24_, n13566 );
not U_inv1997 ( n75212, P2_P2_PHYADDRPOINTER_REG_24_ );
dff P2_P2_PHYADDRPOINTER_REG_25__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_25_, n13571 );
not U_inv1998 ( n74807, P2_P2_PHYADDRPOINTER_REG_25_ );
dff P2_P2_REIP_REG_26__reg ( clk, reset, P2_P2_REIP_REG_26_, n14371 );
not U_inv1999 ( n73295, P2_P2_REIP_REG_26_ );
dff P2_P2_INSTADDRPOINTER_REG_26__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_26_, n13416 );
not U_inv2000 ( n74950, P2_P2_INSTADDRPOINTER_REG_26_ );
dff P2_P2_INSTADDRPOINTER_REG_29__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_29_, n13431 );
not U_inv2001 ( n75008, P2_P2_INSTADDRPOINTER_REG_29_ );
dff P2_P2_PHYADDRPOINTER_REG_26__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_26_, n13576 );
not U_inv2002 ( n75046, P2_P2_PHYADDRPOINTER_REG_26_ );
dff P2_P2_PHYADDRPOINTER_REG_29__reg ( clk, reset, P2_P2_PHYADDRPOINTER_REG_29_, n13591 );
not U_inv2003 ( n74911, P2_P2_PHYADDRPOINTER_REG_29_ );
dff P2_P2_REIP_REG_31__reg ( clk, reset, P2_P2_REIP_REG_31_, n14396 );
not U_inv2004 ( n75177, P2_P2_REIP_REG_31_ );
dff P2_P2_REIP_REG_27__reg ( clk, reset, P2_P2_REIP_REG_27_, n14376 );
not U_inv2005 ( n75000, P2_P2_REIP_REG_27_ );
dff P2_P2_ADDRESS_REG_25__reg ( clk, reset, P2_P2_ADDRESS_REG_25_, n12271 );
dff P2_P2_ADDRESS_REG_26__reg ( clk, reset, P2_P2_ADDRESS_REG_26_, n12266 );
dff P2_P2_ADDRESS_REG_19__reg ( clk, reset, P2_P2_ADDRESS_REG_19_, n12301 );
dff P2_P2_ADDRESS_REG_13__reg ( clk, reset, P2_P2_ADDRESS_REG_13_, n12331 );
not U_inv2006 ( n74385, P2_P2_ADDRESS_REG_13_ );
dff P2_P2_ADDRESS_REG_12__reg ( clk, reset, P2_P2_ADDRESS_REG_12_, n12336 );
not U_inv2007 ( n73069, P2_P2_ADDRESS_REG_12_ );
dff P2_P2_ADDRESS_REG_7__reg ( clk, reset, P2_P2_ADDRESS_REG_7_, n12361 );
not U_inv2008 ( n73528, P2_P2_ADDRESS_REG_7_ );
dff P2_P2_ADDRESS_REG_8__reg ( clk, reset, P2_P2_ADDRESS_REG_8_, n12356 );
not U_inv2009 ( n73061, P2_P2_ADDRESS_REG_8_ );
dff P2_P2_ADDRESS_REG_6__reg ( clk, reset, P2_P2_ADDRESS_REG_6_, n12366 );
not U_inv2010 ( n73056, P2_P2_ADDRESS_REG_6_ );
dff P3_REG2_REG_7__reg ( clk, reset, P3_REG2_REG_7_, n1476 );
not U_inv2011 ( n74336, P3_REG2_REG_7_ );
dff P3_REG1_REG_11__reg ( clk, reset, P3_REG1_REG_11_, n1336 );
not U_inv2012 ( n74379, P3_REG1_REG_11_ );
dff P3_REG0_REG_11__reg ( clk, reset, P3_REG0_REG_11_, n1176 );
dff P3_REG2_REG_6__reg ( clk, reset, P3_REG2_REG_6_, n1471 );
not U_inv2013 ( n74281, P3_REG2_REG_6_ );
dff P3_REG2_REG_1__reg ( clk, reset, P3_REG2_REG_1_, n1446 );
not U_inv2014 ( n73827, P3_REG2_REG_1_ );
dff P3_REG2_REG_0__reg ( clk, reset, P3_REG2_REG_0_, n1441 );
not U_inv2015 ( n73633, P3_REG2_REG_0_ );
dff P3_ADDR_REG_0__reg ( clk, reset, P3_ADDR_REG_0_, n1696 );
dff P3_ADDR_REG_1__reg ( clk, reset, P3_ADDR_REG_1_, n1691 );
dff P3_ADDR_REG_3__reg ( clk, reset, ex_wire245, n1681 );
not U_inv2016 ( n73475, ex_wire245 );
dff P3_ADDR_REG_5__reg ( clk, reset, ex_wire246, n1671 );
not U_inv2017 ( n73501, ex_wire246 );
dff P3_ADDR_REG_6__reg ( clk, reset, ex_wire247, n1666 );
not U_inv2018 ( n73523, ex_wire247 );
dff P3_ADDR_REG_7__reg ( clk, reset, ex_wire248, n1661 );
not U_inv2019 ( n73531, ex_wire248 );
dff P3_ADDR_REG_8__reg ( clk, reset, ex_wire249, n1656 );
not U_inv2020 ( n73551, ex_wire249 );
dff P3_ADDR_REG_2__reg ( clk, reset, P3_ADDR_REG_2_, n1686 );
dff P3_ADDR_REG_4__reg ( clk, reset, P3_ADDR_REG_4_, n1676 );
dff P3_REG3_REG_19__reg ( clk, reset, P3_REG3_REG_19_, n1976 );
not U_inv2021 ( n74462, P3_REG3_REG_19_ );
dff P3_REG3_REG_20__reg ( clk, reset, P3_REG3_REG_20_, n1906 );
dff P3_REG3_REG_21__reg ( clk, reset, P3_REG3_REG_21_, n1956 );
not U_inv2022 ( n74492, P3_REG3_REG_21_ );
dff P3_REG3_REG_22__reg ( clk, reset, P3_REG3_REG_22_, n1896 );
dff P3_REG3_REG_23__reg ( clk, reset, P3_REG3_REG_23_, n1991 );
not U_inv2023 ( n74567, P3_REG3_REG_23_ );
dff P3_REG3_REG_24__reg ( clk, reset, P3_REG3_REG_24_, n1926 );
dff P3_REG3_REG_25__reg ( clk, reset, P3_REG3_REG_25_, n1946 );
not U_inv2024 ( n74674, P3_REG3_REG_25_ );
dff P3_REG3_REG_26__reg ( clk, reset, P3_REG3_REG_26_, n1871 );
dff P3_REG3_REG_27__reg ( clk, reset, P3_REG3_REG_27_, n2001 );
not U_inv2025 ( n74736, P3_REG3_REG_27_ );
dff P3_REG3_REG_28__reg ( clk, reset, P3_REG3_REG_28_, n1971 );
dff P1_P3_EBX_REG_10__reg ( clk, reset, P1_P3_EBX_REG_10_, n5151 );
not U_inv2026 ( n74719, P1_P3_EBX_REG_10_ );
dff P1_P3_EBX_REG_11__reg ( clk, reset, P1_P3_EBX_REG_11_, n5156 );
not U_inv2027 ( n73208, P1_P3_EBX_REG_11_ );
dff P1_P3_EBX_REG_12__reg ( clk, reset, P1_P3_EBX_REG_12_, n5161 );
not U_inv2028 ( n74762, P1_P3_EBX_REG_12_ );
dff P1_P3_EBX_REG_13__reg ( clk, reset, P1_P3_EBX_REG_13_, n5166 );
not U_inv2029 ( n73227, P1_P3_EBX_REG_13_ );
dff P1_P3_EBX_REG_14__reg ( clk, reset, P1_P3_EBX_REG_14_, n5171 );
not U_inv2030 ( n74792, P1_P3_EBX_REG_14_ );
dff P1_P3_EBX_REG_15__reg ( clk, reset, P1_P3_EBX_REG_15_, n5176 );
not U_inv2031 ( n73242, P1_P3_EBX_REG_15_ );
dff P1_P3_EBX_REG_16__reg ( clk, reset, P1_P3_EBX_REG_16_, n5181 );
not U_inv2032 ( n74832, P1_P3_EBX_REG_16_ );
dff P1_P3_EBX_REG_17__reg ( clk, reset, P1_P3_EBX_REG_17_, n5186 );
not U_inv2033 ( n73256, P1_P3_EBX_REG_17_ );
dff P1_P3_EBX_REG_18__reg ( clk, reset, P1_P3_EBX_REG_18_, n5191 );
not U_inv2034 ( n74893, P1_P3_EBX_REG_18_ );
dff P1_P3_EBX_REG_19__reg ( clk, reset, P1_P3_EBX_REG_19_, n5196 );
not U_inv2035 ( n73270, P1_P3_EBX_REG_19_ );
dff P1_P3_EBX_REG_20__reg ( clk, reset, P1_P3_EBX_REG_20_, n5201 );
not U_inv2036 ( n74933, P1_P3_EBX_REG_20_ );
dff P1_P3_EBX_REG_21__reg ( clk, reset, P1_P3_EBX_REG_21_, n5206 );
not U_inv2037 ( n73283, P1_P3_EBX_REG_21_ );
dff P1_P3_EBX_REG_22__reg ( clk, reset, P1_P3_EBX_REG_22_, n5211 );
not U_inv2038 ( n74979, P1_P3_EBX_REG_22_ );
dff P1_P3_EBX_REG_23__reg ( clk, reset, P1_P3_EBX_REG_23_, n5216 );
not U_inv2039 ( n73299, P1_P3_EBX_REG_23_ );
dff P1_P3_EBX_REG_24__reg ( clk, reset, P1_P3_EBX_REG_24_, n5221 );
not U_inv2040 ( n75022, P1_P3_EBX_REG_24_ );
dff P1_P3_EBX_REG_25__reg ( clk, reset, P1_P3_EBX_REG_25_, n5226 );
not U_inv2041 ( n73311, P1_P3_EBX_REG_25_ );
dff P1_P3_EBX_REG_26__reg ( clk, reset, P1_P3_EBX_REG_26_, n5231 );
not U_inv2042 ( n75072, P1_P3_EBX_REG_26_ );
dff P1_P3_EBX_REG_27__reg ( clk, reset, P1_P3_EBX_REG_27_, n5236 );
not U_inv2043 ( n75171, P1_P3_EBX_REG_27_ );
dff P1_P3_EBX_REG_28__reg ( clk, reset, P1_P3_EBX_REG_28_, n5241 );
not U_inv2044 ( n73387, P1_P3_EBX_REG_28_ );
dff P1_P3_EBX_REG_29__reg ( clk, reset, P1_P3_EBX_REG_29_, n5246 );
not U_inv2045 ( n75181, P1_P3_EBX_REG_29_ );
dff P1_P3_EBX_REG_30__reg ( clk, reset, P1_P3_EBX_REG_30_, n5251 );
not U_inv2046 ( n75213, P1_P3_EBX_REG_30_ );
dff P1_P3_EBX_REG_31__reg ( clk, reset, P1_P3_EBX_REG_31_, n5256 );
dff P1_P2_PHYADDRPOINTER_REG_0__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_0_, n6711 );
not U_inv2047 ( n75222, P1_P2_PHYADDRPOINTER_REG_0_ );
dff P1_P2_REIP_REG_1__reg ( clk, reset, P1_P2_REIP_REG_1_, n7511 );
not U_inv2048 ( n72958, P1_P2_REIP_REG_1_ );
dff P1_P2_INSTADDRPOINTER_REG_1__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_1_, n6556 );
not U_inv2049 ( n75056, P1_P2_INSTADDRPOINTER_REG_1_ );
dff P1_P2_PHYADDRPOINTER_REG_1__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_1_, n6716 );
not U_inv2050 ( n74471, P1_P2_PHYADDRPOINTER_REG_1_ );
dff P1_P2_REIP_REG_2__reg ( clk, reset, P1_P2_REIP_REG_2_, n7516 );
not U_inv2051 ( n74620, P1_P2_REIP_REG_2_ );
dff P1_P2_PHYADDRPOINTER_REG_2__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_2_, n6721 );
not U_inv2052 ( n74701, P1_P2_PHYADDRPOINTER_REG_2_ );
dff P1_P2_REIP_REG_4__reg ( clk, reset, P1_P2_REIP_REG_4_, n7526 );
not U_inv2053 ( n74641, P1_P2_REIP_REG_4_ );
dff P1_P2_INSTADDRPOINTER_REG_4__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_4_, n6571 );
not U_inv2054 ( n75938, P1_P2_INSTADDRPOINTER_REG_4_ );
dff P1_P2_PHYADDRPOINTER_REG_4__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_4_, n6731 );
not U_inv2055 ( n74480, P1_P2_PHYADDRPOINTER_REG_4_ );
dff P1_P2_PHYADDRPOINTER_REG_5__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_5_, n6736 );
not U_inv2056 ( n73094, P1_P2_PHYADDRPOINTER_REG_5_ );
dff P1_P2_REIP_REG_5__reg ( clk, reset, P1_P2_REIP_REG_5_, n7531 );
not U_inv2057 ( n74694, P1_P2_REIP_REG_5_ );
dff P1_P2_REIP_REG_6__reg ( clk, reset, ex_wire250, n7536 );
not U_inv2058 ( n74710, ex_wire250 );
dff P1_P2_INSTADDRPOINTER_REG_6__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_6_, n6581 );
not U_inv2059 ( n73067, P1_P2_INSTADDRPOINTER_REG_6_ );
dff P1_P2_INSTADDRPOINTER_REG_7__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_7_, n6586 );
not U_inv2060 ( n74697, P1_P2_INSTADDRPOINTER_REG_7_ );
dff P1_P2_PHYADDRPOINTER_REG_8__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_8_, n6751 );
not U_inv2061 ( n74528, P1_P2_PHYADDRPOINTER_REG_8_ );
dff P1_P2_PHYADDRPOINTER_REG_9__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_9_, n6756 );
not U_inv2062 ( n73113, P1_P2_PHYADDRPOINTER_REG_9_ );
dff P1_P2_PHYADDRPOINTER_REG_10__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_10_, n6761 );
not U_inv2063 ( n74559, P1_P2_PHYADDRPOINTER_REG_10_ );
dff P1_P2_PHYADDRPOINTER_REG_11__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_11_, n6766 );
not U_inv2064 ( n74466, P1_P2_PHYADDRPOINTER_REG_11_ );
dff P1_P2_REIP_REG_11__reg ( clk, reset, P1_P2_REIP_REG_11_, n7561 );
not U_inv2065 ( n74789, P1_P2_REIP_REG_11_ );
dff P1_P2_REIP_REG_12__reg ( clk, reset, ex_wire251, n7566 );
not U_inv2066 ( n74799, ex_wire251 );
dff P1_P2_INSTADDRPOINTER_REG_12__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_12_, n6611 );
not U_inv2067 ( n74439, P1_P2_INSTADDRPOINTER_REG_12_ );
dff P1_P2_INSTADDRPOINTER_REG_15__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_15_, n6626 );
not U_inv2068 ( n74853, P1_P2_INSTADDRPOINTER_REG_15_ );
dff P1_P2_PHYADDRPOINTER_REG_15__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_15_, n6786 );
not U_inv2069 ( n75198, P1_P2_PHYADDRPOINTER_REG_15_ );
dff P1_P2_REIP_REG_15__reg ( clk, reset, P1_P2_REIP_REG_15_, n7581 );
not U_inv2070 ( n74838, P1_P2_REIP_REG_15_ );
dff P1_P2_REIP_REG_16__reg ( clk, reset, P1_P2_REIP_REG_16_, n7586 );
not U_inv2071 ( n73248, P1_P2_REIP_REG_16_ );
dff P1_P2_PHYADDRPOINTER_REG_16__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_16_, n6791 );
dff P1_P2_REIP_REG_17__reg ( clk, reset, P1_P2_REIP_REG_17_, n7591 );
not U_inv2072 ( n74883, P1_P2_REIP_REG_17_ );
dff P1_P2_REIP_REG_18__reg ( clk, reset, P1_P2_REIP_REG_18_, n7596 );
not U_inv2073 ( n74899, P1_P2_REIP_REG_18_ );
dff P1_P2_REIP_REG_19__reg ( clk, reset, P1_P2_REIP_REG_19_, n7601 );
not U_inv2074 ( n73262, P1_P2_REIP_REG_19_ );
dff P1_P2_INSTADDRPOINTER_REG_19__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_19_, n6646 );
not U_inv2075 ( n74575, P1_P2_INSTADDRPOINTER_REG_19_ );
dff P1_P2_INSTADDRPOINTER_REG_21__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_21_, n6656 );
not U_inv2076 ( n73150, P1_P2_INSTADDRPOINTER_REG_21_ );
dff P1_P2_INSTADDRPOINTER_REG_22__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_22_, n6661 );
not U_inv2077 ( n74596, P1_P2_INSTADDRPOINTER_REG_22_ );
dff P1_P2_PHYADDRPOINTER_REG_22__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_22_, n6821 );
not U_inv2078 ( n75241, P1_P2_PHYADDRPOINTER_REG_22_ );
dff P1_P2_REIP_REG_22__reg ( clk, reset, P1_P2_REIP_REG_22_, n7616 );
not U_inv2079 ( n73276, P1_P2_REIP_REG_22_ );
dff P1_P2_REIP_REG_23__reg ( clk, reset, P1_P2_REIP_REG_23_, n7621 );
not U_inv2080 ( n74970, P1_P2_REIP_REG_23_ );
dff P1_P2_REIP_REG_24__reg ( clk, reset, P1_P2_REIP_REG_24_, n7626 );
not U_inv2081 ( n74991, P1_P2_REIP_REG_24_ );
dff P1_P2_REIP_REG_25__reg ( clk, reset, P1_P2_REIP_REG_25_, n7631 );
not U_inv2082 ( n73291, P1_P2_REIP_REG_25_ );
dff P1_P2_INSTADDRPOINTER_REG_28__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_28_, n6691 );
not U_inv2083 ( n74975, P1_P2_INSTADDRPOINTER_REG_28_ );
dff P1_P2_PHYADDRPOINTER_REG_30__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_30_, n6861 );
not U_inv2084 ( n75186, P1_P2_PHYADDRPOINTER_REG_30_ );
dff P1_P2_PHYADDRPOINTER_REG_31__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_31_, n6866 );
dff P1_P2_REIP_REG_3__reg ( clk, reset, P1_P2_REIP_REG_3_, n7521 );
not U_inv2085 ( n72961, P1_P2_REIP_REG_3_ );
dff P1_P2_INSTADDRPOINTER_REG_3__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_3_, n6566 );
not U_inv2086 ( n74409, P1_P2_INSTADDRPOINTER_REG_3_ );
dff P1_P2_INSTADDRPOINTER_REG_5__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_5_, n6576 );
not U_inv2087 ( n74453, P1_P2_INSTADDRPOINTER_REG_5_ );
dff P1_P2_PHYADDRPOINTER_REG_3__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_3_, n6726 );
not U_inv2088 ( n73083, P1_P2_PHYADDRPOINTER_REG_3_ );
dff P1_P2_PHYADDRPOINTER_REG_6__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_6_, n6741 );
not U_inv2089 ( n74504, P1_P2_PHYADDRPOINTER_REG_6_ );
dff P1_P2_REIP_REG_7__reg ( clk, reset, P1_P2_REIP_REG_7_, n7541 );
not U_inv2090 ( n73199, P1_P2_REIP_REG_7_ );
dff P1_P2_PHYADDRPOINTER_REG_7__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_7_, n6746 );
not U_inv2091 ( n73103, P1_P2_PHYADDRPOINTER_REG_7_ );
dff P1_P2_REIP_REG_8__reg ( clk, reset, P1_P2_REIP_REG_8_, n7546 );
not U_inv2092 ( n74748, P1_P2_REIP_REG_8_ );
dff P1_P2_REIP_REG_9__reg ( clk, reset, ex_wire252, n7551 );
not U_inv2093 ( n73215, ex_wire252 );
dff P1_P2_REIP_REG_10__reg ( clk, reset, P1_P2_REIP_REG_10_, n7556 );
not U_inv2094 ( n74744, P1_P2_REIP_REG_10_ );
dff P1_P2_INSTADDRPOINTER_REG_10__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_10_, n6601 );
not U_inv2095 ( n74759, P1_P2_INSTADDRPOINTER_REG_10_ );
dff P1_P2_PHYADDRPOINTER_REG_12__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_12_, n6771 );
not U_inv2096 ( n74617, P1_P2_PHYADDRPOINTER_REG_12_ );
dff P1_P2_PHYADDRPOINTER_REG_13__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_13_, n6776 );
dff P1_P2_REIP_REG_13__reg ( clk, reset, P1_P2_REIP_REG_13_, n7571 );
not U_inv2097 ( n73234, P1_P2_REIP_REG_13_ );
dff P1_P2_REIP_REG_14__reg ( clk, reset, P1_P2_REIP_REG_14_, n7576 );
not U_inv2098 ( n74828, P1_P2_REIP_REG_14_ );
dff P1_P2_INSTADDRPOINTER_REG_14__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_14_, n6621 );
not U_inv2099 ( n74432, P1_P2_INSTADDRPOINTER_REG_14_ );
dff P1_P2_INSTADDRPOINTER_REG_17__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_17_, n6636 );
not U_inv2100 ( n74873, P1_P2_INSTADDRPOINTER_REG_17_ );
dff P1_P2_INSTADDRPOINTER_REG_18__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_18_, n6641 );
not U_inv2101 ( n74547, P1_P2_INSTADDRPOINTER_REG_18_ );
dff P1_P2_INSTADDRPOINTER_REG_23__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_23_, n6666 );
not U_inv2102 ( n74638, P1_P2_INSTADDRPOINTER_REG_23_ );
dff P1_P2_PHYADDRPOINTER_REG_14__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_14_, n6781 );
not U_inv2103 ( n74857, P1_P2_PHYADDRPOINTER_REG_14_ );
dff P1_P2_PHYADDRPOINTER_REG_17__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_17_, n6796 );
not U_inv2104 ( n74565, P1_P2_PHYADDRPOINTER_REG_17_ );
dff P1_P2_PHYADDRPOINTER_REG_18__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_18_, n6801 );
not U_inv2105 ( n75193, P1_P2_PHYADDRPOINTER_REG_18_ );
dff P1_P2_PHYADDRPOINTER_REG_19__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_19_, n6806 );
dff P1_P2_REIP_REG_20__reg ( clk, reset, P1_P2_REIP_REG_20_, n7606 );
not U_inv2106 ( n74926, P1_P2_REIP_REG_20_ );
dff P1_P2_PHYADDRPOINTER_REG_20__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_20_, n6811 );
not U_inv2107 ( n74942, P1_P2_PHYADDRPOINTER_REG_20_ );
dff P1_P2_REIP_REG_21__reg ( clk, reset, P1_P2_REIP_REG_21_, n7611 );
not U_inv2108 ( n74939, P1_P2_REIP_REG_21_ );
dff P1_P2_PHYADDRPOINTER_REG_21__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_21_, n6816 );
not U_inv2109 ( n74689, P1_P2_PHYADDRPOINTER_REG_21_ );
dff P1_P2_PHYADDRPOINTER_REG_23__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_23_, n6826 );
not U_inv2110 ( n74753, P1_P2_PHYADDRPOINTER_REG_23_ );
dff P1_P2_PHYADDRPOINTER_REG_24__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_24_, n6831 );
not U_inv2111 ( n75211, P1_P2_PHYADDRPOINTER_REG_24_ );
dff P1_P2_PHYADDRPOINTER_REG_25__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_25_, n6836 );
not U_inv2112 ( n74806, P1_P2_PHYADDRPOINTER_REG_25_ );
dff P1_P2_REIP_REG_26__reg ( clk, reset, P1_P2_REIP_REG_26_, n7636 );
not U_inv2113 ( n73294, P1_P2_REIP_REG_26_ );
dff P1_P2_INSTADDRPOINTER_REG_26__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_26_, n6681 );
not U_inv2114 ( n74949, P1_P2_INSTADDRPOINTER_REG_26_ );
dff P1_P2_INSTADDRPOINTER_REG_29__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_29_, n6696 );
not U_inv2115 ( n75007, P1_P2_INSTADDRPOINTER_REG_29_ );
dff P1_P2_PHYADDRPOINTER_REG_26__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_26_, n6841 );
not U_inv2116 ( n75043, P1_P2_PHYADDRPOINTER_REG_26_ );
dff P1_P2_PHYADDRPOINTER_REG_29__reg ( clk, reset, P1_P2_PHYADDRPOINTER_REG_29_, n6856 );
not U_inv2117 ( n74910, P1_P2_PHYADDRPOINTER_REG_29_ );
dff P1_P2_REIP_REG_31__reg ( clk, reset, P1_P2_REIP_REG_31_, n7661 );
not U_inv2118 ( n75178, P1_P2_REIP_REG_31_ );
dff P1_P2_REIP_REG_27__reg ( clk, reset, P1_P2_REIP_REG_27_, n7641 );
not U_inv2119 ( n74999, P1_P2_REIP_REG_27_ );
dff P1_P2_REIP_REG_0__reg ( clk, reset, P1_P2_REIP_REG_0_, n7506 );
not U_inv2120 ( n75260, P1_P2_REIP_REG_0_ );
dff P1_P2_BYTEENABLE_REG_0__reg ( clk, reset, P1_P2_BYTEENABLE_REG_0_, n7681 );
dff P1_P2_BE_N_REG_0__reg ( clk, reset, P1_P2_BE_N_REG_0_, n5511 );
dff P1_P2_BYTEENABLE_REG_2__reg ( clk, reset, P1_P2_BYTEENABLE_REG_2_, n7671 );
dff P1_P2_BE_N_REG_2__reg ( clk, reset, P1_P2_BE_N_REG_2_, n5501 );
dff P1_P2_BYTEENABLE_REG_1__reg ( clk, reset, P1_P2_BYTEENABLE_REG_1_, n7676 );
dff P1_P2_BE_N_REG_1__reg ( clk, reset, P1_P2_BE_N_REG_1_, n5506 );
dff P1_P2_BYTEENABLE_REG_3__reg ( clk, reset, P1_P2_BYTEENABLE_REG_3_, n7666 );
dff P4_REG1_REG_2__reg ( clk, reset, P4_REG1_REG_2_, n2516 );
not U_inv2121 ( n73896, P4_REG1_REG_2_ );
dff P4_REG0_REG_2__reg ( clk, reset, P4_REG0_REG_2_, n2356 );
dff P4_REG2_REG_1__reg ( clk, reset, P4_REG2_REG_1_, n2671 );
not U_inv2122 ( n73802, P4_REG2_REG_1_ );
dff P4_REG1_REG_4__reg ( clk, reset, P4_REG1_REG_4_, n2526 );
not U_inv2123 ( n74220, P4_REG1_REG_4_ );
dff P4_REG0_REG_4__reg ( clk, reset, P4_REG0_REG_4_, n2366 );
dff P4_REG2_REG_3__reg ( clk, reset, P4_REG2_REG_3_, n2681 );
not U_inv2124 ( n73997, P4_REG2_REG_3_ );
dff P4_REG1_REG_8__reg ( clk, reset, P4_REG1_REG_8_, n2546 );
not U_inv2125 ( n74372, P4_REG1_REG_8_ );
dff P4_REG0_REG_8__reg ( clk, reset, P4_REG0_REG_8_, n2386 );
dff P4_REG2_REG_7__reg ( clk, reset, P4_REG2_REG_7_, n2701 );
not U_inv2126 ( n74314, P4_REG2_REG_7_ );
dff P4_REG2_REG_5__reg ( clk, reset, P4_REG2_REG_5_, n2691 );
not U_inv2127 ( n74165, P4_REG2_REG_5_ );
dff P4_REG2_REG_6__reg ( clk, reset, P4_REG2_REG_6_, n2696 );
not U_inv2128 ( n74234, P4_REG2_REG_6_ );
dff P4_REG2_REG_9__reg ( clk, reset, P4_REG2_REG_9_, n2711 );
not U_inv2129 ( n74360, P4_REG2_REG_9_ );
dff P4_REG1_REG_9__reg ( clk, reset, P4_REG1_REG_9_, n2551 );
not U_inv2130 ( n74366, P4_REG1_REG_9_ );
dff P4_REG0_REG_9__reg ( clk, reset, P4_REG0_REG_9_, n2391 );
dff P4_REG3_REG_10__reg ( clk, reset, P4_REG3_REG_10_, n3211 );
not U_inv2131 ( n72933, P4_REG3_REG_10_ );
dff P4_REG2_REG_10__reg ( clk, reset, P4_REG2_REG_10_, n2716 );
not U_inv2132 ( n74356, P4_REG2_REG_10_ );
dff P4_REG3_REG_11__reg ( clk, reset, P4_REG3_REG_11_, n3116 );
not U_inv2133 ( n72938, P4_REG3_REG_11_ );
dff P4_REG3_REG_12__reg ( clk, reset, P4_REG3_REG_12_, n3176 );
not U_inv2134 ( n72940, P4_REG3_REG_12_ );
dff P4_REG3_REG_13__reg ( clk, reset, P4_REG3_REG_13_, n3126 );
not U_inv2135 ( n72941, P4_REG3_REG_13_ );
dff P4_REG2_REG_11__reg ( clk, reset, P4_REG2_REG_11_, n2721 );
not U_inv2136 ( n74393, P4_REG2_REG_11_ );
dff P4_REG3_REG_14__reg ( clk, reset, P4_REG3_REG_14_, n3221 );
not U_inv2137 ( n72945, P4_REG3_REG_14_ );
dff P4_REG3_REG_15__reg ( clk, reset, P4_REG3_REG_15_, n3091 );
not U_inv2138 ( n72944, P4_REG3_REG_15_ );
dff P4_REG3_REG_16__reg ( clk, reset, P4_REG3_REG_16_, n3166 );
not U_inv2139 ( n72947, P4_REG3_REG_16_ );
dff P4_REG3_REG_17__reg ( clk, reset, P4_REG3_REG_17_, n3156 );
not U_inv2140 ( n72953, P4_REG3_REG_17_ );
dff P4_REG3_REG_0__reg ( clk, reset, P4_REG3_REG_0_, n3136 );
not U_inv2141 ( n73800, P4_REG3_REG_0_ );
dff P4_REG2_REG_0__reg ( clk, reset, P4_REG2_REG_0_, n2666 );
not U_inv2142 ( n73799, P4_REG2_REG_0_ );
dff P4_ADDR_REG_0__reg ( clk, reset, P4_ADDR_REG_0_, n2921 );
dff P4_ADDR_REG_1__reg ( clk, reset, P4_ADDR_REG_1_, n2916 );
dff P4_ADDR_REG_2__reg ( clk, reset, P4_ADDR_REG_2_, n2911 );
dff P4_ADDR_REG_3__reg ( clk, reset, ex_wire253, n2906 );
not U_inv2143 ( n73484, ex_wire253 );
dff P4_ADDR_REG_4__reg ( clk, reset, P4_ADDR_REG_4_, n2901 );
dff P4_ADDR_REG_5__reg ( clk, reset, ex_wire254, n2896 );
not U_inv2144 ( n73470, ex_wire254 );
dff P4_ADDR_REG_6__reg ( clk, reset, ex_wire255, n2891 );
not U_inv2145 ( n73468, ex_wire255 );
dff P4_ADDR_REG_7__reg ( clk, reset, ex_wire256, n2886 );
not U_inv2146 ( n73459, ex_wire256 );
dff P4_ADDR_REG_8__reg ( clk, reset, ex_wire257, n2881 );
not U_inv2147 ( n73458, ex_wire257 );
dff P4_ADDR_REG_9__reg ( clk, reset, ex_wire258, n2876 );
not U_inv2148 ( n73464, ex_wire258 );
dff P4_ADDR_REG_10__reg ( clk, reset, ex_wire259, n2871 );
not U_inv2149 ( n73452, ex_wire259 );
dff P4_ADDR_REG_11__reg ( clk, reset, ex_wire260, n2866 );
not U_inv2150 ( n73440, ex_wire260 );
dff P4_REG3_REG_18__reg ( clk, reset, P4_REG3_REG_18_, n3106 );
not U_inv2151 ( n72956, P4_REG3_REG_18_ );
dff P4_REG3_REG_19__reg ( clk, reset, P4_REG3_REG_19_, n3201 );
not U_inv2152 ( n74459, P4_REG3_REG_19_ );
dff P4_REG3_REG_20__reg ( clk, reset, P4_REG3_REG_20_, n3131 );
dff P4_REG3_REG_21__reg ( clk, reset, P4_REG3_REG_21_, n3181 );
not U_inv2153 ( n74485, P4_REG3_REG_21_ );
dff P4_REG3_REG_22__reg ( clk, reset, P4_REG3_REG_22_, n3121 );
dff P4_REG3_REG_23__reg ( clk, reset, P4_REG3_REG_23_, n3216 );
not U_inv2154 ( n74578, P4_REG3_REG_23_ );
dff P4_REG3_REG_24__reg ( clk, reset, P4_REG3_REG_24_, n3151 );
dff P4_REG3_REG_25__reg ( clk, reset, P4_REG3_REG_25_, n3171 );
not U_inv2155 ( n74627, P4_REG3_REG_25_ );
dff P4_REG3_REG_26__reg ( clk, reset, P4_REG3_REG_26_, n3096 );
dff P4_REG3_REG_27__reg ( clk, reset, P4_REG3_REG_27_, n3226 );
not U_inv2156 ( n74708, P4_REG3_REG_27_ );
dff P4_REG3_REG_28__reg ( clk, reset, P4_REG3_REG_28_, n3196 );
dff P2_P1_EBX_REG_15__reg ( clk, reset, P2_P1_EBX_REG_15_, n16401 );
not U_inv2157 ( n73241, P2_P1_EBX_REG_15_ );
dff P2_P1_EBX_REG_16__reg ( clk, reset, P2_P1_EBX_REG_16_, n16406 );
not U_inv2158 ( n74831, P2_P1_EBX_REG_16_ );
dff P2_P1_EBX_REG_17__reg ( clk, reset, P2_P1_EBX_REG_17_, n16411 );
not U_inv2159 ( n73255, P2_P1_EBX_REG_17_ );
dff P2_P1_EBX_REG_18__reg ( clk, reset, P2_P1_EBX_REG_18_, n16416 );
not U_inv2160 ( n74892, P2_P1_EBX_REG_18_ );
dff P2_P1_EBX_REG_19__reg ( clk, reset, P2_P1_EBX_REG_19_, n16421 );
not U_inv2161 ( n73269, P2_P1_EBX_REG_19_ );
dff P2_P1_EBX_REG_20__reg ( clk, reset, P2_P1_EBX_REG_20_, n16426 );
not U_inv2162 ( n74932, P2_P1_EBX_REG_20_ );
dff P2_P1_EBX_REG_21__reg ( clk, reset, P2_P1_EBX_REG_21_, n16431 );
not U_inv2163 ( n73282, P2_P1_EBX_REG_21_ );
dff P2_P1_EBX_REG_22__reg ( clk, reset, P2_P1_EBX_REG_22_, n16436 );
not U_inv2164 ( n74978, P2_P1_EBX_REG_22_ );
dff P2_P1_EBX_REG_23__reg ( clk, reset, P2_P1_EBX_REG_23_, n16441 );
not U_inv2165 ( n73298, P2_P1_EBX_REG_23_ );
dff P2_P1_EBX_REG_24__reg ( clk, reset, P2_P1_EBX_REG_24_, n16446 );
not U_inv2166 ( n75021, P2_P1_EBX_REG_24_ );
dff P2_P1_EBX_REG_25__reg ( clk, reset, P2_P1_EBX_REG_25_, n16451 );
not U_inv2167 ( n73310, P2_P1_EBX_REG_25_ );
dff P2_P1_EBX_REG_26__reg ( clk, reset, P2_P1_EBX_REG_26_, n16456 );
not U_inv2168 ( n75071, P2_P1_EBX_REG_26_ );
dff P2_P1_EBX_REG_27__reg ( clk, reset, P2_P1_EBX_REG_27_, n16461 );
not U_inv2169 ( n75175, P2_P1_EBX_REG_27_ );
dff P2_P1_EBX_REG_28__reg ( clk, reset, P2_P1_EBX_REG_28_, n16466 );
not U_inv2170 ( n73385, P2_P1_EBX_REG_28_ );
dff P2_P1_EBX_REG_29__reg ( clk, reset, P2_P1_EBX_REG_29_, n16471 );
not U_inv2171 ( n75190, P2_P1_EBX_REG_29_ );
dff P2_P1_EBX_REG_30__reg ( clk, reset, P2_P1_EBX_REG_30_, n16476 );
not U_inv2172 ( n75220, P2_P1_EBX_REG_30_ );
dff P2_P1_EBX_REG_31__reg ( clk, reset, P2_P1_EBX_REG_31_, n16481 );
not U_inv2173 ( n74992, P2_P1_EBX_REG_31_ );
dff P2_P1_REIP_REG_16__reg ( clk, reset, P2_P1_REIP_REG_16_, n16566 );
not U_inv2174 ( n73253, P2_P1_REIP_REG_16_ );
dff P2_P1_PHYADDRPOINTER_REG_16__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_16_, n15771 );
dff P2_P1_REIP_REG_17__reg ( clk, reset, P2_P1_REIP_REG_17_, n16571 );
not U_inv2175 ( n74904, P2_P1_REIP_REG_17_ );
dff P2_P1_REIP_REG_18__reg ( clk, reset, P2_P1_REIP_REG_18_, n16576 );
not U_inv2176 ( n74914, P2_P1_REIP_REG_18_ );
dff P2_P1_ADDRESS_REG_16__reg ( clk, reset, P2_P1_ADDRESS_REG_16_, n14561 );
not U_inv2177 ( n74445, P2_P1_ADDRESS_REG_16_ );
dff P2_P1_REIP_REG_19__reg ( clk, reset, P2_P1_REIP_REG_19_, n16581 );
not U_inv2178 ( n73267, P2_P1_REIP_REG_19_ );
dff P2_P1_INSTADDRPOINTER_REG_19__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_19_, n15626 );
not U_inv2179 ( n74550, P2_P1_INSTADDRPOINTER_REG_19_ );
dff P2_P1_INSTADDRPOINTER_REG_21__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_21_, n15636 );
not U_inv2180 ( n73148, P2_P1_INSTADDRPOINTER_REG_21_ );
dff P2_P1_INSTADDRPOINTER_REG_22__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_22_, n15641 );
not U_inv2181 ( n74585, P2_P1_INSTADDRPOINTER_REG_22_ );
dff P2_P1_PHYADDRPOINTER_REG_22__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_22_, n15801 );
not U_inv2182 ( n74680, P2_P1_PHYADDRPOINTER_REG_22_ );
dff P2_P1_REIP_REG_22__reg ( clk, reset, P2_P1_REIP_REG_22_, n16596 );
not U_inv2183 ( n73280, P2_P1_REIP_REG_22_ );
dff P2_P1_REIP_REG_23__reg ( clk, reset, P2_P1_REIP_REG_23_, n16601 );
not U_inv2184 ( n74995, P2_P1_REIP_REG_23_ );
dff P2_P1_REIP_REG_24__reg ( clk, reset, P2_P1_REIP_REG_24_, n16606 );
not U_inv2185 ( n75005, P2_P1_REIP_REG_24_ );
dff P2_P1_ADDRESS_REG_22__reg ( clk, reset, P2_P1_ADDRESS_REG_22_, n14531 );
dff P2_P1_REIP_REG_25__reg ( clk, reset, P2_P1_REIP_REG_25_, n16611 );
not U_inv2186 ( n73304, P2_P1_REIP_REG_25_ );
dff P2_P1_PHYADDRPOINTER_REG_26__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_26_, n15821 );
not U_inv2187 ( n74810, P2_P1_PHYADDRPOINTER_REG_26_ );
dff P2_P1_REIP_REG_26__reg ( clk, reset, P2_P1_REIP_REG_26_, n16616 );
not U_inv2188 ( n73308, P2_P1_REIP_REG_26_ );
dff P2_P1_REIP_REG_27__reg ( clk, reset, P2_P1_REIP_REG_27_, n16621 );
not U_inv2189 ( n75014, P2_P1_REIP_REG_27_ );
dff P2_P1_PHYADDRPOINTER_REG_27__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_27_, n15826 );
not U_inv2190 ( n75208, P2_P1_PHYADDRPOINTER_REG_27_ );
dff P2_P1_REIP_REG_28__reg ( clk, reset, P2_P1_REIP_REG_28_, n16626 );
not U_inv2191 ( n75302, P2_P1_REIP_REG_28_ );
dff P2_P1_REIP_REG_29__reg ( clk, reset, P2_P1_REIP_REG_29_, n16631 );
not U_inv2192 ( n73391, P2_P1_REIP_REG_29_ );
dff P2_P1_ADDRESS_REG_27__reg ( clk, reset, P2_P1_ADDRESS_REG_27_, n14506 );
dff P2_P1_REIP_REG_30__reg ( clk, reset, P2_P1_REIP_REG_30_, n16636 );
not U_inv2193 ( n75237, P2_P1_REIP_REG_30_ );
dff P2_P1_ADDRESS_REG_28__reg ( clk, reset, P2_P1_ADDRESS_REG_28_, n14501 );
dff P2_P1_REIP_REG_31__reg ( clk, reset, P2_P1_REIP_REG_31_, n16641 );
not U_inv2194 ( n75328, P2_P1_REIP_REG_31_ );
dff P2_P1_INSTADDRPOINTER_REG_31__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_31_, n15686 );
not U_inv2195 ( n75052, P2_P1_INSTADDRPOINTER_REG_31_ );
dff P2_P1_PHYADDRPOINTER_REG_31__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_31_, n15846 );
not U_inv2196 ( n74967, P2_P1_PHYADDRPOINTER_REG_31_ );
dff P2_P1_REIP_REG_0__reg ( clk, reset, P2_P1_REIP_REG_0_, n16486 );
not U_inv2197 ( n75259, P2_P1_REIP_REG_0_ );
dff P2_P1_PHYADDRPOINTER_REG_0__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_0_, n15691 );
not U_inv2198 ( n75225, P2_P1_PHYADDRPOINTER_REG_0_ );
dff P2_P1_REIP_REG_1__reg ( clk, reset, P2_P1_REIP_REG_1_, n16491 );
not U_inv2199 ( n72962, P2_P1_REIP_REG_1_ );
dff P2_P1_BYTEENABLE_REG_0__reg ( clk, reset, P2_P1_BYTEENABLE_REG_0_, n16661 );
dff P2_P1_BE_N_REG_0__reg ( clk, reset, P2_P1_BE_N_REG_0_, n14491 );
dff P2_P1_BYTEENABLE_REG_1__reg ( clk, reset, P2_P1_BYTEENABLE_REG_1_, n16656 );
dff P2_P1_BE_N_REG_1__reg ( clk, reset, P2_P1_BE_N_REG_1_, n14486 );
dff P2_P1_PHYADDRPOINTER_REG_1__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_1_, n15696 );
not U_inv2200 ( n74467, P2_P1_PHYADDRPOINTER_REG_1_ );
dff P2_P1_BYTEENABLE_REG_3__reg ( clk, reset, P2_P1_BYTEENABLE_REG_3_, n16646 );
dff P2_P1_BE_N_REG_3__reg ( clk, reset, P2_P1_BE_N_REG_3_, n14476 );
dff P2_P1_BYTEENABLE_REG_2__reg ( clk, reset, P2_P1_BYTEENABLE_REG_2_, n16651 );
dff P2_P1_BE_N_REG_2__reg ( clk, reset, P2_P1_BE_N_REG_2_, n14481 );
dff P2_P1_REIP_REG_2__reg ( clk, reset, P2_P1_REIP_REG_2_, n16496 );
not U_inv2201 ( n74655, P2_P1_REIP_REG_2_ );
dff P2_P1_ADDRESS_REG_0__reg ( clk, reset, P2_P1_ADDRESS_REG_0_, n14641 );
dff P2_P1_PHYADDRPOINTER_REG_2__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_2_, n15701 );
not U_inv2202 ( n74717, P2_P1_PHYADDRPOINTER_REG_2_ );
dff P2_P1_REIP_REG_3__reg ( clk, reset, P2_P1_REIP_REG_3_, n16501 );
not U_inv2203 ( n72964, P2_P1_REIP_REG_3_ );
dff P2_P1_ADDRESS_REG_1__reg ( clk, reset, P2_P1_ADDRESS_REG_1_, n14636 );
dff P2_P1_REIP_REG_4__reg ( clk, reset, P2_P1_REIP_REG_4_, n16506 );
not U_inv2204 ( n74672, P2_P1_REIP_REG_4_ );
dff P2_P1_INSTADDRPOINTER_REG_4__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_4_, n15551 );
not U_inv2205 ( n75934, P2_P1_INSTADDRPOINTER_REG_4_ );
dff P2_P1_INSTADDRPOINTER_REG_5__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_5_, n15556 );
not U_inv2206 ( n74443, P2_P1_INSTADDRPOINTER_REG_5_ );
dff P2_P1_INSTADDRPOINTER_REG_6__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_6_, n15561 );
not U_inv2207 ( n73065, P2_P1_INSTADDRPOINTER_REG_6_ );
dff P2_P1_PHYADDRPOINTER_REG_6__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_6_, n15721 );
not U_inv2208 ( n74500, P2_P1_PHYADDRPOINTER_REG_6_ );
dff P2_P1_INSTADDRPOINTER_REG_7__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_7_, n15566 );
not U_inv2209 ( n74659, P2_P1_INSTADDRPOINTER_REG_7_ );
dff P2_P1_PHYADDRPOINTER_REG_7__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_7_, n15726 );
not U_inv2210 ( n73098, P2_P1_PHYADDRPOINTER_REG_7_ );
dff P2_P1_REIP_REG_7__reg ( clk, reset, P2_P1_REIP_REG_7_, n16521 );
not U_inv2211 ( n73206, P2_P1_REIP_REG_7_ );
dff P2_P1_PHYADDRPOINTER_REG_8__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_8_, n15731 );
not U_inv2212 ( n74522, P2_P1_PHYADDRPOINTER_REG_8_ );
dff P2_P1_REIP_REG_8__reg ( clk, reset, P2_P1_REIP_REG_8_, n16526 );
not U_inv2213 ( n75965, P2_P1_REIP_REG_8_ );
dff P2_P1_ADDRESS_REG_6__reg ( clk, reset, P2_P1_ADDRESS_REG_6_, n14611 );
not U_inv2214 ( n73057, P2_P1_ADDRESS_REG_6_ );
dff P2_P1_PHYADDRPOINTER_REG_9__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_9_, n15736 );
not U_inv2215 ( n73108, P2_P1_PHYADDRPOINTER_REG_9_ );
dff P2_P1_REIP_REG_9__reg ( clk, reset, ex_wire261, n16531 );
not U_inv2216 ( n73221, ex_wire261 );
dff P2_P1_ADDRESS_REG_7__reg ( clk, reset, P2_P1_ADDRESS_REG_7_, n14606 );
not U_inv2217 ( n73529, P2_P1_ADDRESS_REG_7_ );
dff P2_P1_PHYADDRPOINTER_REG_10__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_10_, n15741 );
not U_inv2218 ( n74554, P2_P1_PHYADDRPOINTER_REG_10_ );
dff P2_P1_REIP_REG_10__reg ( clk, reset, P2_P1_REIP_REG_10_, n16536 );
not U_inv2219 ( n74769, P2_P1_REIP_REG_10_ );
dff P2_P1_INSTADDRPOINTER_REG_10__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_10_, n15581 );
not U_inv2220 ( n74734, P2_P1_INSTADDRPOINTER_REG_10_ );
dff P2_P1_ADDRESS_REG_8__reg ( clk, reset, P2_P1_ADDRESS_REG_8_, n14601 );
not U_inv2221 ( n73062, P2_P1_ADDRESS_REG_8_ );
dff P2_P1_PHYADDRPOINTER_REG_11__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_11_, n15746 );
not U_inv2222 ( n74451, P2_P1_PHYADDRPOINTER_REG_11_ );
dff P2_P1_REIP_REG_11__reg ( clk, reset, P2_P1_REIP_REG_11_, n16541 );
not U_inv2223 ( n74811, P2_P1_REIP_REG_11_ );
dff P2_P1_ADDRESS_REG_9__reg ( clk, reset, P2_P1_ADDRESS_REG_9_, n14596 );
not U_inv2224 ( n73822, P2_P1_ADDRESS_REG_9_ );
dff P2_P1_REIP_REG_12__reg ( clk, reset, ex_wire262, n16546 );
not U_inv2225 ( n74815, ex_wire262 );
dff P2_P1_INSTADDRPOINTER_REG_12__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_12_, n15591 );
not U_inv2226 ( n74427, P2_P1_INSTADDRPOINTER_REG_12_ );
dff P2_P1_PHYADDRPOINTER_REG_12__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_12_, n15751 );
not U_inv2227 ( n74607, P2_P1_PHYADDRPOINTER_REG_12_ );
dff P2_P1_PHYADDRPOINTER_REG_13__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_13_, n15756 );
dff P2_P1_REIP_REG_13__reg ( clk, reset, P2_P1_REIP_REG_13_, n16551 );
not U_inv2228 ( n73239, P2_P1_REIP_REG_13_ );
dff P2_P1_REIP_REG_14__reg ( clk, reset, P2_P1_REIP_REG_14_, n16556 );
not U_inv2229 ( n74860, P2_P1_REIP_REG_14_ );
dff P2_P1_INSTADDRPOINTER_REG_14__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_14_, n15601 );
not U_inv2230 ( n74417, P2_P1_INSTADDRPOINTER_REG_14_ );
dff P2_P1_PHYADDRPOINTER_REG_14__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_14_, n15761 );
not U_inv2231 ( n74871, P2_P1_PHYADDRPOINTER_REG_14_ );
dff P2_P1_ADDRESS_REG_12__reg ( clk, reset, P2_P1_ADDRESS_REG_12_, n14581 );
not U_inv2232 ( n73070, P2_P1_ADDRESS_REG_12_ );
dff P2_P1_INSTADDRPOINTER_REG_15__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_15_, n15606 );
not U_inv2233 ( n74822, P2_P1_INSTADDRPOINTER_REG_15_ );
dff P2_P1_INSTADDRPOINTER_REG_17__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_17_, n15616 );
not U_inv2234 ( n74841, P2_P1_INSTADDRPOINTER_REG_17_ );
dff P2_P1_INSTADDRPOINTER_REG_18__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_18_, n15621 );
not U_inv2235 ( n74524, P2_P1_INSTADDRPOINTER_REG_18_ );
dff P2_P1_INSTADDRPOINTER_REG_23__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_23_, n15646 );
not U_inv2236 ( n73159, P2_P1_INSTADDRPOINTER_REG_23_ );
dff P2_P1_INSTADDRPOINTER_REG_28__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_28_, n15671 );
not U_inv2237 ( n74974, P2_P1_INSTADDRPOINTER_REG_28_ );
dff P2_P1_INSTADDRPOINTER_REG_29__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_29_, n15676 );
not U_inv2238 ( n74986, P2_P1_INSTADDRPOINTER_REG_29_ );
dff P2_P1_PHYADDRPOINTER_REG_15__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_15_, n15766 );
not U_inv2239 ( n75197, P2_P1_PHYADDRPOINTER_REG_15_ );
dff P2_P1_PHYADDRPOINTER_REG_17__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_17_, n15776 );
not U_inv2240 ( n74515, P2_P1_PHYADDRPOINTER_REG_17_ );
dff P2_P1_PHYADDRPOINTER_REG_18__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_18_, n15781 );
not U_inv2241 ( n74772, P2_P1_PHYADDRPOINTER_REG_18_ );
dff P2_P1_PHYADDRPOINTER_REG_19__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_19_, n15786 );
dff P2_P1_REIP_REG_15__reg ( clk, reset, P2_P1_REIP_REG_15_, n16561 );
not U_inv2242 ( n74868, P2_P1_REIP_REG_15_ );
dff P2_P1_REIP_REG_20__reg ( clk, reset, P2_P1_REIP_REG_20_, n16586 );
not U_inv2243 ( n74951, P2_P1_REIP_REG_20_ );
dff P2_P1_PHYADDRPOINTER_REG_20__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_20_, n15791 );
not U_inv2244 ( n74957, P2_P1_PHYADDRPOINTER_REG_20_ );
dff P2_P1_REIP_REG_21__reg ( clk, reset, P2_P1_REIP_REG_21_, n16591 );
not U_inv2245 ( n74958, P2_P1_REIP_REG_21_ );
dff P2_P1_PHYADDRPOINTER_REG_21__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_21_, n15796 );
not U_inv2246 ( n75202, P2_P1_PHYADDRPOINTER_REG_21_ );
dff P2_P1_PHYADDRPOINTER_REG_23__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_23_, n15806 );
not U_inv2247 ( n74998, P2_P1_PHYADDRPOINTER_REG_23_ );
dff P2_P1_PHYADDRPOINTER_REG_24__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_24_, n15811 );
not U_inv2248 ( n74740, P2_P1_PHYADDRPOINTER_REG_24_ );
dff P2_P1_PHYADDRPOINTER_REG_25__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_25_, n15816 );
not U_inv2249 ( n75236, P2_P1_PHYADDRPOINTER_REG_25_ );
dff P2_P1_PHYADDRPOINTER_REG_28__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_28_, n15831 );
not U_inv2250 ( n74891, P2_P1_PHYADDRPOINTER_REG_28_ );
dff P2_P1_PHYADDRPOINTER_REG_29__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_29_, n15836 );
not U_inv2251 ( n75077, P2_P1_PHYADDRPOINTER_REG_29_ );
dff P2_P1_PHYADDRPOINTER_REG_30__reg ( clk, reset, P2_P1_PHYADDRPOINTER_REG_30_, n15841 );
not U_inv2252 ( n74931, P2_P1_PHYADDRPOINTER_REG_30_ );
dff P2_P1_ADDRESS_REG_19__reg ( clk, reset, P2_P1_ADDRESS_REG_19_, n14546 );
dff P2_P1_ADDRESS_REG_13__reg ( clk, reset, P2_P1_ADDRESS_REG_13_, n14576 );
not U_inv2253 ( n74387, P2_P1_ADDRESS_REG_13_ );
dff P2_P1_ADDRESS_REG_10__reg ( clk, reset, P2_P1_ADDRESS_REG_10_, n14591 );
not U_inv2254 ( n73064, P2_P1_ADDRESS_REG_10_ );
dff P2_P1_ADDRESS_REG_11__reg ( clk, reset, P2_P1_ADDRESS_REG_11_, n14586 );
not U_inv2255 ( n74273, P2_P1_ADDRESS_REG_11_ );
dff P2_P1_ADDRESS_REG_2__reg ( clk, reset, P2_P1_ADDRESS_REG_2_, n14631 );
not U_inv2256 ( n73028, P2_P1_ADDRESS_REG_2_ );
dff P2_P1_ADDRESS_REG_3__reg ( clk, reset, P2_P1_ADDRESS_REG_3_, n14626 );
not U_inv2257 ( n73473, P2_P1_ADDRESS_REG_3_ );
dff P2_P1_ADDRESS_REG_29__reg ( clk, reset, P2_P1_ADDRESS_REG_29_, n14496 );
dff P2_P1_ADDRESS_REG_25__reg ( clk, reset, P2_P1_ADDRESS_REG_25_, n14516 );
dff P2_P1_ADDRESS_REG_26__reg ( clk, reset, P2_P1_ADDRESS_REG_26_, n14511 );
dff P2_P1_ADDRESS_REG_23__reg ( clk, reset, P2_P1_ADDRESS_REG_23_, n14526 );
dff P2_P1_ADDRESS_REG_24__reg ( clk, reset, P2_P1_ADDRESS_REG_24_, n14521 );
dff P2_P1_ADDRESS_REG_20__reg ( clk, reset, P2_P1_ADDRESS_REG_20_, n14541 );
dff P2_P1_ADDRESS_REG_21__reg ( clk, reset, P2_P1_ADDRESS_REG_21_, n14536 );
dff P2_P1_ADDRESS_REG_17__reg ( clk, reset, P2_P1_ADDRESS_REG_17_, n14556 );
not U_inv2258 ( n73125, P2_P1_ADDRESS_REG_17_ );
dff P2_P1_ADDRESS_REG_18__reg ( clk, reset, P2_P1_ADDRESS_REG_18_, n14551 );
not U_inv2259 ( n74494, P2_P1_ADDRESS_REG_18_ );
dff P2_P1_ADDRESS_REG_14__reg ( clk, reset, P2_P1_ADDRESS_REG_14_, n14571 );
not U_inv2260 ( n73096, P2_P1_ADDRESS_REG_14_ );
dff P2_P1_ADDRESS_REG_15__reg ( clk, reset, P2_P1_ADDRESS_REG_15_, n14566 );
not U_inv2261 ( n74436, P2_P1_ADDRESS_REG_15_ );
dff P1_P3_REQUESTPENDING_REG_reg ( clk, reset, P1_P3_REQUESTPENDING_REG, n5461 );
not U_inv2262 ( n75256, P1_P3_REQUESTPENDING_REG );
dff P1_P2_ADDRESS_REG_0__reg ( clk, reset, P1_P2_ADDRESS_REG_0_, n5661 );
not U_inv2263 ( n73514, P1_P2_ADDRESS_REG_0_ );
dff P1_P2_ADDRESS_REG_1__reg ( clk, reset, P1_P2_ADDRESS_REG_1_, n5656 );
not U_inv2264 ( n73488, P1_P2_ADDRESS_REG_1_ );
dff P1_P2_ADDRESS_REG_2__reg ( clk, reset, P1_P2_ADDRESS_REG_2_, n5651 );
not U_inv2265 ( n73489, P1_P2_ADDRESS_REG_2_ );
dff P1_P2_ADDRESS_REG_3__reg ( clk, reset, P1_P2_ADDRESS_REG_3_, n5646 );
not U_inv2266 ( n73043, P1_P2_ADDRESS_REG_3_ );
dff P1_P2_ADDRESS_REG_4__reg ( clk, reset, P1_P2_ADDRESS_REG_4_, n5641 );
not U_inv2267 ( n73476, P1_P2_ADDRESS_REG_4_ );
dff P1_P2_ADDRESS_REG_5__reg ( clk, reset, P1_P2_ADDRESS_REG_5_, n5636 );
not U_inv2268 ( n73040, P1_P2_ADDRESS_REG_5_ );
dff P1_P2_ADDRESS_REG_6__reg ( clk, reset, P1_P2_ADDRESS_REG_6_, n5631 );
not U_inv2269 ( n73466, P1_P2_ADDRESS_REG_6_ );
dff P1_P2_ADDRESS_REG_7__reg ( clk, reset, P1_P2_ADDRESS_REG_7_, n5626 );
not U_inv2270 ( n73036, P1_P2_ADDRESS_REG_7_ );
dff P1_P2_ADDRESS_REG_8__reg ( clk, reset, P1_P2_ADDRESS_REG_8_, n5621 );
not U_inv2271 ( n73037, P1_P2_ADDRESS_REG_8_ );
dff P1_P2_ADDRESS_REG_9__reg ( clk, reset, P1_P2_ADDRESS_REG_9_, n5616 );
not U_inv2272 ( n73460, P1_P2_ADDRESS_REG_9_ );
dff P1_P2_ADDRESS_REG_10__reg ( clk, reset, P1_P2_ADDRESS_REG_10_, n5611 );
not U_inv2273 ( n73450, P1_P2_ADDRESS_REG_10_ );
dff P1_P2_ADDRESS_REG_11__reg ( clk, reset, P1_P2_ADDRESS_REG_11_, n5606 );
not U_inv2274 ( n73029, P1_P2_ADDRESS_REG_11_ );
dff P1_P2_ADDRESS_REG_12__reg ( clk, reset, P1_P2_ADDRESS_REG_12_, n5601 );
not U_inv2275 ( n73031, P1_P2_ADDRESS_REG_12_ );
dff P1_P2_ADDRESS_REG_13__reg ( clk, reset, P1_P2_ADDRESS_REG_13_, n5596 );
not U_inv2276 ( n73444, P1_P2_ADDRESS_REG_13_ );
dff P1_P2_ADDRESS_REG_14__reg ( clk, reset, P1_P2_ADDRESS_REG_14_, n5591 );
not U_inv2277 ( n73033, P1_P2_ADDRESS_REG_14_ );
dff P1_P2_ADDRESS_REG_15__reg ( clk, reset, P1_P2_ADDRESS_REG_15_, n5586 );
not U_inv2278 ( n73454, P1_P2_ADDRESS_REG_15_ );
dff P1_P2_ADDRESS_REG_16__reg ( clk, reset, P1_P2_ADDRESS_REG_16_, n5581 );
not U_inv2279 ( n73482, P1_P2_ADDRESS_REG_16_ );
dff P1_P2_ADDRESS_REG_17__reg ( clk, reset, P1_P2_ADDRESS_REG_17_, n5576 );
not U_inv2280 ( n73048, P1_P2_ADDRESS_REG_17_ );
dff P1_P2_ADDRESS_REG_18__reg ( clk, reset, P1_P2_ADDRESS_REG_18_, n5571 );
not U_inv2281 ( n73507, P1_P2_ADDRESS_REG_18_ );
dff P1_P2_ADDRESS_REG_19__reg ( clk, reset, P1_P2_ADDRESS_REG_19_, n5566 );
dff P1_P2_ADDRESS_REG_20__reg ( clk, reset, P1_P2_ADDRESS_REG_20_, n5561 );
dff P1_P2_ADDRESS_REG_21__reg ( clk, reset, P1_P2_ADDRESS_REG_21_, n5556 );
dff P1_P2_ADDRESS_REG_22__reg ( clk, reset, P1_P2_ADDRESS_REG_22_, n5551 );
dff P1_P2_ADDRESS_REG_23__reg ( clk, reset, P1_P2_ADDRESS_REG_23_, n5546 );
dff P1_P2_ADDRESS_REG_24__reg ( clk, reset, P1_P2_ADDRESS_REG_24_, n5541 );
dff P1_P2_ADDRESS_REG_25__reg ( clk, reset, P1_P2_ADDRESS_REG_25_, n5536 );
dff P1_P2_ADDRESS_REG_26__reg ( clk, reset, P1_P2_ADDRESS_REG_26_, n5531 );
dff P1_P2_ADDRESS_REG_27__reg ( clk, reset, P1_P2_ADDRESS_REG_27_, n5526 );
dff P1_P2_ADDRESS_REG_28__reg ( clk, reset, P1_P2_ADDRESS_REG_28_, n5521 );
dff P1_P1_REIP_REG_2__reg ( clk, reset, P1_P1_REIP_REG_2_, n9761 );
not U_inv2282 ( n74656, P1_P1_REIP_REG_2_ );
dff P1_P1_ADDRESS_REG_0__reg ( clk, reset, P1_P1_ADDRESS_REG_0_, n7906 );
dff P1_P1_PHYADDRPOINTER_REG_2__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_2_, n8966 );
not U_inv2283 ( n74718, P1_P1_PHYADDRPOINTER_REG_2_ );
dff P1_P1_REIP_REG_3__reg ( clk, reset, P1_P1_REIP_REG_3_, n9766 );
not U_inv2284 ( n72965, P1_P1_REIP_REG_3_ );
dff P1_P1_ADDRESS_REG_1__reg ( clk, reset, P1_P1_ADDRESS_REG_1_, n7901 );
dff P1_P1_REIP_REG_4__reg ( clk, reset, P1_P1_REIP_REG_4_, n9771 );
not U_inv2285 ( n74673, P1_P1_REIP_REG_4_ );
dff P1_P1_INSTADDRPOINTER_REG_4__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_4_, n8816 );
not U_inv2286 ( n75941, P1_P1_INSTADDRPOINTER_REG_4_ );
dff P1_P1_INSTADDRPOINTER_REG_5__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_5_, n8821 );
not U_inv2287 ( n74461, P1_P1_INSTADDRPOINTER_REG_5_ );
dff P1_P1_INSTADDRPOINTER_REG_6__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_6_, n8826 );
not U_inv2288 ( n73090, P1_P1_INSTADDRPOINTER_REG_6_ );
dff P1_P1_PHYADDRPOINTER_REG_6__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_6_, n8986 );
not U_inv2289 ( n74506, P1_P1_PHYADDRPOINTER_REG_6_ );
dff P1_P1_INSTADDRPOINTER_REG_7__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_7_, n8831 );
not U_inv2290 ( n74658, P1_P1_INSTADDRPOINTER_REG_7_ );
dff P1_P1_PHYADDRPOINTER_REG_7__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_7_, n8991 );
not U_inv2291 ( n73097, P1_P1_PHYADDRPOINTER_REG_7_ );
dff P1_P1_REIP_REG_7__reg ( clk, reset, P1_P1_REIP_REG_7_, n9786 );
not U_inv2292 ( n73207, P1_P1_REIP_REG_7_ );
dff P1_P1_PHYADDRPOINTER_REG_8__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_8_, n8996 );
not U_inv2293 ( n74541, P1_P1_PHYADDRPOINTER_REG_8_ );
dff P1_P1_REIP_REG_8__reg ( clk, reset, P1_P1_REIP_REG_8_, n9791 );
not U_inv2294 ( n75967, P1_P1_REIP_REG_8_ );
dff P1_P1_ADDRESS_REG_6__reg ( clk, reset, P1_P1_ADDRESS_REG_6_, n7876 );
not U_inv2295 ( n73467, P1_P1_ADDRESS_REG_6_ );
dff P1_P1_PHYADDRPOINTER_REG_9__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_9_, n9001 );
not U_inv2296 ( n73107, P1_P1_PHYADDRPOINTER_REG_9_ );
dff P1_P1_REIP_REG_9__reg ( clk, reset, ex_wire263, n9796 );
not U_inv2297 ( n73222, ex_wire263 );
dff P1_P1_ADDRESS_REG_7__reg ( clk, reset, P1_P1_ADDRESS_REG_7_, n7871 );
not U_inv2298 ( n73038, P1_P1_ADDRESS_REG_7_ );
dff P1_P1_PHYADDRPOINTER_REG_10__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_10_, n9006 );
not U_inv2299 ( n74577, P1_P1_PHYADDRPOINTER_REG_10_ );
dff P1_P1_REIP_REG_10__reg ( clk, reset, P1_P1_REIP_REG_10_, n9801 );
not U_inv2300 ( n74770, P1_P1_REIP_REG_10_ );
dff P1_P1_INSTADDRPOINTER_REG_10__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_10_, n8846 );
not U_inv2301 ( n74735, P1_P1_INSTADDRPOINTER_REG_10_ );
dff P1_P1_ADDRESS_REG_8__reg ( clk, reset, P1_P1_ADDRESS_REG_8_, n7866 );
not U_inv2302 ( n73039, P1_P1_ADDRESS_REG_8_ );
dff P1_P1_PHYADDRPOINTER_REG_11__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_11_, n9011 );
not U_inv2303 ( n74450, P1_P1_PHYADDRPOINTER_REG_11_ );
dff P1_P1_REIP_REG_11__reg ( clk, reset, P1_P1_REIP_REG_11_, n9806 );
not U_inv2304 ( n74812, P1_P1_REIP_REG_11_ );
dff P1_P1_ADDRESS_REG_9__reg ( clk, reset, P1_P1_ADDRESS_REG_9_, n7861 );
not U_inv2305 ( n73463, P1_P1_ADDRESS_REG_9_ );
dff P1_P1_REIP_REG_12__reg ( clk, reset, ex_wire264, n9811 );
not U_inv2306 ( n74816, ex_wire264 );
dff P1_P1_INSTADDRPOINTER_REG_12__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_12_, n8856 );
not U_inv2307 ( n74476, P1_P1_INSTADDRPOINTER_REG_12_ );
dff P1_P1_PHYADDRPOINTER_REG_12__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_12_, n9016 );
not U_inv2308 ( n74644, P1_P1_PHYADDRPOINTER_REG_12_ );
dff P1_P1_PHYADDRPOINTER_REG_13__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_13_, n9021 );
dff P1_P1_REIP_REG_13__reg ( clk, reset, P1_P1_REIP_REG_13_, n9816 );
not U_inv2309 ( n73240, P1_P1_REIP_REG_13_ );
dff P1_P1_INSTADDRPOINTER_REG_14__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_14_, n8866 );
not U_inv2310 ( n73117, P1_P1_INSTADDRPOINTER_REG_14_ );
dff P1_P1_PHYADDRPOINTER_REG_14__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_14_, n9026 );
not U_inv2311 ( n74870, P1_P1_PHYADDRPOINTER_REG_14_ );
dff P1_P1_REIP_REG_14__reg ( clk, reset, P1_P1_REIP_REG_14_, n9821 );
not U_inv2312 ( n74861, P1_P1_REIP_REG_14_ );
dff P1_P1_ADDRESS_REG_12__reg ( clk, reset, P1_P1_ADDRESS_REG_12_, n7846 );
not U_inv2313 ( n73032, P1_P1_ADDRESS_REG_12_ );
dff P1_P1_INSTADDRPOINTER_REG_15__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_15_, n8871 );
not U_inv2314 ( n74823, P1_P1_INSTADDRPOINTER_REG_15_ );
dff P1_P1_INSTADDRPOINTER_REG_17__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_17_, n8881 );
not U_inv2315 ( n74847, P1_P1_INSTADDRPOINTER_REG_17_ );
dff P1_P1_INSTADDRPOINTER_REG_18__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_18_, n8886 );
not U_inv2316 ( n74599, P1_P1_INSTADDRPOINTER_REG_18_ );
dff P1_P1_PHYADDRPOINTER_REG_15__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_15_, n9031 );
not U_inv2317 ( n75200, P1_P1_PHYADDRPOINTER_REG_15_ );
dff P1_P1_PHYADDRPOINTER_REG_17__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_17_, n9041 );
not U_inv2318 ( n74512, P1_P1_PHYADDRPOINTER_REG_17_ );
dff P1_P1_PHYADDRPOINTER_REG_18__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_18_, n9046 );
not U_inv2319 ( n74785, P1_P1_PHYADDRPOINTER_REG_18_ );
dff P1_P1_PHYADDRPOINTER_REG_19__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_19_, n9051 );
dff P1_P1_REIP_REG_15__reg ( clk, reset, P1_P1_REIP_REG_15_, n9826 );
not U_inv2320 ( n74869, P1_P1_REIP_REG_15_ );
dff P1_P1_REIP_REG_20__reg ( clk, reset, P1_P1_REIP_REG_20_, n9851 );
not U_inv2321 ( n74952, P1_P1_REIP_REG_20_ );
dff P1_P1_PHYADDRPOINTER_REG_20__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_20_, n9056 );
not U_inv2322 ( n74956, P1_P1_PHYADDRPOINTER_REG_20_ );
dff P1_P1_REIP_REG_21__reg ( clk, reset, P1_P1_REIP_REG_21_, n9856 );
not U_inv2323 ( n74959, P1_P1_REIP_REG_21_ );
dff P1_P1_PHYADDRPOINTER_REG_21__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_21_, n9061 );
not U_inv2324 ( n75201, P1_P1_PHYADDRPOINTER_REG_21_ );
dff P1_P1_ADDRESS_REG_19__reg ( clk, reset, P1_P1_ADDRESS_REG_19_, n7811 );
dff P1_P1_REIP_REG_22__reg ( clk, reset, P1_P1_REIP_REG_22_, n9861 );
not U_inv2325 ( n73281, P1_P1_REIP_REG_22_ );
dff P1_P1_PHYADDRPOINTER_REG_22__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_22_, n9066 );
not U_inv2326 ( n74677, P1_P1_PHYADDRPOINTER_REG_22_ );
dff P1_P1_REIP_REG_23__reg ( clk, reset, P1_P1_REIP_REG_23_, n9866 );
not U_inv2327 ( n74996, P1_P1_REIP_REG_23_ );
dff P1_P1_INSTADDRPOINTER_REG_23__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_23_, n8911 );
not U_inv2328 ( n74920, P1_P1_INSTADDRPOINTER_REG_23_ );
dff P1_P1_PHYADDRPOINTER_REG_23__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_23_, n9071 );
not U_inv2329 ( n74997, P1_P1_PHYADDRPOINTER_REG_23_ );
dff P1_P1_PHYADDRPOINTER_REG_25__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_25_, n9081 );
not U_inv2330 ( n75235, P1_P1_PHYADDRPOINTER_REG_25_ );
dff P1_P1_REIP_REG_28__reg ( clk, reset, P1_P1_REIP_REG_28_, n9891 );
not U_inv2331 ( n75303, P1_P1_REIP_REG_28_ );
dff P1_P1_INSTADDRPOINTER_REG_29__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_29_, n8941 );
not U_inv2332 ( n73279, P1_P1_INSTADDRPOINTER_REG_29_ );
dff P1_P1_INSTADDRPOINTER_REG_30__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_30_, n8946 );
not U_inv2333 ( n74989, P1_P1_INSTADDRPOINTER_REG_30_ );
dff P1_P1_PHYADDRPOINTER_REG_28__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_28_, n9096 );
not U_inv2334 ( n74880, P1_P1_PHYADDRPOINTER_REG_28_ );
dff P1_P1_PHYADDRPOINTER_REG_29__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_29_, n9101 );
not U_inv2335 ( n75170, P1_P1_PHYADDRPOINTER_REG_29_ );
dff P1_P1_PHYADDRPOINTER_REG_30__reg ( clk, reset, P1_P1_PHYADDRPOINTER_REG_30_, n9106 );
not U_inv2336 ( n74924, P1_P1_PHYADDRPOINTER_REG_30_ );
dff P1_P1_ADDRESS_REG_27__reg ( clk, reset, P1_P1_ADDRESS_REG_27_, n7771 );
dff P1_P1_ADDRESS_REG_22__reg ( clk, reset, P1_P1_ADDRESS_REG_22_, n7796 );
dff P1_P1_ADDRESS_REG_20__reg ( clk, reset, P1_P1_ADDRESS_REG_20_, n7806 );
dff P1_P1_ADDRESS_REG_21__reg ( clk, reset, P1_P1_ADDRESS_REG_21_, n7801 );
dff P1_P1_ADDRESS_REG_13__reg ( clk, reset, P1_P1_ADDRESS_REG_13_, n7841 );
not U_inv2337 ( n73445, P1_P1_ADDRESS_REG_13_ );
dff P1_P1_ADDRESS_REG_10__reg ( clk, reset, P1_P1_ADDRESS_REG_10_, n7856 );
not U_inv2338 ( n73451, P1_P1_ADDRESS_REG_10_ );
dff P1_P1_ADDRESS_REG_11__reg ( clk, reset, P1_P1_ADDRESS_REG_11_, n7851 );
not U_inv2339 ( n73030, P1_P1_ADDRESS_REG_11_ );
dff P1_P1_ADDRESS_REG_2__reg ( clk, reset, P1_P1_ADDRESS_REG_2_, n7896 );
not U_inv2340 ( n73490, P1_P1_ADDRESS_REG_2_ );
dff P1_P1_ADDRESS_REG_3__reg ( clk, reset, P1_P1_ADDRESS_REG_3_, n7891 );
not U_inv2341 ( n73044, P1_P1_ADDRESS_REG_3_ );
dff P1_P1_ADDRESS_REG_29__reg ( clk, reset, P1_P1_ADDRESS_REG_29_, n7761 );
dff P1_P1_ADDRESS_REG_25__reg ( clk, reset, P1_P1_ADDRESS_REG_25_, n7781 );
dff P1_P1_ADDRESS_REG_26__reg ( clk, reset, P1_P1_ADDRESS_REG_26_, n7776 );
dff P1_P1_ADDRESS_REG_23__reg ( clk, reset, P1_P1_ADDRESS_REG_23_, n7791 );
dff P1_P1_ADDRESS_REG_24__reg ( clk, reset, P1_P1_ADDRESS_REG_24_, n7786 );
dff P1_P1_ADDRESS_REG_17__reg ( clk, reset, P1_P1_ADDRESS_REG_17_, n7821 );
not U_inv2342 ( n73049, P1_P1_ADDRESS_REG_17_ );
dff P1_P1_ADDRESS_REG_18__reg ( clk, reset, P1_P1_ADDRESS_REG_18_, n7816 );
not U_inv2343 ( n73508, P1_P1_ADDRESS_REG_18_ );
dff P1_P1_ADDRESS_REG_14__reg ( clk, reset, P1_P1_ADDRESS_REG_14_, n7836 );
not U_inv2344 ( n73034, P1_P1_ADDRESS_REG_14_ );
dff P1_P1_ADDRESS_REG_15__reg ( clk, reset, P1_P1_ADDRESS_REG_15_, n7831 );
not U_inv2345 ( n73455, P1_P1_ADDRESS_REG_15_ );
dff P2_P3_REQUESTPENDING_REG_reg ( clk, reset, P2_P3_REQUESTPENDING_REG, n12196 );
not U_inv2346 ( n75227, P2_P3_REQUESTPENDING_REG );
dff P2_P2_ADDRESS_REG_23__reg ( clk, reset, P2_P2_ADDRESS_REG_23_, n12281 );
dff P2_P2_ADDRESS_REG_24__reg ( clk, reset, P2_P2_ADDRESS_REG_24_, n12276 );
dff P2_P2_ADDRESS_REG_20__reg ( clk, reset, P2_P2_ADDRESS_REG_20_, n12296 );
dff P2_P2_ADDRESS_REG_21__reg ( clk, reset, P2_P2_ADDRESS_REG_21_, n12291 );
dff P2_P2_ADDRESS_REG_17__reg ( clk, reset, P2_P2_ADDRESS_REG_17_, n12311 );
not U_inv2347 ( n73124, P2_P2_ADDRESS_REG_17_ );
dff P2_P2_ADDRESS_REG_18__reg ( clk, reset, P2_P2_ADDRESS_REG_18_, n12306 );
not U_inv2348 ( n74493, P2_P2_ADDRESS_REG_18_ );
dff P2_P2_ADDRESS_REG_14__reg ( clk, reset, P2_P2_ADDRESS_REG_14_, n12326 );
not U_inv2349 ( n73095, P2_P2_ADDRESS_REG_14_ );
dff P2_P2_ADDRESS_REG_15__reg ( clk, reset, P2_P2_ADDRESS_REG_15_, n12321 );
not U_inv2350 ( n74434, P2_P2_ADDRESS_REG_15_ );
dff P2_P2_ADDRESS_REG_10__reg ( clk, reset, P2_P2_ADDRESS_REG_10_, n12346 );
not U_inv2351 ( n73063, P2_P2_ADDRESS_REG_10_ );
dff P2_P2_ADDRESS_REG_11__reg ( clk, reset, P2_P2_ADDRESS_REG_11_, n12341 );
not U_inv2352 ( n74266, P2_P2_ADDRESS_REG_11_ );
dff P2_P2_ADDRESS_REG_4__reg ( clk, reset, P2_P2_ADDRESS_REG_4_, n12376 );
not U_inv2353 ( n73045, P2_P2_ADDRESS_REG_4_ );
dff P2_P2_ADDRESS_REG_5__reg ( clk, reset, P2_P2_ADDRESS_REG_5_, n12371 );
not U_inv2354 ( n73498, P2_P2_ADDRESS_REG_5_ );
dff P2_P1_LWORD_REG_7__reg ( clk, reset, P2_P1_LWORD_REG_7_, n15891 );
not U_inv2355 ( n75652, P2_P1_LWORD_REG_7_ );
dff P2_P1_DATAO_REG_7__reg ( clk, reset, P2_P1_DATAO_REG_7_, n16041 );
dff P2_BUF1_REG_7__reg ( clk, reset, P2_BUF1_REG_7_, n496 );
not U_inv2356 ( n75448, P2_BUF1_REG_7_ );
dff P3_REG2_REG_10__reg ( clk, reset, ex_wire265, n1491 );
not U_inv2357 ( n74381, ex_wire265 );
dff P3_REG1_REG_12__reg ( clk, reset, P3_REG1_REG_12_, n1341 );
not U_inv2358 ( n74397, P3_REG1_REG_12_ );
dff P3_REG0_REG_12__reg ( clk, reset, P3_REG0_REG_12_, n1181 );
dff P3_REG1_REG_14__reg ( clk, reset, P3_REG1_REG_14_, n1351 );
not U_inv2359 ( n74430, P3_REG1_REG_14_ );
dff P3_REG0_REG_14__reg ( clk, reset, P3_REG0_REG_14_, n1191 );
dff P3_REG2_REG_13__reg ( clk, reset, P3_REG2_REG_13_, n1506 );
not U_inv2360 ( n74401, P3_REG2_REG_13_ );
dff P3_REG1_REG_15__reg ( clk, reset, P3_REG1_REG_15_, n1356 );
not U_inv2361 ( n74413, P3_REG1_REG_15_ );
dff P3_REG0_REG_15__reg ( clk, reset, P3_REG0_REG_15_, n1196 );
dff P3_REG1_REG_17__reg ( clk, reset, P3_REG1_REG_17_, n1366 );
not U_inv2362 ( n74449, P3_REG1_REG_17_ );
dff P3_REG0_REG_17__reg ( clk, reset, P3_REG0_REG_17_, n1206 );
dff P3_REG2_REG_16__reg ( clk, reset, P3_REG2_REG_16_, n1521 );
not U_inv2363 ( n74415, P3_REG2_REG_16_ );
dff P3_REG1_REG_18__reg ( clk, reset, P3_REG1_REG_18_, n1371 );
not U_inv2364 ( n74475, P3_REG1_REG_18_ );
dff P3_REG0_REG_18__reg ( clk, reset, P3_REG0_REG_18_, n1211 );
dff P3_REG1_REG_20__reg ( clk, reset, P3_REG1_REG_20_, n1381 );
not U_inv2365 ( n74501, P3_REG1_REG_20_ );
dff P3_REG0_REG_20__reg ( clk, reset, P3_REG0_REG_20_, n1221 );
dff P3_REG2_REG_19__reg ( clk, reset, ex_wire266, n1536 );
not U_inv2366 ( n74497, ex_wire266 );
dff P3_REG1_REG_21__reg ( clk, reset, P3_REG1_REG_21_, n1386 );
not U_inv2367 ( n74521, P3_REG1_REG_21_ );
dff P3_REG0_REG_21__reg ( clk, reset, P3_REG0_REG_21_, n1226 );
dff P3_REG1_REG_22__reg ( clk, reset, P3_REG1_REG_22_, n1391 );
not U_inv2368 ( n74551, P3_REG1_REG_22_ );
dff P3_REG0_REG_22__reg ( clk, reset, P3_REG0_REG_22_, n1231 );
dff P3_REG1_REG_23__reg ( clk, reset, P3_REG1_REG_23_, n1396 );
not U_inv2369 ( n74553, P3_REG1_REG_23_ );
dff P3_REG0_REG_23__reg ( clk, reset, P3_REG0_REG_23_, n1236 );
dff P3_REG1_REG_24__reg ( clk, reset, P3_REG1_REG_24_, n1401 );
not U_inv2370 ( n74647, P3_REG1_REG_24_ );
dff P3_REG0_REG_24__reg ( clk, reset, P3_REG0_REG_24_, n1241 );
dff P3_REG1_REG_25__reg ( clk, reset, P3_REG1_REG_25_, n1406 );
not U_inv2371 ( n74725, P3_REG1_REG_25_ );
dff P3_REG0_REG_25__reg ( clk, reset, P3_REG0_REG_25_, n1246 );
dff P3_REG1_REG_26__reg ( clk, reset, P3_REG1_REG_26_, n1411 );
not U_inv2372 ( n74768, P3_REG1_REG_26_ );
dff P3_REG0_REG_26__reg ( clk, reset, P3_REG0_REG_26_, n1251 );
dff P3_REG2_REG_29__reg ( clk, reset, ex_wire267, n1586 );
not U_inv2373 ( n74862, ex_wire267 );
dff P3_REG1_REG_28__reg ( clk, reset, P3_REG1_REG_28_, n1421 );
not U_inv2374 ( n74813, P3_REG1_REG_28_ );
dff P3_REG0_REG_28__reg ( clk, reset, P3_REG0_REG_28_, n1261 );
dff P3_REG1_REG_27__reg ( clk, reset, P3_REG1_REG_27_, n1416 );
not U_inv2375 ( n74824, P3_REG1_REG_27_ );
dff P3_REG0_REG_27__reg ( clk, reset, P3_REG0_REG_27_, n1256 );
dff P3_REG2_REG_9__reg ( clk, reset, P3_REG2_REG_9_, n1486 );
not U_inv2376 ( n74384, P3_REG2_REG_9_ );
dff P3_ADDR_REG_9__reg ( clk, reset, ex_wire268, n1651 );
not U_inv2377 ( n73828, ex_wire268 );
dff P3_ADDR_REG_10__reg ( clk, reset, ex_wire269, n1646 );
not U_inv2378 ( n74041, ex_wire269 );
dff P3_ADDR_REG_14__reg ( clk, reset, ex_wire270, n1626 );
not U_inv2379 ( n74405, ex_wire270 );
dff P3_ADDR_REG_15__reg ( clk, reset, ex_wire271, n1621 );
not U_inv2380 ( n74441, ex_wire271 );
dff P3_ADDR_REG_16__reg ( clk, reset, ex_wire272, n1616 );
not U_inv2381 ( n74447, ex_wire272 );
dff P3_ADDR_REG_17__reg ( clk, reset, ex_wire273, n1611 );
not U_inv2382 ( n74489, ex_wire273 );
dff P3_ADDR_REG_18__reg ( clk, reset, ex_wire274, n1606 );
not U_inv2383 ( n74496, ex_wire274 );
dff P3_ADDR_REG_11__reg ( clk, reset, ex_wire275, n1641 );
not U_inv2384 ( n74279, ex_wire275 );
dff P3_ADDR_REG_12__reg ( clk, reset, ex_wire276, n1636 );
not U_inv2385 ( n74346, ex_wire276 );
dff P3_ADDR_REG_13__reg ( clk, reset, ex_wire277, n1631 );
not U_inv2386 ( n74389, ex_wire277 );
dff P1_P3_INSTADDRPOINTER_REG_1__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_1_, n4311 );
not U_inv2387 ( n75055, P1_P3_INSTADDRPOINTER_REG_1_ );
dff P1_P3_PHYADDRPOINTER_REG_1__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_1_, n4471 );
not U_inv2388 ( n74470, P1_P3_PHYADDRPOINTER_REG_1_ );
dff P1_P3_REIP_REG_1__reg ( clk, reset, P1_P3_REIP_REG_1_, n5266 );
not U_inv2389 ( n73164, P1_P3_REIP_REG_1_ );
dff P1_P3_BYTEENABLE_REG_0__reg ( clk, reset, P1_P3_BYTEENABLE_REG_0_, n5436 );
dff P1_P3_BYTEENABLE_REG_1__reg ( clk, reset, P1_P3_BYTEENABLE_REG_1_, n5431 );
dff P1_P3_BYTEENABLE_REG_2__reg ( clk, reset, P1_P3_BYTEENABLE_REG_2_, n5426 );
dff P1_P3_PHYADDRPOINTER_REG_2__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_2_, n4476 );
not U_inv2390 ( n74699, P1_P3_PHYADDRPOINTER_REG_2_ );
dff P1_P3_REIP_REG_2__reg ( clk, reset, P1_P3_REIP_REG_2_, n5271 );
not U_inv2391 ( n74622, P1_P3_REIP_REG_2_ );
dff P1_P3_INSTADDRPOINTER_REG_3__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_3_, n4321 );
not U_inv2392 ( n74412, P1_P3_INSTADDRPOINTER_REG_3_ );
dff P1_P3_PHYADDRPOINTER_REG_3__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_3_, n4481 );
not U_inv2393 ( n73082, P1_P3_PHYADDRPOINTER_REG_3_ );
dff P1_P3_REIP_REG_3__reg ( clk, reset, P1_P3_REIP_REG_3_, n5276 );
not U_inv2394 ( n73169, P1_P3_REIP_REG_3_ );
dff P1_P3_PHYADDRPOINTER_REG_4__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_4_, n4486 );
not U_inv2395 ( n74478, P1_P3_PHYADDRPOINTER_REG_4_ );
dff P1_P3_REIP_REG_4__reg ( clk, reset, P1_P3_REIP_REG_4_, n5281 );
not U_inv2396 ( n74643, P1_P3_REIP_REG_4_ );
dff P1_P3_INSTADDRPOINTER_REG_4__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_4_, n4326 );
not U_inv2397 ( n75940, P1_P3_INSTADDRPOINTER_REG_4_ );
dff P1_P3_PHYADDRPOINTER_REG_5__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_5_, n4491 );
not U_inv2398 ( n73093, P1_P3_PHYADDRPOINTER_REG_5_ );
dff P1_P3_REIP_REG_5__reg ( clk, reset, P1_P3_REIP_REG_5_, n5286 );
not U_inv2399 ( n73194, P1_P3_REIP_REG_5_ );
dff P1_P3_INSTADDRPOINTER_REG_5__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_5_, n4331 );
not U_inv2400 ( n74455, P1_P3_INSTADDRPOINTER_REG_5_ );
dff P1_P3_REIP_REG_6__reg ( clk, reset, ex_wire278, n5291 );
not U_inv2401 ( n74712, ex_wire278 );
dff P1_P3_INSTADDRPOINTER_REG_6__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_6_, n4336 );
not U_inv2402 ( n73088, P1_P3_INSTADDRPOINTER_REG_6_ );
dff P1_P3_PHYADDRPOINTER_REG_6__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_6_, n4496 );
not U_inv2403 ( n74503, P1_P3_PHYADDRPOINTER_REG_6_ );
dff P1_P3_INSTADDRPOINTER_REG_7__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_7_, n4341 );
not U_inv2404 ( n74696, P1_P3_INSTADDRPOINTER_REG_7_ );
dff P1_P3_PHYADDRPOINTER_REG_7__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_7_, n4501 );
not U_inv2405 ( n73102, P1_P3_PHYADDRPOINTER_REG_7_ );
dff P1_P3_REIP_REG_7__reg ( clk, reset, P1_P3_REIP_REG_7_, n5296 );
not U_inv2406 ( n72967, P1_P3_REIP_REG_7_ );
dff P1_P3_INSTADDRPOINTER_REG_8__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_8_, n4346 );
not U_inv2407 ( n73197, P1_P3_INSTADDRPOINTER_REG_8_ );
dff P1_P3_PHYADDRPOINTER_REG_8__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_8_, n4506 );
not U_inv2408 ( n74527, P1_P3_PHYADDRPOINTER_REG_8_ );
dff P1_P3_REIP_REG_8__reg ( clk, reset, P1_P3_REIP_REG_8_, n5301 );
not U_inv2409 ( n74750, P1_P3_REIP_REG_8_ );
dff P1_P3_PHYADDRPOINTER_REG_9__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_9_, n4511 );
not U_inv2410 ( n73112, P1_P3_PHYADDRPOINTER_REG_9_ );
dff P1_P3_REIP_REG_9__reg ( clk, reset, ex_wire279, n5306 );
not U_inv2411 ( n73217, ex_wire279 );
dff P1_P3_PHYADDRPOINTER_REG_10__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_10_, n4516 );
not U_inv2412 ( n74557, P1_P3_PHYADDRPOINTER_REG_10_ );
dff P1_P3_REIP_REG_10__reg ( clk, reset, P1_P3_REIP_REG_10_, n5311 );
not U_inv2413 ( n74746, P1_P3_REIP_REG_10_ );
dff P1_P3_INSTADDRPOINTER_REG_10__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_10_, n4356 );
not U_inv2414 ( n73115, P1_P3_INSTADDRPOINTER_REG_10_ );
dff P1_P3_PHYADDRPOINTER_REG_11__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_11_, n4521 );
not U_inv2415 ( n74465, P1_P3_PHYADDRPOINTER_REG_11_ );
dff P1_P3_REIP_REG_11__reg ( clk, reset, P1_P3_REIP_REG_11_, n5316 );
not U_inv2416 ( n74791, P1_P3_REIP_REG_11_ );
dff P1_P3_REIP_REG_12__reg ( clk, reset, ex_wire280, n5321 );
not U_inv2417 ( n74801, ex_wire280 );
dff P1_P3_INSTADDRPOINTER_REG_12__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_12_, n4366 );
not U_inv2418 ( n74458, P1_P3_INSTADDRPOINTER_REG_12_ );
dff P1_P3_PHYADDRPOINTER_REG_12__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_12_, n4526 );
not U_inv2419 ( n74615, P1_P3_PHYADDRPOINTER_REG_12_ );
dff P1_P3_PHYADDRPOINTER_REG_13__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_13_, n4531 );
dff P1_P3_REIP_REG_13__reg ( clk, reset, P1_P3_REIP_REG_13_, n5326 );
not U_inv2420 ( n73235, P1_P3_REIP_REG_13_ );
dff P1_P3_INSTADDRPOINTER_REG_14__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_14_, n4376 );
not U_inv2421 ( n73160, P1_P3_INSTADDRPOINTER_REG_14_ );
dff P1_P3_PHYADDRPOINTER_REG_14__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_14_, n4536 );
not U_inv2422 ( n74859, P1_P3_PHYADDRPOINTER_REG_14_ );
dff P1_P3_REIP_REG_14__reg ( clk, reset, P1_P3_REIP_REG_14_, n5331 );
not U_inv2423 ( n74829, P1_P3_REIP_REG_14_ );
dff P1_P3_REIP_REG_15__reg ( clk, reset, P1_P3_REIP_REG_15_, n5336 );
not U_inv2424 ( n74839, P1_P3_REIP_REG_15_ );
dff P1_P3_INSTADDRPOINTER_REG_15__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_15_, n4381 );
not U_inv2425 ( n74855, P1_P3_INSTADDRPOINTER_REG_15_ );
dff P1_P3_PHYADDRPOINTER_REG_15__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_15_, n4541 );
not U_inv2426 ( n75195, P1_P3_PHYADDRPOINTER_REG_15_ );
dff P1_P3_REIP_REG_16__reg ( clk, reset, P1_P3_REIP_REG_16_, n5341 );
not U_inv2427 ( n73250, P1_P3_REIP_REG_16_ );
dff P1_P3_PHYADDRPOINTER_REG_16__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_16_, n4546 );
dff P1_P3_REIP_REG_17__reg ( clk, reset, P1_P3_REIP_REG_17_, n5346 );
not U_inv2428 ( n74885, P1_P3_REIP_REG_17_ );
dff P1_P3_INSTADDRPOINTER_REG_17__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_17_, n4391 );
not U_inv2429 ( n74879, P1_P3_INSTADDRPOINTER_REG_17_ );
dff P1_P3_PHYADDRPOINTER_REG_17__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_17_, n4551 );
not U_inv2430 ( n74564, P1_P3_PHYADDRPOINTER_REG_17_ );
dff P1_P3_REIP_REG_18__reg ( clk, reset, P1_P3_REIP_REG_18_, n5351 );
not U_inv2431 ( n74901, P1_P3_REIP_REG_18_ );
dff P1_P3_INSTADDRPOINTER_REG_18__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_18_, n4396 );
not U_inv2432 ( n74635, P1_P3_INSTADDRPOINTER_REG_18_ );
dff P1_P3_PHYADDRPOINTER_REG_18__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_18_, n4556 );
not U_inv2433 ( n75191, P1_P3_PHYADDRPOINTER_REG_18_ );
dff P1_P3_REIP_REG_19__reg ( clk, reset, P1_P3_REIP_REG_19_, n5356 );
not U_inv2434 ( n73264, P1_P3_REIP_REG_19_ );
dff P1_P3_INSTADDRPOINTER_REG_19__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_19_, n4401 );
not U_inv2435 ( n74610, P1_P3_INSTADDRPOINTER_REG_19_ );
dff P1_P3_PHYADDRPOINTER_REG_19__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_19_, n4561 );
dff P1_P3_PHYADDRPOINTER_REG_20__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_20_, n4566 );
not U_inv2436 ( n74941, P1_P3_PHYADDRPOINTER_REG_20_ );
dff P1_P3_REIP_REG_20__reg ( clk, reset, P1_P3_REIP_REG_20_, n5361 );
not U_inv2437 ( n74929, P1_P3_REIP_REG_20_ );
dff P1_P3_INSTADDRPOINTER_REG_21__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_21_, n4411 );
not U_inv2438 ( n73167, P1_P3_INSTADDRPOINTER_REG_21_ );
dff P1_P3_PHYADDRPOINTER_REG_21__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_21_, n4571 );
not U_inv2439 ( n74688, P1_P3_PHYADDRPOINTER_REG_21_ );
dff P1_P3_REIP_REG_21__reg ( clk, reset, P1_P3_REIP_REG_21_, n5366 );
not U_inv2440 ( n74945, P1_P3_REIP_REG_21_ );
dff P1_P3_INSTADDRPOINTER_REG_22__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_22_, n4416 );
not U_inv2441 ( n74652, P1_P3_INSTADDRPOINTER_REG_22_ );
dff P1_P3_PHYADDRPOINTER_REG_22__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_22_, n4576 );
not U_inv2442 ( n75239, P1_P3_PHYADDRPOINTER_REG_22_ );
dff P1_P3_REIP_REG_22__reg ( clk, reset, P1_P3_REIP_REG_22_, n5371 );
not U_inv2443 ( n73278, P1_P3_REIP_REG_22_ );
dff P1_P3_INSTADDRPOINTER_REG_23__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_23_, n4421 );
not U_inv2444 ( n75050, P1_P3_INSTADDRPOINTER_REG_23_ );
dff P1_P3_PHYADDRPOINTER_REG_23__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_23_, n4581 );
not U_inv2445 ( n74752, P1_P3_PHYADDRPOINTER_REG_23_ );
dff P1_P3_REIP_REG_23__reg ( clk, reset, P1_P3_REIP_REG_23_, n5376 );
not U_inv2446 ( n74988, P1_P3_REIP_REG_23_ );
dff P1_P3_PHYADDRPOINTER_REG_24__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_24_, n4586 );
not U_inv2447 ( n75209, P1_P3_PHYADDRPOINTER_REG_24_ );
dff P1_P3_REIP_REG_24__reg ( clk, reset, P1_P3_REIP_REG_24_, n5381 );
not U_inv2448 ( n74994, P1_P3_REIP_REG_24_ );
dff P1_P3_REIP_REG_25__reg ( clk, reset, P1_P3_REIP_REG_25_, n5386 );
not U_inv2449 ( n73293, P1_P3_REIP_REG_25_ );
dff P1_P3_PHYADDRPOINTER_REG_25__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_25_, n4591 );
not U_inv2450 ( n74804, P1_P3_PHYADDRPOINTER_REG_25_ );
dff P1_P3_INSTADDRPOINTER_REG_26__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_26_, n4436 );
not U_inv2451 ( n74948, P1_P3_INSTADDRPOINTER_REG_26_ );
dff P1_P3_PHYADDRPOINTER_REG_26__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_26_, n4596 );
not U_inv2452 ( n75044, P1_P3_PHYADDRPOINTER_REG_26_ );
dff P1_P3_REIP_REG_26__reg ( clk, reset, P1_P3_REIP_REG_26_, n5391 );
not U_inv2453 ( n73297, P1_P3_REIP_REG_26_ );
dff P1_P3_REIP_REG_27__reg ( clk, reset, P1_P3_REIP_REG_27_, n5396 );
not U_inv2454 ( n75004, P1_P3_REIP_REG_27_ );
dff P1_P3_INSTADDRPOINTER_REG_28__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_28_, n4446 );
not U_inv2455 ( n74973, P1_P3_INSTADDRPOINTER_REG_28_ );
dff P1_P3_INSTADDRPOINTER_REG_29__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_29_, n4451 );
not U_inv2456 ( n75010, P1_P3_INSTADDRPOINTER_REG_29_ );
dff P1_P3_PHYADDRPOINTER_REG_29__reg ( clk, reset, P1_P3_PHYADDRPOINTER_REG_29_, n4611 );
not U_inv2457 ( n74912, P1_P3_PHYADDRPOINTER_REG_29_ );
dff P1_P3_REIP_REG_31__reg ( clk, reset, P1_P3_REIP_REG_31_, n5416 );
not U_inv2458 ( n75180, P1_P3_REIP_REG_31_ );
dff P1_P3_BE_N_REG_0__reg ( clk, reset, P1_P3_BE_N_REG_0_, n3266 );
dff P1_P3_BE_N_REG_1__reg ( clk, reset, P1_P3_BE_N_REG_1_, n3261 );
dff P1_P3_BE_N_REG_2__reg ( clk, reset, P1_P3_BE_N_REG_2_, n3256 );
dff P1_P3_ADDRESS_REG_0__reg ( clk, reset, P1_P3_ADDRESS_REG_0_, n3416 );
not U_inv2459 ( n73513, P1_P3_ADDRESS_REG_0_ );
dff P1_P3_ADDRESS_REG_1__reg ( clk, reset, P1_P3_ADDRESS_REG_1_, n3411 );
not U_inv2460 ( n73486, P1_P3_ADDRESS_REG_1_ );
dff P1_P3_ADDRESS_REG_2__reg ( clk, reset, P1_P3_ADDRESS_REG_2_, n3406 );
not U_inv2461 ( n73491, P1_P3_ADDRESS_REG_2_ );
dff P1_P3_ADDRESS_REG_3__reg ( clk, reset, P1_P3_ADDRESS_REG_3_, n3401 );
not U_inv2462 ( n73485, P1_P3_ADDRESS_REG_3_ );
dff P1_P3_ADDRESS_REG_4__reg ( clk, reset, P1_P3_ADDRESS_REG_4_, n3396 );
not U_inv2463 ( n73478, P1_P3_ADDRESS_REG_4_ );
dff P1_P3_ADDRESS_REG_5__reg ( clk, reset, P1_P3_ADDRESS_REG_5_, n3391 );
not U_inv2464 ( n73471, P1_P3_ADDRESS_REG_5_ );
dff P1_P3_ADDRESS_REG_6__reg ( clk, reset, P1_P3_ADDRESS_REG_6_, n3386 );
not U_inv2465 ( n73469, P1_P3_ADDRESS_REG_6_ );
dff P1_P3_ADDRESS_REG_7__reg ( clk, reset, P1_P3_ADDRESS_REG_7_, n3381 );
not U_inv2466 ( n73461, P1_P3_ADDRESS_REG_7_ );
dff P1_P3_ADDRESS_REG_8__reg ( clk, reset, P1_P3_ADDRESS_REG_8_, n3376 );
not U_inv2467 ( n73462, P1_P3_ADDRESS_REG_8_ );
dff P1_P3_ADDRESS_REG_9__reg ( clk, reset, P1_P3_ADDRESS_REG_9_, n3371 );
not U_inv2468 ( n73465, P1_P3_ADDRESS_REG_9_ );
dff P1_P3_ADDRESS_REG_10__reg ( clk, reset, P1_P3_ADDRESS_REG_10_, n3366 );
not U_inv2469 ( n73453, P1_P3_ADDRESS_REG_10_ );
dff P1_P3_ADDRESS_REG_11__reg ( clk, reset, P1_P3_ADDRESS_REG_11_, n3361 );
not U_inv2470 ( n73441, P1_P3_ADDRESS_REG_11_ );
dff P1_P3_ADDRESS_REG_12__reg ( clk, reset, P1_P3_ADDRESS_REG_12_, n3356 );
not U_inv2471 ( n73443, P1_P3_ADDRESS_REG_12_ );
dff P1_P3_ADDRESS_REG_13__reg ( clk, reset, P1_P3_ADDRESS_REG_13_, n3351 );
not U_inv2472 ( n73447, P1_P3_ADDRESS_REG_13_ );
dff P1_P3_ADDRESS_REG_14__reg ( clk, reset, P1_P3_ADDRESS_REG_14_, n3346 );
not U_inv2473 ( n73449, P1_P3_ADDRESS_REG_14_ );
dff P1_P3_ADDRESS_REG_15__reg ( clk, reset, P1_P3_ADDRESS_REG_15_, n3341 );
not U_inv2474 ( n73457, P1_P3_ADDRESS_REG_15_ );
dff P1_P3_ADDRESS_REG_16__reg ( clk, reset, P1_P3_ADDRESS_REG_16_, n3336 );
not U_inv2475 ( n73481, P1_P3_ADDRESS_REG_16_ );
dff P1_P3_ADDRESS_REG_17__reg ( clk, reset, P1_P3_ADDRESS_REG_17_, n3331 );
not U_inv2476 ( n73493, P1_P3_ADDRESS_REG_17_ );
dff P1_P3_ADDRESS_REG_18__reg ( clk, reset, P1_P3_ADDRESS_REG_18_, n3326 );
not U_inv2477 ( n73510, P1_P3_ADDRESS_REG_18_ );
dff P4_REG1_REG_14__reg ( clk, reset, P4_REG1_REG_14_, n2576 );
not U_inv2478 ( n74414, P4_REG1_REG_14_ );
dff P4_REG0_REG_14__reg ( clk, reset, P4_REG0_REG_14_, n2416 );
dff P4_REG2_REG_13__reg ( clk, reset, P4_REG2_REG_13_, n2731 );
not U_inv2479 ( n74402, P4_REG2_REG_13_ );
dff P4_REG1_REG_21__reg ( clk, reset, P4_REG1_REG_21_, n2611 );
not U_inv2480 ( n74545, P4_REG1_REG_21_ );
dff P4_REG0_REG_21__reg ( clk, reset, P4_REG0_REG_21_, n2451 );
dff P4_REG2_REG_20__reg ( clk, reset, ex_wire281, n2766 );
not U_inv2481 ( n74518, ex_wire281 );
dff P4_REG2_REG_19__reg ( clk, reset, ex_wire282, n2761 );
not U_inv2482 ( n74508, ex_wire282 );
dff P4_REG2_REG_18__reg ( clk, reset, ex_wire283, n2756 );
not U_inv2483 ( n74482, ex_wire283 );
dff P4_REG2_REG_16__reg ( clk, reset, P4_REG2_REG_16_, n2746 );
not U_inv2484 ( n74419, P4_REG2_REG_16_ );
dff P4_REG1_REG_15__reg ( clk, reset, P4_REG1_REG_15_, n2581 );
not U_inv2485 ( n74422, P4_REG1_REG_15_ );
dff P4_REG0_REG_15__reg ( clk, reset, P4_REG0_REG_15_, n2421 );
dff P4_REG2_REG_17__reg ( clk, reset, P4_REG2_REG_17_, n2751 );
not U_inv2486 ( n74456, P4_REG2_REG_17_ );
dff P4_REG1_REG_22__reg ( clk, reset, P4_REG1_REG_22_, n2616 );
not U_inv2487 ( n74530, P4_REG1_REG_22_ );
dff P4_REG0_REG_22__reg ( clk, reset, P4_REG0_REG_22_, n2456 );
dff P4_REG1_REG_23__reg ( clk, reset, P4_REG1_REG_23_, n2621 );
not U_inv2488 ( n74600, P4_REG1_REG_23_ );
dff P4_REG0_REG_23__reg ( clk, reset, P4_REG0_REG_23_, n2461 );
dff P4_REG1_REG_25__reg ( clk, reset, P4_REG1_REG_25_, n2631 );
not U_inv2489 ( n74706, P4_REG1_REG_25_ );
dff P4_REG0_REG_25__reg ( clk, reset, P4_REG0_REG_25_, n2471 );
dff P4_REG2_REG_24__reg ( clk, reset, ex_wire284, n2786 );
not U_inv2490 ( n74692, ex_wire284 );
dff P4_REG2_REG_29__reg ( clk, reset, ex_wire285, n2811 );
not U_inv2491 ( n74782, ex_wire285 );
dff P4_REG1_REG_28__reg ( clk, reset, P4_REG1_REG_28_, n2646 );
not U_inv2492 ( n74783, P4_REG1_REG_28_ );
dff P4_REG0_REG_28__reg ( clk, reset, P4_REG0_REG_28_, n2486 );
dff P4_REG1_REG_27__reg ( clk, reset, P4_REG1_REG_27_, n2641 );
not U_inv2493 ( n74781, P4_REG1_REG_27_ );
dff P4_REG0_REG_27__reg ( clk, reset, P4_REG0_REG_27_, n2481 );
dff P4_REG2_REG_26__reg ( clk, reset, ex_wire286, n2796 );
not U_inv2494 ( n74715, ex_wire286 );
dff P4_REG2_REG_12__reg ( clk, reset, P4_REG2_REG_12_, n2726 );
not U_inv2495 ( n74398, P4_REG2_REG_12_ );
dff P4_ADDR_REG_12__reg ( clk, reset, ex_wire287, n2861 );
not U_inv2496 ( n73442, ex_wire287 );
dff P4_ADDR_REG_13__reg ( clk, reset, ex_wire288, n2856 );
not U_inv2497 ( n73446, ex_wire288 );
dff P4_ADDR_REG_14__reg ( clk, reset, ex_wire289, n2851 );
not U_inv2498 ( n73448, ex_wire289 );
dff P4_ADDR_REG_15__reg ( clk, reset, ex_wire290, n2846 );
not U_inv2499 ( n73456, ex_wire290 );
dff P4_ADDR_REG_16__reg ( clk, reset, ex_wire291, n2841 );
not U_inv2500 ( n73480, ex_wire291 );
dff P4_ADDR_REG_17__reg ( clk, reset, ex_wire292, n2836 );
not U_inv2501 ( n73492, ex_wire292 );
dff P4_ADDR_REG_18__reg ( clk, reset, ex_wire293, n2831 );
not U_inv2502 ( n73509, ex_wire293 );
dff P2_P3_INSTADDRPOINTER_REG_1__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_1_, n11046 );
not U_inv2503 ( n75054, P2_P3_INSTADDRPOINTER_REG_1_ );
dff P2_P3_PHYADDRPOINTER_REG_1__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_1_, n11206 );
not U_inv2504 ( n74469, P2_P3_PHYADDRPOINTER_REG_1_ );
dff P2_P3_REIP_REG_1__reg ( clk, reset, P2_P3_REIP_REG_1_, n12001 );
not U_inv2505 ( n73163, P2_P3_REIP_REG_1_ );
dff P2_P3_PHYADDRPOINTER_REG_2__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_2_, n11211 );
not U_inv2506 ( n74700, P2_P3_PHYADDRPOINTER_REG_2_ );
dff P2_P3_REIP_REG_2__reg ( clk, reset, P2_P3_REIP_REG_2_, n12006 );
not U_inv2507 ( n74621, P2_P3_REIP_REG_2_ );
dff P2_P3_INSTADDRPOINTER_REG_3__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_3_, n11056 );
not U_inv2508 ( n74408, P2_P3_INSTADDRPOINTER_REG_3_ );
dff P2_P3_PHYADDRPOINTER_REG_3__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_3_, n11216 );
not U_inv2509 ( n73080, P2_P3_PHYADDRPOINTER_REG_3_ );
dff P2_P3_REIP_REG_3__reg ( clk, reset, P2_P3_REIP_REG_3_, n12011 );
not U_inv2510 ( n73168, P2_P3_REIP_REG_3_ );
dff P2_P3_PHYADDRPOINTER_REG_4__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_4_, n11221 );
not U_inv2511 ( n74479, P2_P3_PHYADDRPOINTER_REG_4_ );
dff P2_P3_REIP_REG_4__reg ( clk, reset, P2_P3_REIP_REG_4_, n12016 );
not U_inv2512 ( n74642, P2_P3_REIP_REG_4_ );
dff P2_P3_INSTADDRPOINTER_REG_4__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_4_, n11061 );
not U_inv2513 ( n75937, P2_P3_INSTADDRPOINTER_REG_4_ );
dff P2_P3_PHYADDRPOINTER_REG_5__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_5_, n11226 );
not U_inv2514 ( n73091, P2_P3_PHYADDRPOINTER_REG_5_ );
dff P2_P3_REIP_REG_5__reg ( clk, reset, P2_P3_REIP_REG_5_, n12021 );
not U_inv2515 ( n73193, P2_P3_REIP_REG_5_ );
dff P2_P3_INSTADDRPOINTER_REG_5__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_5_, n11066 );
not U_inv2516 ( n74452, P2_P3_INSTADDRPOINTER_REG_5_ );
dff P2_P3_REIP_REG_6__reg ( clk, reset, ex_wire294, n12026 );
not U_inv2517 ( n74711, ex_wire294 );
dff P2_P3_INSTADDRPOINTER_REG_6__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_6_, n11071 );
not U_inv2518 ( n73066, P2_P3_INSTADDRPOINTER_REG_6_ );
dff P2_P3_PHYADDRPOINTER_REG_6__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_6_, n11231 );
not U_inv2519 ( n74502, P2_P3_PHYADDRPOINTER_REG_6_ );
dff P2_P3_INSTADDRPOINTER_REG_7__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_7_, n11076 );
not U_inv2520 ( n74695, P2_P3_INSTADDRPOINTER_REG_7_ );
dff P2_P3_PHYADDRPOINTER_REG_7__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_7_, n11236 );
not U_inv2521 ( n73100, P2_P3_PHYADDRPOINTER_REG_7_ );
dff P2_P3_REIP_REG_7__reg ( clk, reset, P2_P3_REIP_REG_7_, n12031 );
not U_inv2522 ( n72966, P2_P3_REIP_REG_7_ );
dff P2_P3_PHYADDRPOINTER_REG_8__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_8_, n11241 );
not U_inv2523 ( n74526, P2_P3_PHYADDRPOINTER_REG_8_ );
dff P2_P3_REIP_REG_8__reg ( clk, reset, P2_P3_REIP_REG_8_, n12036 );
not U_inv2524 ( n74749, P2_P3_REIP_REG_8_ );
dff P2_P3_PHYADDRPOINTER_REG_9__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_9_, n11246 );
not U_inv2525 ( n73110, P2_P3_PHYADDRPOINTER_REG_9_ );
dff P2_P3_REIP_REG_9__reg ( clk, reset, ex_wire295, n12041 );
not U_inv2526 ( n73216, ex_wire295 );
dff P2_P3_PHYADDRPOINTER_REG_10__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_10_, n11251 );
not U_inv2527 ( n74558, P2_P3_PHYADDRPOINTER_REG_10_ );
dff P2_P3_REIP_REG_10__reg ( clk, reset, P2_P3_REIP_REG_10_, n12046 );
not U_inv2528 ( n74745, P2_P3_REIP_REG_10_ );
dff P2_P3_INSTADDRPOINTER_REG_10__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_10_, n11091 );
not U_inv2529 ( n74758, P2_P3_INSTADDRPOINTER_REG_10_ );
dff P2_P3_PHYADDRPOINTER_REG_11__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_11_, n11256 );
not U_inv2530 ( n74463, P2_P3_PHYADDRPOINTER_REG_11_ );
dff P2_P3_REIP_REG_11__reg ( clk, reset, P2_P3_REIP_REG_11_, n12051 );
not U_inv2531 ( n74790, P2_P3_REIP_REG_11_ );
dff P2_P3_REIP_REG_12__reg ( clk, reset, ex_wire296, n12056 );
not U_inv2532 ( n74800, ex_wire296 );
dff P2_P3_INSTADDRPOINTER_REG_12__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_12_, n11101 );
not U_inv2533 ( n74438, P2_P3_INSTADDRPOINTER_REG_12_ );
dff P2_P3_PHYADDRPOINTER_REG_12__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_12_, n11261 );
not U_inv2534 ( n74616, P2_P3_PHYADDRPOINTER_REG_12_ );
dff P2_P3_PHYADDRPOINTER_REG_13__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_13_, n11266 );
dff P2_P3_REIP_REG_13__reg ( clk, reset, P2_P3_REIP_REG_13_, n12061 );
not U_inv2535 ( n73236, P2_P3_REIP_REG_13_ );
dff P2_P3_REIP_REG_14__reg ( clk, reset, P2_P3_REIP_REG_14_, n12066 );
not U_inv2536 ( n74830, P2_P3_REIP_REG_14_ );
dff P2_P3_INSTADDRPOINTER_REG_14__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_14_, n11111 );
not U_inv2537 ( n74431, P2_P3_INSTADDRPOINTER_REG_14_ );
dff P2_P3_PHYADDRPOINTER_REG_14__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_14_, n11271 );
not U_inv2538 ( n74856, P2_P3_PHYADDRPOINTER_REG_14_ );
dff P2_P3_INSTADDRPOINTER_REG_15__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_15_, n11116 );
not U_inv2539 ( n74852, P2_P3_INSTADDRPOINTER_REG_15_ );
dff P2_P3_PHYADDRPOINTER_REG_15__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_15_, n11276 );
not U_inv2540 ( n75196, P2_P3_PHYADDRPOINTER_REG_15_ );
dff P2_P3_REIP_REG_15__reg ( clk, reset, P2_P3_REIP_REG_15_, n12071 );
not U_inv2541 ( n74840, P2_P3_REIP_REG_15_ );
dff P2_P3_REIP_REG_16__reg ( clk, reset, P2_P3_REIP_REG_16_, n12076 );
not U_inv2542 ( n73249, P2_P3_REIP_REG_16_ );
dff P2_P3_PHYADDRPOINTER_REG_16__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_16_, n11281 );
dff P2_P3_REIP_REG_17__reg ( clk, reset, P2_P3_REIP_REG_17_, n12081 );
not U_inv2543 ( n74884, P2_P3_REIP_REG_17_ );
dff P2_P3_INSTADDRPOINTER_REG_17__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_17_, n11126 );
not U_inv2544 ( n74872, P2_P3_INSTADDRPOINTER_REG_17_ );
dff P2_P3_PHYADDRPOINTER_REG_17__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_17_, n11286 );
not U_inv2545 ( n74563, P2_P3_PHYADDRPOINTER_REG_17_ );
dff P2_P3_REIP_REG_18__reg ( clk, reset, P2_P3_REIP_REG_18_, n12086 );
not U_inv2546 ( n74900, P2_P3_REIP_REG_18_ );
dff P2_P3_INSTADDRPOINTER_REG_18__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_18_, n11131 );
not U_inv2547 ( n74546, P2_P3_INSTADDRPOINTER_REG_18_ );
dff P2_P3_PHYADDRPOINTER_REG_18__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_18_, n11291 );
not U_inv2548 ( n75192, P2_P3_PHYADDRPOINTER_REG_18_ );
dff P2_P3_REIP_REG_19__reg ( clk, reset, P2_P3_REIP_REG_19_, n12091 );
not U_inv2549 ( n73263, P2_P3_REIP_REG_19_ );
dff P2_P3_INSTADDRPOINTER_REG_19__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_19_, n11136 );
not U_inv2550 ( n74574, P2_P3_INSTADDRPOINTER_REG_19_ );
dff P2_P3_PHYADDRPOINTER_REG_19__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_19_, n11296 );
dff P2_P3_PHYADDRPOINTER_REG_20__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_20_, n11301 );
not U_inv2551 ( n74940, P2_P3_PHYADDRPOINTER_REG_20_ );
dff P2_P3_REIP_REG_20__reg ( clk, reset, P2_P3_REIP_REG_20_, n12096 );
not U_inv2552 ( n74928, P2_P3_REIP_REG_20_ );
dff P2_P3_INSTADDRPOINTER_REG_21__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_21_, n11146 );
not U_inv2553 ( n73149, P2_P3_INSTADDRPOINTER_REG_21_ );
dff P2_P3_PHYADDRPOINTER_REG_21__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_21_, n11306 );
not U_inv2554 ( n74687, P2_P3_PHYADDRPOINTER_REG_21_ );
dff P2_P3_REIP_REG_21__reg ( clk, reset, P2_P3_REIP_REG_21_, n12101 );
not U_inv2555 ( n74944, P2_P3_REIP_REG_21_ );
dff P2_P3_INSTADDRPOINTER_REG_22__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_22_, n11151 );
not U_inv2556 ( n74595, P2_P3_INSTADDRPOINTER_REG_22_ );
dff P2_P3_PHYADDRPOINTER_REG_22__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_22_, n11311 );
not U_inv2557 ( n75240, P2_P3_PHYADDRPOINTER_REG_22_ );
dff P2_P3_REIP_REG_22__reg ( clk, reset, P2_P3_REIP_REG_22_, n12106 );
not U_inv2558 ( n73277, P2_P3_REIP_REG_22_ );
dff P2_P3_REIP_REG_23__reg ( clk, reset, P2_P3_REIP_REG_23_, n12111 );
not U_inv2559 ( n74987, P2_P3_REIP_REG_23_ );
dff P2_P3_INSTADDRPOINTER_REG_23__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_23_, n11156 );
not U_inv2560 ( n74637, P2_P3_INSTADDRPOINTER_REG_23_ );
dff P2_P3_PHYADDRPOINTER_REG_23__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_23_, n11316 );
not U_inv2561 ( n74751, P2_P3_PHYADDRPOINTER_REG_23_ );
dff P2_P3_REIP_REG_24__reg ( clk, reset, P2_P3_REIP_REG_24_, n12116 );
not U_inv2562 ( n74993, P2_P3_REIP_REG_24_ );
dff P2_P3_PHYADDRPOINTER_REG_24__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_24_, n11321 );
not U_inv2563 ( n75210, P2_P3_PHYADDRPOINTER_REG_24_ );
dff P2_P3_REIP_REG_25__reg ( clk, reset, P2_P3_REIP_REG_25_, n12121 );
not U_inv2564 ( n73292, P2_P3_REIP_REG_25_ );
dff P2_P3_PHYADDRPOINTER_REG_25__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_25_, n11326 );
not U_inv2565 ( n74805, P2_P3_PHYADDRPOINTER_REG_25_ );
dff P2_P3_INSTADDRPOINTER_REG_26__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_26_, n11171 );
not U_inv2566 ( n74947, P2_P3_INSTADDRPOINTER_REG_26_ );
dff P2_P3_PHYADDRPOINTER_REG_26__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_26_, n11331 );
not U_inv2567 ( n75045, P2_P3_PHYADDRPOINTER_REG_26_ );
dff P2_P3_REIP_REG_26__reg ( clk, reset, P2_P3_REIP_REG_26_, n12126 );
not U_inv2568 ( n73296, P2_P3_REIP_REG_26_ );
dff P2_P3_REIP_REG_27__reg ( clk, reset, P2_P3_REIP_REG_27_, n12131 );
not U_inv2569 ( n75003, P2_P3_REIP_REG_27_ );
dff P2_P3_INSTADDRPOINTER_REG_28__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_28_, n11181 );
not U_inv2570 ( n74976, P2_P3_INSTADDRPOINTER_REG_28_ );
dff P2_P3_INSTADDRPOINTER_REG_29__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_29_, n11186 );
not U_inv2571 ( n75009, P2_P3_INSTADDRPOINTER_REG_29_ );
dff P2_P3_PHYADDRPOINTER_REG_29__reg ( clk, reset, P2_P3_PHYADDRPOINTER_REG_29_, n11346 );
not U_inv2572 ( n74913, P2_P3_PHYADDRPOINTER_REG_29_ );
dff P2_P3_REIP_REG_31__reg ( clk, reset, P2_P3_REIP_REG_31_, n12151 );
not U_inv2573 ( n75179, P2_P3_REIP_REG_31_ );
dff P2_P3_DATAWIDTH_REG_31__reg ( clk, reset, ex_wire297, n10326 );
not U_inv2574 ( n75134, ex_wire297 );
dff P2_P3_DATAWIDTH_REG_30__reg ( clk, reset, ex_wire298, n10321 );
not U_inv2575 ( n73334, ex_wire298 );
dff P2_P3_DATAWIDTH_REG_29__reg ( clk, reset, ex_wire299, n10316 );
not U_inv2576 ( n73322, ex_wire299 );
dff P2_P3_DATAWIDTH_REG_28__reg ( clk, reset, ex_wire300, n10311 );
not U_inv2577 ( n75078, ex_wire300 );
dff P2_P3_DATAWIDTH_REG_27__reg ( clk, reset, ex_wire301, n10306 );
not U_inv2578 ( n73348, ex_wire301 );
dff P2_P3_DATAWIDTH_REG_26__reg ( clk, reset, ex_wire302, n10301 );
not U_inv2579 ( n75122, ex_wire302 );
dff P2_P3_DATAWIDTH_REG_25__reg ( clk, reset, ex_wire303, n10296 );
not U_inv2580 ( n73329, ex_wire303 );
dff P2_P3_DATAWIDTH_REG_24__reg ( clk, reset, ex_wire304, n10291 );
not U_inv2581 ( n75087, ex_wire304 );
dff P2_P3_DATAWIDTH_REG_23__reg ( clk, reset, ex_wire305, n10286 );
not U_inv2582 ( n73376, ex_wire305 );
dff P2_P3_DATAWIDTH_REG_22__reg ( clk, reset, ex_wire306, n10281 );
not U_inv2583 ( n75158, ex_wire306 );
dff P2_P3_DATAWIDTH_REG_21__reg ( clk, reset, ex_wire307, n10276 );
not U_inv2584 ( n73354, ex_wire307 );
dff P2_P3_DATAWIDTH_REG_20__reg ( clk, reset, ex_wire308, n10271 );
not U_inv2585 ( n75128, ex_wire308 );
dff P2_P3_DATAWIDTH_REG_19__reg ( clk, reset, ex_wire309, n10266 );
not U_inv2586 ( n73382, ex_wire309 );
dff P2_P3_DATAWIDTH_REG_18__reg ( clk, reset, ex_wire310, n10261 );
not U_inv2587 ( n75164, ex_wire310 );
dff P2_P3_DATAWIDTH_REG_17__reg ( clk, reset, ex_wire311, n10256 );
not U_inv2588 ( n73366, ex_wire311 );
dff P2_P3_DATAWIDTH_REG_16__reg ( clk, reset, ex_wire312, n10251 );
not U_inv2589 ( n75140, ex_wire312 );
dff P2_P3_DATAWIDTH_REG_15__reg ( clk, reset, ex_wire313, n10246 );
not U_inv2590 ( n73346, ex_wire313 );
dff P2_P3_DATAWIDTH_REG_14__reg ( clk, reset, ex_wire314, n10241 );
not U_inv2591 ( n75116, ex_wire314 );
dff P2_P3_DATAWIDTH_REG_13__reg ( clk, reset, ex_wire315, n10236 );
not U_inv2592 ( n73328, ex_wire315 );
dff P2_P3_DATAWIDTH_REG_12__reg ( clk, reset, ex_wire316, n10231 );
not U_inv2593 ( n75086, ex_wire316 );
dff P2_P3_DATAWIDTH_REG_11__reg ( clk, reset, ex_wire317, n10226 );
not U_inv2594 ( n73332, ex_wire317 );
dff P2_P3_DATAWIDTH_REG_10__reg ( clk, reset, ex_wire318, n10221 );
not U_inv2595 ( n75098, ex_wire318 );
dff P2_P3_DATAWIDTH_REG_9__reg ( clk, reset, ex_wire319, n10216 );
not U_inv2596 ( n73368, ex_wire319 );
dff P2_P3_DATAWIDTH_REG_8__reg ( clk, reset, ex_wire320, n10211 );
not U_inv2597 ( n75146, ex_wire320 );
dff P2_P3_DATAWIDTH_REG_7__reg ( clk, reset, ex_wire321, n10206 );
not U_inv2598 ( n73340, ex_wire321 );
dff P2_P3_DATAWIDTH_REG_6__reg ( clk, reset, ex_wire322, n10201 );
not U_inv2599 ( n75110, ex_wire322 );
dff P2_P3_DATAWIDTH_REG_5__reg ( clk, reset, ex_wire323, n10196 );
not U_inv2600 ( n73370, ex_wire323 );
dff P2_P3_DATAWIDTH_REG_4__reg ( clk, reset, ex_wire324, n10191 );
not U_inv2601 ( n75152, ex_wire324 );
dff P2_P3_DATAWIDTH_REG_3__reg ( clk, reset, ex_wire325, n10186 );
not U_inv2602 ( n73360, ex_wire325 );
dff P2_P3_DATAWIDTH_REG_2__reg ( clk, reset, ex_wire326, n10181 );
not U_inv2603 ( n75104, ex_wire326 );
dff P2_P3_DATAWIDTH_REG_1__reg ( clk, reset, P2_P3_DATAWIDTH_REG_1_, n10176 );
dff P2_P3_BYTEENABLE_REG_0__reg ( clk, reset, P2_P3_BYTEENABLE_REG_0_, n12171 );
dff P2_P3_BYTEENABLE_REG_1__reg ( clk, reset, P2_P3_BYTEENABLE_REG_1_, n12166 );
dff P2_P3_BYTEENABLE_REG_2__reg ( clk, reset, P2_P3_BYTEENABLE_REG_2_, n12161 );
dff P2_P3_BE_N_REG_1__reg ( clk, reset, P2_P3_BE_N_REG_1_, n9996 );
dff P2_P3_BE_N_REG_2__reg ( clk, reset, P2_P3_BE_N_REG_2_, n9991 );
dff P2_P3_M_IO_N_REG_reg ( clk, reset, P2_P3_M_IO_N_REG, n12206 );
dff P2_P3_D_C_N_REG_reg ( clk, reset, P2_P3_D_C_N_REG, n12201 );
dff P2_P3_W_R_N_REG_reg ( clk, reset, P2_P3_W_R_N_REG, n12176 );
dff P2_P3_BE_N_REG_0__reg ( clk, reset, P2_P3_BE_N_REG_0_, n10001 );
dff P2_P3_ADDRESS_REG_0__reg ( clk, reset, P2_P3_ADDRESS_REG_0_, n10151 );
not U_inv2604 ( n73434, P2_P3_ADDRESS_REG_0_ );
dff P2_P3_ADDRESS_REG_1__reg ( clk, reset, P2_P3_ADDRESS_REG_1_, n10146 );
not U_inv2605 ( n73438, P2_P3_ADDRESS_REG_1_ );
dff P2_P3_ADDRESS_REG_2__reg ( clk, reset, P2_P3_ADDRESS_REG_2_, n10141 );
not U_inv2606 ( n73439, P2_P3_ADDRESS_REG_2_ );
dff P2_P3_ADDRESS_REG_3__reg ( clk, reset, P2_P3_ADDRESS_REG_3_, n10136 );
not U_inv2607 ( n73474, P2_P3_ADDRESS_REG_3_ );
dff P2_P3_ADDRESS_REG_4__reg ( clk, reset, P2_P3_ADDRESS_REG_4_, n10131 );
not U_inv2608 ( n73487, P2_P3_ADDRESS_REG_4_ );
dff P2_P3_ADDRESS_REG_5__reg ( clk, reset, P2_P3_ADDRESS_REG_5_, n10126 );
not U_inv2609 ( n73500, P2_P3_ADDRESS_REG_5_ );
dff P2_P3_ADDRESS_REG_6__reg ( clk, reset, P2_P3_ADDRESS_REG_6_, n10121 );
not U_inv2610 ( n73522, P2_P3_ADDRESS_REG_6_ );
dff P2_P3_ADDRESS_REG_7__reg ( clk, reset, P2_P3_ADDRESS_REG_7_, n10116 );
not U_inv2611 ( n73530, P2_P3_ADDRESS_REG_7_ );
dff P2_P3_ADDRESS_REG_8__reg ( clk, reset, P2_P3_ADDRESS_REG_8_, n10111 );
not U_inv2612 ( n73544, P2_P3_ADDRESS_REG_8_ );
dff P2_P3_ADDRESS_REG_9__reg ( clk, reset, P2_P3_ADDRESS_REG_9_, n10106 );
not U_inv2613 ( n73824, P2_P3_ADDRESS_REG_9_ );
dff P2_P3_ADDRESS_REG_10__reg ( clk, reset, P2_P3_ADDRESS_REG_10_, n10101 );
not U_inv2614 ( n74020, P2_P3_ADDRESS_REG_10_ );
dff P2_P3_ADDRESS_REG_11__reg ( clk, reset, P2_P3_ADDRESS_REG_11_, n10096 );
not U_inv2615 ( n74274, P2_P3_ADDRESS_REG_11_ );
dff P2_P3_ADDRESS_REG_12__reg ( clk, reset, P2_P3_ADDRESS_REG_12_, n10091 );
not U_inv2616 ( n74342, P2_P3_ADDRESS_REG_12_ );
dff P2_P3_ADDRESS_REG_13__reg ( clk, reset, P2_P3_ADDRESS_REG_13_, n10086 );
not U_inv2617 ( n74388, P2_P3_ADDRESS_REG_13_ );
dff P2_P3_ADDRESS_REG_14__reg ( clk, reset, P2_P3_ADDRESS_REG_14_, n10081 );
not U_inv2618 ( n74403, P2_P3_ADDRESS_REG_14_ );
dff P2_P3_ADDRESS_REG_15__reg ( clk, reset, P2_P3_ADDRESS_REG_15_, n10076 );
not U_inv2619 ( n74437, P2_P3_ADDRESS_REG_15_ );
dff P2_P3_ADDRESS_REG_16__reg ( clk, reset, P2_P3_ADDRESS_REG_16_, n10071 );
not U_inv2620 ( n74446, P2_P3_ADDRESS_REG_16_ );
dff P2_P3_ADDRESS_REG_17__reg ( clk, reset, P2_P3_ADDRESS_REG_17_, n10066 );
not U_inv2621 ( n74486, P2_P3_ADDRESS_REG_17_ );
dff P2_P3_ADDRESS_REG_18__reg ( clk, reset, P2_P3_ADDRESS_REG_18_, n10061 );
not U_inv2622 ( n74495, P2_P3_ADDRESS_REG_18_ );
not U67951 ( n2040, n36481 );
dff P2_P3_INSTADDRPOINTER_REG_30__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_30_, n11191 );
not U_inv2623 ( n75039, P2_P3_INSTADDRPOINTER_REG_30_ );
dff P1_P3_INSTADDRPOINTER_REG_30__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_30_, n4456 );
not U_inv2624 ( n75042, P1_P3_INSTADDRPOINTER_REG_30_ );
dff P2_P2_INSTADDRPOINTER_REG_30__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_30_, n13436 );
not U_inv2625 ( n75040, P2_P2_INSTADDRPOINTER_REG_30_ );
dff P1_P2_INSTADDRPOINTER_REG_30__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_30_, n6701 );
not U_inv2626 ( n75038, P1_P2_INSTADDRPOINTER_REG_30_ );
dff P2_P1_INSTADDRPOINTER_REG_30__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_30_, n15681 );
not U_inv2627 ( n75016, P2_P1_INSTADDRPOINTER_REG_30_ );
dff P1_P1_INSTADDRPOINTER_REG_28__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_28_, n8936 );
not U_inv2628 ( n74946, P1_P1_INSTADDRPOINTER_REG_28_ );
dff P1_P1_INSTADDRPOINTER_REG_26__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_26_, n8926 );
not U_inv2629 ( n74886, P1_P1_INSTADDRPOINTER_REG_26_ );
dff P2_P1_INSTADDRPOINTER_REG_26__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_26_, n15661 );
not U_inv2630 ( n74919, P2_P1_INSTADDRPOINTER_REG_26_ );
dff P1_P1_INSTADDRPOINTER_REG_25__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_25_, n8921 );
not U_inv2631 ( n74774, P1_P1_INSTADDRPOINTER_REG_25_ );
dff P2_P2_INSTADDRPOINTER_REG_25__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_25_, n13411 );
not U_inv2632 ( n73225, P2_P2_INSTADDRPOINTER_REG_25_ );
dff P1_P2_INSTADDRPOINTER_REG_25__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_25_, n6676 );
not U_inv2633 ( n73224, P1_P2_INSTADDRPOINTER_REG_25_ );
dff P2_P3_INSTADDRPOINTER_REG_25__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_25_, n11166 );
not U_inv2634 ( n73223, P2_P3_INSTADDRPOINTER_REG_25_ );
dff P1_P3_INSTADDRPOINTER_REG_25__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_25_, n4431 );
not U_inv2635 ( n73232, P1_P3_INSTADDRPOINTER_REG_25_ );
dff P2_P1_INSTADDRPOINTER_REG_25__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_25_, n15656 );
not U_inv2636 ( n73220, P2_P1_INSTADDRPOINTER_REG_25_ );
dff P2_P2_INSTADDRPOINTER_REG_24__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_24_, n13406 );
not U_inv2637 ( n74918, P2_P2_INSTADDRPOINTER_REG_24_ );
dff P1_P2_INSTADDRPOINTER_REG_24__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_24_, n6671 );
not U_inv2638 ( n74917, P1_P2_INSTADDRPOINTER_REG_24_ );
dff P2_P3_INSTADDRPOINTER_REG_24__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_24_, n11161 );
not U_inv2639 ( n74916, P2_P3_INSTADDRPOINTER_REG_24_ );
dff P2_P1_INSTADDRPOINTER_REG_24__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_24_, n15651 );
not U_inv2640 ( n74881, P2_P1_INSTADDRPOINTER_REG_24_ );
dff P1_P1_INSTADDRPOINTER_REG_24__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_24_, n8916 );
not U_inv2641 ( n74653, P1_P1_INSTADDRPOINTER_REG_24_ );
dff P1_P3_INSTADDRPOINTER_REG_24__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_24_, n4426 );
not U_inv2642 ( n74671, P1_P3_INSTADDRPOINTER_REG_24_ );
dff P1_P1_INSTADDRPOINTER_REG_20__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_20_, n8896 );
not U_inv2643 ( n75053, P1_P1_INSTADDRPOINTER_REG_20_ );
dff P1_P1_STATE2_REG_2__reg ( clk, reset, P1_P1_STATE2_REG_2_, n8091 );
not U_inv2644 ( n73191, P1_P1_STATE2_REG_2_ );
dff P2_P1_STATE2_REG_2__reg ( clk, reset, P2_P1_STATE2_REG_2_, n14826 );
not U_inv2645 ( n73190, P2_P1_STATE2_REG_2_ );
dff P2_P1_STATE2_REG_1__reg ( clk, reset, P2_P1_STATE2_REG_1_, n14831 );
not U_inv2646 ( n74686, P2_P1_STATE2_REG_1_ );
dff P1_P1_STATE2_REG_1__reg ( clk, reset, P1_P1_STATE2_REG_1_, n8096 );
not U_inv2647 ( n74685, P1_P1_STATE2_REG_1_ );
dff P1_P3_INSTADDRPOINTER_REG_20__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_20_, n4406 );
not U_inv2648 ( n75060, P1_P3_INSTADDRPOINTER_REG_20_ );
dff P1_P1_STATE2_REG_0__reg ( clk, reset, P1_P1_STATE2_REG_0_, n8101 );
not U_inv2649 ( n74649, P1_P1_STATE2_REG_0_ );
dff P2_P1_STATE2_REG_0__reg ( clk, reset, P2_P1_STATE2_REG_0_, n14836 );
not U_inv2650 ( n74648, P2_P1_STATE2_REG_0_ );
dff P2_P3_STATE2_REG_2__reg ( clk, reset, P2_P3_STATE2_REG_2_, n10336 );
not U_inv2651 ( n74660, P2_P3_STATE2_REG_2_ );
dff P2_P2_STATE2_REG_2__reg ( clk, reset, P2_P2_STATE2_REG_2_, n12581 );
not U_inv2652 ( n74661, P2_P2_STATE2_REG_2_ );
dff P1_P2_STATE2_REG_2__reg ( clk, reset, P1_P2_STATE2_REG_2_, n5846 );
not U_inv2653 ( n74663, P1_P2_STATE2_REG_2_ );
dff P1_P3_STATE2_REG_2__reg ( clk, reset, P1_P3_STATE2_REG_2_, n3601 );
not U_inv2654 ( n74662, P1_P3_STATE2_REG_2_ );
dff P2_P3_STATE2_REG_1__reg ( clk, reset, P2_P3_STATE2_REG_1_, n10341 );
not U_inv2655 ( n73183, P2_P3_STATE2_REG_1_ );
dff P1_P2_STATE2_REG_1__reg ( clk, reset, P1_P2_STATE2_REG_1_, n5851 );
not U_inv2656 ( n73181, P1_P2_STATE2_REG_1_ );
dff P2_P2_STATE2_REG_1__reg ( clk, reset, P2_P2_STATE2_REG_1_, n12586 );
not U_inv2657 ( n73180, P2_P2_STATE2_REG_1_ );
dff P2_P2_INSTADDRPOINTER_REG_20__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_20_, n13386 );
not U_inv2658 ( n75019, P2_P2_INSTADDRPOINTER_REG_20_ );
dff P1_P2_INSTADDRPOINTER_REG_20__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_20_, n6651 );
not U_inv2659 ( n75018, P1_P2_INSTADDRPOINTER_REG_20_ );
dff P2_P3_INSTADDRPOINTER_REG_20__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_20_, n11141 );
not U_inv2660 ( n75017, P2_P3_INSTADDRPOINTER_REG_20_ );
dff P1_P3_STATE2_REG_1__reg ( clk, reset, P1_P3_STATE2_REG_1_, n3606 );
not U_inv2661 ( n73182, P1_P3_STATE2_REG_1_ );
dff P2_P1_INSTADDRPOINTER_REG_20__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_20_, n15631 );
not U_inv2662 ( n75020, P2_P1_INSTADDRPOINTER_REG_20_ );
dff P2_P1_EBX_REG_1__reg ( clk, reset, P2_P1_EBX_REG_1_, n16331 );
dff P1_P1_EBX_REG_1__reg ( clk, reset, P1_P1_EBX_REG_1_, n9596 );
dff P2_P2_INSTADDRPOINTER_REG_16__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_16_, n13366 );
not U_inv2663 ( n73132, P2_P2_INSTADDRPOINTER_REG_16_ );
dff P1_P2_INSTADDRPOINTER_REG_16__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_16_, n6631 );
not U_inv2664 ( n73131, P1_P2_INSTADDRPOINTER_REG_16_ );
dff P2_P3_INSTADDRPOINTER_REG_16__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_16_, n11121 );
not U_inv2665 ( n73130, P2_P3_INSTADDRPOINTER_REG_16_ );
dff P2_P2_EBX_REG_1__reg ( clk, reset, P2_P2_EBX_REG_1_, n14086 );
dff P2_P3_EBX_REG_1__reg ( clk, reset, P2_P3_EBX_REG_1_, n11841 );
dff P1_P2_EBX_REG_1__reg ( clk, reset, P1_P2_EBX_REG_1_, n7351 );
dff P1_P3_EBX_REG_1__reg ( clk, reset, P1_P3_EBX_REG_1_, n5106 );
dff P2_P1_INSTADDRPOINTER_REG_16__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_16_, n15611 );
not U_inv2666 ( n73118, P2_P1_INSTADDRPOINTER_REG_16_ );
dff P1_P1_INSTADDRPOINTER_REG_13__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_13_, n8861 );
not U_inv2667 ( n74468, P1_P1_INSTADDRPOINTER_REG_13_ );
dff P2_P3_STATE2_REG_0__reg ( clk, reset, P2_P3_STATE2_REG_0_, n10346 );
not U_inv2668 ( n74593, P2_P3_STATE2_REG_0_ );
dff P2_P2_STATE2_REG_0__reg ( clk, reset, P2_P2_STATE2_REG_0_, n12591 );
not U_inv2669 ( n74594, P2_P2_STATE2_REG_0_ );
dff P1_P2_STATE2_REG_0__reg ( clk, reset, P1_P2_STATE2_REG_0_, n5856 );
not U_inv2670 ( n74592, P1_P2_STATE2_REG_0_ );
dff P1_P3_STATE2_REG_0__reg ( clk, reset, P1_P3_STATE2_REG_0_, n3611 );
not U_inv2671 ( n74591, P1_P3_STATE2_REG_0_ );
dff P1_P1_INSTADDRPOINTER_REG_11__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_11_, n8851 );
not U_inv2672 ( n73116, P1_P1_INSTADDRPOINTER_REG_11_ );
dff P2_P1_INSTQUEUEWR_ADDR_REG_2__reg ( clk, reset, P2_P1_INSTQUEUEWR_ADDR_REG_2_, n15516 );
not U_inv2673 ( n73133, P2_P1_INSTQUEUEWR_ADDR_REG_2_ );
dff P1_P1_INSTQUEUEWR_ADDR_REG_2__reg ( clk, reset, P1_P1_INSTQUEUEWR_ADDR_REG_2_, n8781 );
not U_inv2674 ( n73134, P1_P1_INSTQUEUEWR_ADDR_REG_2_ );
dff P1_P1_INSTADDRPOINTER_REG_8__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_8_, n8836 );
not U_inv2675 ( n73176, P1_P1_INSTADDRPOINTER_REG_8_ );
dff P1_P3_INSTADDRPOINTER_REG_13__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_13_, n4371 );
not U_inv2676 ( n74460, P1_P3_INSTADDRPOINTER_REG_13_ );
dff P1_P1_INSTADDRPOINTER_REG_9__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_9_, n8841 );
not U_inv2677 ( n73109, P1_P1_INSTADDRPOINTER_REG_9_ );
dff P1_P3_INSTADDRPOINTER_REG_9__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_9_, n4351 );
not U_inv2678 ( n73114, P1_P3_INSTADDRPOINTER_REG_9_ );
dff P2_P2_INSTADDRPOINTER_REG_13__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_13_, n13351 );
not U_inv2679 ( n73106, P2_P2_INSTADDRPOINTER_REG_13_ );
dff P1_P2_INSTADDRPOINTER_REG_13__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_13_, n6616 );
not U_inv2680 ( n73105, P1_P2_INSTADDRPOINTER_REG_13_ );
dff P2_P3_INSTADDRPOINTER_REG_13__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_13_, n11106 );
not U_inv2681 ( n73104, P2_P3_INSTADDRPOINTER_REG_13_ );
dff P2_P1_INSTADDRPOINTER_REG_13__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_13_, n15596 );
not U_inv2682 ( n73099, P2_P1_INSTADDRPOINTER_REG_13_ );
dff P2_P2_INSTADDRPOINTER_REG_11__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_11_, n13341 );
not U_inv2683 ( n72952, P2_P2_INSTADDRPOINTER_REG_11_ );
dff P1_P2_INSTADDRPOINTER_REG_11__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_11_, n6606 );
not U_inv2684 ( n72951, P1_P2_INSTADDRPOINTER_REG_11_ );
dff P2_P3_INSTADDRPOINTER_REG_11__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_11_, n11096 );
not U_inv2685 ( n72950, P2_P3_INSTADDRPOINTER_REG_11_ );
dff P2_P1_INSTADDRPOINTER_REG_11__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_11_, n15586 );
not U_inv2686 ( n72948, P2_P1_INSTADDRPOINTER_REG_11_ );
dff P1_P3_INSTQUEUEWR_ADDR_REG_2__reg ( clk, reset, P1_P3_INSTQUEUEWR_ADDR_REG_2_, n4291 );
not U_inv2687 ( n74513, P1_P3_INSTQUEUEWR_ADDR_REG_2_ );
dff P2_P3_INSTQUEUEWR_ADDR_REG_2__reg ( clk, reset, P2_P3_INSTQUEUEWR_ADDR_REG_2_, n11026 );
not U_inv2688 ( n74514, P2_P3_INSTQUEUEWR_ADDR_REG_2_ );
dff P1_P2_INSTQUEUEWR_ADDR_REG_2__reg ( clk, reset, P1_P2_INSTQUEUEWR_ADDR_REG_2_, n6536 );
not U_inv2689 ( n74516, P1_P2_INSTQUEUEWR_ADDR_REG_2_ );
dff P2_P2_INSTQUEUEWR_ADDR_REG_2__reg ( clk, reset, P2_P2_INSTQUEUEWR_ADDR_REG_2_, n13271 );
not U_inv2690 ( n74517, P2_P2_INSTQUEUEWR_ADDR_REG_2_ );
dff P2_P2_INSTADDRPOINTER_REG_8__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_8_, n13326 );
not U_inv2691 ( n73189, P2_P2_INSTADDRPOINTER_REG_8_ );
dff P1_P2_INSTADDRPOINTER_REG_8__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_8_, n6591 );
not U_inv2692 ( n73188, P1_P2_INSTADDRPOINTER_REG_8_ );
dff P2_P3_INSTADDRPOINTER_REG_8__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_8_, n11081 );
not U_inv2693 ( n73187, P2_P3_INSTADDRPOINTER_REG_8_ );
dff P2_P1_INSTADDRPOINTER_REG_8__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_8_, n15571 );
not U_inv2694 ( n73178, P2_P1_INSTADDRPOINTER_REG_8_ );
dff P2_P2_INSTADDRPOINTER_REG_9__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_9_, n13331 );
not U_inv2695 ( n73086, P2_P2_INSTADDRPOINTER_REG_9_ );
dff P1_P2_INSTADDRPOINTER_REG_9__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_9_, n6596 );
not U_inv2696 ( n73085, P1_P2_INSTADDRPOINTER_REG_9_ );
dff P2_P3_INSTADDRPOINTER_REG_9__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_9_, n11086 );
not U_inv2697 ( n73084, P2_P3_INSTADDRPOINTER_REG_9_ );
dff P2_P1_INSTADDRPOINTER_REG_9__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_9_, n15576 );
not U_inv2698 ( n73078, P2_P1_INSTADDRPOINTER_REG_9_ );
dff P1_P1_INSTADDRPOINTER_REG_2__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_2_, n8806 );
not U_inv2699 ( n74579, P1_P1_INSTADDRPOINTER_REG_2_ );
dff P1_P3_INSTADDRPOINTER_REG_2__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_2_, n4316 );
not U_inv2700 ( n74588, P1_P3_INSTADDRPOINTER_REG_2_ );
dff P1_P1_INSTADDRPOINTER_REG_0__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_0_, n8796 );
not U_inv2701 ( n73079, P1_P1_INSTADDRPOINTER_REG_0_ );
dff P1_P3_INSTADDRPOINTER_REG_0__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_0_, n4306 );
not U_inv2702 ( n73077, P1_P3_INSTADDRPOINTER_REG_0_ );
dff P2_P2_INSTADDRPOINTER_REG_2__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_2_, n13296 );
not U_inv2703 ( n74590, P2_P2_INSTADDRPOINTER_REG_2_ );
dff P1_P2_INSTADDRPOINTER_REG_2__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_2_, n6561 );
not U_inv2704 ( n74589, P1_P2_INSTADDRPOINTER_REG_2_ );
dff P2_P3_INSTADDRPOINTER_REG_2__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_2_, n11051 );
not U_inv2705 ( n74587, P2_P3_INSTADDRPOINTER_REG_2_ );
dff P2_P1_INSTADDRPOINTER_REG_2__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_2_, n15541 );
not U_inv2706 ( n74580, P2_P1_INSTADDRPOINTER_REG_2_ );
dff P2_P3_INSTADDRPOINTER_REG_0__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_0_, n11041 );
not U_inv2707 ( n73076, P2_P3_INSTADDRPOINTER_REG_0_ );
dff P2_P2_INSTADDRPOINTER_REG_0__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_0_, n13286 );
not U_inv2708 ( n73074, P2_P2_INSTADDRPOINTER_REG_0_ );
dff P1_P2_INSTADDRPOINTER_REG_0__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_0_, n6551 );
not U_inv2709 ( n73075, P1_P2_INSTADDRPOINTER_REG_0_ );
dff P2_P1_INSTADDRPOINTER_REG_0__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_0_, n15531 );
not U_inv2710 ( n73071, P2_P1_INSTADDRPOINTER_REG_0_ );
dff P1_P1_INSTQUEUERD_ADDR_REG_1__reg ( clk, reset, P1_P1_INSTQUEUERD_ADDR_REG_1_, n8761 );
not U_inv2711 ( n73060, P1_P1_INSTQUEUERD_ADDR_REG_1_ );
dff P1_P1_INSTQUEUERD_ADDR_REG_3__reg ( clk, reset, P1_P1_INSTQUEUERD_ADDR_REG_3_, n8751 );
not U_inv2712 ( n73525, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
dff P1_P3_INSTQUEUERD_ADDR_REG_1__reg ( clk, reset, P1_P3_INSTQUEUERD_ADDR_REG_1_, n4271 );
not U_inv2713 ( n73059, P1_P3_INSTQUEUERD_ADDR_REG_1_ );
dff P1_P3_INSTQUEUERD_ADDR_REG_3__reg ( clk, reset, P1_P3_INSTQUEUERD_ADDR_REG_3_, n4261 );
not U_inv2714 ( n73524, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
dff P2_P2_INSTQUEUERD_ADDR_REG_1__reg ( clk, reset, P2_P2_INSTQUEUERD_ADDR_REG_1_, n13251 );
not U_inv2715 ( n73054, P2_P2_INSTQUEUERD_ADDR_REG_1_ );
dff P1_P2_INSTQUEUERD_ADDR_REG_1__reg ( clk, reset, P1_P2_INSTQUEUERD_ADDR_REG_1_, n6516 );
not U_inv2716 ( n73055, P1_P2_INSTQUEUERD_ADDR_REG_1_ );
dff P2_P3_INSTQUEUERD_ADDR_REG_1__reg ( clk, reset, P2_P3_INSTQUEUERD_ADDR_REG_1_, n11006 );
not U_inv2717 ( n73053, P2_P3_INSTQUEUERD_ADDR_REG_1_ );
dff P2_P1_INSTQUEUERD_ADDR_REG_1__reg ( clk, reset, P2_P1_INSTQUEUERD_ADDR_REG_1_, n15496 );
not U_inv2718 ( n73052, P2_P1_INSTQUEUERD_ADDR_REG_1_ );
dff P2_P2_INSTQUEUERD_ADDR_REG_3__reg ( clk, reset, P2_P2_INSTQUEUERD_ADDR_REG_3_, n13241 );
not U_inv2719 ( n73504, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
dff P1_P2_INSTQUEUERD_ADDR_REG_3__reg ( clk, reset, P1_P2_INSTQUEUERD_ADDR_REG_3_, n6506 );
not U_inv2720 ( n73503, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
dff P2_P3_INSTQUEUERD_ADDR_REG_3__reg ( clk, reset, P2_P3_INSTQUEUERD_ADDR_REG_3_, n10996 );
not U_inv2721 ( n73502, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
dff P2_P1_INSTQUEUERD_ADDR_REG_3__reg ( clk, reset, P2_P1_INSTQUEUERD_ADDR_REG_3_, n15486 );
not U_inv2722 ( n73497, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
dff P3_DATAO_REG_0__reg ( clk, reset, P3_DATAO_REG_0_, n1701 );
dff P4_DATAO_REG_0__reg ( clk, reset, P4_DATAO_REG_0_, n2926 );
not U_inv2723 ( n74955, P4_DATAO_REG_0_ );
dff P3_DATAO_REG_4__reg ( clk, reset, P3_DATAO_REG_4_, n1721 );
not U_inv2724 ( n73021, P3_DATAO_REG_4_ );
dff P3_DATAO_REG_5__reg ( clk, reset, P3_DATAO_REG_5_, n1726 );
not U_inv2725 ( n73421, P3_DATAO_REG_5_ );
dff P3_DATAO_REG_6__reg ( clk, reset, P3_DATAO_REG_6_, n1731 );
not U_inv2726 ( n73019, P3_DATAO_REG_6_ );
dff P4_DATAO_REG_5__reg ( clk, reset, P4_DATAO_REG_5_, n2951 );
not U_inv2727 ( n73020, P4_DATAO_REG_5_ );
dff P3_DATAO_REG_22__reg ( clk, reset, P3_DATAO_REG_22_, n1811 );
not U_inv2728 ( n73411, P3_DATAO_REG_22_ );
dff P4_DATAO_REG_6__reg ( clk, reset, P4_DATAO_REG_6_, n2956 );
not U_inv2729 ( n73420, P4_DATAO_REG_6_ );
dff P3_DATAO_REG_8__reg ( clk, reset, P3_DATAO_REG_8_, n1741 );
not U_inv2730 ( n73017, P3_DATAO_REG_8_ );
dff P3_DATAO_REG_9__reg ( clk, reset, P3_DATAO_REG_9_, n1746 );
not U_inv2731 ( n73413, P3_DATAO_REG_9_ );
dff P3_DATAO_REG_10__reg ( clk, reset, P3_DATAO_REG_10_, n1751 );
not U_inv2732 ( n73412, P3_DATAO_REG_10_ );
dff P3_DATAO_REG_12__reg ( clk, reset, P3_DATAO_REG_12_, n1761 );
not U_inv2733 ( n73410, P3_DATAO_REG_12_ );
dff P3_DATAO_REG_11__reg ( clk, reset, P3_DATAO_REG_11_, n1756 );
not U_inv2734 ( n73008, P3_DATAO_REG_11_ );
dff P4_DATAO_REG_8__reg ( clk, reset, P4_DATAO_REG_8_, n2966 );
not U_inv2735 ( n73418, P4_DATAO_REG_8_ );
dff P3_DATAO_REG_13__reg ( clk, reset, P3_DATAO_REG_13_, n1766 );
not U_inv2736 ( n73003, P3_DATAO_REG_13_ );
dff P3_DATAO_REG_16__reg ( clk, reset, P3_DATAO_REG_16_, n1781 );
not U_inv2737 ( n73397, P3_DATAO_REG_16_ );
dff P3_DATAO_REG_15__reg ( clk, reset, P3_DATAO_REG_15_, n1776 );
not U_inv2738 ( n72999, P3_DATAO_REG_15_ );
dff P4_DATAO_REG_18__reg ( clk, reset, P4_DATAO_REG_18_, n3016 );
not U_inv2739 ( n73007, P4_DATAO_REG_18_ );
dff P4_DATAO_REG_9__reg ( clk, reset, P4_DATAO_REG_9_, n2971 );
not U_inv2740 ( n73015, P4_DATAO_REG_9_ );
dff P4_DATAO_REG_10__reg ( clk, reset, P4_DATAO_REG_10_, n2976 );
not U_inv2741 ( n73414, P4_DATAO_REG_10_ );
dff P4_DATAO_REG_13__reg ( clk, reset, P4_DATAO_REG_13_, n2991 );
not U_inv2742 ( n73009, P4_DATAO_REG_13_ );
dff P4_DATAO_REG_12__reg ( clk, reset, P4_DATAO_REG_12_, n2986 );
not U_inv2743 ( n75913, P4_DATAO_REG_12_ );
dff P4_DATAO_REG_11__reg ( clk, reset, P4_DATAO_REG_11_, n2981 );
not U_inv2744 ( n73012, P4_DATAO_REG_11_ );
dff P4_DATAO_REG_16__reg ( clk, reset, P4_DATAO_REG_16_, n3006 );
not U_inv2745 ( n73406, P4_DATAO_REG_16_ );
dff P4_DATAO_REG_15__reg ( clk, reset, P4_DATAO_REG_15_, n3001 );
not U_inv2746 ( n75911, P4_DATAO_REG_15_ );
dff P2_P2_INSTADDRPOINTER_REG_27__reg ( clk, reset, P2_P2_INSTADDRPOINTER_REG_27_, n13421 );
not U_inv2747 ( n74963, P2_P2_INSTADDRPOINTER_REG_27_ );
dff P2_P3_INSTADDRPOINTER_REG_27__reg ( clk, reset, P2_P3_INSTADDRPOINTER_REG_27_, n11176 );
not U_inv2748 ( n74962, P2_P3_INSTADDRPOINTER_REG_27_ );
dff P1_P3_INSTADDRPOINTER_REG_27__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_27_, n4441 );
not U_inv2749 ( n74961, P1_P3_INSTADDRPOINTER_REG_27_ );
dff P1_P2_INSTADDRPOINTER_REG_27__reg ( clk, reset, P1_P2_INSTADDRPOINTER_REG_27_, n6686 );
not U_inv2750 ( n74960, P1_P2_INSTADDRPOINTER_REG_27_ );
dff P2_P1_INSTADDRPOINTER_REG_27__reg ( clk, reset, P2_P1_INSTADDRPOINTER_REG_27_, n15666 );
not U_inv2751 ( n74930, P2_P1_INSTADDRPOINTER_REG_27_ );
dff P1_P3_INSTADDRPOINTER_REG_16__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_16_, n4386 );
not U_inv2752 ( n74845, P1_P3_INSTADDRPOINTER_REG_16_ );
dff P1_P1_INSTADDRPOINTER_REG_16__reg ( clk, reset, P1_P1_INSTADDRPOINTER_REG_16_, n8876 );
not U_inv2753 ( n74818, P1_P1_INSTADDRPOINTER_REG_16_ );
dff P1_P3_INSTADDRPOINTER_REG_11__reg ( clk, reset, P1_P3_INSTADDRPOINTER_REG_11_, n4361 );
not U_inv2754 ( n74755, P1_P3_INSTADDRPOINTER_REG_11_ );
dff P2_P1_INSTQUEUEWR_ADDR_REG_0__reg ( clk, reset, P2_P1_INSTQUEUEWR_ADDR_REG_0_, n15526 );
not U_inv2755 ( n74442, P2_P1_INSTQUEUEWR_ADDR_REG_0_ );
dff P1_P1_INSTQUEUEWR_ADDR_REG_0__reg ( clk, reset, P1_P1_INSTQUEUEWR_ADDR_REG_0_, n8791 );
not U_inv2756 ( n74435, P1_P1_INSTQUEUEWR_ADDR_REG_0_ );
dff P1_P3_INSTQUEUEWR_ADDR_REG_0__reg ( clk, reset, P1_P3_INSTQUEUEWR_ADDR_REG_0_, n4301 );
not U_inv2757 ( n74426, P1_P3_INSTQUEUEWR_ADDR_REG_0_ );
dff P2_P3_INSTQUEUEWR_ADDR_REG_0__reg ( clk, reset, P2_P3_INSTQUEUEWR_ADDR_REG_0_, n11036 );
not U_inv2758 ( n74425, P2_P3_INSTQUEUEWR_ADDR_REG_0_ );
dff P2_P2_INSTQUEUEWR_ADDR_REG_0__reg ( clk, reset, P2_P2_INSTQUEUEWR_ADDR_REG_0_, n13281 );
not U_inv2759 ( n74424, P2_P2_INSTQUEUEWR_ADDR_REG_0_ );
dff P1_P2_INSTQUEUEWR_ADDR_REG_0__reg ( clk, reset, P1_P2_INSTQUEUEWR_ADDR_REG_0_, n6546 );
not U_inv2760 ( n74423, P1_P2_INSTQUEUEWR_ADDR_REG_0_ );
dff P1_P1_INSTQUEUERD_ADDR_REG_0__reg ( clk, reset, P1_P1_INSTQUEUERD_ADDR_REG_0_, n8766 );
not U_inv2761 ( n73533, P1_P1_INSTQUEUERD_ADDR_REG_0_ );
dff P1_P3_INSTQUEUERD_ADDR_REG_0__reg ( clk, reset, P1_P3_INSTQUEUERD_ADDR_REG_0_, n4276 );
not U_inv2762 ( n73532, P1_P3_INSTQUEUERD_ADDR_REG_0_ );
dff P1_P1_INSTQUEUERD_ADDR_REG_2__reg ( clk, reset, P1_P1_INSTQUEUERD_ADDR_REG_2_, n8756 );
not U_inv2763 ( n73527, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
dff P1_P3_INSTQUEUERD_ADDR_REG_2__reg ( clk, reset, P1_P3_INSTQUEUERD_ADDR_REG_2_, n4266 );
not U_inv2764 ( n73526, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
dff P2_P2_INSTQUEUERD_ADDR_REG_0__reg ( clk, reset, P2_P2_INSTQUEUERD_ADDR_REG_0_, n13256 );
not U_inv2765 ( n73521, P2_P2_INSTQUEUERD_ADDR_REG_0_ );
dff P1_P2_INSTQUEUERD_ADDR_REG_0__reg ( clk, reset, P1_P2_INSTQUEUERD_ADDR_REG_0_, n6521 );
not U_inv2766 ( n73520, P1_P2_INSTQUEUERD_ADDR_REG_0_ );
dff P2_P3_INSTQUEUERD_ADDR_REG_0__reg ( clk, reset, P2_P3_INSTQUEUERD_ADDR_REG_0_, n11011 );
not U_inv2767 ( n73518, P2_P3_INSTQUEUERD_ADDR_REG_0_ );
dff P2_P2_INSTQUEUERD_ADDR_REG_2__reg ( clk, reset, P2_P2_INSTQUEUERD_ADDR_REG_2_, n13246 );
not U_inv2768 ( n73517, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
dff P1_P2_INSTQUEUERD_ADDR_REG_2__reg ( clk, reset, P1_P2_INSTQUEUERD_ADDR_REG_2_, n6511 );
not U_inv2769 ( n73516, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
dff P2_P3_INSTQUEUERD_ADDR_REG_2__reg ( clk, reset, P2_P3_INSTQUEUERD_ADDR_REG_2_, n11001 );
not U_inv2770 ( n73515, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
dff P2_P1_INSTQUEUERD_ADDR_REG_0__reg ( clk, reset, P2_P1_INSTQUEUERD_ADDR_REG_0_, n15501 );
not U_inv2771 ( n73512, P2_P1_INSTQUEUERD_ADDR_REG_0_ );
dff P2_P1_INSTQUEUERD_ADDR_REG_2__reg ( clk, reset, P2_P1_INSTQUEUERD_ADDR_REG_2_, n15491 );
not U_inv2772 ( n73511, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
dff P3_DATAO_REG_2__reg ( clk, reset, P3_DATAO_REG_2_, n1711 );
not U_inv2773 ( n73426, P3_DATAO_REG_2_ );
dff P3_DATAO_REG_1__reg ( clk, reset, P3_DATAO_REG_1_, n1706 );
not U_inv2774 ( n73425, P3_DATAO_REG_1_ );
dff P3_DATAO_REG_3__reg ( clk, reset, P3_DATAO_REG_3_, n1716 );
not U_inv2775 ( n73424, P3_DATAO_REG_3_ );
dff P4_DATAO_REG_2__reg ( clk, reset, P4_DATAO_REG_2_, n2936 );
not U_inv2776 ( n73423, P4_DATAO_REG_2_ );
dff P4_DATAO_REG_1__reg ( clk, reset, P4_DATAO_REG_1_, n2931 );
not U_inv2777 ( n73422, P4_DATAO_REG_1_ );
dff P4_DATAO_REG_4__reg ( clk, reset, P4_DATAO_REG_4_, n2946 );
not U_inv2778 ( n75919, P4_DATAO_REG_4_ );
dff P3_DATAO_REG_7__reg ( clk, reset, P3_DATAO_REG_7_, n1736 );
not U_inv2779 ( n73419, P3_DATAO_REG_7_ );
dff P4_DATAO_REG_3__reg ( clk, reset, P4_DATAO_REG_3_, n2941 );
not U_inv2780 ( n73022, P4_DATAO_REG_3_ );
dff P4_DATAO_REG_7__reg ( clk, reset, P4_DATAO_REG_7_, n2961 );
not U_inv2781 ( n73018, P4_DATAO_REG_7_ );
dff P3_IR_REG_31__reg ( clk, reset, P3_IR_REG_31_, n956 );
dff P4_IR_REG_31__reg ( clk, reset, P4_IR_REG_31_, n2181 );
nand U72950 ( n50496, DIN_7_, n76930 );
nand U72951 ( n16966, DIN_7_, n76927 );
nand U72952 ( n17035, DIN_19_, n76928 );
nand U72953 ( n16943, DIN_3_, n76927 );
nand U72954 ( n17014, DIN_11_, n76928 );
nand U72955 ( n17525, DIN_10_, n76928 );
nand U72956 ( n17047, DIN_20_, n76928 );
nand U72957 ( n49898, DIN_3_, n76930 );
nand U72958 ( n49989, DIN_19_, n76929 );
nand U72959 ( n50320, DIN_11_, n76930 );
nand U72960 ( n50543, DIN_10_, n76930 );
nand U72961 ( n50001, DIN_20_, n76929 );
nand U72962 ( n50508, DIN_5_, n76929 );
nand U72963 ( n49982, DIN_17_, n76929 );
nand U72964 ( n17028, DIN_17_, n76928 );
nand U72965 ( n16861, DIN_15_, n76928 );
nand U72966 ( n49816, DIN_15_, n76930 );
nand U72967 ( n38866, n76804, n37303 );
xnor U72968 ( n31517, n73059, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
xnor U72969 ( n65767, n73053, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
xnor U72970 ( n57345, n73054, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
xnor U72971 ( n44902, n73052, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
xnor U72972 ( n24223, n73055, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
xnor U72973 ( n11194, n73060, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U72974 ( n48133, n47945, n73190 );
nand U72975 ( n61624, n839, n829 );
nand U72976 ( n61618, n67222, n842 );
nand U72977 ( n62272, n67224, n845 );
not U72978 ( n832, n61612 );
nand U72979 ( n14947, n14729, n73191 );
nand U72980 ( n38872, n2007, n2083 );
nand U72981 ( n38865, n40326, n37303 );
nor U72982 ( n38861, n37776, n2069 );
not U72983 ( n1239, n71327 );
nand U72984 ( n27124, n26965, n74663 );
xnor U72985 ( n27384, n26946, P1_P2_INSTQUEUEWR_ADDR_REG_2_ );
xnor U72986 ( n34629, n34191, P1_P3_INSTQUEUEWR_ADDR_REG_2_ );
nand U72987 ( n34369, n34210, n74662 );
xnor U72988 ( n15273, n14705, P1_P1_INSTQUEUEWR_ADDR_REG_2_ );
nand U72989 ( n69121, n68964, n74660 );
xnor U72990 ( n69375, n68945, P2_P3_INSTQUEUEWR_ADDR_REG_2_ );
xnor U72991 ( n48413, n47926, P2_P1_INSTQUEUEWR_ADDR_REG_2_ );
xnor U72992 ( n60532, n60086, P2_P2_INSTQUEUEWR_ADDR_REG_2_ );
nand U72993 ( n60268, n60105, n74661 );
not U72994 ( n593, n40826 );
not U72995 ( n833, n61613 );
not U72996 ( n2039, n38861 );
nand U72997 ( n37513, n40327, n37303 );
nand U72998 ( n38764, n40336, n2083 );
nand U72999 ( n38822, n2082, n37080 );
not U73000 ( n2033, n38764 );
not U73001 ( n1205, n71259 );
not U73002 ( n1222, n71096 );
xnor U73003 ( n63460, n66830, P2_P3_PHYADDRPOINTER_REG_19_ );
xor U73004 ( n63557, n6164, P2_P3_PHYADDRPOINTER_REG_15_ );
xnor U73005 ( n63616, n66950, P2_P3_PHYADDRPOINTER_REG_13_ );
xor U73006 ( n63731, n66989, n74463 );
xor U73007 ( n63775, n67057, n73110 );
xor U73008 ( n63827, n67099, n73100 );
xor U73009 ( n63887, n67138, n73091 );
nand U73010 ( n63953, n64984, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
xor U73011 ( n63940, n67166, n73080 );
xnor U73012 ( n29557, n32184, P1_P3_PHYADDRPOINTER_REG_19_ );
xor U73013 ( n29658, n3549, P1_P3_PHYADDRPOINTER_REG_15_ );
xnor U73014 ( n29717, n32311, P1_P3_PHYADDRPOINTER_REG_13_ );
xor U73015 ( n29771, n32350, n74465 );
xor U73016 ( n29815, n32394, n73112 );
xor U73017 ( n29871, n32443, n73102 );
xor U73018 ( n29931, n32482, n73093 );
nand U73019 ( n29997, n30782, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
xor U73020 ( n29984, n32510, n73082 );
xor U73021 ( n8637, P1_P1_PHYADDRPOINTER_REG_23_, n11993 );
xor U73022 ( n8708, P1_P1_PHYADDRPOINTER_REG_21_, n5307 );
xor U73023 ( n8884, P1_P1_PHYADDRPOINTER_REG_15_, n5297 );
xnor U73024 ( n8958, n12327, P1_P1_PHYADDRPOINTER_REG_13_ );
xor U73025 ( n9025, n12375, n74450 );
xor U73026 ( n9080, n12437, n73107 );
xor U73027 ( n9145, n12489, n73097 );
nand U73028 ( n9303, n10273, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
xor U73029 ( n42764, P2_P1_PHYADDRPOINTER_REG_21_, n7962 );
xor U73030 ( n42905, P2_P1_PHYADDRPOINTER_REG_15_, n7952 );
xnor U73031 ( n42978, n46010, P2_P1_PHYADDRPOINTER_REG_13_ );
xor U73032 ( n43032, n46049, n74451 );
xor U73033 ( n43076, n46093, n73108 );
xor U73034 ( n43128, n46135, n73098 );
nand U73035 ( n43268, n44142, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
xor U73036 ( n42582, P2_P1_PHYADDRPOINTER_REG_27_, n45640 );
xor U73037 ( n42628, P2_P1_PHYADDRPOINTER_REG_25_, n45694 );
xor U73038 ( n42703, P2_P1_PHYADDRPOINTER_REG_23_, n45727 );
xnor U73039 ( n42808, n45879, P2_P1_PHYADDRPOINTER_REG_19_ );
xor U73040 ( n42863, n45894, n74515 );
xnor U73041 ( n22396, n25074, P1_P2_PHYADDRPOINTER_REG_13_ );
xor U73042 ( n22548, n25201, n73103 );
xor U73043 ( n22661, n25268, n73083 );
xnor U73044 ( n22240, n24954, P1_P2_PHYADDRPOINTER_REG_19_ );
xor U73045 ( n22337, n4387, P1_P2_PHYADDRPOINTER_REG_15_ );
xor U73046 ( n22450, n25113, n74466 );
xor U73047 ( n22496, n25157, n73113 );
xor U73048 ( n22608, n25240, n73094 );
nand U73049 ( n22674, n23475, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
xnor U73050 ( n55508, n58209, P2_P2_PHYADDRPOINTER_REG_13_ );
xor U73051 ( n55661, n58337, n73101 );
nand U73052 ( n55787, n56597, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U73053 ( n34735, n35515, P1_BUF2_REG_25_ );
nand U73054 ( n34771, n35515, P1_BUF2_REG_29_ );
nand U73055 ( n34780, n35515, P1_BUF2_REG_30_ );
nand U73056 ( n34796, n35515, P1_BUF2_REG_31_ );
not U73057 ( n85, n27125 );
not U73058 ( n65, n27037 );
nand U73059 ( n34753, n35515, P1_BUF2_REG_27_ );
not U73060 ( n74, n27073 );
nand U73061 ( n34762, n35515, P1_BUF2_REG_28_ );
not U73062 ( n77, n27084 );
nand U73063 ( n34724, n35515, P1_BUF2_REG_24_ );
nand U73064 ( n28127, n28196, n26934 );
not U73065 ( n71, n27062 );
nand U73066 ( n27642, n27467, n27379 );
nand U73067 ( n15317, n16450, n10114 );
nand U73068 ( n14858, n16450, n10628 );
nand U73069 ( n15328, n16450, n10058 );
nand U73070 ( n14872, n16450, n10573 );
not U73071 ( n80, n27095 );
nand U73072 ( n15357, n16450, n9954 );
nand U73073 ( n14899, n16450, n10467 );
nand U73074 ( n15290, n16450, n10235 );
nand U73075 ( n14829, n16450, n10694 );
nand U73076 ( n16240, n16225, n15058 );
nand U73077 ( n16038, n15809, n15278 );
nand U73078 ( n15930, n15809, n15167 );
nand U73079 ( n15825, n15809, n15058 );
nand U73080 ( n15613, n15395, n15278 );
nand U73081 ( n69479, n70243, P2_BUF2_REG_25_ );
nand U73082 ( n69497, n70243, P2_BUF2_REG_27_ );
nand U73083 ( n69524, n70243, P2_BUF2_REG_30_ );
nand U73084 ( n69540, n70243, P2_BUF2_REG_31_ );
nand U73085 ( n69515, n70243, P2_BUF2_REG_29_ );
not U73086 ( n344, n60239 );
not U73087 ( n348, n60250 );
not U73088 ( n329, n60192 );
not U73089 ( n325, n60178 );
not U73090 ( n333, n60203 );
nand U73091 ( n69506, n70243, P2_BUF2_REG_28_ );
not U73092 ( n340, n60225 );
nand U73093 ( n48465, n49451, n44019 );
nand U73094 ( n48054, n49451, n44440 );
nand U73095 ( n69468, n70243, P2_BUF2_REG_24_ );
nand U73096 ( n48428, n49451, n44112 );
nand U73097 ( n48031, n49451, n44493 );
nand U73098 ( n48440, n49451, n44065 );
nand U73099 ( n48043, n49451, n44482 );
nand U73100 ( n49279, n49251, n48237 );
nand U73101 ( n48994, n48882, n48319 );
nand U73102 ( n48895, n48882, n48237 );
nand U73103 ( n48474, n49451, n43974 );
nand U73104 ( n48065, n49451, n44382 );
nand U73105 ( n48492, n49451, n43845 );
nand U73106 ( n48101, n49451, n44297 );
not U73107 ( n337, n60214 );
nand U73108 ( n61282, n61360, n60074 );
nand U73109 ( n60795, n60616, n60527 );
nand U73110 ( n48722, n48522, n48417 );
nand U73111 ( n49089, n48882, n48417 );
nand U73112 ( n48136, n49451, n44210 );
nand U73113 ( n48139, n76325, n45424 );
nand U73114 ( n15305, n16450, n10177 );
nand U73115 ( n14844, n16450, n10680 );
not U73116 ( n68, n27051 );
xor U73117 ( n28913, n28914, n28643 );
not U73118 ( n83, n27106 );
nand U73119 ( n69488, n70243, P2_BUF2_REG_26_ );
nand U73120 ( n48483, n49451, n43893 );
nand U73121 ( n49357, n49251, n48319 );
nand U73122 ( n48090, n49451, n44305 );
nand U73123 ( n49450, n49251, n48417 );
nand U73124 ( n48112, n49451, n44253 );
nand U73125 ( n34744, n35515, P1_BUF2_REG_26_ );
nand U73126 ( n15339, n16450, n9970 );
nand U73127 ( n16345, n16225, n15167 );
nand U73128 ( n14885, n16450, n10477 );
nand U73129 ( n15368, n16450, n9893 );
nand U73130 ( n14913, n16450, n10412 );
xor U73131 ( n62218, n62219, n61948 );
xor U73132 ( n36092, n36093, n35822 );
xor U73133 ( n8515, P1_P1_PHYADDRPOINTER_REG_27_, n11865 );
xor U73134 ( n8573, P1_P1_PHYADDRPOINTER_REG_25_, n11928 );
xnor U73135 ( n8763, n12165, P1_P1_PHYADDRPOINTER_REG_19_ );
xnor U73136 ( n55352, n58089, P2_P2_PHYADDRPOINTER_REG_19_ );
xor U73137 ( n55449, n7019, P2_P2_PHYADDRPOINTER_REG_15_ );
xor U73138 ( n55565, n58251, n74464 );
xor U73139 ( n55609, n58295, n73111 );
xor U73140 ( n55721, n58376, n73092 );
xor U73141 ( n55774, n58404, n73081 );
not U73142 ( n350, n60269 );
xor U73143 ( n54590, n54591, n54320 );
xor U73144 ( n43188, n46174, n73089 );
xor U73145 ( n43255, n46202, n73073 );
nor U73146 ( n45754, n41472, n45363 );
nand U73147 ( n61443, n76010, n842 );
nand U73148 ( n41487, n67224, n41908 );
nand U73149 ( n36167, P1_P3_STATE_REG_2_, n76501 );
xor U73150 ( n21607, n21608, n21337 );
xor U73151 ( n9220, n12537, n73087 );
xor U73152 ( n9287, n12573, n73072 );
nand U73153 ( n14950, n16450, n10358 );
nand U73154 ( n16449, n16225, n15278 );
nand U73155 ( n14954, n76591, n11638 );
xor U73156 ( n70818, n70819, n70548 );
nand U73157 ( n70876, P2_P3_STATE_REG_2_, n76647 );
not U73158 ( n1218, n71098 );
nand U73159 ( n27133, n76518, n24559 );
nand U73160 ( n27043, n76517, n24531 );
nand U73161 ( n27099, n76518, n24551 );
nand U73162 ( n34287, n76461, P1_BUF2_REG_0_ );
nand U73163 ( n27110, n76518, n24555 );
nand U73164 ( n60243, n76260, n57682 );
nand U73165 ( n60184, n76259, n57659 );
nand U73166 ( n69039, n76193, P2_BUF2_REG_0_ );
nand U73167 ( n49276, n49244, n47908 );
nand U73168 ( n48892, n48982, n47908 );
nand U73169 ( n48531, n48515, n47908 );
nand U73170 ( n60254, n76260, n57686 );
nand U73171 ( n60277, n76260, n57690 );
nand U73172 ( n31646, P1_P3_STATE2_REG_0_, n31619 );
nand U73173 ( n24390, P1_P2_STATE2_REG_0_, n24323 );
nand U73174 ( n57515, P2_P2_STATE2_REG_0_, n57446 );
nand U73175 ( n45111, P2_P1_STATE2_REG_0_, n45317 );
buf U73176 ( n76555, n75707 );
buf U73177 ( n76645, n75709 );
buf U73178 ( n76301, n75706 );
nand U73179 ( n28291, n28111, n27379 );
nand U73180 ( n11410, P1_P1_STATE2_REG_0_, n11494 );
nand U73181 ( n66054, P2_P3_STATE2_REG_0_, n65905 );
nand U73182 ( n61513, n61266, n60527 );
buf U73183 ( n76373, n75708 );
and U73184 ( n75011, n70842, n70843 );
and U73185 ( n75027, n36122, n36123 );
and U73186 ( n75029, n62405, n62406 );
and U73187 ( n75047, n21639, n21640 );
and U73188 ( n75048, n54661, n54662 );
and U73189 ( n75049, n28949, n28950 );
buf U73190 ( n76366, n75713 );
buf U73191 ( n76492, n75711 );
buf U73192 ( n76545, n75715 );
buf U73193 ( n76225, n75712 );
buf U73194 ( n76287, n75716 );
buf U73195 ( n76636, n75714 );
buf U73196 ( n76365, n75713 );
buf U73197 ( n76491, n75711 );
buf U73198 ( n76224, n75712 );
buf U73199 ( n76544, n75715 );
buf U73200 ( n76286, n75716 );
buf U73201 ( n76635, n75714 );
buf U73202 ( n76843, n615 );
buf U73203 ( n76824, n2023 );
buf U73204 ( n76343, n75700 );
buf U73205 ( n76199, n75701 );
buf U73206 ( n76523, n75702 );
buf U73207 ( n76265, n75703 );
buf U73208 ( n76473, n75704 );
buf U73209 ( n76604, n76601 );
buf U73210 ( n76853, n570 );
buf U73211 ( n76216, n75757 );
buf U73212 ( n76483, n75758 );
buf U73213 ( n76540, n75756 );
buf U73214 ( n76282, n75755 );
buf U73215 ( n76614, n11508 );
buf U73216 ( n76528, n24466 );
buf U73217 ( n76270, n57595 );
buf U73218 ( n76204, n66168 );
buf U73219 ( n76348, n45328 );
buf U73220 ( n76627, n75759 );
buf U73221 ( n76799, n2065 );
buf U73222 ( n76390, n75765 );
buf U73223 ( n76459, n75766 );
and U73224 ( n75700, n7564, n46277 );
and U73225 ( n75701, n5777, n67338 );
and U73226 ( n75702, n4018, n25331 );
and U73227 ( n75703, n6650, n58470 );
and U73228 ( n75704, n3178, n32573 );
buf U73229 ( n76601, n12218 );
not U73230 ( n568, n54923 );
buf U73231 ( n76337, n45748 );
buf U73232 ( n76290, n76291 );
buf U73233 ( n76289, n76291 );
not U73234 ( n2002, n37100 );
buf U73235 ( n76423, n75774 );
buf U73236 ( n76424, n75774 );
buf U73237 ( n76375, n76377 );
buf U73238 ( n76450, n76452 );
buf U73239 ( n76408, n75777 );
buf U73240 ( n76485, n30427 );
buf U73241 ( n76218, n64586 );
buf U73242 ( n76359, n43743 );
buf U73243 ( n76629, n9827 );
buf U73244 ( n76396, n40471 );
buf U73245 ( n76392, n40477 );
nand U73246 ( n38956, n40327, n2042 );
nor U73247 ( n37266, n1928, n36286 );
nor U73248 ( n37500, n36572, n1975 );
nor U73249 ( n39495, n2175, n1982 );
buf U73250 ( n76381, n75705 );
not U73251 ( n76385, n76387 );
nor U73252 ( n62465, n40913, n76387 );
nor U73253 ( n37402, n2113, n2183 );
nand U73254 ( n40708, n41446, n41447 );
buf U73255 ( n76740, n4760 );
buf U73256 ( n76673, n7405 );
buf U73257 ( n76437, n38146 );
buf U73258 ( n76441, n38129 );
buf U73259 ( n76445, n38127 );
nor U73260 ( n61612, n42291, n67217 );
nor U73261 ( n61613, n42291, n842 );
buf U73262 ( n76257, n76258 );
buf U73263 ( n76256, n76258 );
buf U73264 ( n76454, n76453 );
buf U73265 ( n76455, n76453 );
buf U73266 ( n76427, n76428 );
buf U73267 ( n76426, n76428 );
nand U73268 ( n38604, n2082, n2153 );
buf U73269 ( n76346, n45532 );
buf U73270 ( n76480, n31833 );
buf U73271 ( n76526, n24619 );
buf U73272 ( n76202, n66456 );
buf U73273 ( n76268, n57751 );
buf U73274 ( n76607, n11762 );
nand U73275 ( n28208, n27952, n27462 );
nand U73276 ( n61372, n61105, n60611 );
nand U73277 ( n27887, n27952, n27127 );
nand U73278 ( n61034, n61105, n60271 );
nand U73279 ( n28045, n27792, n27462 );
nand U73280 ( n61204, n60940, n60611 );
nand U73281 ( n27720, n27792, n27127 );
nand U73282 ( n60871, n60940, n60271 );
nor U73283 ( n35514, n34213, n3430 );
nor U73284 ( n70242, n68967, n6045 );
nand U73285 ( n27566, n27296, n27462 );
nand U73286 ( n60716, n60439, n60611 );
nand U73287 ( n15184, n14953, n15278 );
nand U73288 ( n14973, n15058, n14953 );
nand U73289 ( n48154, n48237, n48138 );
nand U73290 ( n48349, n48138, n48417 );
nand U73291 ( n15410, n15058, n15395 );
nand U73292 ( n48534, n48237, n48522 );
nand U73293 ( n27311, n27136, n27379 );
nand U73294 ( n60454, n60280, n60527 );
nand U73295 ( n27147, n27214, n27136 );
nand U73296 ( n60289, n60359, n60280 );
buf U73297 ( n76591, n14747 );
buf U73298 ( n76325, n47970 );
nand U73299 ( n28128, n28112, n4295 );
nand U73300 ( n61283, n61267, n6928 );
buf U73301 ( n76231, n75011 );
buf U73302 ( n76498, n75027 );
buf U73303 ( n76297, n75029 );
buf U73304 ( n76369, n75048 );
buf U73305 ( n76641, n75047 );
buf U73306 ( n76551, n75049 );
and U73307 ( n71265, n76043, n71274 );
buf U73308 ( n76247, n61294 );
or U73309 ( n61295, n67248, n783 );
buf U73310 ( n76240, n61595 );
buf U73311 ( n76251, n61291 );
buf U73312 ( n76413, n38756 );
buf U73313 ( n76402, n38843 );
or U73314 ( n38757, n40353, n2195 );
buf U73315 ( n76417, n38753 );
and U73316 ( n71247, n72692, n72693 );
nor U73317 ( n37273, n2160, n36655 );
buf U73318 ( n76835, n76833 );
buf U73319 ( n76790, n76792 );
buf U73320 ( n76836, n76838 );
and U73321 ( n71196, n72820, n72821 );
nor U73322 ( n42049, n41323, n700 );
buf U73323 ( n76387, n76384 );
buf U73324 ( n76388, n76384 );
and U73325 ( n75705, n829, n41908 );
nand U73326 ( n61617, n67223, n41908 );
nand U73327 ( n38875, n40324, n76804 );
buf U73328 ( n76453, n36287 );
buf U73329 ( n76547, n21935 );
buf U73330 ( n76494, n29252 );
buf U73331 ( n76227, n63019 );
buf U73332 ( n76293, n55047 );
buf U73333 ( n76226, n63019 );
buf U73334 ( n76493, n29252 );
buf U73335 ( n76546, n21935 );
buf U73336 ( n76292, n55047 );
nand U73337 ( n61441, n830, n41449 );
nand U73338 ( n14735, n15385, n5204 );
nand U73339 ( n47941, n48515, n7865 );
nand U73340 ( n34215, n34709, n3460 );
nand U73341 ( n68969, n69453, n6075 );
nand U73342 ( n26970, n27464, n4298 );
nand U73343 ( n60110, n60613, n6930 );
nand U73344 ( n27969, n27874, n26955 );
nand U73345 ( n61118, n61021, n60095 );
nand U73346 ( n27805, n27874, n26934 );
nand U73347 ( n60953, n61021, n60074 );
buf U73348 ( n76597, n12687 );
nor U73349 ( n48417, n74442, n47916 );
buf U73350 ( n76331, n46298 );
buf U73351 ( n76594, n76593 );
buf U73352 ( n76595, n76593 );
buf U73353 ( n76211, n65910 );
buf U73354 ( n76277, n57451 );
buf U73355 ( n76535, n24328 );
buf U73356 ( n76355, n45025 );
nor U73357 ( n15278, n74435, n21114 );
buf U73358 ( n76328, n76327 );
buf U73359 ( n76329, n76327 );
nand U73360 ( n34725, n34797, n34179 );
nand U73361 ( n69469, n69541, n68933 );
nand U73362 ( n27480, n27552, n26934 );
nand U73363 ( n60629, n60704, n60074 );
buf U73364 ( n76621, n11324 );
nor U73365 ( n27379, n74423, n28413 );
nor U73366 ( n60527, n74424, n61722 );
nor U73367 ( n34624, n74426, n35594 );
nor U73368 ( n69370, n74425, n70322 );
nor U73369 ( n15058, n5207, n74435 );
nand U73370 ( n15715, n15809, n14952 );
nand U73371 ( n48814, n48882, n48137 );
nand U73372 ( n16134, n16225, n14952 );
nand U73373 ( n49183, n49251, n48137 );
nor U73374 ( n26935, n27297, n27214 );
nor U73375 ( n60075, n60440, n60359 );
nor U73376 ( n44507, n44136, n44544 );
nor U73377 ( n31128, n30776, n31165 );
nor U73378 ( n65382, n64978, n65419 );
nor U73379 ( n23836, n23469, n23873 );
nor U73380 ( n56960, n56591, n56997 );
nor U73381 ( n10712, n10265, n10758 );
nand U73382 ( n15295, n14952, n15395 );
nand U73383 ( n14828, n14952, n14953 );
nand U73384 ( n15077, n15167, n14953 );
nand U73385 ( n48432, n48137, n48522 );
nand U73386 ( n48030, n48137, n48138 );
nand U73387 ( n48252, n48319, n48138 );
nor U73388 ( n34180, n34542, n34459 );
nor U73389 ( n68934, n69290, n69209 );
nand U73390 ( n15517, n15167, n15395 );
nand U73391 ( n48628, n48319, n48522 );
nand U73392 ( n27229, n27297, n27136 );
nand U73393 ( n60374, n60440, n60280 );
nand U73394 ( n27044, n27135, n27136 );
nand U73395 ( n60185, n60279, n60280 );
nand U73396 ( n34474, n34542, n34381 );
nand U73397 ( n69224, n69290, n69133 );
nand U73398 ( n34288, n34380, n34381 );
nand U73399 ( n69040, n69132, n69133 );
nand U73400 ( n27397, n27135, n27467 );
nand U73401 ( n60545, n60279, n60616 );
nand U73402 ( n34642, n34380, n34712 );
nand U73403 ( n69388, n69132, n69456 );
buf U73404 ( n76429, n38306 );
buf U73405 ( n76433, n38305 );
buf U73406 ( n76477, n76479 );
buf U73407 ( n76509, n27751 );
buf U73408 ( n76513, n27750 );
buf U73409 ( n76612, n76609 );
nand U73410 ( n60218, n76260, n57671 );
nand U73411 ( n60207, n76260, n57667 );
nand U73412 ( n60196, n76260, n57663 );
nand U73413 ( n60229, n76260, n57675 );
nand U73414 ( n27066, n76518, n24539 );
nand U73415 ( n27077, n76518, n24543 );
nand U73416 ( n27055, n76518, n24535 );
nand U73417 ( n27088, n76518, n24547 );
nand U73418 ( n48155, n48238, n47908 );
nand U73419 ( n15407, n15385, n5210 );
nand U73420 ( n48625, n48711, n48515 );
nand U73421 ( n15513, n15600, n15385 );
nand U73422 ( n49354, n48711, n49244 );
nand U73423 ( n16034, n15915, n5204 );
nand U73424 ( n15185, n15059, n5204 );
nand U73425 ( n16342, n15600, n16217 );
nand U73426 ( n15822, n15915, n5210 );
nand U73427 ( n14974, n15059, n5210 );
nand U73428 ( n49086, n48982, n7865 );
nand U73429 ( n48350, n48238, n7865 );
nand U73430 ( n27481, n27464, n4295 );
nand U73431 ( n34726, n34709, n3458 );
nand U73432 ( n60630, n60613, n6928 );
nand U73433 ( n69470, n69453, n6073 );
nand U73434 ( n27567, n27631, n27464 );
nand U73435 ( n34810, n34876, n34709 );
nand U73436 ( n60717, n60784, n60613 );
nand U73437 ( n69554, n69618, n69453 );
nand U73438 ( n61373, n60784, n61267 );
nand U73439 ( n28209, n27631, n28112 );
nand U73440 ( n70172, n69618, n70079 );
nand U73441 ( n35442, n34876, n35347 );
nand U73442 ( n27393, n27463, n27464 );
nand U73443 ( n60541, n60612, n60613 );
nand U73444 ( n34638, n34708, n34709 );
nand U73445 ( n69384, n69452, n69453 );
nand U73446 ( n28042, n27463, n28112 );
nand U73447 ( n61201, n60612, n61267 );
nand U73448 ( n27314, n27220, n4298 );
nand U73449 ( n34559, n34465, n3460 );
nand U73450 ( n69307, n69215, n6075 );
nand U73451 ( n60457, n60365, n6930 );
nand U73452 ( n27970, n27875, n4298 );
nand U73453 ( n35205, n35114, n3460 );
nand U73454 ( n61119, n61022, n6930 );
nand U73455 ( n69941, n69850, n6075 );
nand U73456 ( n27150, n27220, n4295 );
nand U73457 ( n60292, n60365, n6928 );
nand U73458 ( n27806, n27875, n4295 );
nand U73459 ( n60954, n61022, n6928 );
nand U73460 ( n35279, n34708, n35347 );
nand U73461 ( n70013, n69452, n70079 );
nand U73462 ( n15927, n16023, n14940 );
nand U73463 ( n34393, n34465, n3458 );
nand U73464 ( n69145, n69215, n6073 );
nand U73465 ( n35047, n35114, n3458 );
nand U73466 ( n69785, n69850, n6073 );
nand U73467 ( n48991, n49077, n48127 );
nand U73468 ( n27888, n27953, n27130 );
nand U73469 ( n35127, n35192, n34374 );
nand U73470 ( n61035, n61106, n60274 );
nand U73471 ( n69863, n69928, n69126 );
buf U73472 ( n76235, n75982 );
buf U73473 ( n76504, n75983 );
buf U73474 ( n76304, n75984 );
buf U73475 ( n76563, n75985 );
buf U73476 ( n76236, n62480 );
buf U73477 ( n76505, n28968 );
buf U73478 ( n76305, n54696 );
buf U73479 ( n76564, n21658 );
buf U73480 ( n76560, n76556 );
buf U73481 ( n76559, n76556 );
buf U73482 ( n76467, n76463 );
buf U73483 ( n76466, n76463 );
buf U73484 ( n76927, SEL );
buf U73485 ( n76574, n16974 );
buf U73486 ( n76585, n16956 );
buf U73487 ( n76584, n16957 );
nand U73488 ( n71274, n72795, n72796 );
nand U73489 ( n40697, n66119, n66120 );
and U73490 ( n21935, n22774, P1_P2_STATE2_REG_1_ );
and U73491 ( n29252, n30095, P1_P3_STATE2_REG_1_ );
and U73492 ( n63019, n64112, P2_P3_STATE2_REG_1_ );
and U73493 ( n55047, n55888, P2_P2_STATE2_REG_1_ );
nor U73494 ( n47908, n74442, P2_P1_INSTQUEUEWR_ADDR_REG_1_ );
buf U73495 ( n76593, n12689 );
buf U73496 ( n76327, n46300 );
not U73497 ( n8208, HOLD );
nor U73498 ( n48319, P2_P1_INSTQUEUEWR_ADDR_REG_0_, n47916 );
nor U73499 ( n47920, n7859, P2_P1_INSTQUEUEWR_ADDR_REG_0_ );
nor U73500 ( n14690, n5205, P1_P1_INSTQUEUEWR_ADDR_REG_0_ );
nor U73501 ( n15167, P1_P1_INSTQUEUEWR_ADDR_REG_0_, n21114 );
nor U73502 ( n60074, n6924, P2_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U73503 ( n26934, n4292, P1_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U73504 ( n34179, n3454, P1_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U73505 ( n68933, n6069, P2_P3_INSTQUEUEWR_ADDR_REG_0_ );
and U73506 ( n44882, n54249, n54250 );
and U73507 ( n31497, n35751, n35752 );
and U73508 ( n24203, n28572, n28573 );
and U73509 ( n65747, n70477, n70478 );
and U73510 ( n57325, n61877, n61878 );
and U73511 ( n11169, n21243, n21244 );
buf U73512 ( n76912, n76913 );
buf U73513 ( n76916, n76917 );
buf U73514 ( n76918, n76919 );
buf U73515 ( n76914, n76915 );
buf U73516 ( n76923, n76924 );
nand U73517 ( n34343, n76462, P1_BUF2_REG_5_ );
nand U73518 ( n34354, n76462, P1_BUF2_REG_6_ );
nand U73519 ( n34321, n76462, P1_BUF2_REG_3_ );
nand U73520 ( n34332, n76462, P1_BUF2_REG_4_ );
nand U73521 ( n69073, n76194, P2_BUF2_REG_3_ );
nand U73522 ( n69106, n76194, P2_BUF2_REG_6_ );
nand U73523 ( n69095, n76194, P2_BUF2_REG_5_ );
nand U73524 ( n69084, n76194, P2_BUF2_REG_4_ );
nand U73525 ( n69062, n76194, P2_BUF2_REG_2_ );
nand U73526 ( n34310, n76462, P1_BUF2_REG_2_ );
nand U73527 ( n34377, n76462, P1_BUF2_REG_7_ );
nand U73528 ( n34299, n76462, P1_BUF2_REG_1_ );
nand U73529 ( n69129, n76194, P2_BUF2_REG_7_ );
nand U73530 ( n69051, n76194, P2_BUF2_REG_1_ );
nand U73531 ( n15078, n15168, n14940 );
nand U73532 ( n48253, n48320, n48127 );
nand U73533 ( n14823, n14939, n14940 );
nand U73534 ( n48026, n48126, n48127 );
nand U73535 ( n27232, n27302, n27130 );
nand U73536 ( n34477, n34547, n34374 );
nand U73537 ( n69227, n69295, n69126 );
nand U73538 ( n60377, n60445, n60274 );
nand U73539 ( n27717, n27789, n27130 );
nand U73540 ( n34962, n35030, n34374 );
nand U73541 ( n69702, n69768, n69126 );
nand U73542 ( n60868, n60937, n60274 );
nand U73543 ( n27038, n27129, n27130 );
nand U73544 ( n34282, n34373, n34374 );
nand U73545 ( n69034, n69125, n69126 );
nand U73546 ( n60179, n60273, n60274 );
and U73547 ( n75706, P2_P2_STATE_REG_1_, n74683 );
and U73548 ( n75707, P1_P2_STATE_REG_1_, n74691 );
and U73549 ( n75708, P2_P1_STATE_REG_1_, n74684 );
and U73550 ( n75709, P1_P1_STATE_REG_1_, n74713 );
not U73551 ( n4827, n13214 );
not U73552 ( n5685, n67503 );
not U73553 ( n7470, n46439 );
not U73554 ( n3928, n25498 );
not U73555 ( n6560, n58635 );
not U73556 ( n3084, n32738 );
buf U73557 ( n76774, n3102 );
buf U73558 ( n76754, n3945 );
buf U73559 ( n76708, n5703 );
buf U73560 ( n76687, n6578 );
buf U73561 ( n76660, n7489 );
buf U73562 ( n76727, n4847 );
not U73563 ( n5723, n67395 );
not U73564 ( n3123, n32630 );
not U73565 ( n7509, n46331 );
not U73566 ( n3965, n25390 );
not U73567 ( n6598, n58527 );
not U73568 ( n4864, n12732 );
nand U73569 ( n13214, n4832, n4864 );
not U73570 ( n5708, n67826 );
not U73571 ( n3107, n33070 );
not U73572 ( n3950, n25823 );
not U73573 ( n6583, n58961 );
not U73574 ( n7494, n46779 );
not U73575 ( n5684, n67396 );
not U73576 ( n3083, n32631 );
not U73577 ( n3927, n25391 );
not U73578 ( n6559, n58528 );
not U73579 ( n4850, n12828 );
not U73580 ( n4825, n12733 );
not U73581 ( n7469, n46332 );
nand U73582 ( n67503, n5689, n5723 );
nand U73583 ( n46439, n7474, n7509 );
nand U73584 ( n25498, n3932, n3965 );
nand U73585 ( n58635, n6564, n6598 );
nand U73586 ( n32738, n3088, n3123 );
buf U73587 ( n76661, n7489 );
buf U73588 ( n76755, n3945 );
buf U73589 ( n76775, n3102 );
buf U73590 ( n76709, n5703 );
buf U73591 ( n76688, n6578 );
buf U73592 ( n76728, n4847 );
buf U73593 ( n76816, n2029 );
buf U73594 ( n76815, n2029 );
buf U73595 ( n76817, n2029 );
not U73596 ( n3102, n32712 );
not U73597 ( n3945, n25472 );
not U73598 ( n5703, n67477 );
not U73599 ( n6578, n58609 );
not U73600 ( n7489, n46413 );
not U73601 ( n4847, n13055 );
nand U73602 ( n46331, n7517, n7518 );
nand U73603 ( n67395, n5732, n5733 );
nand U73604 ( n32630, n3130, n3132 );
nand U73605 ( n25390, n3974, n3975 );
nand U73606 ( n58527, n6607, n6608 );
not U73607 ( n7518, n46349 );
not U73608 ( n3975, n25408 );
not U73609 ( n6608, n58545 );
not U73610 ( n3132, n32648 );
not U73611 ( n5733, n67413 );
not U73612 ( n76489, n76491 );
not U73613 ( n76363, n76365 );
not U73614 ( n76222, n76224 );
not U73615 ( n76633, n76635 );
not U73616 ( n76284, n76286 );
not U73617 ( n76542, n76544 );
not U73618 ( n76490, n76491 );
nand U73619 ( n12732, n4872, n4873 );
not U73620 ( n76634, n76635 );
not U73621 ( n76223, n76224 );
not U73622 ( n76364, n76365 );
not U73623 ( n76543, n76544 );
not U73624 ( n76285, n76286 );
not U73625 ( n4873, n12777 );
buf U73626 ( n76023, n76492 );
buf U73627 ( n75991, n76225 );
buf U73628 ( n76028, n76545 );
buf U73629 ( n75999, n76287 );
buf U73630 ( n76007, n76366 );
buf U73631 ( n76036, n76636 );
buf U73632 ( n76024, n76492 );
buf U73633 ( n76029, n76545 );
buf U73634 ( n76037, n76636 );
buf U73635 ( n75992, n76225 );
buf U73636 ( n76000, n76287 );
buf U73637 ( n76008, n76366 );
buf U73638 ( n76025, n76492 );
buf U73639 ( n76030, n76545 );
buf U73640 ( n75993, n76225 );
buf U73641 ( n76001, n76287 );
buf U73642 ( n76009, n76366 );
buf U73643 ( n76038, n76636 );
not U73644 ( n4832, n12999 );
nand U73645 ( n12733, n4855, n4832 );
nand U73646 ( n46332, n7500, n7474 );
nand U73647 ( n67396, n5714, n5689 );
nand U73648 ( n32631, n3113, n3088 );
nand U73649 ( n25391, n3957, n3932 );
nand U73650 ( n58528, n6589, n6564 );
nand U73651 ( n67826, n5714, n5723 );
nand U73652 ( n33070, n3113, n3123 );
nand U73653 ( n25823, n3957, n3965 );
nand U73654 ( n58961, n6589, n6598 );
not U73655 ( n7474, n46438 );
nor U73656 ( n47867, n7519, n47869 );
nand U73657 ( n46779, n7500, n7509 );
nand U73658 ( n12828, n4855, n4864 );
not U73659 ( n5689, n67502 );
not U73660 ( n3932, n25497 );
not U73661 ( n6564, n58634 );
nor U73662 ( n68887, n5734, n68889 );
nor U73663 ( n26888, n3977, n26890 );
nor U73664 ( n60028, n6609, n60030 );
not U73665 ( n3088, n32737 );
nor U73666 ( n34133, n3133, n34135 );
nor U73667 ( n35825, n34135, n3100 );
nor U73668 ( n28646, n26890, n3944 );
nor U73669 ( n70551, n68889, n5702 );
nor U73670 ( n61951, n60030, n6577 );
nor U73671 ( n54323, n47869, n7488 );
nor U73672 ( n21340, n14635, n4845 );
not U73673 ( n76134, n76131 );
not U73674 ( n76135, n76131 );
not U73675 ( n76137, n76132 );
not U73676 ( n76136, n76131 );
not U73677 ( n76138, n76132 );
not U73678 ( n76139, n76133 );
not U73679 ( n76140, n76133 );
not U73680 ( n76141, n76131 );
buf U73681 ( n76844, n76843 );
buf U73682 ( n76845, n76843 );
buf U73683 ( n76828, n76824 );
buf U73684 ( n76827, n76824 );
nand U73685 ( n72270, n72367, n72368 );
nand U73686 ( n72368, n72369, n1112 );
nor U73687 ( n72367, n72370, n72371 );
nor U73688 ( n72370, n1108, n72378 );
and U73689 ( n71927, n72042, n72043 );
nand U73690 ( n72043, n72044, n1087 );
nor U73691 ( n72042, n72045, n72046 );
nor U73692 ( n72045, n1085, n72053 );
and U73693 ( n72361, n72430, n72431 );
nand U73694 ( n72431, n72432, n1185 );
nor U73695 ( n72430, n72433, n72434 );
nor U73696 ( n72433, n1184, n72441 );
nor U73697 ( n46216, n573, n46221 );
not U73698 ( n76342, n76343 );
not U73699 ( n76198, n76199 );
not U73700 ( n76522, n76523 );
not U73701 ( n76264, n76265 );
buf U73702 ( n76846, n76843 );
nor U73703 ( n46933, n573, n46938 );
not U73704 ( n1099, n71212 );
not U73705 ( n76472, n76473 );
not U73706 ( n76341, n76343 );
not U73707 ( n76197, n76199 );
not U73708 ( n76521, n76523 );
not U73709 ( n76263, n76265 );
not U73710 ( n76471, n76473 );
not U73711 ( n749, n42017 );
buf U73712 ( n76006, n76344 );
buf U73713 ( n76027, n76524 );
buf U73714 ( n75998, n76266 );
buf U73715 ( n75990, n76200 );
buf U73716 ( n76005, n76344 );
buf U73717 ( n76026, n76524 );
buf U73718 ( n75997, n76266 );
buf U73719 ( n75989, n76200 );
buf U73720 ( n76035, n76605 );
buf U73721 ( n76022, n76474 );
buf U73722 ( n76021, n76474 );
not U73723 ( n7562, n47300 );
not U73724 ( n5774, n68331 );
not U73725 ( n4015, n26330 );
not U73726 ( n6648, n59469 );
not U73727 ( n76602, n76604 );
nor U73728 ( n62756, n727, n820 );
nor U73729 ( n40102, n2000, n1855 );
buf U73730 ( n76857, n76853 );
not U73731 ( n76335, n75753 );
buf U73732 ( n76826, n76824 );
nor U73733 ( n66361, n819, n54754 );
not U73734 ( n3175, n33575 );
not U73735 ( n4912, n13930 );
buf U73736 ( n76856, n76853 );
buf U73737 ( n76855, n76853 );
not U73738 ( n76603, n76604 );
not U73739 ( n2029, n38108 );
not U73740 ( n2034, n38792 );
not U73741 ( n76470, n76473 );
nand U73742 ( n60030, n58604, n57738 );
nand U73743 ( n26890, n25467, n24606 );
not U73744 ( n76281, n76282 );
not U73745 ( n76539, n76540 );
nand U73746 ( n68889, n67472, n66414 );
not U73747 ( n76215, n76216 );
nand U73748 ( n34135, n32707, n31822 );
not U73749 ( n76482, n76483 );
not U73750 ( n6689, n55882 );
not U73751 ( n4057, n22768 );
not U73752 ( n5828, n64106 );
not U73753 ( n3229, n30089 );
nor U73754 ( n58545, n61859, n55882 );
nor U73755 ( n25408, n28554, n22768 );
nand U73756 ( n32712, n35781, n3230 );
nor U73757 ( n67413, n70459, n64106 );
nor U73758 ( n32648, n35733, n30089 );
nand U73759 ( n67477, n70507, n5829 );
nand U73760 ( n46413, n54279, n7617 );
nand U73761 ( n25472, n28602, n4058 );
nand U73762 ( n58609, n61907, n6690 );
not U73763 ( n823, n61410 );
nand U73764 ( n13055, n21287, n4963 );
not U73765 ( n2000, n38819 );
buf U73766 ( n76034, n76605 );
nor U73767 ( n57444, n55882, n56203 );
nor U73768 ( n24321, n22768, n23082 );
nor U73769 ( n65903, n64106, n64572 );
nor U73770 ( n31617, n30089, n30413 );
not U73771 ( n819, n61439 );
not U73772 ( n4008, n28560 );
not U73773 ( n6640, n61865 );
not U73774 ( n5767, n70465 );
not U73775 ( n3168, n35739 );
nand U73776 ( n35685, n35713, n34061 );
nand U73777 ( n28506, n28534, n26816 );
nand U73778 ( n70411, n70439, n68815 );
nand U73779 ( n61811, n61839, n59956 );
nand U73780 ( n54183, n54211, n47795 );
not U73781 ( n7517, n43731 );
not U73782 ( n3130, n30414 );
not U73783 ( n3974, n23083 );
not U73784 ( n5732, n64573 );
not U73785 ( n6607, n56204 );
not U73786 ( n4845, n14634 );
nor U73787 ( n46349, n54231, n43362 );
not U73788 ( n4878, n12835 );
not U73789 ( n7488, n47868 );
nand U73790 ( n21199, n21248, n14543 );
not U73791 ( n7523, n46407 );
not U73792 ( n4872, n9812 );
nor U73793 ( n12777, n21233, n9419 );
nand U73794 ( n14635, n12837, n11748 );
nand U73795 ( n47869, n46408, n45521 );
and U73796 ( n21258, n14543, n21248 );
not U73797 ( n4962, n9419 );
not U73798 ( n3100, n34134 );
not U73799 ( n3944, n26889 );
not U73800 ( n5702, n68888 );
not U73801 ( n6577, n60029 );
not U73802 ( n7615, n43362 );
not U73803 ( n3137, n32706 );
not U73804 ( n3980, n25466 );
not U73805 ( n5738, n67471 );
not U73806 ( n6613, n58603 );
buf U73807 ( n76866, n495 );
buf U73808 ( n76892, n224 );
buf U73809 ( n76893, n224 );
buf U73810 ( n76867, n495 );
or U73811 ( n21198, n21199, n4903 );
buf U73812 ( n76616, n76614 );
buf U73813 ( n76615, n76614 );
buf U73814 ( n76617, n76614 );
not U73815 ( n4858, n21287 );
not U73816 ( n3117, n35781 );
not U73817 ( n5718, n70507 );
not U73818 ( n3960, n28602 );
not U73819 ( n6593, n61907 );
not U73820 ( n7504, n54279 );
buf U73821 ( n76272, n76270 );
buf U73822 ( n76530, n76528 );
buf U73823 ( n76529, n76528 );
buf U73824 ( n76271, n76270 );
buf U73825 ( n76206, n76204 );
buf U73826 ( n76205, n76204 );
buf U73827 ( n76207, n76204 );
buf U73828 ( n76531, n76528 );
buf U73829 ( n76273, n76270 );
not U73830 ( n4904, n21239 );
not U73831 ( n7553, n54237 );
buf U73832 ( n76350, n76348 );
buf U73833 ( n76349, n76348 );
or U73834 ( n35684, n35685, n3167 );
or U73835 ( n28505, n28506, n4007 );
or U73836 ( n70410, n70411, n5765 );
or U73837 ( n61810, n61811, n6639 );
or U73838 ( n54182, n54183, n7552 );
buf U73839 ( n76351, n76348 );
not U73840 ( n3097, n32707 );
not U73841 ( n3940, n25467 );
not U73842 ( n5698, n67472 );
not U73843 ( n6573, n58604 );
not U73844 ( n7484, n46408 );
buf U73845 ( n76891, n224 );
buf U73846 ( n76865, n495 );
not U73847 ( n4842, n12837 );
not U73848 ( n76626, n76627 );
nand U73849 ( n12999, n14633, n14634 );
nor U73850 ( n14633, n4874, n14635 );
not U73851 ( n4855, n12775 );
not U73852 ( n7500, n46365 );
nor U73853 ( n54904, n6689, n6693 );
nor U73854 ( n21828, n4057, n4060 );
nor U73855 ( n29143, n3229, n3233 );
nor U73856 ( n62810, n5828, n5832 );
nor U73857 ( n42322, n7615, n7619 );
nor U73858 ( n11317, n9419, n9810 );
nor U73859 ( n44995, n43362, n43730 );
not U73860 ( n76625, n76627 );
not U73861 ( n5714, n67429 );
not U73862 ( n3113, n32664 );
not U73863 ( n3957, n25424 );
not U73864 ( n6589, n58561 );
nand U73865 ( n46438, n47867, n47868 );
nor U73866 ( n8262, n4962, n4965 );
not U73867 ( n4874, n14637 );
nand U73868 ( n67502, n68887, n68888 );
nand U73869 ( n25497, n26888, n26889 );
nand U73870 ( n58634, n60028, n60029 );
nand U73871 ( n32737, n34133, n34134 );
not U73872 ( n7519, n47870 );
buf U73873 ( n76772, n3104 );
buf U73874 ( n76705, n5705 );
buf U73875 ( n76751, n3948 );
buf U73876 ( n76684, n6580 );
buf U73877 ( n76724, n4849 );
buf U73878 ( n76657, n7492 );
buf U73879 ( n76756, n3915 );
buf U73880 ( n76689, n6548 );
not U73881 ( n5734, n68890 );
not U73882 ( n3133, n34136 );
not U73883 ( n3977, n26891 );
not U73884 ( n6609, n60031 );
buf U73885 ( n76757, n3915 );
buf U73886 ( n76690, n6548 );
buf U73887 ( n76773, n3104 );
nand U73888 ( n76100, n47867, n47868 );
nand U73889 ( n76057, n68887, n68888 );
nand U73890 ( n76127, n34133, n34134 );
nand U73891 ( n76155, n26888, n26889 );
nand U73892 ( n76083, n60028, n60029 );
buf U73893 ( n76706, n5705 );
buf U73894 ( n76752, n3948 );
buf U73895 ( n76685, n6580 );
buf U73896 ( n76725, n4849 );
buf U73897 ( n76658, n7492 );
buf U73898 ( n76707, n5705 );
buf U73899 ( n76753, n3948 );
buf U73900 ( n76686, n6580 );
buf U73901 ( n76726, n4849 );
nand U73902 ( n76058, n68887, n68888 );
nand U73903 ( n76101, n47867, n47868 );
nand U73904 ( n76156, n26888, n26889 );
nand U73905 ( n76084, n60028, n60029 );
nand U73906 ( n76128, n34133, n34134 );
buf U73907 ( n76659, n7492 );
nor U73908 ( n12823, n4877, n4874 );
not U73909 ( n4877, n11748 );
nor U73910 ( n46393, n7522, n7519 );
not U73911 ( n7522, n45521 );
nor U73912 ( n67457, n5737, n5734 );
not U73913 ( n5737, n66414 );
nor U73914 ( n32692, n3135, n3133 );
not U73915 ( n3135, n31822 );
nor U73916 ( n25452, n3979, n3977 );
not U73917 ( n3979, n24606 );
nor U73918 ( n58589, n6612, n6609 );
not U73919 ( n6612, n57738 );
not U73920 ( n4848, n13060 );
not U73921 ( n5704, n67479 );
not U73922 ( n3103, n32714 );
not U73923 ( n3947, n25474 );
not U73924 ( n6579, n58611 );
not U73925 ( n7490, n46415 );
not U73926 ( n76131, n31728 );
not U73927 ( n76132, n31728 );
not U73928 ( n76133, n31728 );
not U73929 ( n1755, n49885 );
not U73930 ( n1362, n49713 );
not U73931 ( n1738, n49952 );
not U73932 ( n1717, n49962 );
not U73933 ( n1278, n49693 );
nand U73934 ( n50278, n49885, n50273 );
not U73935 ( n1749, n50273 );
nand U73936 ( n50231, n49962, n49960 );
nand U73937 ( n50254, n49952, n49950 );
not U73938 ( n2478, n16757 );
not U73939 ( n2855, n16997 );
not U73940 ( n2834, n17007 );
not U73941 ( n2393, n16737 );
not U73942 ( n8229, n49930 );
not U73943 ( n2639, n20421 );
not U73944 ( n2485, n18185 );
nand U73945 ( n17285, n17007, n17005 );
nand U73946 ( n17308, n16997, n16995 );
not U73947 ( n1729, n49950 );
not U73948 ( n1369, n51141 );
not U73949 ( n1517, n53275 );
not U73950 ( n1539, n53395 );
not U73951 ( n1407, n52638 );
not U73952 ( n1542, n53417 );
not U73953 ( n2527, n19682 );
not U73954 ( n2847, n16995 );
not U73955 ( n2662, n20535 );
not U73956 ( n2664, n20244 );
not U73957 ( n1728, n50258 );
not U73958 ( n1707, n49960 );
not U73959 ( n1628, n51957 );
not U73960 ( n1645, n52855 );
or U73961 ( n51632, n51633, n51634 );
not U73962 ( n2824, n17005 );
not U73963 ( n1648, n52413 );
not U73964 ( n1660, n51573 );
or U73965 ( n18676, n18677, n18678 );
not U73966 ( n2768, n19324 );
not U73967 ( n2782, n18621 );
not U73968 ( n1658, n50180 );
not U73969 ( n1650, n51422 );
not U73970 ( n2770, n18466 );
not U73971 ( n1507, n49754 );
not U73972 ( n2629, n16799 );
not U73973 ( n76389, n76390 );
nor U73974 ( n40820, n40831, n40819 );
nor U73975 ( n40831, n515, n40817 );
not U73976 ( n515, n40706 );
not U73977 ( n76457, n76459 );
nor U73978 ( n36833, n36834, n2013 );
nor U73979 ( n36834, n2015, n36548 );
nor U73980 ( n36830, n36831, n36832 );
nor U73981 ( n36831, n36837, n36836 );
nor U73982 ( n36832, n2011, n36833 );
nor U73983 ( n36837, n36839, n2015 );
not U73984 ( n76458, n76459 );
buf U73985 ( n76801, n76799 );
buf U73986 ( n76807, n2037 );
nand U73987 ( n36545, n36550, n36548 );
nand U73988 ( n36550, n36436, n36438 );
nand U73989 ( n38785, n1902, n2038 );
nand U73990 ( n38813, n38814, n38815 );
not U73991 ( n564, n61438 );
nand U73992 ( n61403, n837, n564 );
nor U73993 ( n61399, n41597, n61400 );
nor U73994 ( n61400, n61401, n61402 );
nand U73995 ( n61401, n61405, n61406 );
nand U73996 ( n61402, n61403, n61404 );
nand U73997 ( n61433, n61434, n61435 );
nand U73998 ( n61421, n61422, n61423 );
nand U73999 ( n61422, n61439, n61440 );
nand U74000 ( n61423, n778, n61424 );
nand U74001 ( n61424, n61425, n61426 );
nand U74002 ( n61434, n837, n61438 );
nand U74003 ( n61406, n825, n564 );
nor U74004 ( n38922, n2132, n1900 );
nand U74005 ( n40892, n40893, n40703 );
nand U74006 ( n40893, n40894, n76850 );
nor U74007 ( n40894, n40895, n40896 );
nor U74008 ( n40896, n598, n40897 );
nand U74009 ( n40897, n40898, n40899 );
nand U74010 ( n40899, n608, n40900 );
not U74011 ( n1843, n36509 );
not U74012 ( n540, n62254 );
nor U74013 ( n61626, n832, n61609 );
nand U74014 ( n62282, n62283, n41517 );
nand U74015 ( n62283, n563, n62284 );
nand U74016 ( n62284, n765, n61410 );
not U74017 ( n563, n62285 );
and U74018 ( n62339, n62275, n825 );
and U74019 ( n62342, n62275, n837 );
nor U74020 ( n72504, n1124, n1140 );
nor U74021 ( n71532, n1037, n1043 );
not U74022 ( n1179, n72523 );
not U74023 ( n1107, n72409 );
not U74024 ( n1083, n72282 );
not U74025 ( n1062, n71955 );
not U74026 ( n1043, n71530 );
nand U74027 ( n72174, n72273, n72274 );
nand U74028 ( n72274, n72275, n1083 );
nor U74029 ( n72273, n72276, n72277 );
nor U74030 ( n72276, n1083, n72283 );
nor U74031 ( n72730, n72731, n72524 );
nor U74032 ( n72731, n72732, n72525 );
nor U74033 ( n72732, n1165, n72523 );
nor U74034 ( n72404, n72405, n72406 );
nor U74035 ( n72405, n72407, n72408 );
nor U74036 ( n72407, n1095, n72409 );
nor U74037 ( n72277, n72278, n72279 );
nor U74038 ( n72278, n72280, n72281 );
nor U74039 ( n72280, n1073, n72282 );
nand U74040 ( n71653, n72077, n72078 );
nand U74041 ( n72078, n71955, n71952 );
nor U74042 ( n72077, n71954, n71948 );
nand U74043 ( n72519, n72727, n72728 );
nand U74044 ( n72728, n72526, n1179 );
nor U74045 ( n72727, n72729, n72730 );
nor U74046 ( n72729, n1179, n72734 );
and U74047 ( n72494, n72647, n72648 );
nand U74048 ( n72648, n72505, n1140 );
nor U74049 ( n72647, n72650, n72651 );
nor U74050 ( n72650, n1140, n72654 );
and U74051 ( n72382, n72400, n72401 );
nand U74052 ( n72401, n72402, n1107 );
nor U74053 ( n72400, n72403, n72404 );
nor U74054 ( n72403, n1107, n72410 );
and U74055 ( n71658, n71935, n71936 );
nand U74056 ( n71936, n71533, n1043 );
nor U74057 ( n71935, n71938, n71939 );
nor U74058 ( n71938, n1043, n71942 );
not U74059 ( n1059, n71646 );
not U74060 ( n1044, n71361 );
nand U74061 ( n71641, n72304, n72305 );
nand U74062 ( n72305, n72282, n72279 );
nor U74063 ( n72304, n72281, n72275 );
buf U74064 ( n76847, n613 );
nand U74065 ( n71051, n71052, n71053 );
nor U74066 ( n71950, n71951, n71952 );
nor U74067 ( n71951, n71953, n71954 );
nor U74068 ( n71953, n1053, n71955 );
and U74069 ( n71934, n71946, n71947 );
nand U74070 ( n71947, n71948, n1062 );
nor U74071 ( n71946, n71949, n71950 );
nor U74072 ( n71949, n1062, n71956 );
nor U74073 ( n38930, n2039, n38879 );
not U74074 ( n1180, n72683 );
nand U74075 ( n72517, n72705, n72706 );
nand U74076 ( n72706, n72683, n72680 );
nor U74077 ( n72705, n72682, n72676 );
nand U74078 ( n38938, n2005, n38877 );
nor U74079 ( n71579, n1127, n1147 );
not U74080 ( n1188, n71590 );
not U74081 ( n1082, n71550 );
not U74082 ( n1109, n71563 );
nand U74083 ( n71637, n72484, n72485 );
nand U74084 ( n72485, n71566, n1109 );
nor U74085 ( n72484, n72486, n72487 );
nor U74086 ( n72486, n1109, n72491 );
nand U74087 ( n71625, n72527, n72528 );
nand U74088 ( n72528, n71593, n1188 );
nor U74089 ( n72527, n72529, n72530 );
nor U74090 ( n72529, n1188, n72534 );
nand U74091 ( n71631, n72506, n72507 );
nand U74092 ( n72507, n71580, n1147 );
nor U74093 ( n72506, n72509, n72510 );
nor U74094 ( n72509, n1147, n72513 );
nor U74095 ( n72530, n72531, n71591 );
nor U74096 ( n72531, n72532, n71592 );
nor U74097 ( n72532, n1174, n71590 );
nor U74098 ( n72392, n72393, n71551 );
nor U74099 ( n72393, n72394, n71552 );
nor U74100 ( n72394, n1072, n71550 );
nor U74101 ( n72487, n72488, n71564 );
nor U74102 ( n72488, n72489, n71565 );
nor U74103 ( n72489, n1097, n71563 );
and U74104 ( n71643, n72389, n72390 );
nand U74105 ( n72390, n71553, n1082 );
nor U74106 ( n72389, n72391, n72392 );
nor U74107 ( n72391, n1082, n72396 );
not U74108 ( n1060, n71375 );
nor U74109 ( n71544, n71543, n71546 );
xor U74110 ( n71546, n1060, n1068 );
and U74111 ( n71488, n71541, n71542 );
nand U74112 ( n71542, n71376, n1060 );
nor U74113 ( n71541, n71544, n71545 );
and U74114 ( n71545, n1068, n71377 );
nand U74115 ( n71635, n72555, n72556 );
nand U74116 ( n72556, n72409, n72406 );
nor U74117 ( n72555, n72408, n72402 );
not U74118 ( n538, n61628 );
nor U74119 ( n62262, n62264, n62265 );
nor U74120 ( n62264, n538, n833 );
nor U74121 ( n62265, n538, n832 );
nand U74122 ( n62665, n62462, n62466 );
nand U74123 ( n62550, n62558, n62559 );
nand U74124 ( n62558, n62570, n41919 );
nand U74125 ( n62559, n748, n62560 );
nand U74126 ( n62570, n62571, n62572 );
nand U74127 ( n62560, n62561, n62562 );
nor U74128 ( n62561, n62568, n62569 );
nor U74129 ( n62562, n62563, n62564 );
nor U74130 ( n62568, n832, n62473 );
and U74131 ( n72676, n1167, n72680 );
nand U74132 ( n71623, n72521, n72522 );
nand U74133 ( n72522, n72523, n72524 );
nor U74134 ( n72521, n72525, n72526 );
not U74135 ( n1878, n38130 );
nand U74136 ( n71140, n71372, n71373 );
nand U74137 ( n71373, n71374, n71375 );
nor U74138 ( n71372, n71376, n71377 );
not U74139 ( n1034, n71350 );
nor U74140 ( n72678, n72679, n72680 );
nor U74141 ( n72679, n72681, n72682 );
nor U74142 ( n72681, n1167, n72683 );
nand U74143 ( n72612, n72674, n72675 );
nand U74144 ( n72675, n72676, n1180 );
nor U74145 ( n72674, n72677, n72678 );
nor U74146 ( n72677, n1180, n72684 );
nor U74147 ( n72161, n1129, n1154 );
not U74148 ( n1193, n72260 );
not U74149 ( n1118, n71979 );
not U74150 ( n1089, n71926 );
not U74151 ( n1067, n71691 );
nand U74152 ( n71982, n72153, n72154 );
nand U74153 ( n72154, n72155, n1154 );
nor U74154 ( n72153, n72156, n72157 );
nor U74155 ( n72156, n1153, n72164 );
nand U74156 ( n72149, n72249, n72250 );
nand U74157 ( n72250, n72251, n1193 );
nor U74158 ( n72249, n72252, n72253 );
nor U74159 ( n72252, n1192, n72259 );
and U74160 ( n71914, n71968, n71969 );
nand U74161 ( n71969, n71970, n1118 );
nor U74162 ( n71968, n71971, n71972 );
nor U74163 ( n71971, n1117, n71978 );
not U74164 ( n542, n62308 );
nor U74165 ( n62377, n62381, n62382 );
nor U74166 ( n62381, n542, n833 );
nor U74167 ( n62382, n542, n832 );
and U74168 ( n72526, n1165, n72524 );
nor U74169 ( n39162, n2112, n39194 );
nor U74170 ( n72467, n1125, n1144 );
not U74171 ( n1182, n72644 );
nand U74172 ( n72593, n72635, n72636 );
nand U74173 ( n72636, n72637, n1182 );
nor U74174 ( n72635, n72638, n72639 );
nor U74175 ( n72638, n1182, n72645 );
nand U74176 ( n72363, n72459, n72460 );
nand U74177 ( n72460, n72461, n1144 );
nor U74178 ( n72459, n72462, n72463 );
nor U74179 ( n72462, n1144, n72470 );
nor U74180 ( n72371, n72372, n72373 );
nor U74181 ( n72372, n72374, n72375 );
nor U74182 ( n72374, n72376, n72377 );
nor U74183 ( n72639, n72640, n72641 );
nor U74184 ( n72640, n72642, n72643 );
nor U74185 ( n72642, n1168, n72644 );
and U74186 ( n72375, n72376, n72377 );
and U74187 ( n72275, n1073, n72279 );
nand U74188 ( n71483, n71548, n71549 );
nand U74189 ( n71549, n71550, n71551 );
nor U74190 ( n71548, n71552, n71553 );
not U74191 ( n1068, n71374 );
nand U74192 ( n62312, n62313, n62314 );
nand U74193 ( n62313, n62318, n62316 );
nand U74194 ( n62314, n62315, n62316 );
nor U74195 ( n62318, n832, n62317 );
nor U74196 ( n71556, n71558, n71559 );
xor U74197 ( n71559, n71388, n71387 );
nor U74198 ( n62383, n62384, n62385 );
nand U74199 ( n62384, n62390, n62391 );
nand U74200 ( n62385, n62386, n62387 );
nor U74201 ( n62391, n62392, n62393 );
nor U74202 ( n62390, n62396, n62397 );
nor U74203 ( n62396, n833, n62308 );
nor U74204 ( n62397, n832, n62308 );
not U74205 ( n1084, n72091 );
nand U74206 ( n72414, n72597, n72598 );
nand U74207 ( n72598, n72599, n1143 );
nor U74208 ( n72597, n72600, n72601 );
nor U74209 ( n72600, n1142, n72608 );
and U74210 ( n72402, n1095, n72406 );
and U74211 ( n71948, n1053, n71952 );
not U74212 ( n1113, n72208 );
nand U74213 ( n72056, n72094, n72095 );
nand U74214 ( n72095, n72048, n72052 );
nor U74215 ( n72094, n72044, n72050 );
nor U74216 ( n72203, n72204, n72205 );
nor U74217 ( n72204, n72206, n72207 );
nor U74218 ( n72206, n1102, n72208 );
and U74219 ( n72044, n72051, n72048 );
and U74220 ( n72172, n72199, n72200 );
nand U74221 ( n72200, n72201, n1113 );
nor U74222 ( n72199, n72202, n72203 );
nor U74223 ( n72202, n1113, n72209 );
nand U74224 ( n62263, n822, n61628 );
nor U74225 ( n72224, n1128, n1152 );
not U74226 ( n1190, n72358 );
nand U74227 ( n72261, n72347, n72348 );
nand U74228 ( n72348, n72349, n1190 );
nor U74229 ( n72347, n72350, n72351 );
nor U74230 ( n72350, n1187, n72357 );
nor U74231 ( n72046, n72047, n72048 );
nor U74232 ( n72047, n72049, n72050 );
nor U74233 ( n72049, n72051, n72052 );
and U74234 ( n72050, n72051, n72052 );
and U74235 ( n71800, n71819, n71820 );
nand U74236 ( n71820, n71821, n1064 );
nor U74237 ( n71819, n71822, n71823 );
nor U74238 ( n71822, n1063, n71830 );
and U74239 ( n72168, n72216, n72217 );
nand U74240 ( n72217, n72218, n1152 );
nor U74241 ( n72216, n72219, n72220 );
nor U74242 ( n72219, n1150, n72227 );
nand U74243 ( n39117, n1903, n2038 );
not U74244 ( n1183, n72590 );
nand U74245 ( n72595, n72619, n72620 );
nand U74246 ( n72620, n72590, n72587 );
nor U74247 ( n72619, n72589, n72583 );
and U74248 ( n71553, n1072, n71551 );
not U74249 ( n1087, n72052 );
or U74250 ( n72053, n72051, n1087 );
not U74251 ( n1112, n72377 );
or U74252 ( n72378, n72376, n1112 );
and U74253 ( n62392, n62351, n825 );
nand U74254 ( n72271, n72309, n72310 );
nand U74255 ( n72310, n72208, n72205 );
nor U74256 ( n72309, n72207, n72201 );
nor U74257 ( n71381, n71380, n71383 );
xor U74258 ( n71383, n71155, n71156 );
not U74259 ( n1064, n71829 );
not U74260 ( n1119, n71908 );
not U74261 ( n1092, n71792 );
not U74262 ( n1090, n71787 );
nand U74263 ( n71933, n71958, n71959 );
nand U74264 ( n71959, n71825, n71829 );
nor U74265 ( n71958, n71821, n71827 );
nor U74266 ( n45492, n61444, n61440 );
or U74267 ( n61444, n61447, n61448 );
nor U74268 ( n61447, n61450, n61451 );
nor U74269 ( n61448, n778, n61449 );
and U74270 ( n71593, n1174, n71591 );
nand U74271 ( n71117, n71118, n71119 );
nand U74272 ( n71119, n1038, n71120 );
not U74273 ( n1038, n71121 );
not U74274 ( n1088, n71921 );
not U74275 ( n1065, n71686 );
not U74276 ( n1085, n72048 );
nor U74277 ( n72034, n1130, n1157 );
not U74278 ( n1195, n72148 );
and U74279 ( n72583, n1169, n72587 );
nand U74280 ( n72380, n72412, n72413 );
nand U74281 ( n72413, n72373, n72377 );
nor U74282 ( n72412, n72375, n72369 );
nand U74283 ( n71124, n71118, n71121 );
not U74284 ( n1194, n72143 );
nand U74285 ( n72614, n72658, n72659 );
nand U74286 ( n72659, n72644, n72641 );
nor U74287 ( n72658, n72643, n72637 );
nand U74288 ( n71895, n72026, n72027 );
nand U74289 ( n72027, n72028, n1157 );
nor U74290 ( n72026, n72029, n72030 );
nor U74291 ( n72029, n1155, n72037 );
nor U74292 ( n71557, n71388, n71390 );
nand U74293 ( n62387, n837, n62351 );
nand U74294 ( n71477, n71561, n71562 );
nand U74295 ( n71562, n71563, n71564 );
nor U74296 ( n71561, n71565, n71566 );
and U74297 ( n71566, n1097, n71564 );
not U74298 ( n1114, n72105 );
nor U74299 ( n72028, n1130, n1155 );
nor U74300 ( n62443, n62447, n62448 );
nor U74301 ( n62447, n540, n833 );
nor U74302 ( n62448, n540, n832 );
not U74303 ( n1192, n72255 );
and U74304 ( n71376, n71543, n71374 );
nor U74305 ( n72585, n72586, n72587 );
nor U74306 ( n72586, n72588, n72589 );
nor U74307 ( n72588, n1169, n72590 );
nand U74308 ( n72423, n72581, n72582 );
nand U74309 ( n72582, n72583, n1183 );
nor U74310 ( n72581, n72584, n72585 );
nor U74311 ( n72584, n1183, n72591 );
nor U74312 ( n71570, n71569, n71572 );
xor U74313 ( n71572, n71402, n71401 );
and U74314 ( n71479, n71567, n71568 );
nand U74315 ( n71568, n71403, n1110 );
nor U74316 ( n71567, n71570, n71571 );
not U74317 ( n1110, n71402 );
nor U74318 ( n72155, n1129, n1153 );
nand U74319 ( n71390, n71558, n71387 );
and U74320 ( n72369, n72376, n72373 );
not U74321 ( n1063, n71825 );
and U74322 ( n72637, n1168, n72641 );
and U74323 ( n72264, n72331, n72332 );
nand U74324 ( n72332, n72255, n72260 );
nor U74325 ( n72331, n72251, n72257 );
not U74326 ( n1108, n72373 );
nor U74327 ( n71394, n71393, n71397 );
xor U74328 ( n71397, n71178, n71179 );
nor U74329 ( n72434, n72435, n72436 );
nor U74330 ( n72435, n72437, n72438 );
nor U74331 ( n72437, n72439, n72440 );
and U74332 ( n72268, n72314, n72315 );
nand U74333 ( n72315, n72316, n1149 );
nor U74334 ( n72314, n72317, n72318 );
nor U74335 ( n72317, n1145, n72325 );
and U74336 ( n72438, n72439, n72440 );
nor U74337 ( n62449, n62450, n62451 );
nand U74338 ( n62450, n62456, n62457 );
nand U74339 ( n62451, n62452, n62453 );
nor U74340 ( n62457, n62458, n62459 );
nor U74341 ( n62456, n62469, n62470 );
nor U74342 ( n62469, n833, n62254 );
nor U74343 ( n62470, n832, n62254 );
not U74344 ( n1187, n72353 );
nor U74345 ( n72218, n1128, n1150 );
and U74346 ( n72201, n1102, n72205 );
not U74347 ( n1185, n72440 );
or U74348 ( n72441, n72439, n1185 );
xor U74349 ( n45753, n61586, n61450 );
nand U74350 ( n61584, n61585, n810 );
nand U74351 ( n61585, n45753, n827 );
and U74352 ( n72362, n72442, n72443 );
nand U74353 ( n72443, n72353, n72358 );
nor U74354 ( n72442, n72349, n72355 );
nor U74355 ( n62745, n62746, n41917 );
nor U74356 ( n62746, n62747, n62748 );
nand U74357 ( n62748, n62749, n62750 );
nand U74358 ( n62747, n62751, n62752 );
nand U74359 ( n72425, n72565, n72566 );
nand U74360 ( n72566, n72436, n72440 );
nor U74361 ( n72565, n72432, n72438 );
not U74362 ( n1197, n72004 );
xor U74363 ( n71148, n71149, n71150 );
nand U74364 ( n71149, n71157, n71158 );
nor U74365 ( n71150, n71151, n71152 );
nand U74366 ( n71158, n1069, n71159 );
nand U74367 ( n71154, n71380, n71156 );
nand U74368 ( n46221, n62305, n62306 );
nand U74369 ( n62305, n758, n62307 );
or U74370 ( n62307, n62308, n760 );
nor U74371 ( n71133, n71137, n71138 );
nor U74372 ( n71137, n1054, n71139 );
not U74373 ( n1054, n71140 );
and U74374 ( n72432, n72439, n72436 );
nor U74375 ( n71854, n1158, n1132 );
and U74376 ( n71764, n71846, n71847 );
nand U74377 ( n71847, n71848, n1158 );
nor U74378 ( n71846, n71849, n71850 );
nor U74379 ( n71849, n1158, n71857 );
nor U74380 ( n71408, n71407, n71411 );
xor U74381 ( n71411, n71201, n71202 );
and U74382 ( n71403, n71569, n71401 );
nand U74383 ( n62664, n62586, n837 );
not U74384 ( n559, n62462 );
nor U74385 ( n71314, n71138, n71140 );
xor U74386 ( n46551, n62308, n757 );
nand U74387 ( n62357, n62358, n810 );
nand U74388 ( n62358, n46551, n827 );
nand U74389 ( n45744, n45751, n45752 );
nand U74390 ( n45751, n45753, n45754 );
and U74391 ( n71151, n71155, n71156 );
xor U74392 ( n45999, n41926, n61589 );
not U74393 ( n740, n41581 );
nand U74394 ( n71177, n71393, n71179 );
not U74395 ( n1184, n72436 );
nor U74396 ( n71712, n1133, n1159 );
and U74397 ( n71893, n71998, n71999 );
nand U74398 ( n71999, n72000, n1198 );
nor U74399 ( n71998, n72001, n72002 );
nor U74400 ( n72001, n1197, n72008 );
nand U74401 ( n71465, n71588, n71589 );
nand U74402 ( n71589, n71590, n71591 );
nor U74403 ( n71588, n71592, n71593 );
nor U74404 ( n71718, n1133, n1160 );
nand U74405 ( n62774, n559, n825 );
nor U74406 ( n62564, n833, n62473 );
nand U74407 ( n46545, n46550, n45752 );
nand U74408 ( n46550, n46551, n45754 );
nor U74409 ( n71597, n71596, n71599 );
xor U74410 ( n71599, n71433, n71432 );
nand U74411 ( n71467, n71594, n71595 );
nand U74412 ( n71595, n71434, n1189 );
nor U74413 ( n71594, n71597, n71598 );
not U74414 ( n1189, n71433 );
not U74415 ( n534, n62757 );
nand U74416 ( n71200, n71407, n71202 );
nand U74417 ( n39282, n39283, n2103 );
nor U74418 ( n39283, n2058, n39284 );
nor U74419 ( n39284, n39285, n39286 );
nor U74420 ( n39285, n2052, n2002 );
not U74421 ( n7564, n47281 );
not U74422 ( n7610, n47602 );
not U74423 ( n1882, n39286 );
nand U74424 ( n71159, n71160, n71161 );
nand U74425 ( n71161, n1075, n71162 );
not U74426 ( n1075, n71163 );
nand U74427 ( n57542, n62820, n62821 );
nor U74428 ( n62821, n62822, n62823 );
nor U74429 ( n62820, n62834, n48210 );
nand U74430 ( n62823, n62824, n810 );
nand U74431 ( n62749, n837, n62462 );
xor U74432 ( n46938, n62254, n41920 );
nand U74433 ( n48206, n48207, n48208 );
or U74434 ( n48208, n48209, n573 );
nand U74435 ( n48207, n76857, n48210 );
nor U74436 ( n38262, n39287, n39288 );
nor U74437 ( n39288, n39289, n39290 );
nor U74438 ( n39287, n39259, n2103 );
nand U74439 ( n39289, n2103, n39293 );
not U74440 ( n5777, n68312 );
not U74441 ( n4018, n26311 );
not U74442 ( n6650, n59450 );
not U74443 ( n5823, n68623 );
not U74444 ( n4054, n26622 );
not U74445 ( n6687, n59764 );
nand U74446 ( n62837, n62849, n62850 );
nand U74447 ( n62849, n62854, n62852 );
nand U74448 ( n62850, n62851, n62852 );
nor U74449 ( n62854, n832, n62853 );
nand U74450 ( n71306, n71436, n71437 );
nand U74451 ( n71437, n71300, n1204 );
nor U74452 ( n71436, n71439, n71440 );
not U74453 ( n1204, n71299 );
not U74454 ( n537, n62577 );
nor U74455 ( n62668, n62672, n62673 );
nor U74456 ( n62672, n537, n833 );
nor U74457 ( n62673, n537, n832 );
nor U74458 ( n62744, n833, n62741 );
nand U74459 ( n62741, n48075, n48074 );
and U74460 ( n71434, n71596, n71432 );
not U74461 ( n1845, n36530 );
nand U74462 ( n39585, n39595, n39596 );
nand U74463 ( n39595, n39606, n1977 );
nand U74464 ( n39596, n39581, n39597 );
nand U74465 ( n39606, n39607, n39608 );
not U74466 ( n519, n40928 );
nand U74467 ( n62572, n822, n62473 );
not U74468 ( n589, n41100 );
nand U74469 ( n71181, n1078, n71182 );
not U74470 ( n1078, n71187 );
nand U74471 ( n71182, n71183, n71184 );
nand U74472 ( n71184, n1098, n71185 );
xnor U74473 ( n47416, n62473, n748 );
nor U74474 ( n46452, n76341, n7493 );
nor U74475 ( n67516, n76197, n5707 );
nor U74476 ( n25511, n76521, n3949 );
nor U74477 ( n58648, n76263, n6582 );
nand U74478 ( n71180, n71187, n71188 );
nand U74479 ( n71188, n71185, n71189 );
nand U74480 ( n71189, n71183, n71186 );
not U74481 ( n1098, n71186 );
not U74482 ( n1964, n36716 );
nor U74483 ( n39533, n39536, n1978 );
nor U74484 ( n39536, n1979, n1865 );
nand U74485 ( n39474, n2038, n39430 );
not U74486 ( n727, n62686 );
xor U74487 ( n47960, n62577, n744 );
nand U74488 ( n62632, n62633, n810 );
nand U74489 ( n62633, n47960, n827 );
buf U74490 ( n76829, n76825 );
buf U74491 ( n76825, n2023 );
nor U74492 ( n64018, n64020, n64021 );
nor U74493 ( n64020, n533, n833 );
nor U74494 ( n64021, n533, n832 );
and U74495 ( n71511, n71710, n71711 );
nand U74496 ( n71711, n71712, n1160 );
nor U74497 ( n71710, n71713, n71714 );
nor U74498 ( n71713, n1159, n71721 );
xor U74499 ( n71212, n71217, n71218 );
nor U74500 ( n71218, n71219, n71220 );
xor U74501 ( n71217, n71223, n71224 );
nor U74502 ( n71219, n1162, n1163 );
nand U74503 ( n71203, n71205, n71206 );
nand U74504 ( n71205, n71212, n71213 );
nand U74505 ( n71206, n1099, n71207 );
nand U74506 ( n71213, n71210, n71214 );
nand U74507 ( n41515, n41516, n41517 );
nand U74508 ( n41516, n41518, n41519 );
nand U74509 ( n41519, n41520, n41521 );
nand U74510 ( n41520, n41522, n41523 );
nor U74511 ( n64217, n698, n64219 );
nor U74512 ( n64219, n64220, n64221 );
nand U74513 ( n64221, n64222, n64223 );
nand U74514 ( n64220, n64224, n64225 );
nand U74515 ( n47954, n47959, n45752 );
nand U74516 ( n47959, n47960, n45754 );
not U74517 ( n3178, n33556 );
not U74518 ( n3224, n33867 );
nand U74519 ( n71207, n71208, n71209 );
nand U74520 ( n71209, n1134, n71210 );
not U74521 ( n1134, n71211 );
nand U74522 ( n71214, n71208, n71211 );
nand U74523 ( n64222, n64032, n837 );
or U74524 ( n42066, n770, n41597 );
not U74525 ( n530, n64513 );
nand U74526 ( n64505, n64506, n64507 );
nand U74527 ( n64506, n825, n64518 );
nand U74528 ( n64507, n49026, n64216 );
nand U74529 ( n42017, n41522, n41518 );
nor U74530 ( n42073, n42017, n42051 );
and U74531 ( n41985, n42073, n42088 );
nor U74532 ( n42088, n41579, n649 );
nand U74533 ( n41527, n41528, n41529 );
nor U74534 ( n32751, n76470, n3105 );
nor U74535 ( n39708, n39709, n39710 );
nor U74536 ( n39710, n2039, n39668 );
nor U74537 ( n39709, n2002, n39678 );
not U74538 ( n1863, n39773 );
and U74539 ( n42046, n41529, n41528 );
nor U74540 ( n39834, n2039, n39835 );
xor U74541 ( n39835, n1955, n1864 );
nor U74542 ( n64795, n64801, n682 );
nor U74543 ( n64801, n64802, n64803 );
nor U74544 ( n64802, n555, n64800 );
nor U74545 ( n64803, n819, n530 );
nand U74546 ( n41915, n41919, n41920 );
nand U74547 ( n41935, n41936, n41937 );
nor U74548 ( n37503, n2105, n2112 );
not U74549 ( n1993, n37454 );
buf U74550 ( n76344, n75700 );
nand U74551 ( n41916, n41917, n41918 );
nand U74552 ( n41929, n41933, n773 );
xor U74553 ( n38381, n39668, n1968 );
not U74554 ( n598, n40901 );
not U74555 ( n529, n65823 );
nor U74556 ( n65817, n819, n65801 );
buf U74557 ( n76524, n75702 );
buf U74558 ( n76266, n75703 );
buf U74559 ( n76200, n75701 );
and U74560 ( n39935, n39930, n75710 );
and U74561 ( n75710, n39931, n38819 );
and U74562 ( n47517, n47601, n47480 );
nand U74563 ( n47601, n7595, n47602 );
not U74564 ( n763, n41937 );
not U74565 ( n725, n62845 );
and U74566 ( n26537, n26621, n26500 );
nand U74567 ( n26621, n4042, n26622 );
and U74568 ( n59679, n59763, n59639 );
nand U74569 ( n59763, n6674, n59764 );
and U74570 ( n68538, n68622, n68501 );
nand U74571 ( n68622, n5808, n68623 );
nor U74572 ( n41212, n40847, n40842 );
not U74573 ( n739, n41917 );
buf U74574 ( n76345, n75700 );
not U74575 ( n528, n65801 );
buf U74576 ( n76525, n75702 );
buf U74577 ( n76267, n75703 );
buf U74578 ( n76201, n75701 );
buf U74579 ( n76802, n76799 );
nor U74580 ( n62555, n748, n747 );
not U74581 ( n748, n41919 );
nand U74582 ( n38441, n39930, n39931 );
not U74583 ( n4914, n13907 );
not U74584 ( n4957, n14293 );
buf U74585 ( n76605, n76601 );
buf U74586 ( n76474, n75704 );
and U74587 ( n39983, n38819, n38459 );
not U74588 ( n758, n62321 );
xnor U74589 ( n47483, n47480, n7583 );
not U74590 ( n757, n41936 );
nand U74591 ( n47330, n47431, n47297 );
nand U74592 ( n47431, n7572, n47432 );
nand U74593 ( n45406, n45752, n45758 );
nand U74594 ( n45758, n48080, n568 );
nand U74595 ( n61426, n41597, n61410 );
nand U74596 ( n26361, n26451, n26327 );
nand U74597 ( n26451, n4023, n26452 );
nand U74598 ( n59500, n59590, n59466 );
nand U74599 ( n59590, n6655, n59591 );
nand U74600 ( n68362, n68452, n68328 );
nand U74601 ( n68452, n5784, n68453 );
xnor U74602 ( n68504, n68501, n5795 );
xnor U74603 ( n26503, n26500, n4032 );
xnor U74604 ( n59642, n59639, n6664 );
xor U74605 ( n49569, n529, n665 );
not U74606 ( n744, n41918 );
not U74607 ( n2019, n36502 );
xnor U74608 ( n47300, n47297, n7563 );
nor U74609 ( n42002, n747, n692 );
xnor U74610 ( n68331, n68328, n5775 );
xnor U74611 ( n26330, n26327, n4017 );
xnor U74612 ( n59469, n59466, n6649 );
buf U74613 ( n76808, n2037 );
nand U74614 ( n37407, n37467, n37468 );
nor U74615 ( n37434, n37407, n37455 );
buf U74616 ( n76848, n613 );
buf U74617 ( n76475, n75704 );
not U74618 ( n773, n61586 );
not U74619 ( n1855, n38509 );
buf U74620 ( n76606, n76601 );
and U74621 ( n33782, n33866, n33745 );
nand U74622 ( n33866, n3209, n33867 );
nand U74623 ( n40017, n40014, n38792 );
not U74624 ( n655, n42059 );
not U74625 ( n1924, n37382 );
nor U74626 ( n37502, n2115, n2120 );
and U74627 ( n14187, n14292, n14140 );
nand U74628 ( n14292, n4942, n14293 );
nor U74629 ( n37452, n1985, n37454 );
nor U74630 ( n38885, n2132, n2137 );
nand U74631 ( n54629, n527, n45754 );
nand U74632 ( n33606, n33696, n33572 );
nand U74633 ( n33696, n3185, n33697 );
xnor U74634 ( n33748, n33745, n3197 );
not U74635 ( n569, n54915 );
buf U74636 ( n76858, n76854 );
buf U74637 ( n76854, n570 );
xor U74638 ( n54754, n66293, n41938 );
xnor U74639 ( n33575, n33572, n3177 );
and U74640 ( n40190, n38819, n38540 );
not U74641 ( n2013, n36436 );
not U74642 ( n1977, n39581 );
nand U74643 ( n13984, n14079, n13927 );
nand U74644 ( n14079, n4920, n14080 );
xnor U74645 ( n14144, n14140, n4929 );
or U74646 ( n37335, n37336, n1945 );
xnor U74647 ( n13930, n13927, n4913 );
nor U74648 ( n40225, n2000, n38555 );
nor U74649 ( n66434, n819, n54813 );
not U74650 ( n644, n41579 );
nor U74651 ( n66745, n820, n524 );
not U74652 ( n2015, n36438 );
not U74653 ( n2125, n38989 );
nor U74654 ( n39590, n1974, n39581 );
nor U74655 ( n66748, n833, n54868 );
not U74656 ( n630, n41959 );
buf U74657 ( n76336, n75753 );
not U74658 ( n577, n42198 );
nand U74659 ( n39887, n1944, n38792 );
not U74660 ( n2011, n36836 );
not U74661 ( n2050, n39349 );
nor U74662 ( n67008, n819, n54914 );
nor U74663 ( n40271, n1905, n2034 );
and U74664 ( n40309, n38819, n38585 );
buf U74665 ( n76811, n76813 );
buf U74666 ( n76819, n2028 );
buf U74667 ( n76818, n2028 );
nand U74668 ( n38108, n76811, n76409 );
nand U74669 ( n38791, n2144, n38792 );
buf U74670 ( n76820, n2028 );
nor U74671 ( n66741, n553, n823 );
buf U74672 ( n76338, n76337 );
buf U74673 ( n76339, n76337 );
nand U74674 ( n38568, n38570, n76444 );
buf U74675 ( n76340, n76337 );
not U74676 ( n2078, n37690 );
buf U74677 ( n76830, n2004 );
buf U74678 ( n76831, n2004 );
buf U74679 ( n76832, n2004 );
not U74680 ( n573, n45754 );
xor U74681 ( n47521, n47443, n7583 );
buf U74682 ( n76803, n76799 );
nor U74683 ( n47332, n47443, n7583 );
xor U74684 ( n33786, n33708, n3197 );
xor U74685 ( n26541, n26463, n4032 );
xor U74686 ( n59683, n59602, n6664 );
nand U74687 ( n38792, n37104, n37098 );
xor U74688 ( n68542, n68464, n5795 );
not U74689 ( n76374, n76375 );
nor U74690 ( n33608, n33708, n3197 );
nor U74691 ( n68364, n68464, n5795 );
nor U74692 ( n26363, n26463, n4032 );
nor U74693 ( n59502, n59602, n6664 );
not U74694 ( n578, n40884 );
xor U74695 ( n14192, n14094, n4929 );
not U74696 ( n76288, n76289 );
not U74697 ( n76449, n76450 );
nor U74698 ( n13963, n14094, n4929 );
not U74699 ( n76422, n76423 );
not U74700 ( n76421, n76423 );
xor U74701 ( n47293, n47240, n7563 );
buf U74702 ( n76812, n76813 );
buf U74703 ( n76809, n76814 );
buf U74704 ( n76810, n76814 );
xor U74705 ( n33568, n33516, n3177 );
xor U74706 ( n26323, n26270, n4017 );
xor U74707 ( n59462, n59409, n6649 );
xor U74708 ( n68324, n68271, n5775 );
not U74709 ( n76637, n75775 );
buf U74710 ( n76004, n76290 );
buf U74711 ( n76003, n76290 );
buf U74712 ( n76002, n76290 );
nand U74713 ( n25467, n28651, n4057 );
nor U74714 ( n28651, n4047, n28485 );
nand U74715 ( n58604, n61956, n6689 );
nor U74716 ( n61956, n6679, n61790 );
nand U74717 ( n67472, n70556, n5828 );
nor U74718 ( n70556, n5815, n70390 );
nand U74719 ( n32707, n35830, n3229 );
nor U74720 ( n35830, n3217, n35664 );
nand U74721 ( n22768, n4059, n4067 );
nand U74722 ( n55882, n6692, n6699 );
nand U74723 ( n64106, n5830, n5842 );
nand U74724 ( n30089, n3232, n3242 );
buf U74725 ( n76849, n613 );
buf U74726 ( n76014, n76424 );
buf U74727 ( n76012, n76424 );
buf U74728 ( n76013, n76424 );
buf U74729 ( n76805, n2062 );
buf U74730 ( n76806, n2062 );
buf U74731 ( n76850, n585 );
xor U74732 ( n13922, n13857, n4913 );
buf U74733 ( n76851, n585 );
not U74734 ( n76400, n75776 );
buf U74735 ( n76852, n585 );
nand U74736 ( n24606, n4060, n28565 );
nand U74737 ( n57738, n6693, n61870 );
nand U74738 ( n66414, n5832, n70470 );
nand U74739 ( n31822, n3233, n35744 );
nand U74740 ( n61859, n61939, n6639 );
nor U74741 ( n61939, n6659, n61940 );
nand U74742 ( n28554, n28634, n4007 );
nor U74743 ( n28634, n4027, n28635 );
nand U74744 ( n61940, n61942, n6679 );
nor U74745 ( n61942, n6610, n6668 );
nand U74746 ( n28635, n28637, n4047 );
nor U74747 ( n28637, n3978, n4035 );
not U74748 ( n3230, n29177 );
nand U74749 ( n70459, n70539, n5765 );
nor U74750 ( n70539, n5790, n70540 );
nand U74751 ( n70540, n70542, n5815 );
nor U74752 ( n70542, n5735, n5802 );
nand U74753 ( n35733, n35813, n3167 );
nor U74754 ( n35813, n3192, n35814 );
nand U74755 ( n35814, n35816, n3217 );
nor U74756 ( n35816, n3134, n3203 );
not U74757 ( n4058, n21864 );
not U74758 ( n7617, n42390 );
not U74759 ( n5829, n62899 );
not U74760 ( n6690, n54955 );
not U74761 ( n4007, n24316 );
not U74762 ( n6639, n57439 );
not U74763 ( n5765, n65898 );
not U74764 ( n3167, n31612 );
nor U74765 ( n35781, n35815, n35814 );
nand U74766 ( n35815, n3165, n3192 );
nor U74767 ( n70507, n70541, n70540 );
nand U74768 ( n70541, n5764, n5790 );
nor U74769 ( n28602, n28636, n28635 );
nand U74770 ( n28636, n4005, n4027 );
nor U74771 ( n61907, n61941, n61940 );
nand U74772 ( n61941, n6638, n6659 );
nor U74773 ( n54279, n54313, n54312 );
nand U74774 ( n54313, n7550, n7578 );
nand U74775 ( n54312, n54314, n7603 );
nor U74776 ( n54314, n7520, n7589 );
buf U74777 ( n76821, n2027 );
buf U74778 ( n76822, n2027 );
nand U74779 ( n61410, n41473, n41467 );
not U74780 ( n4963, n8304 );
buf U74781 ( n76823, n2027 );
nor U74782 ( n21287, n21330, n21329 );
nand U74783 ( n21330, n4902, n4925 );
nand U74784 ( n21329, n21331, n4949 );
nor U74785 ( n21331, n4875, n4935 );
not U74786 ( n4060, n22756 );
not U74787 ( n6693, n55870 );
not U74788 ( n5832, n64094 );
not U74789 ( n3233, n30077 );
not U74790 ( n3165, n34149 );
not U74791 ( n4005, n26904 );
not U74792 ( n5764, n68903 );
not U74793 ( n6638, n60044 );
not U74794 ( n7550, n47883 );
nand U74795 ( n47194, n47239, n47240 );
nor U74796 ( n47239, n7530, n7563 );
nand U74797 ( n38819, n2002, n2039 );
not U74798 ( n4902, n14653 );
not U74799 ( n3060, n32562 );
not U74800 ( n5662, n67327 );
not U74801 ( n3904, n25320 );
not U74802 ( n6537, n58459 );
not U74803 ( n7435, n46266 );
not U74804 ( n4792, n12638 );
nand U74805 ( n33474, n33515, n33516 );
nor U74806 ( n33515, n3143, n3177 );
nand U74807 ( n68225, n68270, n68271 );
nor U74808 ( n68270, n5744, n5775 );
nand U74809 ( n26224, n26269, n26270 );
nor U74810 ( n26269, n3987, n4017 );
nand U74811 ( n59363, n59408, n59409 );
nor U74812 ( n59408, n6619, n6649 );
not U74813 ( n76407, n76408 );
not U74814 ( n76406, n76408 );
nand U74815 ( n61439, n820, n833 );
not U74816 ( n820, n41469 );
nand U74817 ( n56203, n6610, n6659 );
nand U74818 ( n23082, n3978, n4027 );
nand U74819 ( n64572, n5735, n5790 );
nand U74820 ( n30413, n3134, n3192 );
nand U74821 ( n13807, n13855, n13857 );
nor U74822 ( n13855, n4885, n4913 );
nand U74823 ( n28560, n28568, n28569 );
nand U74824 ( n61865, n61873, n61874 );
nand U74825 ( n70465, n70473, n70474 );
nand U74826 ( n35739, n35747, n35748 );
nor U74827 ( n35780, n34149, n30089 );
nor U74828 ( n28601, n26904, n22768 );
nor U74829 ( n70506, n68903, n64106 );
nor U74830 ( n61906, n60044, n55882 );
and U74831 ( n34061, n35756, n35757 );
nor U74832 ( n35757, n35758, n35759 );
nor U74833 ( n35756, n35766, n35767 );
nand U74834 ( n35759, n35760, n35761 );
and U74835 ( n26816, n28577, n28578 );
nor U74836 ( n28578, n28579, n28580 );
nor U74837 ( n28577, n28587, n28588 );
nand U74838 ( n28580, n28581, n28582 );
and U74839 ( n68815, n70482, n70483 );
nor U74840 ( n70483, n70484, n70485 );
nor U74841 ( n70482, n70492, n70493 );
nand U74842 ( n70485, n70486, n70487 );
and U74843 ( n59956, n61882, n61883 );
nor U74844 ( n61883, n61884, n61885 );
nor U74845 ( n61882, n61892, n61893 );
nand U74846 ( n61885, n61886, n61887 );
nand U74847 ( n43362, n7618, n7629 );
nor U74848 ( n54278, n47883, n43362 );
and U74849 ( n47795, n54254, n54255 );
nor U74850 ( n54255, n54256, n54257 );
nor U74851 ( n54254, n54264, n54265 );
nand U74852 ( n54257, n54258, n54259 );
nor U74853 ( n30414, n35733, n30077 );
nor U74854 ( n23083, n28554, n22756 );
nor U74855 ( n64573, n70459, n64094 );
nor U74856 ( n56204, n61859, n55870 );
nor U74857 ( n43731, n54231, n43350 );
nand U74858 ( n54231, n54311, n7552 );
nor U74859 ( n54311, n7578, n54312 );
nor U74860 ( n35779, n29177, n31612 );
nor U74861 ( n28600, n21864, n24316 );
nor U74862 ( n70505, n62899, n65898 );
nor U74863 ( n61905, n54955, n57439 );
nor U74864 ( n54277, n42390, n44990 );
not U74865 ( n4967, n9420 );
nor U74866 ( n14634, n4878, n12833 );
nand U74867 ( n12835, n21290, n4963 );
not U74868 ( n7620, n43363 );
nor U74869 ( n47868, n7523, n46405 );
nand U74870 ( n9419, n4964, n4975 );
nor U74871 ( n21286, n14653, n9419 );
and U74872 ( n14543, n21261, n21262 );
nor U74873 ( n21262, n21263, n21264 );
nor U74874 ( n21261, n21272, n21273 );
nand U74875 ( n21264, n21265, n21266 );
nand U74876 ( n46407, n54242, n7617 );
buf U74877 ( n76781, n3042 );
buf U74878 ( n76763, n3885 );
buf U74879 ( n76715, n5643 );
buf U74880 ( n76696, n6518 );
buf U74881 ( n76667, n7418 );
buf U74882 ( n76782, n3042 );
buf U74883 ( n76716, n5643 );
buf U74884 ( n76668, n7418 );
buf U74885 ( n76764, n3885 );
buf U74886 ( n76697, n6518 );
buf U74887 ( n76669, n7418 );
buf U74888 ( n76765, n3885 );
buf U74889 ( n76698, n6518 );
and U74890 ( n75711, n3075, n3134 );
buf U74891 ( n76783, n3042 );
buf U74892 ( n76717, n5643 );
nor U74893 ( n9812, n21233, n9404 );
nand U74894 ( n21233, n21328, n4903 );
nor U74895 ( n21328, n4925, n21329 );
and U74896 ( n75712, n5677, n5735 );
and U74897 ( n75713, n7462, n7520 );
and U74898 ( n75714, n4818, n4875 );
and U74899 ( n75715, n3919, n3978 );
and U74900 ( n75716, n6552, n6610 );
nor U74901 ( n21285, n8304, n11310 );
not U74902 ( n4903, n11310 );
not U74903 ( n7552, n44990 );
buf U74904 ( n76734, n4774 );
buf U74905 ( n76735, n4774 );
buf U74906 ( n76736, n4774 );
nand U74907 ( n12837, n21345, n4962 );
nor U74908 ( n21345, n4949, n21179 );
nand U74909 ( n46408, n54328, n7615 );
nor U74910 ( n54328, n7603, n54162 );
not U74911 ( n3234, n30090 );
not U74912 ( n4062, n22769 );
not U74913 ( n5833, n64107 );
not U74914 ( n6694, n55883 );
nor U74915 ( n68888, n5738, n67469 );
nor U74916 ( n34134, n3137, n32704 );
nor U74917 ( n26889, n3980, n25464 );
nor U74918 ( n60029, n6613, n58601 );
and U74919 ( n64800, n41467, n41473 );
nand U74920 ( n32706, n35744, n3230 );
nand U74921 ( n25466, n28565, n4058 );
nand U74922 ( n67471, n70470, n5829 );
nand U74923 ( n58603, n61870, n6690 );
nand U74924 ( n35764, n3167, n3192 );
nand U74925 ( n28585, n4007, n4027 );
nand U74926 ( n70490, n5765, n5790 );
nand U74927 ( n61890, n6639, n6659 );
nand U74928 ( n35758, n35763, n35764 );
nand U74929 ( n35763, n35765, n3183 );
nor U74930 ( n35765, n3169, n35748 );
nand U74931 ( n28579, n28584, n28585 );
nand U74932 ( n28584, n28586, n4020 );
nor U74933 ( n28586, n4009, n28569 );
nand U74934 ( n70484, n70489, n70490 );
nand U74935 ( n70489, n70491, n5782 );
nor U74936 ( n70491, n5768, n70474 );
nand U74937 ( n61884, n61889, n61890 );
nand U74938 ( n61889, n61891, n6653 );
nor U74939 ( n61891, n6642, n61874 );
nand U74940 ( n54262, n7552, n7578 );
nand U74941 ( n54256, n54261, n54262 );
nand U74942 ( n54261, n54263, n7569 );
nor U74943 ( n54263, n7554, n54246 );
nand U74944 ( n26910, n28611, n28612 );
nand U74945 ( n28612, n4007, n4058 );
nor U74946 ( n28611, n28613, n28614 );
nor U74947 ( n28614, n4047, n28615 );
nand U74948 ( n60050, n61916, n61917 );
nand U74949 ( n61917, n6639, n6690 );
nor U74950 ( n61916, n61918, n61919 );
nor U74951 ( n61919, n6679, n61920 );
nor U74952 ( n28619, n28568, n28621 );
nor U74953 ( n28621, n4027, n4007 );
nor U74954 ( n61924, n61873, n61926 );
nor U74955 ( n61926, n6659, n6639 );
nand U74956 ( n34155, n35790, n35791 );
nand U74957 ( n35791, n3167, n3230 );
nor U74958 ( n35790, n35792, n35793 );
nor U74959 ( n35793, n3217, n35794 );
nor U74960 ( n35798, n35747, n35800 );
nor U74961 ( n35800, n3192, n3167 );
nand U74962 ( n68909, n70516, n70517 );
nand U74963 ( n70517, n5765, n5829 );
nor U74964 ( n70516, n70518, n70519 );
nor U74965 ( n70519, n5815, n70520 );
nor U74966 ( n70524, n70473, n70526 );
nor U74967 ( n70526, n5790, n5765 );
not U74968 ( n224, n9908 );
not U74969 ( n495, n43808 );
buf U74970 ( n76283, n75755 );
buf U74971 ( n76541, n75756 );
buf U74972 ( n76484, n75758 );
buf U74973 ( n76217, n75757 );
nor U74974 ( n35713, n34062, n35781 );
nor U74975 ( n28534, n26817, n28602 );
nor U74976 ( n70439, n68816, n70507 );
nor U74977 ( n61839, n59957, n61907 );
nor U74978 ( n54211, n47796, n54279 );
nand U74979 ( n47889, n54288, n54289 );
nand U74980 ( n54289, n7552, n7617 );
nor U74981 ( n54288, n54290, n54291 );
nor U74982 ( n54291, n7603, n54292 );
nor U74983 ( n54296, n54245, n54298 );
nor U74984 ( n54298, n7578, n7552 );
nand U74985 ( n21269, n4903, n4925 );
nand U74986 ( n21263, n21268, n21269 );
nand U74987 ( n21268, n21270, n4918 );
nor U74988 ( n21270, n4905, n21271 );
nand U74989 ( n11748, n4965, n21290 );
nand U74990 ( n14660, n21305, n21306 );
nand U74991 ( n21306, n4903, n4963 );
nor U74992 ( n21305, n21307, n21308 );
nor U74993 ( n21308, n4949, n21309 );
nor U74994 ( n21313, n21293, n21315 );
nor U74995 ( n21315, n4925, n4903 );
nand U74996 ( n45521, n7619, n54242 );
nor U74997 ( n35766, n3165, n30090 );
nor U74998 ( n28587, n4005, n22769 );
nor U74999 ( n70492, n5764, n64107 );
nor U75000 ( n61892, n6638, n55883 );
nor U75001 ( n54264, n7550, n43363 );
nor U75002 ( n21248, n14544, n21287 );
nand U75003 ( n11508, n76619, n4964 );
nor U75004 ( n12679, n4858, n9404 );
nor U75005 ( n32588, n3117, n30077 );
nor U75006 ( n67353, n5718, n64094 );
nor U75007 ( n25346, n3960, n22756 );
nor U75008 ( n58485, n6593, n55870 );
nor U75009 ( n46292, n7504, n43350 );
nor U75010 ( n30412, n30077, n30413 );
nand U75011 ( n24466, n76533, n4059 );
nand U75012 ( n57595, n76275, n6692 );
nand U75013 ( n43730, n7520, n7578 );
nand U75014 ( n9810, n4875, n4925 );
nor U75015 ( n64571, n64094, n64572 );
nor U75016 ( n43729, n43350, n43730 );
nor U75017 ( n9809, n9404, n9810 );
nand U75018 ( n66168, n76209, n5830 );
nor U75019 ( n23081, n22756, n23082 );
nor U75020 ( n56202, n55870, n56203 );
nand U75021 ( n21239, n21293, n21271 );
nand U75022 ( n54237, n54245, n54246 );
nand U75023 ( n45328, n76353, n7618 );
nor U75024 ( n21272, n4902, n9420 );
nor U75025 ( n28622, n4035, n4062 );
nor U75026 ( n61927, n6668, n6694 );
nor U75027 ( n35801, n3203, n3234 );
nor U75028 ( n70527, n5802, n5833 );
not U75029 ( n478, n63068 );
not U75030 ( n207, n29301 );
not U75031 ( n445, n55096 );
not U75032 ( n173, n21986 );
nor U75033 ( n54299, n7589, n7620 );
nor U75034 ( n40321, n76797, n76409 );
not U75035 ( n4965, n9404 );
not U75036 ( n7619, n43350 );
nor U75037 ( n21316, n4935, n4967 );
not U75038 ( n76618, n76619 );
not U75039 ( n76274, n76275 );
not U75040 ( n76532, n76533 );
not U75041 ( n76208, n76209 );
not U75042 ( n76352, n76353 );
nand U75043 ( n34136, n35738, n3168 );
nor U75044 ( n35738, n3134, n30089 );
nand U75045 ( n26891, n28559, n4008 );
nor U75046 ( n28559, n3978, n22768 );
nand U75047 ( n68890, n70464, n5767 );
nor U75048 ( n70464, n5735, n64106 );
nand U75049 ( n60031, n61864, n6640 );
nor U75050 ( n61864, n6610, n55882 );
nand U75051 ( n47870, n54236, n7553 );
nor U75052 ( n54236, n7520, n43362 );
nand U75053 ( n28620, n4067, n4027 );
nand U75054 ( n61925, n6699, n6659 );
nand U75055 ( n35799, n3242, n3192 );
nand U75056 ( n70525, n5842, n5790 );
nand U75057 ( n54297, n7629, n7578 );
not U75058 ( n4045, n26906 );
not U75059 ( n6678, n60046 );
not U75060 ( n3215, n34151 );
not U75061 ( n5814, n68905 );
nand U75062 ( n21314, n4975, n4925 );
nand U75063 ( n12775, n14542, n14543 );
nor U75064 ( n14542, n14544, n14545 );
nor U75065 ( n14545, n4858, n9420 );
nand U75066 ( n46365, n47794, n47795 );
nor U75067 ( n47794, n47796, n47797 );
nor U75068 ( n47797, n7504, n43363 );
nand U75069 ( n14637, n21238, n4904 );
nor U75070 ( n21238, n4875, n9419 );
buf U75071 ( n76399, n76396 );
buf U75072 ( n76395, n76392 );
buf U75073 ( n76398, n76396 );
buf U75074 ( n76397, n76396 );
nand U75075 ( n67429, n68814, n68815 );
nor U75076 ( n68814, n68816, n68817 );
nor U75077 ( n68817, n5718, n64107 );
nand U75078 ( n32664, n34060, n34061 );
nor U75079 ( n34060, n34062, n34063 );
nor U75080 ( n34063, n3117, n30090 );
nand U75081 ( n25424, n26815, n26816 );
nor U75082 ( n26815, n26817, n26818 );
nor U75083 ( n26818, n3960, n22769 );
nand U75084 ( n58561, n59955, n59956 );
nor U75085 ( n59955, n59957, n59958 );
nor U75086 ( n59958, n6593, n55883 );
not U75087 ( n3095, n32911 );
not U75088 ( n5697, n67672 );
not U75089 ( n3939, n25667 );
not U75090 ( n6572, n58807 );
not U75091 ( n4828, n13239 );
not U75092 ( n4839, n13095 );
not U75093 ( n7482, n46625 );
not U75094 ( n174, n22036 );
not U75095 ( n446, n55146 );
not U75096 ( n479, n63118 );
not U75097 ( n208, n29355 );
nor U75098 ( n31611, n3244, n76486 );
nor U75099 ( n65897, n5844, n76219 );
buf U75100 ( n76486, n76485 );
buf U75101 ( n76219, n76218 );
nor U75102 ( n31542, n3143, n76486 );
nor U75103 ( n65792, n5744, n76219 );
nor U75104 ( n31553, n3177, n76486 );
nor U75105 ( n31574, n3197, n76486 );
nor U75106 ( n65843, n5775, n76219 );
nor U75107 ( n65864, n5795, n76219 );
nor U75108 ( n31563, n3185, n76486 );
nor U75109 ( n31587, n3209, n76486 );
nor U75110 ( n65853, n5784, n76219 );
nor U75111 ( n65873, n5808, n76219 );
nor U75112 ( n31598, n3223, n76486 );
nor U75113 ( n65884, n5822, n76219 );
buf U75114 ( n76487, n76485 );
buf U75115 ( n76220, n76218 );
nor U75116 ( n30755, n30184, n76487 );
nor U75117 ( n64957, n64250, n76220 );
buf U75118 ( n76488, n76485 );
buf U75119 ( n76221, n76218 );
nor U75120 ( n30484, n30129, n76488 );
nor U75121 ( n30527, n30139, n76488 );
nor U75122 ( n30572, n30147, n76488 );
nor U75123 ( n30617, n30155, n76488 );
nor U75124 ( n30662, n30165, n76488 );
nor U75125 ( n30706, n30174, n76488 );
nor U75126 ( n64643, n64142, n76221 );
nor U75127 ( n64686, n64152, n76221 );
nor U75128 ( n64731, n64160, n76221 );
nor U75129 ( n64823, n64168, n76221 );
nor U75130 ( n64868, n64178, n76221 );
nor U75131 ( n64912, n64240, n76221 );
nor U75132 ( n11309, n4978, n76630 );
nor U75133 ( n44989, n7632, n76360 );
buf U75134 ( n76360, n76359 );
buf U75135 ( n76630, n76629 );
not U75136 ( n3094, n33137 );
not U75137 ( n5695, n67893 );
not U75138 ( n3938, n25890 );
not U75139 ( n6570, n59028 );
nor U75140 ( n44927, n7530, n76360 );
nor U75141 ( n11225, n4885, n76630 );
nor U75142 ( n44938, n7563, n76360 );
nor U75143 ( n11239, n4913, n76630 );
nor U75144 ( n44957, n7583, n76360 );
nor U75145 ( n11269, n4929, n76630 );
nor U75146 ( n11257, n4920, n76630 );
nor U75147 ( n11283, n4942, n76630 );
nor U75148 ( n44947, n7572, n76360 );
nor U75149 ( n44968, n7595, n76360 );
nor U75150 ( n11293, n4955, n76630 );
nor U75151 ( n44976, n7609, n76360 );
buf U75152 ( n76631, n76629 );
buf U75153 ( n76361, n76359 );
buf U75154 ( n76632, n76629 );
buf U75155 ( n76362, n76359 );
not U75156 ( n4838, n13385 );
not U75157 ( n7480, n46846 );
not U75158 ( n5687, n67774 );
not U75159 ( n7472, n46727 );
not U75160 ( n3929, n25771 );
not U75161 ( n6562, n58909 );
not U75162 ( n3085, n33018 );
not U75163 ( n505, n42577 );
not U75164 ( n234, n8509 );
not U75165 ( n3120, n33181 );
not U75166 ( n3104, n32604 );
not U75167 ( n5705, n67369 );
not U75168 ( n3948, n25364 );
not U75169 ( n6580, n58501 );
not U75170 ( n4862, n13440 );
not U75171 ( n4849, n12887 );
not U75172 ( n7492, n46453 );
not U75173 ( n7832, n48719 );
not U75174 ( n3915, n22798 );
not U75175 ( n6548, n55912 );
not U75176 ( n164, n23096 );
not U75177 ( n437, n56217 );
nor U75178 ( n28483, n28484, n28485 );
nor U75179 ( n28484, n4062, n4057 );
nor U75180 ( n61788, n61789, n61790 );
nor U75181 ( n61789, n6694, n6689 );
nor U75182 ( n35662, n35663, n35664 );
nor U75183 ( n35663, n3234, n3229 );
nor U75184 ( n70388, n70389, n70390 );
nor U75185 ( n70389, n5833, n5828 );
nor U75186 ( n21177, n21178, n21179 );
nor U75187 ( n21178, n4967, n4962 );
nor U75188 ( n54156, n54157, n54158 );
nor U75189 ( n54157, n7619, n7617 );
nor U75190 ( n12824, n12833, n12834 );
nand U75191 ( n12834, n12835, n12837 );
nor U75192 ( n46394, n46405, n46406 );
nand U75193 ( n46406, n46407, n46408 );
not U75194 ( n7602, n47885 );
not U75195 ( n4948, n14655 );
nand U75196 ( n31181, n31116, n31612 );
nand U75197 ( n65435, n65370, n65898 );
nand U75198 ( n57007, n56949, n57439 );
nand U75199 ( n23883, n23825, n24316 );
nand U75200 ( n23152, n23825, n4020 );
nand U75201 ( n56273, n56949, n6653 );
nand U75202 ( n30481, n31116, n3183 );
nand U75203 ( n64640, n65370, n5782 );
nand U75204 ( n10785, n10695, n11310 );
nand U75205 ( n44561, n44494, n44990 );
nor U75206 ( n67458, n67469, n67470 );
nand U75207 ( n67470, n67471, n67472 );
nor U75208 ( n32693, n32704, n32705 );
nand U75209 ( n32705, n32706, n32707 );
nor U75210 ( n25453, n25464, n25465 );
nand U75211 ( n25465, n25466, n25467 );
nor U75212 ( n58590, n58601, n58602 );
nand U75213 ( n58602, n58603, n58604 );
nand U75214 ( n43799, n44494, n7569 );
nand U75215 ( n9897, n10695, n4918 );
not U75216 ( n4869, n13003 );
not U75217 ( n5729, n67634 );
not U75218 ( n3972, n25629 );
not U75219 ( n6604, n58766 );
not U75220 ( n3128, n32873 );
nor U75221 ( n23251, n22822, n23096 );
nor U75222 ( n56375, n55936, n56217 );
nor U75223 ( n56518, n55966, n56217 );
nor U75224 ( n23396, n22849, n23096 );
buf U75225 ( n76628, n75759 );
not U75226 ( n5724, n67913 );
not U75227 ( n7510, n46866 );
not U75228 ( n3967, n25910 );
not U75229 ( n6599, n59048 );
nand U75230 ( n13060, n4885, n12679 );
buf U75231 ( n76393, n76392 );
buf U75232 ( n76394, n76392 );
not U75233 ( n4867, n13152 );
not U75234 ( n7513, n46663 );
not U75235 ( n5727, n67710 );
not U75236 ( n3125, n32956 );
not U75237 ( n3969, n25705 );
not U75238 ( n6602, n58845 );
nand U75239 ( n67479, n5744, n67353 );
nand U75240 ( n32714, n3143, n32588 );
nand U75241 ( n25474, n3987, n25346 );
nand U75242 ( n58611, n6619, n58485 );
nand U75243 ( n46415, n7530, n46292 );
nand U75244 ( n31728, n217, n3232 );
not U75245 ( n3072, n30123 );
not U75246 ( n5673, n64136 );
not U75247 ( n7458, n43392 );
not U75248 ( n4814, n9457 );
nand U75249 ( n14482, n13060, n12887 );
nand U75250 ( n68767, n67479, n67369 );
nand U75251 ( n34011, n32714, n32604 );
nand U75252 ( n26768, n25474, n25364 );
nand U75253 ( n59908, n58611, n58501 );
nand U75254 ( n47746, n46415, n46453 );
not U75255 ( n933, n13650 );
not U75256 ( n4756, n14854 );
not U75257 ( n7400, n48051 );
nand U75258 ( n16519, n5195, n4756 );
nand U75259 ( n49507, n7850, n7400 );
not U75260 ( n4755, n14868 );
not U75261 ( n7399, n48062 );
nand U75262 ( n16555, n5195, n4755 );
nand U75263 ( n49536, n7850, n7399 );
not U75264 ( n7402, n48040 );
not U75265 ( n4757, n14840 );
nand U75266 ( n49474, n7850, n7402 );
nand U75267 ( n16478, n5195, n4757 );
not U75268 ( n4754, n14882 );
not U75269 ( n7398, n48087 );
nand U75270 ( n16593, n5195, n4754 );
nand U75271 ( n49582, n7850, n7398 );
not U75272 ( n4753, n14895 );
not U75273 ( n7397, n48098 );
nand U75274 ( n16629, n5195, n4753 );
nand U75275 ( n49610, n7850, n7397 );
not U75276 ( n4758, n14824 );
not U75277 ( n7403, n48027 );
nand U75278 ( n16440, n5195, n4758 );
nand U75279 ( n49443, n7850, n7403 );
not U75280 ( n7395, n48109 );
not U75281 ( n4752, n14909 );
nand U75282 ( n49639, n7850, n7395 );
nand U75283 ( n16665, n5195, n4752 );
nand U75284 ( n49885, n50283, n50284 );
nand U75285 ( n50284, n1757, n50285 );
nand U75286 ( n50283, n50288, n49914 );
not U75287 ( n1757, n49914 );
nand U75288 ( n49713, n50066, n50067 );
nand U75289 ( n50067, n1363, n50068 );
nand U75290 ( n50066, n50071, n50037 );
not U75291 ( n1363, n50037 );
nand U75292 ( n49952, n50259, n50260 );
nand U75293 ( n50259, n50263, n49878 );
nand U75294 ( n50260, n1739, n50261 );
nand U75295 ( n50263, n49875, n49877 );
nand U75296 ( n49962, n50236, n50237 );
nand U75297 ( n50236, n50241, n49956 );
nand U75298 ( n50237, n1718, n50238 );
nand U75299 ( n50241, n49953, n49955 );
nor U75300 ( n49858, n1717, n1712 );
nor U75301 ( n49768, n1575, n1573 );
nand U75302 ( n49755, n50094, n50095 );
nand U75303 ( n50095, n1532, n50096 );
nand U75304 ( n50094, n50099, n50000 );
not U75305 ( n1532, n50000 );
not U75306 ( n1639, n49797 );
not U75307 ( n1674, n49822 );
not U75308 ( n1607, n49780 );
not U75309 ( n1575, n49996 );
nor U75310 ( n50229, n50230, n49960 );
nor U75311 ( n50230, n49858, n49859 );
nor U75312 ( n50158, n50159, n50156 );
nor U75313 ( n50159, n50160, n49803 );
nor U75314 ( n50160, n1639, n1637 );
nor U75315 ( n50182, n50183, n50180 );
nor U75316 ( n50183, n50184, n49828 );
nor U75317 ( n50184, n1674, n1670 );
nor U75318 ( n50134, n50135, n50132 );
nor U75319 ( n50135, n50136, n49786 );
nor U75320 ( n50136, n1607, n1604 );
nor U75321 ( n50058, n50059, n50056 );
nor U75322 ( n50059, n50060, n49718 );
nor U75323 ( n50060, n1362, n1357 );
nand U75324 ( n49693, n50042, n50043 );
nand U75325 ( n50042, n50046, n49703 );
nand U75326 ( n50043, n1279, n50044 );
nand U75327 ( n50046, n49700, n49702 );
not U75328 ( n1745, n50270 );
not U75329 ( n1320, n50053 );
not U75330 ( n1760, n49908 );
nand U75331 ( n50071, n50035, n50038 );
nand U75332 ( n50288, n49912, n49915 );
nand U75333 ( n50099, n49997, n49999 );
nand U75334 ( n50207, n49844, n49973 );
nand U75335 ( n49699, n49700, n49701 );
nand U75336 ( n49701, n49702, n49703 );
nand U75337 ( n50273, n50279, n50280 );
nand U75338 ( n50280, n50281, n50282 );
not U75339 ( n76323, n75778 );
nand U75340 ( n50061, n49713, n50056 );
not U75341 ( n1693, n49844 );
nand U75342 ( n50137, n49780, n50132 );
nand U75343 ( n50161, n49797, n50156 );
nand U75344 ( n50185, n49822, n50180 );
nand U75345 ( n16757, n17112, n17113 );
nand U75346 ( n17112, n17116, n17083 );
nand U75347 ( n17113, n2479, n17114 );
nand U75348 ( n17116, n17081, n17084 );
nand U75349 ( n16997, n17313, n17314 );
nand U75350 ( n17313, n17317, n16923 );
nand U75351 ( n17314, n2857, n17315 );
nand U75352 ( n17317, n16920, n16922 );
nand U75353 ( n17007, n17290, n17291 );
nand U75354 ( n17290, n17295, n17001 );
nand U75355 ( n17291, n2835, n17292 );
nand U75356 ( n17295, n16998, n17000 );
nor U75357 ( n16903, n2834, n2829 );
nor U75358 ( n16813, n2697, n2694 );
nand U75359 ( n16800, n17148, n17149 );
nand U75360 ( n17149, n2653, n17150 );
nand U75361 ( n17148, n17153, n17046 );
not U75362 ( n2653, n17046 );
not U75363 ( n2608, n17057 );
not U75364 ( n2870, n16930 );
not U75365 ( n2763, n16842 );
not U75366 ( n2793, n16867 );
not U75367 ( n2728, n16825 );
not U75368 ( n2697, n17042 );
nor U75369 ( n17283, n17284, n17005 );
nor U75370 ( n17284, n16903, n16904 );
nor U75371 ( n17329, n17330, n17327 );
nor U75372 ( n17330, n17331, n16935 );
nor U75373 ( n17331, n2870, n2868 );
nor U75374 ( n17212, n17213, n17210 );
nor U75375 ( n17213, n17214, n16848 );
nor U75376 ( n17214, n2763, n2760 );
nor U75377 ( n17236, n17237, n17234 );
nor U75378 ( n17237, n17238, n16873 );
nor U75379 ( n17238, n2793, n2790 );
nor U75380 ( n17188, n17189, n17186 );
nor U75381 ( n17189, n17190, n16831 );
nor U75382 ( n17190, n2728, n2725 );
nor U75383 ( n17104, n17105, n17102 );
nor U75384 ( n17105, n17106, n16762 );
nor U75385 ( n17106, n2478, n2474 );
nand U75386 ( n16737, n17088, n17089 );
nand U75387 ( n17088, n17092, n16747 );
nand U75388 ( n17089, n2394, n17090 );
nand U75389 ( n17092, n16744, n16746 );
not U75390 ( n2514, n17123 );
not U75391 ( n2863, n17324 );
not U75392 ( n2438, n17099 );
not U75393 ( n2877, n16953 );
nand U75394 ( n17153, n17043, n17045 );
nand U75395 ( n17261, n16889, n17019 );
nand U75396 ( n50268, n50515, n50516 );
nand U75397 ( n50515, n50520, n50282 );
nand U75398 ( n50516, n1748, n50517 );
nand U75399 ( n50520, n50279, n50281 );
not U75400 ( n1739, n49878 );
nand U75401 ( n49930, n76653, n76648 );
nand U75402 ( n50297, n49903, n49905 );
nand U75403 ( n16743, n16744, n16745 );
nand U75404 ( n16745, n16746, n16747 );
nand U75405 ( n17332, n16930, n17327 );
not U75406 ( n2864, n17327 );
nor U75407 ( n16931, n2868, n2864 );
not U75408 ( n76589, n75779 );
nand U75409 ( n16659, n17402, n17403 );
nand U75410 ( n17403, n17381, n17384 );
nor U75411 ( n17402, n17405, n17406 );
nor U75412 ( n17405, n17384, n17408 );
xnor U75413 ( n20421, n20528, n20448 );
xor U75414 ( n20528, n20449, n2648 );
nand U75415 ( n18203, n18561, n18562 );
nor U75416 ( n18561, n18563, n18564 );
nor U75417 ( n20419, n2622, n2639 );
nor U75418 ( n19843, n2542, n2554 );
not U75419 ( n2688, n20626 );
nand U75420 ( n18185, n18200, n18201 );
nand U75421 ( n18201, n18202, n18203 );
nor U75422 ( n18204, n2510, n18209 );
nand U75423 ( n20452, n20453, n20454 );
nor U75424 ( n20453, n20419, n20413 );
nor U75425 ( n20707, n2693, n2702 );
not U75426 ( n2812, n16889 );
nand U75427 ( n17239, n16867, n17234 );
nand U75428 ( n17191, n16825, n17186 );
nand U75429 ( n17215, n16842, n17210 );
or U75430 ( n18209, n2520, n18203 );
not U75431 ( n2520, n18208 );
nand U75432 ( n17107, n16757, n17102 );
not U75433 ( n1748, n50282 );
nand U75434 ( n49950, n50255, n50256 );
nand U75435 ( n50256, n50257, n50258 );
not U75436 ( n2397, n17683 );
nor U75437 ( n20706, n2693, n2689 );
and U75438 ( n20699, n20757, n20758 );
nand U75439 ( n20758, n20707, n2689 );
nor U75440 ( n20757, n20759, n20760 );
nor U75441 ( n20759, n2702, n20764 );
nor U75442 ( n50350, n1247, n50351 );
nor U75443 ( n52672, n1423, n1435 );
not U75444 ( n1567, n53497 );
not U75445 ( n1435, n52674 );
not U75446 ( n1282, n50862 );
not U75447 ( n1518, n53385 );
nand U75448 ( n51141, n51156, n51157 );
nor U75449 ( n51156, n51160, n51161 );
nor U75450 ( n51160, n1393, n51165 );
nand U75451 ( n53310, n53311, n53312 );
nand U75452 ( n51159, n51517, n51518 );
nor U75453 ( n51517, n51519, n51520 );
nand U75454 ( n52789, n52928, n52929 );
nand U75455 ( n52929, n52674, n52670 );
nor U75456 ( n52928, n52672, n52666 );
nand U75457 ( n49560, n50598, n50599 );
not U75458 ( n1400, n51164 );
not U75459 ( n1325, n50909 );
not U75460 ( n1434, n53057 );
nand U75461 ( n52787, n53045, n53046 );
nand U75462 ( n53046, n53047, n1434 );
nor U75463 ( n53045, n53048, n53049 );
and U75464 ( n53049, n1464, n53050 );
nor U75465 ( n52648, n1389, n1405 );
nor U75466 ( n52177, n1309, n1332 );
nor U75467 ( n51823, n1265, n1288 );
nand U75468 ( n52333, n52640, n52641 );
nand U75469 ( n52641, n52642, n1405 );
nor U75470 ( n52640, n52643, n52644 );
nor U75471 ( n52643, n1405, n52651 );
nand U75472 ( n50620, n51849, n51850 );
nand U75473 ( n51850, n1252, n50882 );
nor U75474 ( n51849, n51851, n51852 );
not U75475 ( n1252, n50879 );
nor U75476 ( n20804, n2669, n2687 );
not U75477 ( n2640, n20527 );
nand U75478 ( n20512, n20846, n20847 );
nand U75479 ( n20847, n20805, n2687 );
nor U75480 ( n20846, n20849, n20850 );
nor U75481 ( n20849, n2687, n20853 );
nor U75482 ( n17395, n16620, n16622 );
nand U75483 ( n16587, n17643, n17644 );
nor U75484 ( n17643, n17645, n17646 );
nand U75485 ( n19831, n20089, n20090 );
nand U75486 ( n20090, n20091, n2555 );
nor U75487 ( n20089, n20092, n20093 );
and U75488 ( n20093, n2587, n20094 );
xor U75489 ( n53386, n1527, n53387 );
nor U75490 ( n53273, n1500, n1517 );
not U75491 ( n2443, n17952 );
nor U75492 ( n51901, n1479, n1487 );
nand U75493 ( n51890, n52370, n52371 );
nand U75494 ( n52371, n51902, n1487 );
nor U75495 ( n52370, n52373, n52374 );
nor U75496 ( n52373, n1487, n52377 );
not U75497 ( n1538, n52393 );
not U75498 ( n1614, n53702 );
nand U75499 ( n52920, n53055, n53056 );
nand U75500 ( n53056, n53053, n53057 );
nor U75501 ( n53055, n53047, n53050 );
nand U75502 ( n49634, n50357, n50358 );
nand U75503 ( n50358, n50336, n50339 );
nor U75504 ( n50357, n50360, n50361 );
nor U75505 ( n50360, n50339, n50363 );
nand U75506 ( n53396, n53309, n53308 );
nor U75507 ( n19716, n2543, n2557 );
nor U75508 ( n20643, n2709, n2717 );
nand U75509 ( n20637, n20708, n20709 );
nand U75510 ( n20709, n20644, n2717 );
nor U75511 ( n20708, n20711, n20712 );
nor U75512 ( n20711, n2717, n20715 );
not U75513 ( n2442, n18188 );
or U75514 ( n17959, n2482, n17900 );
not U75515 ( n2482, n17901 );
nor U75516 ( n20203, n2598, n2615 );
not U75517 ( n2615, n20207 );
nand U75518 ( n20215, n20332, n20333 );
nand U75519 ( n20333, n20207, n20211 );
nor U75520 ( n20332, n20209, n20203 );
not U75521 ( n1565, n53561 );
not U75522 ( n1544, n53380 );
nor U75523 ( n53643, n53644, n53645 );
nand U75524 ( n19696, n19835, n19836 );
nand U75525 ( n19836, n19837, n2554 );
nor U75526 ( n19835, n19838, n19839 );
nor U75527 ( n19838, n2554, n19846 );
nor U75528 ( n53159, n1478, n1492 );
not U75529 ( n1492, n53163 );
nand U75530 ( n53171, n53186, n53187 );
nand U75531 ( n53187, n53163, n53167 );
nor U75532 ( n53186, n53165, n53159 );
not U75533 ( n2523, n18700 );
xor U75534 ( n52831, n52393, n52392 );
nand U75535 ( n53395, n53408, n53409 );
nand U75536 ( n53409, n53410, n1542 );
nor U75537 ( n53408, n53411, n53412 );
nor U75538 ( n53412, n53413, n1540 );
not U75539 ( n1464, n53053 );
not U75540 ( n2857, n16923 );
nor U75541 ( n52342, n1350, n1370 );
or U75542 ( n49717, n49718, n1322 );
xor U75543 ( n50638, n1282, n1249 );
not U75544 ( n1247, n49603 );
nor U75545 ( n20209, n2598, n2589 );
not U75546 ( n2617, n20410 );
not U75547 ( n2589, n20211 );
and U75548 ( n20072, n20201, n20202 );
nand U75549 ( n20202, n20203, n2589 );
nor U75550 ( n20201, n20204, n20205 );
nor U75551 ( n20204, n2615, n20212 );
and U75552 ( n20395, n20500, n20501 );
nand U75553 ( n20501, n20502, n2643 );
nor U75554 ( n20500, n20503, n20504 );
nor U75555 ( n20503, n2668, n20511 );
nand U75556 ( n52912, n53506, n53507 );
nand U75557 ( n53507, n53413, n53417 );
nor U75558 ( n53506, n53410, n53414 );
nand U75559 ( n52638, n52664, n52665 );
nand U75560 ( n52665, n52666, n1435 );
nor U75561 ( n52664, n52667, n52668 );
nor U75562 ( n52667, n1435, n52675 );
nor U75563 ( n52183, n1309, n1289 );
nor U75564 ( n51829, n1265, n1254 );
nand U75565 ( n51819, n52175, n52176 );
nand U75566 ( n52176, n52177, n1289 );
nor U75567 ( n52175, n52178, n52179 );
nor U75568 ( n52178, n1332, n52186 );
nand U75569 ( n20213, n20411, n20412 );
nand U75570 ( n20412, n20413, n2639 );
nor U75571 ( n20411, n20414, n20415 );
nor U75572 ( n20414, n2639, n20422 );
nand U75573 ( n52187, n52334, n52335 );
nand U75574 ( n52335, n52336, n1370 );
nor U75575 ( n52334, n52337, n52338 );
nor U75576 ( n52337, n1370, n52345 );
not U75577 ( n1534, n53400 );
not U75578 ( n1270, n50601 );
not U75579 ( n1459, n51513 );
not U75580 ( n1462, n51652 );
nor U75581 ( n52526, n1390, n1408 );
nand U75582 ( n52639, n52676, n52677 );
nand U75583 ( n52677, n52530, n52534 );
nor U75584 ( n52676, n52526, n52532 );
not U75585 ( n1408, n52530 );
nand U75586 ( n52651, n1389, n52646 );
nand U75587 ( n50246, n50497, n50498 );
nand U75588 ( n50497, n50502, n50258 );
nand U75589 ( n50498, n1728, n50499 );
nand U75590 ( n50502, n50255, n50257 );
not U75591 ( n1718, n49956 );
nand U75592 ( n53173, n53282, n53283 );
nand U75593 ( n53283, n53284, n1512 );
nor U75594 ( n53282, n53286, n53287 );
not U75595 ( n1512, n53285 );
nor U75596 ( n19692, n2505, n2525 );
nand U75597 ( n53169, n53265, n53266 );
nand U75598 ( n53266, n53267, n1517 );
nor U75599 ( n53265, n53268, n53269 );
nor U75600 ( n53268, n1517, n53276 );
nand U75601 ( n50781, n50810, n50811 );
nand U75602 ( n50811, n50812, n50813 );
nand U75603 ( n50258, n50503, n50504 );
nand U75604 ( n50503, n50505, n50506 );
not U75605 ( n1735, n51045 );
nor U75606 ( n20348, n2623, n2644 );
and U75607 ( n18214, n18901, n18902 );
nand U75608 ( n18902, n18564, n2519 );
nor U75609 ( n18901, n18906, n18907 );
not U75610 ( n2519, n18903 );
not U75611 ( n1601, n53631 );
nand U75612 ( n52652, n52791, n52792 );
nor U75613 ( n52791, n52794, n52795 );
or U75614 ( n50917, n1365, n50855 );
not U75615 ( n1365, n50856 );
nor U75616 ( n20446, n20449, n20448 );
nand U75617 ( n20217, n20428, n20429 );
nand U75618 ( n20429, n20323, n2634 );
nor U75619 ( n20428, n20433, n20434 );
not U75620 ( n2634, n20430 );
nand U75621 ( n20534, n20451, n20450 );
nor U75622 ( n51158, n1393, n51164 );
nand U75623 ( n53417, n53428, n53508 );
nand U75624 ( n53508, n53429, n53426 );
not U75625 ( n1540, n53414 );
nor U75626 ( n53165, n1478, n1467 );
nand U75627 ( n53250, n53358, n53359 );
nand U75628 ( n53359, n53360, n1520 );
nor U75629 ( n53358, n53361, n53362 );
nor U75630 ( n53362, n53363, n53364 );
not U75631 ( n1493, n53264 );
not U75632 ( n1467, n53167 );
and U75633 ( n53028, n53157, n53158 );
nand U75634 ( n53158, n53159, n1467 );
nor U75635 ( n53157, n53160, n53161 );
nor U75636 ( n53160, n1492, n53168 );
not U75637 ( n1515, n53387 );
not U75638 ( n1557, n52392 );
not U75639 ( n2865, n17336 );
nand U75640 ( n51174, n51345, n51346 );
nand U75641 ( n51346, n1425, n50937 );
nor U75642 ( n51345, n51348, n51349 );
not U75643 ( n1425, n50940 );
not U75644 ( n1287, n51846 );
nand U75645 ( n19682, n19708, n19709 );
nand U75646 ( n19709, n19710, n2557 );
nor U75647 ( n19708, n19711, n19712 );
nor U75648 ( n19711, n2557, n19719 );
nand U75649 ( n49710, n49711, n49712 );
nand U75650 ( n49711, n1322, n1357 );
or U75651 ( n49712, n49713, n49714 );
not U75652 ( n1522, n53206 );
nor U75653 ( n17381, n2389, n17385 );
nor U75654 ( n52532, n1390, n1373 );
not U75655 ( n1437, n52777 );
not U75656 ( n1373, n52534 );
and U75657 ( n52316, n52524, n52525 );
nand U75658 ( n52525, n52526, n1373 );
nor U75659 ( n52524, n52527, n52528 );
nor U75660 ( n52527, n1408, n52535 );
nand U75661 ( n19539, n19684, n19685 );
nand U75662 ( n19685, n19686, n2525 );
nor U75663 ( n19684, n19687, n19688 );
nor U75664 ( n19687, n2525, n19695 );
nor U75665 ( n51175, n51158, n51515 );
nand U75666 ( n51516, n51164, n1393 );
nor U75667 ( n52946, n1449, n1438 );
not U75668 ( n1495, n53211 );
not U75669 ( n1409, n52782 );
not U75670 ( n1470, n52961 );
not U75671 ( n1438, n52948 );
and U75672 ( n52770, n52938, n52939 );
nand U75673 ( n52939, n52940, n1438 );
nor U75674 ( n52938, n52941, n52942 );
nor U75675 ( n52941, n1468, n52949 );
nand U75676 ( n53302, n53422, n53423 );
nand U75677 ( n53422, n53427, n53426 );
nand U75678 ( n53423, n1543, n53424 );
nand U75679 ( n53427, n53428, n53429 );
not U75680 ( n1543, n53426 );
not U75681 ( n1514, n53309 );
and U75682 ( n51170, n51857, n51858 );
nand U75683 ( n51858, n51520, n1399 );
nor U75684 ( n51857, n51862, n51863 );
not U75685 ( n1399, n51859 );
nand U75686 ( n52821, n53295, n53293 );
nor U75687 ( n53295, n53291, n53284 );
nor U75688 ( n20354, n2623, n2619 );
nand U75689 ( n52377, n1479, n51900 );
nor U75690 ( n50336, n1274, n50340 );
nor U75691 ( n51348, n1424, n51351 );
or U75692 ( n51351, n1429, n50937 );
nand U75693 ( n16995, n17309, n17310 );
nand U75694 ( n17310, n17311, n17312 );
not U75695 ( n2854, n17557 );
not U75696 ( n2638, n20451 );
nor U75697 ( n18219, n18202, n18559 );
and U75698 ( n18559, n18560, n18203 );
nand U75699 ( n18560, n18208, n2510 );
nor U75700 ( n19570, n2507, n2528 );
nor U75701 ( n52065, n1310, n1334 );
not U75702 ( n1520, n53368 );
nand U75703 ( n53644, n53704, n53705 );
nand U75704 ( n53704, n53710, n53709 );
nand U75705 ( n53705, n1599, n53706 );
nand U75706 ( n53710, n53711, n53712 );
not U75707 ( n1599, n53709 );
nand U75708 ( n18218, n18389, n18390 );
nand U75709 ( n18390, n2547, n17979 );
nor U75710 ( n18389, n18392, n18393 );
not U75711 ( n2547, n17982 );
nand U75712 ( n52332, n52520, n52329 );
nor U75713 ( n52520, n52320, n52327 );
not U75714 ( n2642, n20405 );
nor U75715 ( n18945, n2603, n2610 );
nand U75716 ( n18934, n19261, n19262 );
nand U75717 ( n19262, n18946, n2610 );
nor U75718 ( n19261, n19264, n19265 );
nor U75719 ( n19264, n2610, n19268 );
not U75720 ( n2659, n19289 );
nor U75721 ( n51807, n1267, n1290 );
not U75722 ( n2558, n19821 );
not U75723 ( n1463, n52381 );
nand U75724 ( n20535, n20537, n20538 );
nand U75725 ( n20538, n20245, n2664 );
nor U75726 ( n20537, n20540, n20541 );
and U75727 ( n20541, n2683, n20246 );
not U75728 ( n2683, n20243 );
nor U75729 ( n19549, n2468, n2487 );
nor U75730 ( n19221, n2427, n2449 );
nor U75731 ( n18867, n2382, n2404 );
nand U75732 ( n17664, n18893, n18894 );
nand U75733 ( n18894, n2367, n17926 );
nor U75734 ( n18893, n18895, n18896 );
not U75735 ( n2367, n17923 );
not U75736 ( n1600, n53718 );
nor U75737 ( n18392, n2545, n18395 );
or U75738 ( n18395, n2550, n17979 );
not U75739 ( n1329, n50899 );
nand U75740 ( n53276, n1500, n53271 );
nor U75741 ( n19984, n2568, n2590 );
nand U75742 ( n20069, n20122, n20123 );
nand U75743 ( n20123, n19988, n19992 );
nor U75744 ( n20122, n19984, n19990 );
not U75745 ( n2590, n19988 );
nand U75746 ( n20443, n20619, n20620 );
nand U75747 ( n20619, n20623, n20614 );
nand U75748 ( n20620, n2660, n20621 );
nand U75749 ( n20623, n20611, n20613 );
not U75750 ( n2660, n20614 );
not U75751 ( n2448, n18175 );
not U75752 ( n1519, n53259 );
nand U75753 ( n53372, n53451, n53452 );
nand U75754 ( n53452, n53364, n53368 );
nor U75755 ( n53451, n53360, n53366 );
nor U75756 ( n20554, n20262, n20265 );
nor U75757 ( n19227, n2427, n2405 );
nor U75758 ( n18873, n2382, n2369 );
and U75759 ( n18864, n19219, n19220 );
nand U75760 ( n19220, n19221, n2405 );
nor U75761 ( n19219, n19222, n19223 );
nor U75762 ( n19222, n2449, n19230 );
nand U75763 ( n17351, n16948, n16950 );
not U75764 ( n1497, n53106 );
and U75765 ( n53024, n53083, n53084 );
nand U75766 ( n53084, n53085, n1469 );
nor U75767 ( n53083, n53086, n53087 );
nor U75768 ( n53086, n1494, n53094 );
not U75769 ( n1498, n53228 );
not U75770 ( n1440, n52966 );
not U75771 ( n1473, n52978 );
nand U75772 ( n49594, n51821, n51822 );
nand U75773 ( n51822, n51823, n1254 );
nor U75774 ( n51821, n51824, n51825 );
nor U75775 ( n51824, n1288, n51832 );
xor U75776 ( n19869, n19289, n19288 );
not U75777 ( n1330, n52351 );
nand U75778 ( n19231, n19541, n19542 );
nand U75779 ( n19542, n19543, n2487 );
nor U75780 ( n19541, n19544, n19545 );
nor U75781 ( n19544, n2487, n19552 );
nand U75782 ( n20212, n2598, n20211 );
nor U75783 ( n49694, n50336, n50337 );
and U75784 ( n50337, n50338, n50339 );
nand U75785 ( n50338, n50340, n1274 );
nand U75786 ( n20422, n2622, n20417 );
not U75787 ( n1410, n52547 );
nor U75788 ( n18202, n2510, n18208 );
nand U75789 ( n17300, n17548, n17549 );
nand U75790 ( n17548, n17552, n17312 );
nand U75791 ( n17549, n2845, n17550 );
nand U75792 ( n17552, n17309, n17311 );
not U75793 ( n2835, n17001 );
nor U75794 ( n52940, n1449, n1468 );
nand U75795 ( n53025, n53078, n53079 );
nand U75796 ( n53079, n52944, n52948 );
nor U75797 ( n53078, n52940, n52946 );
not U75798 ( n1468, n52944 );
nor U75799 ( n16738, n17381, n17382 );
and U75800 ( n17382, n17383, n17384 );
nand U75801 ( n17383, n17385, n2389 );
not U75802 ( n2657, n20226 );
not U75803 ( n1469, n53093 );
nand U75804 ( n49998, n49999, n50000 );
nand U75805 ( n52675, n1423, n52670 );
nand U75806 ( n19958, n20320, n20321 );
nor U75807 ( n20320, n20322, n20323 );
or U75808 ( n16761, n16762, n2439 );
nand U75809 ( n51642, n52026, n52027 );
nand U75810 ( n52027, n52028, n52029 );
nand U75811 ( n20244, n20611, n20612 );
nand U75812 ( n20612, n20613, n20614 );
nand U75813 ( n50245, n50492, n50493 );
nand U75814 ( n50493, n50494, n50495 );
nand U75815 ( n50779, n50506, n50504 );
nand U75816 ( n50775, n51034, n51035 );
nand U75817 ( n51034, n51038, n50813 );
nand U75818 ( n51035, n1727, n51036 );
nand U75819 ( n51038, n50810, n50812 );
nand U75820 ( n19950, n20241, n20242 );
nand U75821 ( n20242, n20243, n20244 );
nor U75822 ( n20241, n20245, n20246 );
nand U75823 ( n52315, n52536, n52537 );
nand U75824 ( n52537, n52218, n52222 );
nor U75825 ( n52536, n52214, n52220 );
nor U75826 ( n52214, n1352, n1374 );
not U75827 ( n1374, n52218 );
not U75828 ( n1429, n51341 );
not U75829 ( n2582, n18557 );
not U75830 ( n2584, n18696 );
nand U75831 ( n53752, n53765, n53749 );
nor U75832 ( n53765, n53747, n53740 );
nand U75833 ( n19695, n2505, n19690 );
nand U75834 ( n49960, n50232, n50233 );
nand U75835 ( n50233, n50234, n50235 );
nor U75836 ( n49961, n1712, n1707 );
not U75837 ( n1472, n53111 );
not U75838 ( n2403, n18890 );
nor U75839 ( n20441, n20445, n20446 );
nor U75840 ( n20445, n20447, n2648 );
and U75841 ( n20447, n20448, n20449 );
nand U75842 ( n51914, n52384, n52385 );
nand U75843 ( n52384, n52389, n52029 );
nand U75844 ( n52385, n52386, n1537 );
nand U75845 ( n52389, n52026, n52028 );
not U75846 ( n1537, n52029 );
nand U75847 ( n20262, n20557, n20558 );
nand U75848 ( n20557, n20561, n20319 );
nand U75849 ( n20558, n2719, n20559 );
nand U75850 ( n20561, n20316, n20318 );
not U75851 ( n2733, n20568 );
xor U75852 ( n18184, n18185, n18181 );
nor U75853 ( n19109, n2428, n2452 );
nand U75854 ( n52768, n52950, n52951 );
nand U75855 ( n52951, n52692, n52696 );
nor U75856 ( n52950, n52688, n52694 );
nor U75857 ( n19576, n2507, n2489 );
nand U75858 ( n20197, n20341, n20342 );
nand U75859 ( n20342, n20133, n20137 );
nor U75860 ( n20341, n20129, n20135 );
nand U75861 ( n50606, n1277, n1272 );
nand U75862 ( n53168, n1478, n53167 );
not U75863 ( n2719, n20319 );
not U75864 ( n1442, n52709 );
not U75865 ( n2678, n19288 );
nand U75866 ( n51634, n52018, n52019 );
nand U75867 ( n52019, n52020, n52021 );
nand U75868 ( n51957, n52468, n52469 );
nand U75869 ( n52469, n52470, n52471 );
nand U75870 ( n51643, n51917, n51918 );
nand U75871 ( n51917, n51921, n51638 );
nand U75872 ( n51918, n1559, n51919 );
nand U75873 ( n51921, n51635, n51637 );
not U75874 ( n1629, n52856 );
not U75875 ( n1579, n51928 );
nand U75876 ( n19268, n2603, n18944 );
nand U75877 ( n53153, n53195, n53196 );
nand U75878 ( n53196, n53089, n53093 );
nor U75879 ( n53195, n53085, n53091 );
not U75880 ( n2718, n20567 );
nand U75881 ( n52429, n52864, n52865 );
nand U75882 ( n52864, n52869, n52467 );
nand U75883 ( n52865, n1659, n52866 );
nand U75884 ( n52869, n52464, n52466 );
not U75885 ( n1510, n51648 );
not U75886 ( n1279, n49703 );
nand U75887 ( n52855, n53810, n53811 );
nand U75888 ( n53810, n53815, n52863 );
nand U75889 ( n53811, n1647, n53812 );
nand U75890 ( n53815, n52860, n52862 );
and U75891 ( n20196, n20346, n20347 );
nand U75892 ( n20347, n20348, n2619 );
nor U75893 ( n20346, n20349, n20350 );
nor U75894 ( n20349, n2644, n20357 );
nand U75895 ( n52535, n1390, n52534 );
nand U75896 ( n52949, n1449, n52948 );
not U75897 ( n8220, n18105 );
nor U75898 ( n53300, n53304, n53305 );
nor U75899 ( n53304, n53306, n1527 );
not U75900 ( n1737, n50505 );
nor U75901 ( n52220, n1352, n1335 );
nand U75902 ( n52625, n52698, n52699 );
nand U75903 ( n52699, n52564, n52568 );
nor U75904 ( n52698, n52560, n52566 );
nor U75905 ( n52560, n1392, n1413 );
not U75906 ( n1375, n52552 );
not U75907 ( n1413, n52564 );
not U75908 ( n1335, n52222 );
nand U75909 ( n50489, n50765, n50766 );
nand U75910 ( n50765, n50770, n50495 );
nand U75911 ( n50766, n1715, n50767 );
nand U75912 ( n50770, n50492, n50494 );
not U75913 ( n1443, n52983 );
nor U75914 ( n20146, n2599, n2620 );
nand U75915 ( n52902, n53711, n53715 );
nand U75916 ( n53715, n53712, n53709 );
and U75917 ( n16609, n18865, n18866 );
nand U75918 ( n18866, n18867, n2369 );
nor U75919 ( n18865, n18868, n18869 );
nor U75920 ( n18868, n2404, n18876 );
nor U75921 ( n52071, n1310, n1292 );
and U75922 ( n52170, n52212, n52213 );
nand U75923 ( n52213, n52214, n1335 );
nor U75924 ( n52212, n52215, n52216 );
nor U75925 ( n52215, n1374, n52223 );
not U75926 ( n1715, n50495 );
nor U75927 ( n51813, n1267, n1255 );
nor U75928 ( n51699, n1268, n1293 );
nor U75929 ( n52566, n1392, n1378 );
nor U75930 ( n52163, n1312, n1294 );
nor U75931 ( n51705, n1268, n1257 );
not U75932 ( n1415, n52581 );
not U75933 ( n1339, n52091 );
not U75934 ( n1378, n52568 );
not U75935 ( n1294, n52165 );
and U75936 ( n51798, n52155, n52156 );
nand U75937 ( n52156, n52157, n1294 );
nor U75938 ( n52155, n52158, n52159 );
nor U75939 ( n52158, n1337, n52166 );
and U75940 ( n52308, n52558, n52559 );
nand U75941 ( n52559, n52560, n1378 );
nor U75942 ( n52558, n52561, n52562 );
nor U75943 ( n52561, n1413, n52569 );
nor U75944 ( n18851, n2383, n2407 );
not U75945 ( n2480, n17962 );
nand U75946 ( n16754, n16755, n16756 );
nand U75947 ( n16755, n2439, n2474 );
or U75948 ( n16756, n16757, n16758 );
nor U75949 ( n19990, n2568, n2559 );
not U75950 ( n2593, n20005 );
not U75951 ( n2559, n19992 );
not U75952 ( n1414, n52714 );
not U75953 ( n1444, n52726 );
nand U75954 ( n51973, n52432, n52433 );
nand U75955 ( n52433, n1677, n52434 );
nand U75956 ( n52432, n52437, n52013 );
not U75957 ( n1677, n52013 );
nand U75958 ( n52413, n52419, n52420 );
nand U75959 ( n52420, n1649, n52421 );
nand U75960 ( n52419, n52424, n52017 );
not U75961 ( n1649, n52017 );
nand U75962 ( n52437, n52010, n52012 );
nand U75963 ( n52424, n52014, n52016 );
nor U75964 ( n52157, n1312, n1337 );
not U75965 ( n1337, n52161 );
and U75966 ( n52168, n52224, n52225 );
nand U75967 ( n52225, n52161, n52165 );
nor U75968 ( n52224, n52157, n52163 );
not U75969 ( n2394, n16747 );
not U75970 ( n1494, n53089 );
not U75971 ( n2529, n19826 );
and U75972 ( n19814, n19982, n19983 );
nand U75973 ( n19983, n19984, n2559 );
nor U75974 ( n19982, n19985, n19986 );
nor U75975 ( n19985, n2590, n19993 );
not U75976 ( n2445, n19402 );
and U75977 ( n52627, n52686, n52687 );
nand U75978 ( n52687, n52688, n1412 );
nor U75979 ( n52686, n52689, n52690 );
nor U75980 ( n52689, n1439, n52697 );
nand U75981 ( n51972, n52464, n52465 );
nand U75982 ( n52465, n52466, n52467 );
nor U75983 ( n20018, n2569, n2595 );
not U75984 ( n2562, n20010 );
nand U75985 ( n49752, n49750, n49753 );
nand U75986 ( n49753, n49748, n49754 );
nand U75987 ( n50490, n50814, n50815 );
nand U75988 ( n50815, n50816, n50817 );
not U75989 ( n1412, n52696 );
nand U75990 ( n19540, n19564, n19536 );
nor U75991 ( n19564, n19527, n19534 );
nand U75992 ( n50776, n51030, n51031 );
nand U75993 ( n51031, n51032, n51033 );
nand U75994 ( n51633, n51948, n51949 );
nand U75995 ( n51948, n51953, n51628 );
nand U75996 ( n51949, n1623, n51950 );
nand U75997 ( n51953, n51625, n51627 );
nand U75998 ( n51962, n52014, n52015 );
nand U75999 ( n52015, n52016, n52017 );
nand U76000 ( n51960, n51572, n51571 );
nand U76001 ( n51941, n52399, n52400 );
nand U76002 ( n52399, n52404, n52021 );
nand U76003 ( n52400, n1610, n52401 );
nand U76004 ( n52404, n52018, n52020 );
not U76005 ( n1598, n51561 );
and U76006 ( n51804, n52063, n52064 );
nand U76007 ( n52064, n52065, n1292 );
nor U76008 ( n52063, n52066, n52067 );
nor U76009 ( n52066, n1334, n52074 );
nor U76010 ( n16778, n2575, n2608 );
not U76011 ( n2575, n17056 );
nor U76012 ( n52254, n1353, n1340 );
not U76013 ( n1417, n52731 );
not U76014 ( n1297, n52096 );
not U76015 ( n1382, n52269 );
not U76016 ( n1340, n52256 );
and U76017 ( n52149, n52246, n52247 );
nand U76018 ( n52247, n52248, n1340 );
nor U76019 ( n52246, n52249, n52250 );
nor U76020 ( n52249, n1379, n52257 );
not U76021 ( n1499, n53126 );
not U76022 ( n1647, n52863 );
nand U76023 ( n50224, n50479, n50480 );
nand U76024 ( n50480, n1705, n50481 );
nand U76025 ( n50479, n50484, n50235 );
not U76026 ( n1705, n50235 );
nand U76027 ( n50484, n50232, n50234 );
and U76028 ( n20068, n20127, n20128 );
nand U76029 ( n20128, n20129, n2592 );
nor U76030 ( n20127, n20130, n20131 );
nor U76031 ( n20130, n2618, n20138 );
not U76032 ( n1659, n52467 );
nand U76033 ( n19891, n20316, n20317 );
nand U76034 ( n20317, n20318, n20319 );
not U76035 ( n2592, n20137 );
not U76036 ( n1380, n52586 );
not U76037 ( n1460, n51332 );
xor U76038 ( n53809, n52856, n52855 );
nor U76039 ( n19421, n2469, n2490 );
not U76040 ( n2845, n17312 );
nand U76041 ( n17299, n17544, n17545 );
nand U76042 ( n17545, n17546, n17547 );
nand U76043 ( n17824, n17556, n17554 );
xor U76044 ( n49559, n49560, n49561 );
not U76045 ( n1623, n51628 );
and U76046 ( n52154, n52229, n52230 );
nand U76047 ( n52230, n52231, n1338 );
nor U76048 ( n52229, n52232, n52233 );
nor U76049 ( n52232, n1377, n52240 );
nand U76050 ( n52428, n52860, n52861 );
nand U76051 ( n52861, n52862, n52863 );
nor U76052 ( n20152, n2599, n2594 );
nand U76053 ( n17005, n17286, n17287 );
nand U76054 ( n17287, n17288, n17289 );
not U76055 ( n2833, n17542 );
and U76056 ( n20064, n20144, n20145 );
nand U76057 ( n20145, n20146, n2594 );
nor U76058 ( n20144, n20147, n20148 );
nor U76059 ( n20147, n2620, n20155 );
nor U76060 ( n17006, n2829, n2824 );
nand U76061 ( n52311, n52553, n52554 );
nand U76062 ( n52554, n52235, n52239 );
nor U76063 ( n52553, n52231, n52237 );
not U76064 ( n2530, n19591 );
nand U76065 ( n50548, n50752, n50753 );
nand U76066 ( n50753, n1698, n50754 );
nand U76067 ( n50752, n50757, n50478 );
not U76068 ( n1698, n50478 );
nand U76069 ( n50757, n50475, n50477 );
nand U76070 ( n20573, n20677, n20678 );
nor U76071 ( n20677, n20679, n20680 );
nand U76072 ( n18678, n19062, n19063 );
nand U76073 ( n19063, n19064, n19065 );
not U76074 ( n2750, n19001 );
not U76075 ( n2767, n19909 );
nand U76076 ( n51573, n51964, n51965 );
nand U76077 ( n51964, n51968, n51578 );
nand U76078 ( n51965, n1662, n51966 );
nand U76079 ( n51968, n51575, n51577 );
nand U76080 ( n51588, n52010, n52011 );
nand U76081 ( n52011, n52012, n52013 );
not U76082 ( n1678, n51975 );
not U76083 ( n1559, n51638 );
nand U76084 ( n51027, n51269, n51270 );
nand U76085 ( n51270, n1714, n51271 );
nand U76086 ( n51269, n51274, n51033 );
not U76087 ( n1714, n51033 );
nand U76088 ( n51274, n51030, n51032 );
nor U76089 ( n52137, n1313, n1342 );
nand U76090 ( n52147, n52258, n52259 );
nand U76091 ( n52259, n52141, n52145 );
nor U76092 ( n52258, n52137, n52143 );
not U76093 ( n1342, n52141 );
nand U76094 ( n50225, n50475, n50476 );
nand U76095 ( n50476, n50477, n50478 );
nor U76096 ( n52248, n1353, n1379 );
nand U76097 ( n52306, n52570, n52571 );
nand U76098 ( n52571, n52252, n52256 );
nor U76099 ( n52570, n52248, n52254 );
not U76100 ( n1379, n52252 );
not U76101 ( n1322, n50056 );
nor U76102 ( n49714, n1357, n1322 );
nor U76103 ( n19115, n2428, n2408 );
nand U76104 ( n19669, n19742, n19743 );
nand U76105 ( n19743, n19608, n19612 );
nor U76106 ( n19742, n19604, n19610 );
nor U76107 ( n19604, n2508, n2533 );
nor U76108 ( n19201, n2429, n2454 );
not U76109 ( n2492, n19596 );
not U76110 ( n2533, n19608 );
nor U76111 ( n52143, n1313, n1299 );
not U76112 ( n1384, n52615 );
not U76113 ( n1343, n52274 );
not U76114 ( n1299, n52145 );
not U76115 ( n2752, n19910 );
not U76116 ( n2439, n17102 );
nor U76117 ( n16758, n2474, n2439 );
nor U76118 ( n19427, n2469, n2453 );
and U76119 ( n19214, n19419, n19420 );
nand U76120 ( n19420, n19421, n2453 );
nor U76121 ( n19419, n19422, n19423 );
nor U76122 ( n19422, n2490, n19430 );
not U76123 ( n2658, n19073 );
not U76124 ( n2550, n18385 );
not U76125 ( n1439, n52692 );
not U76126 ( n1338, n52239 );
nor U76127 ( n20024, n2569, n2564 );
nand U76128 ( n17044, n17045, n17046 );
not U76129 ( n2633, n18692 );
nand U76130 ( n50762, n51017, n51018 );
nand U76131 ( n51017, n51022, n50817 );
nand U76132 ( n51018, n1704, n51019 );
nand U76133 ( n51022, n50814, n50816 );
nor U76134 ( n16777, n17057, n17056 );
not U76135 ( n2618, n20133 );
nand U76136 ( n19812, n19994, n19995 );
nand U76137 ( n19995, n19736, n19740 );
nor U76138 ( n19994, n19732, n19738 );
nand U76139 ( n17540, n17810, n17811 );
nand U76140 ( n17810, n17815, n17547 );
nand U76141 ( n17811, n2832, n17812 );
nand U76142 ( n17815, n17544, n17546 );
nor U76143 ( n18857, n2383, n2370 );
nor U76144 ( n18743, n2384, n2409 );
nand U76145 ( n52223, n1352, n52222 );
nand U76146 ( n52852, n52468, n52470 );
nand U76147 ( n52569, n1392, n52568 );
and U76148 ( n19671, n19730, n19731 );
nand U76149 ( n19731, n19732, n2532 );
nor U76150 ( n19730, n19733, n19734 );
nor U76151 ( n19733, n2560, n19741 );
nand U76152 ( n51071, n51252, n51253 );
nand U76153 ( n51253, n1697, n51254 );
nand U76154 ( n51252, n51257, n51066 );
not U76155 ( n1697, n51066 );
nand U76156 ( n51257, n51063, n51065 );
xnor U76157 ( n16584, n16585, n16587 );
nand U76158 ( n17278, n17531, n17532 );
nand U76159 ( n17531, n17535, n17289 );
nand U76160 ( n17532, n2823, n17533 );
nand U76161 ( n17535, n17286, n17288 );
not U76162 ( n1627, n52471 );
and U76163 ( n18848, n19107, n19108 );
nand U76164 ( n19108, n19109, n2408 );
nor U76165 ( n19107, n19110, n19111 );
nor U76166 ( n19110, n2452, n19118 );
not U76167 ( n2532, n19740 );
not U76168 ( n1727, n50813 );
nand U76169 ( n52166, n1312, n52165 );
nand U76170 ( n51026, n51265, n51266 );
nand U76171 ( n51266, n51267, n51268 );
not U76172 ( n2563, n19753 );
nand U76173 ( n19324, n19330, n19331 );
nand U76174 ( n19331, n2769, n19332 );
nand U76175 ( n19330, n19335, n19061 );
not U76176 ( n2769, n19061 );
nand U76177 ( n19335, n19058, n19060 );
nand U76178 ( n51799, n52080, n52081 );
nand U76179 ( n52081, n51721, n51725 );
nor U76180 ( n52080, n51717, n51723 );
not U76181 ( n1298, n51787 );
nand U76182 ( n19993, n2568, n19992 );
not U76183 ( n1662, n51578 );
not U76184 ( n1377, n52235 );
nor U76185 ( n19610, n2508, n2494 );
not U76186 ( n2534, n19758 );
not U76187 ( n2494, n19612 );
and U76188 ( n19806, n20016, n20017 );
nand U76189 ( n20017, n20018, n2564 );
nor U76190 ( n20016, n20019, n20020 );
nor U76191 ( n20019, n2595, n20027 );
nand U76192 ( n18677, n18992, n18993 );
nand U76193 ( n18992, n18997, n18611 );
nand U76194 ( n18993, n2745, n18994 );
nand U76195 ( n18997, n18608, n18610 );
nand U76196 ( n19006, n19058, n19059 );
nand U76197 ( n19059, n19060, n19061 );
nand U76198 ( n19004, n18620, n18619 );
nand U76199 ( n50932, n50940, n51339 );
nand U76200 ( n51339, n51340, n50937 );
nand U76201 ( n51340, n51341, n1424 );
not U76202 ( n2734, n19893 );
and U76203 ( n20272, n2767, n19912 );
nor U76204 ( n19766, n2544, n2565 );
nand U76205 ( n52257, n1353, n52256 );
nand U76206 ( n18985, n19310, n19311 );
nand U76207 ( n19310, n19315, n19065 );
nand U76208 ( n19311, n2735, n19312 );
nand U76209 ( n19315, n19062, n19064 );
not U76210 ( n2714, n18605 );
not U76211 ( n1259, n51792 );
and U76212 ( n51778, n52135, n52136 );
nand U76213 ( n52136, n52137, n1299 );
nor U76214 ( n52135, n52138, n52139 );
nor U76215 ( n52138, n1342, n52146 );
nand U76216 ( n51589, n51977, n51978 );
nand U76217 ( n51977, n51981, n51624 );
nand U76218 ( n51978, n1687, n51979 );
nand U76219 ( n51981, n51621, n51623 );
not U76220 ( n1687, n51624 );
nand U76221 ( n51395, n51635, n51636 );
nand U76222 ( n51636, n51637, n51638 );
not U76223 ( n2535, n19625 );
not U76224 ( n1418, n52610 );
not U76225 ( n1344, n52116 );
xor U76226 ( n20274, n19910, n19909 );
nor U76227 ( n19207, n2429, n2410 );
nor U76228 ( n18749, n2384, n2372 );
not U76229 ( n2457, n19135 );
and U76230 ( n18842, n19199, n19200 );
nand U76231 ( n19200, n19201, n2410 );
nor U76232 ( n19199, n19202, n19203 );
nor U76233 ( n19202, n2454, n19210 );
and U76234 ( n19516, n19602, n19603 );
nand U76235 ( n19603, n19604, n2494 );
nor U76236 ( n19602, n19605, n19606 );
nor U76237 ( n19605, n2533, n19613 );
not U76238 ( n2773, n19946 );
and U76239 ( n49520, n51805, n51806 );
nand U76240 ( n51806, n51807, n1255 );
nor U76241 ( n51805, n51808, n51809 );
nor U76242 ( n51808, n1290, n51816 );
not U76243 ( n2832, n17547 );
not U76244 ( n1458, n50952 );
nand U76245 ( n17541, n17806, n17807 );
nand U76246 ( n17807, n17808, n17809 );
nor U76247 ( n19772, n2544, n2537 );
nand U76248 ( n17974, n17982, n18383 );
nand U76249 ( n18383, n18384, n17979 );
nand U76250 ( n18384, n18385, n2545 );
not U76251 ( n2745, n18611 );
not U76252 ( n2680, n18682 );
nand U76253 ( n17523, n17793, n17794 );
nand U76254 ( n17793, n17797, n17530 );
nand U76255 ( n17794, n2814, n17795 );
nand U76256 ( n17797, n17527, n17529 );
not U76257 ( n2822, n17804 );
nor U76258 ( n19461, n2470, n2458 );
not U76259 ( n2413, n19140 );
not U76260 ( n2498, n19476 );
not U76261 ( n2458, n19463 );
and U76262 ( n19663, n19764, n19765 );
nand U76263 ( n19765, n19766, n2537 );
nor U76264 ( n19764, n19767, n19768 );
nor U76265 ( n19767, n2565, n19775 );
and U76266 ( n19194, n19453, n19454 );
nand U76267 ( n19454, n19455, n2458 );
nor U76268 ( n19453, n19456, n19457 );
nor U76269 ( n19456, n2495, n19464 );
not U76270 ( n2497, n19630 );
not U76271 ( n2483, n17620 );
nand U76272 ( n50761, n51063, n51064 );
nand U76273 ( n51064, n51065, n51066 );
nor U76274 ( n19656, n2509, n2499 );
nor U76275 ( n19187, n2430, n2415 );
nand U76276 ( n19192, n19465, n19466 );
nand U76277 ( n19466, n19185, n19189 );
nor U76278 ( n19465, n19181, n19187 );
not U76279 ( n2462, n19481 );
not U76280 ( n2415, n19189 );
and U76281 ( n19485, n19648, n19649 );
nand U76282 ( n19649, n19650, n2499 );
nor U76283 ( n19648, n19651, n19652 );
nor U76284 ( n19651, n2538, n19659 );
nand U76285 ( n16797, n16795, n16798 );
nand U76286 ( n16798, n16793, n16799 );
not U76287 ( n1704, n50817 );
not U76288 ( n1367, n50577 );
nand U76289 ( n51070, n51248, n51249 );
nand U76290 ( n51249, n51250, n51251 );
nand U76291 ( n51261, n51453, n51454 );
nand U76292 ( n51453, n51458, n51268 );
nand U76293 ( n51454, n1703, n51455 );
nand U76294 ( n51458, n51265, n51267 );
and U76295 ( n19518, n19597, n19598 );
nand U76296 ( n19598, n19442, n19446 );
nor U76297 ( n19597, n19438, n19444 );
nor U76298 ( n19181, n2430, n2459 );
not U76299 ( n2459, n19185 );
not U76300 ( n1347, n52295 );
not U76301 ( n1610, n52021 );
not U76302 ( n1560, n51324 );
not U76303 ( n2800, n19024 );
not U76304 ( n2583, n18376 );
and U76305 ( n19198, n19436, n19437 );
nand U76306 ( n19437, n19438, n2455 );
nor U76307 ( n19436, n19439, n19440 );
nor U76308 ( n19439, n2493, n19447 );
not U76309 ( n2560, n19736 );
nand U76310 ( n18621, n19008, n19009 );
nand U76311 ( n19009, n2783, n19010 );
nand U76312 ( n19008, n19013, n18672 );
not U76313 ( n2783, n18672 );
nand U76314 ( n19013, n18669, n18671 );
not U76315 ( n2823, n17289 );
nor U76316 ( n51741, n1269, n1300 );
nand U76317 ( n51779, n52102, n52103 );
nand U76318 ( n52103, n51745, n51749 );
nor U76319 ( n52102, n51741, n51747 );
not U76320 ( n1300, n51745 );
nand U76321 ( n19514, n19614, n19615 );
nand U76322 ( n19615, n19459, n19463 );
nor U76323 ( n19614, n19455, n19461 );
nor U76324 ( n19455, n2470, n2495 );
not U76325 ( n2495, n19459 );
not U76326 ( n1385, n52290 );
not U76327 ( n2455, n19446 );
not U76328 ( n1360, n50376 );
nand U76329 ( n17279, n17527, n17528 );
nand U76330 ( n17528, n17529, n17530 );
nand U76331 ( n51262, n51449, n51450 );
nand U76332 ( n51450, n51451, n51452 );
nand U76333 ( n51597, n51449, n51451 );
nand U76334 ( n51446, n51592, n51593 );
nand U76335 ( n51593, n1695, n51594 );
nand U76336 ( n51592, n51597, n51452 );
not U76337 ( n1695, n51452 );
nand U76338 ( n18118, n18296, n18297 );
nand U76339 ( n18297, n2813, n18298 );
nand U76340 ( n18296, n18301, n18113 );
not U76341 ( n2813, n18113 );
nand U76342 ( n18301, n18110, n18112 );
nand U76343 ( n17802, n18063, n18064 );
nand U76344 ( n18064, n2820, n18065 );
nand U76345 ( n18063, n18068, n17809 );
not U76346 ( n2820, n17809 );
nand U76347 ( n18068, n17806, n17808 );
not U76348 ( n2493, n19442 );
not U76349 ( n2848, n17858 );
not U76350 ( n2814, n17530 );
not U76351 ( n2517, n17896 );
not U76352 ( n2374, n18836 );
nand U76353 ( n18821, n19179, n19180 );
nand U76354 ( n19180, n19181, n2415 );
nor U76355 ( n19179, n19182, n19183 );
nor U76356 ( n19182, n2459, n19190 );
and U76357 ( n16535, n18849, n18850 );
nand U76358 ( n18850, n18851, n2370 );
nor U76359 ( n18849, n18852, n18853 );
nor U76360 ( n18852, n2407, n18860 );
nand U76361 ( n52146, n1313, n52145 );
not U76362 ( n1694, n51988 );
nor U76363 ( n19650, n2509, n2538 );
not U76364 ( n2463, n19160 );
nor U76365 ( n51747, n1269, n1260 );
not U76366 ( n1260, n51749 );
nand U76367 ( n50180, n50186, n50187 );
nand U76368 ( n50187, n50188, n50189 );
nor U76369 ( n49823, n1670, n1658 );
not U76370 ( n2677, n18372 );
not U76371 ( n1305, n52299 );
not U76372 ( n1703, n51268 );
nand U76373 ( n19613, n2508, n19612 );
nor U76374 ( n19499, n2472, n2464 );
nand U76375 ( n19464, n2470, n19463 );
nor U76376 ( n18785, n2385, n2417 );
not U76377 ( n2417, n18789 );
and U76378 ( n18824, n19146, n19147 );
nand U76379 ( n19147, n18789, n18793 );
nor U76380 ( n19146, n18785, n18791 );
not U76381 ( n2414, n18831 );
nand U76382 ( n50749, n51073, n51074 );
nand U76383 ( n51074, n51075, n51076 );
not U76384 ( n2808, n18668 );
nand U76385 ( n18117, n18345, n18346 );
nand U76386 ( n18346, n18347, n18348 );
and U76387 ( n49458, n51697, n51698 );
nand U76388 ( n51698, n51699, n1257 );
nor U76389 ( n51697, n51700, n51701 );
nor U76390 ( n51700, n1293, n51708 );
nand U76391 ( n17801, n18110, n18111 );
nand U76392 ( n18111, n18112, n18113 );
not U76393 ( n2735, n19065 );
not U76394 ( n2580, n17994 );
not U76395 ( n1485, n51096 );
nand U76396 ( n51246, n51436, n51437 );
nand U76397 ( n51437, n1688, n51438 );
nand U76398 ( n51436, n51441, n51251 );
not U76399 ( n1688, n51251 );
nand U76400 ( n51231, n51423, n51424 );
nand U76401 ( n51423, n51427, n51304 );
nand U76402 ( n51424, n1663, n51425 );
nand U76403 ( n51427, n51301, n51303 );
not U76404 ( n1680, n51434 );
nand U76405 ( n51441, n51248, n51250 );
nor U76406 ( n19493, n2472, n2500 );
not U76407 ( n1303, n51769 );
nand U76408 ( n50176, n50456, n50457 );
nand U76409 ( n50456, n50460, n50189 );
nand U76410 ( n50457, n1657, n50458 );
nand U76411 ( n50460, n50186, n50188 );
not U76412 ( n1643, n49813 );
not U76413 ( n1430, n50394 );
not U76414 ( n1345, n52298 );
or U76415 ( n49779, n49780, n49781 );
not U76416 ( n1683, n50472 );
and U76417 ( n19173, n19491, n19492 );
nand U76418 ( n19492, n19493, n2464 );
nor U76419 ( n19491, n19494, n19495 );
nor U76420 ( n19494, n2500, n19502 );
nand U76421 ( n51232, n51419, n51420 );
nand U76422 ( n51420, n51421, n51422 );
nand U76423 ( n51432, n51579, n51580 );
nand U76424 ( n51580, n1679, n51581 );
nand U76425 ( n51579, n51584, n51486 );
not U76426 ( n1679, n51486 );
nand U76427 ( n51584, n51483, n51485 );
nand U76428 ( n51245, n51483, n51484 );
nand U76429 ( n51484, n51485, n51486 );
not U76430 ( n2779, n17234 );
nor U76431 ( n16868, n2790, n2779 );
not U76432 ( n2479, n17083 );
nand U76433 ( n19190, n2430, n19189 );
nor U76434 ( n18791, n2385, n2375 );
not U76435 ( n2375, n18793 );
not U76436 ( n1619, n50156 );
nor U76437 ( n49798, n1637, n1619 );
not U76438 ( n1657, n50189 );
nor U76439 ( n19508, n2423, n2420 );
nand U76440 ( n51012, n51235, n51236 );
nand U76441 ( n51236, n1682, n51237 );
nand U76442 ( n51235, n51240, n51076 );
not U76443 ( n1682, n51076 );
nand U76444 ( n51240, n51073, n51075 );
nand U76445 ( n50175, n50550, n50551 );
nand U76446 ( n50551, n50552, n50553 );
xor U76447 ( n18229, n17994, n17993 );
not U76448 ( n2825, n18312 );
nand U76449 ( n51416, n51564, n51565 );
nand U76450 ( n51564, n51569, n51422 );
nand U76451 ( n51565, n1650, n51566 );
nand U76452 ( n51569, n51419, n51421 );
not U76453 ( n1508, n50696 );
not U76454 ( n1663, n51304 );
nand U76455 ( n18293, n18480, n18481 );
nand U76456 ( n18480, n18485, n18348 );
nand U76457 ( n18481, n2805, n18482 );
nand U76458 ( n18485, n18345, n18347 );
nand U76459 ( n18279, n18467, n18468 );
nand U76460 ( n18467, n18471, n18352 );
nand U76461 ( n18468, n2784, n18469 );
nand U76462 ( n18471, n18349, n18351 );
not U76463 ( n2797, n18478 );
nand U76464 ( n17790, n18057, n18058 );
nand U76465 ( n18058, n18059, n18060 );
not U76466 ( n2807, n18294 );
nand U76467 ( n50453, n50726, n50727 );
nand U76468 ( n50726, n50731, n50553 );
nand U76469 ( n50727, n1642, n50728 );
nand U76470 ( n50731, n50550, n50552 );
not U76471 ( n2764, n16858 );
nand U76472 ( n51415, n51625, n51626 );
nand U76473 ( n51626, n51627, n51628 );
nand U76474 ( n18280, n18463, n18464 );
nand U76475 ( n18464, n18465, n18466 );
nand U76476 ( n18476, n18623, n18624 );
nand U76477 ( n18624, n2795, n18625 );
nand U76478 ( n18623, n18628, n18530 );
not U76479 ( n2795, n18530 );
nand U76480 ( n18628, n18527, n18529 );
nor U76481 ( n19507, n2423, n2460 );
not U76482 ( n2419, n18813 );
not U76483 ( n2552, n17439 );
and U76484 ( n16459, n18741, n18742 );
nand U76485 ( n18742, n18743, n2372 );
nor U76486 ( n18741, n18744, n18745 );
nor U76487 ( n18744, n2409, n18752 );
nand U76488 ( n51011, n51301, n51302 );
nand U76489 ( n51302, n51303, n51304 );
not U76490 ( n1609, n49981 );
nand U76491 ( n51431, n51575, n51576 );
nand U76492 ( n51576, n51577, n51578 );
nand U76493 ( n18292, n18527, n18528 );
nand U76494 ( n18528, n18529, n18530 );
nand U76495 ( n18054, n18283, n18284 );
nand U76496 ( n18283, n18287, n18060 );
nand U76497 ( n18284, n2798, n18285 );
nand U76498 ( n18287, n18057, n18059 );
nand U76499 ( n45502, n51727, n51728 );
nand U76500 ( n51727, n45481, n45483 );
nand U76501 ( n51728, n45484, n51729 );
or U76502 ( n51729, n45483, n45481 );
nand U76503 ( n45483, n51730, n51731 );
nand U76504 ( n51730, n45474, n45472 );
nand U76505 ( n51731, n45473, n51732 );
or U76506 ( n51732, n45472, n45474 );
not U76507 ( n2799, n17517 );
nand U76508 ( n51445, n51621, n51622 );
nand U76509 ( n51622, n51623, n51624 );
not U76510 ( n2805, n18348 );
nand U76511 ( n51422, n51570, n51571 );
nand U76512 ( n51570, n51572, n51573 );
not U76513 ( n2515, n17128 );
not U76514 ( n1455, n50324 );
nand U76515 ( n18460, n18612, n18613 );
nand U76516 ( n18612, n18617, n18466 );
nand U76517 ( n18613, n2770, n18614 );
nand U76518 ( n18617, n18463, n18465 );
or U76519 ( n16824, n16825, n16826 );
not U76520 ( n1642, n50553 );
and U76521 ( n45504, n51715, n51716 );
nand U76522 ( n51716, n51717, n1258 );
nor U76523 ( n51715, n51718, n51719 );
nor U76524 ( n51718, n1295, n51726 );
not U76525 ( n2784, n18352 );
not U76526 ( n2742, n17210 );
nor U76527 ( n16843, n2760, n2742 );
nand U76528 ( n50452, n50828, n50829 );
nand U76529 ( n50829, n50830, n50831 );
not U76530 ( n1640, n51000 );
not U76531 ( n1258, n51725 );
not U76532 ( n1263, n53943 );
nand U76533 ( n50086, n50409, n50410 );
nand U76534 ( n50409, n50413, n50093 );
nand U76535 ( n50410, n1505, n50411 );
nand U76536 ( n50413, n50090, n50092 );
not U76537 ( n1530, n50420 );
not U76538 ( n1594, n50132 );
nor U76539 ( n49781, n1604, n1594 );
nand U76540 ( n50406, n50680, n50681 );
nand U76541 ( n50680, n50684, n50573 );
nand U76542 ( n50681, n1484, n50682 );
nand U76543 ( n50684, n50570, n50572 );
not U76544 ( n1504, n50691 );
nand U76545 ( n19170, n21026, n21027 );
nand U76546 ( n21027, n19507, n2420 );
nor U76547 ( n21026, n21028, n21029 );
nor U76548 ( n21028, n2460, n21033 );
not U76549 ( n1304, n53938 );
not U76550 ( n2630, n17888 );
nand U76551 ( n18459, n18608, n18609 );
nand U76552 ( n18609, n18610, n18611 );
or U76553 ( n49796, n49797, n49798 );
not U76554 ( n2798, n18060 );
nand U76555 ( n18475, n18669, n18670 );
nand U76556 ( n18670, n18671, n18672 );
nand U76557 ( n18053, n18349, n18350 );
nand U76558 ( n18350, n18351, n18352 );
not U76559 ( n2730, n17027 );
nand U76560 ( n18466, n18618, n18619 );
nand U76561 ( n18618, n18620, n18621 );
not U76562 ( n2765, n17596 );
not U76563 ( n1484, n50573 );
not U76564 ( n1578, n49986 );
nand U76565 ( n50085, n50570, n50571 );
nand U76566 ( n50571, n50572, n50573 );
not U76567 ( n1652, n51080 );
nand U76568 ( n50722, n50989, n50990 );
nand U76569 ( n50989, n50993, n50831 );
nand U76570 ( n50990, n1620, n50991 );
nand U76571 ( n50993, n50828, n50830 );
not U76572 ( n1295, n51721 );
not U76573 ( n1613, n50557 );
not U76574 ( n2578, n17135 );
nand U76575 ( n17141, n17454, n17455 );
nand U76576 ( n17454, n17458, n17147 );
nand U76577 ( n17455, n2628, n17456 );
nand U76578 ( n17458, n17144, n17146 );
not U76579 ( n2652, n17465 );
and U76580 ( n11727, n18759, n18760 );
nand U76581 ( n18760, n18761, n2373 );
nor U76582 ( n18759, n18762, n18763 );
nor U76583 ( n18762, n2412, n18770 );
not U76584 ( n1505, n50093 );
not U76585 ( n2712, n17186 );
nor U76586 ( n16826, n2725, n2712 );
nand U76587 ( n17451, n17725, n17726 );
nand U76588 ( n17726, n2607, n17727 );
nand U76589 ( n17725, n17730, n17616 );
not U76590 ( n2607, n17616 );
nand U76591 ( n17730, n17613, n17615 );
nor U76592 ( n20984, n2380, n2378 );
not U76593 ( n1620, n50831 );
nor U76594 ( n20978, n2380, n2422 );
not U76595 ( n2699, n17032 );
nand U76596 ( n49754, n50090, n50091 );
nand U76597 ( n50091, n50092, n50093 );
or U76598 ( n16841, n16842, n16843 );
nor U76599 ( n49995, n1573, n1555 );
nand U76600 ( n17140, n17613, n17614 );
nand U76601 ( n17614, n17615, n17616 );
not U76602 ( n2628, n17147 );
not U76603 ( n2772, n18123 );
and U76604 ( n45453, n51739, n51740 );
nand U76605 ( n51740, n51741, n1260 );
nor U76606 ( n51739, n51742, n51743 );
nor U76607 ( n51742, n1300, n51750 );
not U76608 ( n2732, n17600 );
not U76609 ( n2744, n17872 );
nand U76610 ( n49832, n49835, n49836 );
nand U76611 ( n49835, n49845, n49846 );
nand U76612 ( n49836, n49837, n49838 );
nor U76613 ( n49845, n49843, n49971 );
or U76614 ( n49821, n49822, n49823 );
nand U76615 ( n45452, n51751, n51752 );
or U76616 ( n51751, n45441, n45444 );
nand U76617 ( n51752, n45443, n51753 );
nand U76618 ( n51753, n45444, n45441 );
nand U76619 ( n16799, n17144, n17145 );
nand U76620 ( n17145, n17146, n17147 );
nor U76621 ( n17041, n2694, n2675 );
nand U76622 ( n51750, n1269, n51749 );
and U76623 ( n11677, n18783, n18784 );
nor U76624 ( n18783, n18786, n18787 );
nand U76625 ( n18784, n18785, n2375 );
nor U76626 ( n18787, n18788, n18789 );
and U76627 ( n45444, n51754, n51755 );
nand U76628 ( n51754, n45431, n45433 );
nand U76629 ( n51755, n45434, n51756 );
or U76630 ( n51756, n45433, n45431 );
nor U76631 ( n18786, n2417, n18794 );
nand U76632 ( n18794, n2385, n18793 );
nor U76633 ( n49971, n1693, n49842 );
nor U76634 ( n49854, n49855, n1719 );
not U76635 ( n1719, n49856 );
nor U76636 ( n49855, n49857, n49858 );
nor U76637 ( n49857, n1707, n49859 );
nand U76638 ( n11674, n18795, n18796 );
nand U76639 ( n18795, n11660, n11663 );
nand U76640 ( n18796, n11664, n18797 );
or U76641 ( n18797, n11663, n11660 );
nor U76642 ( n49837, n49841, n49842 );
nor U76643 ( n49841, n49843, n49844 );
or U76644 ( n16866, n16867, n16868 );
nand U76645 ( n11663, n18798, n18799 );
nand U76646 ( n18798, n11648, n11650 );
nand U76647 ( n18799, n11652, n18800 );
or U76648 ( n18800, n11650, n11648 );
nand U76649 ( n49954, n49955, n49956 );
nor U76650 ( n17017, n2812, n16887 );
nand U76651 ( n51761, n53890, n53891 );
nand U76652 ( n53890, n49645, n49646 );
nand U76653 ( n53891, n49647, n53892 );
or U76654 ( n53892, n49646, n49645 );
nor U76655 ( n16899, n16900, n2837 );
not U76656 ( n2837, n16901 );
nor U76657 ( n16900, n16902, n16903 );
nor U76658 ( n16902, n2824, n16904 );
nor U76659 ( n16882, n16886, n16887 );
nor U76660 ( n16886, n16888, n16889 );
nand U76661 ( n16999, n17000, n17001 );
nand U76662 ( n16673, n20976, n20977 );
nand U76663 ( n20977, n20978, n2378 );
nor U76664 ( n20976, n20979, n20980 );
nor U76665 ( n20979, n2422, n20987 );
nand U76666 ( n18805, n20934, n20935 );
or U76667 ( n20934, n16673, n16675 );
nand U76668 ( n20935, n16674, n20936 );
nand U76669 ( n20936, n16675, n16673 );
nand U76670 ( n49617, n53896, n53897 );
or U76671 ( n53896, n49587, n49590 );
nand U76672 ( n53897, n49589, n53898 );
nand U76673 ( n53898, n49590, n49587 );
nand U76674 ( n49874, n49875, n49876 );
nand U76675 ( n49876, n49877, n49878 );
nand U76676 ( n49778, n1594, n1604 );
nand U76677 ( n16919, n16920, n16921 );
nand U76678 ( n16921, n16922, n16923 );
nand U76679 ( n16823, n2712, n2725 );
nand U76680 ( n49894, n49912, n49913 );
nand U76681 ( n49913, n49914, n49915 );
nand U76682 ( n49906, n49905, n49907 );
nand U76683 ( n49907, n49903, n49908 );
nand U76684 ( n49820, n1658, n1670 );
nand U76685 ( n16918, n16924, n16925 );
nand U76686 ( n16924, n2860, n16932 );
nand U76687 ( n16925, n16926, n16927 );
not U76688 ( n2860, n16926 );
nand U76689 ( n16927, n16928, n16929 );
nand U76690 ( n16928, n2864, n2868 );
or U76691 ( n16929, n16930, n16931 );
nand U76692 ( n16865, n2779, n2790 );
nand U76693 ( n16951, n16950, n16952 );
nand U76694 ( n16952, n16948, n16953 );
nand U76695 ( n40845, n41234, n41235 );
nand U76696 ( n41234, n40739, n40741 );
nand U76697 ( n41235, n41236, n40742 );
or U76698 ( n41236, n40741, n40739 );
nand U76699 ( n40706, n40837, n40838 );
nor U76700 ( n40837, n40846, n40847 );
nor U76701 ( n40838, n40839, n40840 );
nor U76702 ( n40840, n610, n40841 );
nand U76703 ( n40862, n40681, n41348 );
nand U76704 ( n41348, n40687, n40684 );
nand U76705 ( n40725, n41330, n41331 );
nand U76706 ( n41330, n41417, n41418 );
nand U76707 ( n41331, n41332, n589 );
nand U76708 ( n41417, n41419, n41102 );
nand U76709 ( n40741, n41238, n41239 );
nand U76710 ( n41238, n41126, n41128 );
nand U76711 ( n41239, n41240, n41129 );
or U76712 ( n41240, n41128, n41126 );
nand U76713 ( n40810, n40811, n40703 );
nand U76714 ( n40811, n76851, n40812 );
nand U76715 ( n40812, n40813, n40814 );
nand U76716 ( n40813, n40820, n40816 );
nand U76717 ( n40781, n41161, n40777 );
nand U76718 ( n41003, n40964, n40966 );
nand U76719 ( n40687, n40683, n41349 );
nand U76720 ( n41349, n40685, n41194 );
nor U76721 ( n40839, n40842, n40843 );
nand U76722 ( n40843, n40844, n40845 );
nand U76723 ( n40844, n610, n40841 );
nand U76724 ( n41128, n41242, n41243 );
nor U76725 ( n41242, n41289, n41290 );
nor U76726 ( n41243, n41244, n41245 );
nor U76727 ( n41290, n40908, n40907 );
nand U76728 ( n40814, n40815, n602 );
not U76729 ( n602, n40816 );
nor U76730 ( n40815, n40817, n40818 );
nor U76731 ( n40818, n40819, n40706 );
nor U76732 ( n41332, n41111, n41110 );
nand U76733 ( n40701, n40702, n40703 );
nand U76734 ( n40702, n76850, n40704 );
xor U76735 ( n40704, n600, n40705 );
xor U76736 ( n40705, n40706, n40707 );
nand U76737 ( n40944, n41230, n41231 );
nand U76738 ( n41230, n595, n40845 );
nand U76739 ( n41231, n41232, n41019 );
or U76740 ( n41232, n40845, n595 );
and U76741 ( n41211, n41220, n41221 );
xnor U76742 ( n41221, n41215, n41216 );
nor U76743 ( n41220, n41225, n40846 );
and U76744 ( n41225, n41214, n40944 );
nand U76745 ( n41206, n41217, n40703 );
nand U76746 ( n41217, n41218, n41219 );
nor U76747 ( n41218, n41229, n40944 );
nor U76748 ( n41219, n41211, n40846 );
nand U76749 ( n36304, n36431, n36432 );
nand U76750 ( n36432, n2012, n36433 );
nand U76751 ( n36433, n36434, n36435 );
nand U76752 ( n36434, n36436, n36437 );
nand U76753 ( n36460, n36277, n36983 );
nand U76754 ( n36983, n36283, n36280 );
nand U76755 ( n36745, n36861, n36862 );
nand U76756 ( n36861, n36894, n36895 );
nand U76757 ( n36862, n36863, n2019 );
nand U76758 ( n36894, n36896, n36504 );
nand U76759 ( n36629, n36851, n36852 );
nand U76760 ( n36851, n36335, n36337 );
nand U76761 ( n36852, n36853, n36338 );
or U76762 ( n36853, n36337, n36335 );
nand U76763 ( n36378, n36778, n36374 );
nand U76764 ( n36610, n36569, n36571 );
nand U76765 ( n36283, n36279, n36984 );
nand U76766 ( n36984, n36281, n36813 );
or U76767 ( n36431, n75717, n36835 );
or U76768 ( n75717, n36838, n2013 );
nand U76769 ( n36835, n36629, n36632 );
nor U76770 ( n36863, n36397, n36700 );
nand U76771 ( n36337, n36856, n36857 );
nand U76772 ( n36856, n36743, n36745 );
nand U76773 ( n36857, n36858, n36746 );
or U76774 ( n36858, n36745, n36743 );
nand U76775 ( n36411, n36418, n36414 );
nor U76776 ( n36418, n36417, n36430 );
nor U76777 ( n36430, n1838, n36415 );
not U76778 ( n1838, n36304 );
nand U76779 ( n36320, n36962, n36963 );
nand U76780 ( n36962, n37050, n37051 );
nand U76781 ( n36963, n36964, n1964 );
nand U76782 ( n37050, n37052, n36718 );
and U76783 ( n36964, n36727, n36726 );
nand U76784 ( n36412, n36413, n2022 );
not U76785 ( n2022, n36414 );
nor U76786 ( n36413, n36415, n36416 );
nor U76787 ( n36416, n36417, n36304 );
nand U76788 ( n40939, n40940, n40703 );
nand U76789 ( n40940, n76851, n40941 );
xor U76790 ( n40941, n40942, n40943 );
xor U76791 ( n40943, n40944, n40945 );
xor U76792 ( n36302, n36303, n36304 );
nand U76793 ( n36548, n36439, n36835 );
not U76794 ( n2035, n36424 );
not U76795 ( n2037, n37766 );
nand U76796 ( n41015, n41016, n40703 );
nand U76797 ( n41016, n76851, n41017 );
xor U76798 ( n41017, n40841, n41018 );
xor U76799 ( n41018, n40845, n610 );
nor U76800 ( n36842, n2010, n36431 );
not U76801 ( n2010, n36435 );
nand U76802 ( n37178, n37179, n37180 );
nand U76803 ( n37180, n37181, n37182 );
nor U76804 ( n37179, n37183, n37184 );
and U76805 ( n37184, n37185, n37186 );
nand U76806 ( n37125, n37126, n37127 );
nor U76807 ( n37126, n37289, n37290 );
nor U76808 ( n37127, n37128, n37129 );
nor U76809 ( n37290, n37291, n37292 );
nand U76810 ( n37145, n37146, n37147 );
nand U76811 ( n37147, n37148, n37149 );
nor U76812 ( n37146, n37150, n37151 );
and U76813 ( n37151, n37152, n37153 );
or U76814 ( n36546, n75718, n36548 );
xnor U76815 ( n75718, n36549, n2014 );
not U76816 ( n1900, n38886 );
not U76817 ( n1903, n39104 );
nand U76818 ( n39430, n37498, n39481 );
or U76819 ( n39481, n39482, n37551 );
not U76820 ( n1904, n37591 );
not U76821 ( n1905, n40273 );
nor U76822 ( n40014, n40068, n37266 );
and U76823 ( n40068, n40069, n37592 );
nor U76824 ( n40069, n1922, n40072 );
nor U76825 ( n40072, n1904, n40073 );
nand U76826 ( n38916, n38924, n38925 );
nand U76827 ( n38924, n38936, n37331 );
nand U76828 ( n38925, n2135, n38926 );
nand U76829 ( n38936, n38937, n38938 );
and U76830 ( n39847, n39848, n1943 );
nor U76831 ( n39011, n1900, n38956 );
not U76832 ( n590, n40778 );
not U76833 ( n1902, n38818 );
nand U76834 ( n38786, n1902, n2043 );
nor U76835 ( n38781, n37390, n38782 );
nor U76836 ( n38782, n38783, n38784 );
nand U76837 ( n38783, n38787, n38788 );
nand U76838 ( n38784, n38785, n38786 );
nand U76839 ( n38815, n2043, n38818 );
nand U76840 ( n38802, n38803, n38804 );
nand U76841 ( n38803, n38819, n38766 );
nand U76842 ( n38804, n2147, n38805 );
nand U76843 ( n38805, n38806, n38807 );
nand U76844 ( n38814, n2038, n38818 );
nand U76845 ( n38788, n2045, n1902 );
nand U76846 ( n38812, n38816, n38817 );
nand U76847 ( n38816, n2044, n38818 );
nand U76848 ( n38817, n2045, n38818 );
nand U76849 ( n38787, n2044, n1902 );
not U76850 ( n1912, n36375 );
nor U76851 ( n38850, n38867, n2142 );
nor U76852 ( n38867, n38868, n38869 );
nand U76853 ( n38869, n38810, n38814 );
nand U76854 ( n38868, n38880, n38815 );
nand U76855 ( n36626, n36631, n36629 );
nand U76856 ( n36631, n36439, n36632 );
nand U76857 ( n38877, n38900, n38941 );
nand U76858 ( n38941, n38942, n38903 );
nor U76859 ( n38942, n2119, n1884 );
not U76860 ( n1884, n39072 );
not U76861 ( n1887, n39369 );
nand U76862 ( n39678, n39734, n39740 );
nand U76863 ( n39740, n39741, n39737 );
and U76864 ( n39741, n39738, n39742 );
nand U76865 ( n40231, n40282, n40283 );
and U76866 ( n38810, n38870, n38871 );
or U76867 ( n38871, n38857, n38872 );
nor U76868 ( n38870, n38873, n38874 );
nor U76869 ( n38873, n2039, n38860 );
nor U76870 ( n38852, n38853, n38854 );
nand U76871 ( n38854, n1873, n38785 );
nand U76872 ( n38853, n38862, n38786 );
not U76873 ( n1873, n38793 );
nand U76874 ( n40736, n40737, n40703 );
nand U76875 ( n40737, n76852, n40738 );
xnor U76876 ( n40738, n40739, n40740 );
xnor U76877 ( n40740, n40741, n40742 );
nand U76878 ( n62462, n42016, n62775 );
nand U76879 ( n62775, n62776, n41528 );
nand U76880 ( n61438, n42067, n61632 );
nand U76881 ( n61632, n61633, n772 );
not U76882 ( n772, n42062 );
nand U76883 ( n61633, n62273, n62274 );
nand U76884 ( n62274, n62275, n41517 );
nand U76885 ( n62275, n42100, n62350 );
nand U76886 ( n62350, n62351, n41521 );
nand U76887 ( n62351, n42102, n62394 );
nand U76888 ( n62394, n62395, n41529 );
nand U76889 ( n61396, n61397, n61398 );
nand U76890 ( n61397, n41952, n61407 );
nand U76891 ( n61398, n61399, n41952 );
nand U76892 ( n61407, n61408, n61409 );
nand U76893 ( n61404, n564, n835 );
nand U76894 ( n61435, n835, n61438 );
nor U76895 ( n61425, n61427, n61428 );
nor U76896 ( n61428, n61429, n61430 );
nor U76897 ( n61427, n42061, n61431 );
nor U76898 ( n61431, n61432, n61433 );
nand U76899 ( n61432, n61436, n61437 );
nand U76900 ( n61436, n824, n61438 );
nand U76901 ( n61437, n825, n61438 );
nand U76902 ( n38793, n38855, n38856 );
nand U76903 ( n38856, n2005, n38857 );
nor U76904 ( n38855, n38858, n38859 );
and U76905 ( n38858, n38860, n38861 );
and U76906 ( n38859, n38857, n2047 );
nand U76907 ( n61405, n824, n564 );
xnor U76908 ( n36336, n36337, n36338 );
nor U76909 ( n61602, n61619, n773 );
nor U76910 ( n61619, n61620, n61621 );
nand U76911 ( n61621, n61430, n61434 );
nand U76912 ( n61620, n61629, n61435 );
nand U76913 ( n55954, n61581, n61582 );
nor U76914 ( n61582, n61583, n61584 );
nor U76915 ( n61581, n61599, n45759 );
nor U76916 ( n61583, n779, n76061 );
nand U76917 ( n45756, n45757, n45758 );
nand U76918 ( n45757, n76858, n45759 );
nand U76919 ( n38879, n38900, n38943 );
nand U76920 ( n38943, n38944, n38903 );
nor U76921 ( n38944, n2119, n1874 );
not U76922 ( n1874, n38905 );
nand U76923 ( n39739, n39892, n39894 );
nand U76924 ( n39894, n39895, n39891 );
or U76925 ( n39895, n39890, n1949 );
nand U76926 ( n39259, n39292, n39295 );
nand U76927 ( n39295, n2052, n39291 );
nand U76928 ( n39668, n39734, n39735 );
nand U76929 ( n39735, n39736, n39737 );
and U76930 ( n39736, n39738, n39739 );
nor U76931 ( n61604, n61605, n61606 );
nand U76932 ( n61606, n539, n61403 );
nand U76933 ( n61605, n61614, n61404 );
not U76934 ( n539, n61411 );
nand U76935 ( n38951, n38952, n38953 );
nand U76936 ( n38952, n38955, n38921 );
nand U76937 ( n38953, n38954, n38921 );
nor U76938 ( n38955, n38922, n38956 );
nand U76939 ( n40898, n517, n40905 );
not U76940 ( n517, n40904 );
nor U76941 ( n40895, n40901, n40902 );
nand U76942 ( n40902, n40903, n40900 );
nand U76943 ( n40903, n40898, n40906 );
or U76944 ( n40073, n37274, n1927 );
nand U76945 ( n38188, n38977, n38978 );
nor U76946 ( n38978, n38979, n38980 );
nor U76947 ( n38977, n39001, n39002 );
nor U76948 ( n38979, n2039, n38995 );
nand U76949 ( n39002, n39003, n39004 );
nand U76950 ( n39003, n39012, n37343 );
nand U76951 ( n39004, n39005, n38933 );
nand U76952 ( n39012, n39013, n39014 );
nand U76953 ( n40900, n597, n40904 );
not U76954 ( n597, n40905 );
nor U76955 ( n37104, n2043, n2038 );
not U76956 ( n615, n40825 );
nand U76957 ( n41123, n41124, n40703 );
nand U76958 ( n41124, n76850, n41125 );
xnor U76959 ( n41125, n41126, n41127 );
xnor U76960 ( n41127, n41128, n41129 );
nand U76961 ( n36509, n36698, n36699 );
or U76962 ( n36699, n36700, n36397 );
nor U76963 ( n36501, n36502, n36503 );
nand U76964 ( n36503, n36504, n36505 );
nand U76965 ( n36505, n1843, n2018 );
nand U76966 ( n62473, n62575, n62576 );
nand U76967 ( n62576, n62577, n62578 );
nand U76968 ( n62254, n62471, n62472 );
nand U76969 ( n62472, n62473, n62474 );
nand U76970 ( n61609, n61587, n61627 );
nand U76971 ( n61627, n61628, n61590 );
nand U76972 ( n61628, n62249, n62286 );
nand U76973 ( n62286, n62287, n62252 );
nor U76974 ( n62287, n753, n540 );
not U76975 ( n753, n62253 );
nand U76976 ( n62577, n62674, n62675 );
and U76977 ( n62674, n62681, n62682 );
nand U76978 ( n62675, n62676, n62677 );
nand U76979 ( n62682, n62683, n62679 );
nand U76980 ( n66203, n66204, n66205 );
and U76981 ( n66204, n66206, n66207 );
and U76982 ( n64379, n64804, n64805 );
and U76983 ( n61430, n61622, n61623 );
or U76984 ( n61623, n61609, n61624 );
nor U76985 ( n61622, n61625, n61626 );
nor U76986 ( n61625, n833, n61609 );
nand U76987 ( n41079, n41080, n40703 );
nand U76988 ( n41080, n76850, n41081 );
xor U76989 ( n41081, n40905, n41082 );
xor U76990 ( n41082, n40904, n608 );
not U76991 ( n1922, n37271 );
xnor U76992 ( n36744, n36745, n36746 );
not U76993 ( n2038, n38956 );
nor U76994 ( n62258, n767, n62259 );
not U76995 ( n767, n41926 );
nor U76996 ( n62259, n62260, n62261 );
nand U76997 ( n62261, n62262, n62263 );
nand U76998 ( n56052, n62238, n62239 );
nor U76999 ( n62239, n62240, n62241 );
nor U77000 ( n62238, n61296, n46003 );
nor U77001 ( n62241, n775, n76060 );
nor U77002 ( n62271, n62272, n61633 );
nor U77003 ( n62268, n61618, n61633 );
and U77004 ( n40109, n40113, n40114 );
nor U77005 ( n39043, n2124, n39044 );
nor U77006 ( n39044, n39045, n39046 );
nand U77007 ( n39045, n39051, n39052 );
nand U77008 ( n39046, n39047, n39048 );
nand U77009 ( n62285, n62337, n62338 );
nor U77010 ( n62337, n62341, n62342 );
nor U77011 ( n62338, n62339, n62340 );
and U77012 ( n62341, n62275, n835 );
nor U77013 ( n62276, n62277, n62278 );
nand U77014 ( n62278, n62279, n62280 );
nand U77015 ( n62277, n62281, n62282 );
or U77016 ( n62279, n61628, n61624 );
and U77017 ( n62340, n62275, n824 );
nor U77018 ( n38935, n38872, n38877 );
nand U77019 ( n61411, n61607, n61608 );
nand U77020 ( n61608, n822, n61609 );
nor U77021 ( n61607, n61610, n61611 );
and U77022 ( n61610, n61609, n61613 );
and U77023 ( n61611, n61609, n61612 );
not U77024 ( n1885, n38990 );
and U77025 ( n38937, n75719, n75720 );
nand U77026 ( n75719, n38879, n38861 );
nand U77027 ( n75720, n38877, n2047 );
nand U77028 ( n39243, n39127, n37546 );
nor U77029 ( n39169, n2112, n39171 );
nor U77030 ( n39171, n39172, n39173 );
and U77031 ( n39172, n38792, n37402 );
nand U77032 ( n39173, n39229, n39230 );
nor U77033 ( n39229, n39233, n39234 );
nor U77034 ( n39230, n39231, n39232 );
nor U77035 ( n39234, n39194, n38956 );
nand U77036 ( n39156, n39164, n39165 );
nand U77037 ( n39164, n39176, n37326 );
nand U77038 ( n39165, n2114, n39166 );
nand U77039 ( n39176, n39177, n39178 );
xor U77040 ( n71530, n71655, n72070 );
xor U77041 ( n72070, n71653, n71654 );
xnor U77042 ( n72523, n72539, n72757 );
xnor U77043 ( n72757, n72540, n72537 );
xnor U77044 ( n72282, n72379, n72380 );
xnor U77045 ( n72379, n72381, n72382 );
xnor U77046 ( n71955, n72173, n72174 );
xnor U77047 ( n72173, n72175, n72176 );
nor U77048 ( n72408, n72411, n1107 );
nor U77049 ( n72281, n72284, n1083 );
nor U77050 ( n72525, n72733, n1179 );
nor U77051 ( n71954, n71957, n1062 );
not U77052 ( n1140, n72502 );
xnor U77053 ( n72409, n72609, n72496 );
xnor U77054 ( n72609, n72497, n72494 );
not U77055 ( n1030, n71345 );
nand U77056 ( n71340, n71521, n71522 );
nand U77057 ( n71522, n71346, n1030 );
nor U77058 ( n71521, n71524, n71525 );
and U77059 ( n71525, n1032, n71347 );
nand U77060 ( n71053, n71057, n71056 );
nor U77061 ( n71524, n71523, n71526 );
xor U77062 ( n71526, n1030, n1032 );
nor U77063 ( n72651, n72652, n72503 );
nor U77064 ( n72652, n72653, n72504 );
nor U77065 ( n72653, n72649, n72502 );
nor U77066 ( n71939, n71940, n71531 );
nor U77067 ( n71940, n71941, n71532 );
nor U77068 ( n71941, n71937, n71530 );
nand U77069 ( MUL_1411_U378, n71074, n71075 );
nand U77070 ( n71074, n71079, n71078 );
nand U77071 ( n71075, n1018, n71076 );
nand U77072 ( n71079, n71053, n71328 );
xnor U77073 ( n71646, n71643, n72297 );
xnor U77074 ( n72297, n71641, n71642 );
nand U77075 ( n71497, n71534, n71535 );
nand U77076 ( n71535, n71362, n1044 );
nor U77077 ( n71534, n71537, n71538 );
nor U77078 ( n71537, n71536, n71539 );
nand U77079 ( n71086, n71348, n71349 );
nand U77080 ( n71349, n71114, n1034 );
nor U77081 ( n71348, n71352, n71353 );
nor U77082 ( n71353, n71351, n71113 );
nor U77083 ( n71538, n71360, n1039 );
not U77084 ( n1039, n71363 );
nor U77085 ( n71352, n71354, n71355 );
xor U77086 ( n71355, n71351, n71350 );
nor U77087 ( n72186, n72187, n71647 );
nor U77088 ( n72187, n72188, n71648 );
nor U77089 ( n72188, n1052, n71646 );
nand U77090 ( n71655, n72183, n72184 );
nand U77091 ( n72184, n71649, n1059 );
nor U77092 ( n72183, n72185, n72186 );
nor U77093 ( n72185, n1059, n72190 );
nand U77094 ( n71361, n71650, n71651 );
or U77095 ( n71650, n71655, n71654 );
nand U77096 ( n71651, n71652, n71653 );
nand U77097 ( n71652, n71654, n71655 );
nand U77098 ( n71328, n1022, n71052 );
or U77099 ( n71052, n71056, n71057 );
nand U77100 ( n71495, n71528, n71529 );
nand U77101 ( n71529, n71530, n71531 );
nor U77102 ( n71528, n71532, n71533 );
not U77103 ( n1032, n71344 );
nand U77104 ( n36692, n36697, n36509 );
nand U77105 ( n36697, n2018, n36510 );
not U77106 ( n613, n40830 );
nor U77107 ( n39057, n39058, n39059 );
nand U77108 ( n39059, n39060, n39061 );
nand U77109 ( n39058, n39064, n39065 );
nand U77110 ( n39061, n2038, n39020 );
and U77111 ( n39065, n75721, n75722 );
nand U77112 ( n75721, n39020, n2045 );
nand U77113 ( n75722, n39020, n2044 );
nor U77114 ( n39060, n39062, n39063 );
nor U77115 ( n39062, n38872, n38990 );
and U77116 ( n39063, n39020, n2043 );
not U77117 ( n1033, n71351 );
nor U77118 ( n71110, n71111, n71112 );
nor U77119 ( n71111, n1033, n1034 );
nand U77120 ( n71112, n71113, n1028 );
not U77121 ( n1028, n71114 );
not U77122 ( n1018, n71078 );
not U77123 ( n840, n67226 );
nand U77124 ( n61408, n61411, n61412 );
and U77125 ( n71090, n71342, n71343 );
nand U77126 ( n71343, n71344, n71345 );
nor U77127 ( n71342, n71346, n71347 );
not U77128 ( n643, n42092 );
or U77129 ( n39048, n39020, n38956 );
nand U77130 ( n71660, n71814, n71815 );
nand U77131 ( n71815, n71807, n71811 );
nor U77132 ( n71814, n71803, n71809 );
and U77133 ( n71803, n71810, n71807 );
xor U77134 ( n71350, n71126, n71356 );
xor U77135 ( n71356, n71121, n71125 );
nand U77136 ( n71121, n71358, n71359 );
nand U77137 ( n71359, n71360, n71361 );
nor U77138 ( n71358, n71362, n71363 );
xnor U77139 ( n72683, n72717, n72718 );
xnor U77140 ( n72718, n72719, n72720 );
nor U77141 ( n72682, n72685, n1180 );
not U77142 ( n1875, n38975 );
xor U77143 ( n71563, n71631, n72498 );
xor U77144 ( n72498, n71629, n71630 );
xnor U77145 ( n71590, n71618, n72541 );
xnor U77146 ( n72541, n71619, n71616 );
xnor U77147 ( n71550, n72483, n71637 );
xnor U77148 ( n72483, n71636, n71635 );
nor U77149 ( n71565, n72490, n1109 );
nor U77150 ( n71552, n72395, n1082 );
nor U77151 ( n71592, n72533, n1188 );
not U77152 ( n1147, n71577 );
nor U77153 ( n72510, n72511, n71578 );
nor U77154 ( n72511, n72512, n71579 );
nor U77155 ( n72512, n72508, n71577 );
nand U77156 ( n71647, n72191, n72192 );
or U77157 ( n72191, n72174, n72176 );
nand U77158 ( n72192, n72193, n72175 );
nand U77159 ( n72193, n72176, n72174 );
xor U77160 ( n71539, n71361, n71360 );
nor U77161 ( n38984, n38987, n38988 );
nor U77162 ( n38987, n38990, n38991 );
nor U77163 ( n38988, n1885, n38989 );
nand U77164 ( n38991, n38948, n37343 );
nand U77165 ( n46225, n62309, n62310 );
nor U77166 ( n62310, n62311, n62312 );
nor U77167 ( n62309, n62332, n62333 );
nor U77168 ( n62311, n833, n62326 );
nand U77169 ( n56148, n62294, n62295 );
nor U77170 ( n62295, n62296, n62297 );
nor U77171 ( n62294, n61296, n46225 );
nor U77172 ( n62297, n768, n76059 );
nand U77173 ( n62333, n62334, n62335 );
nand U77174 ( n62335, n62336, n62285 );
nand U77175 ( n62334, n62343, n41937 );
nand U77176 ( n62336, n41517, n62273 );
nor U77177 ( n38130, n38765, n38766 );
or U77178 ( n38765, n38767, n38768 );
nor U77179 ( n38767, n38770, n38772 );
nor U77180 ( n38768, n2147, n38769 );
and U77181 ( n71533, n71937, n71531 );
nand U77182 ( n71113, n71354, n71350 );
and U77183 ( n71339, n71662, n71663 );
nand U77184 ( n71662, n71045, n71047 );
nand U77185 ( n71663, n71048, n71664 );
or U77186 ( n71664, n71047, n71045 );
nor U77187 ( n62349, n62272, n62275 );
nand U77188 ( n71375, n71638, n71639 );
nand U77189 ( n71638, n71643, n71642 );
nand U77190 ( n71639, n71640, n71641 );
or U77191 ( n71640, n71642, n71643 );
nor U77192 ( n62346, n61618, n62275 );
nor U77193 ( n39098, n2118, n39099 );
nor U77194 ( n39099, n39100, n39101 );
nand U77195 ( n39100, n39107, n39108 );
nand U77196 ( n39101, n39102, n39103 );
not U77197 ( n2023, n36423 );
nand U77198 ( n71082, n71083, n71084 );
nand U77199 ( n71084, n71085, n71086 );
and U77200 ( n71362, n71536, n71360 );
nor U77201 ( n71377, n1060, n1057 );
and U77202 ( n71346, n71523, n71344 );
nand U77203 ( n62657, n42014, n62665 );
nand U77204 ( n62567, n62651, n62652 );
nor U77205 ( n62651, n62655, n62656 );
nor U77206 ( n62652, n62653, n62654 );
nor U77207 ( n62656, n62586, n62272 );
nor U77208 ( n62563, n62465, n62565 );
nor U77209 ( n62565, n62566, n62567 );
nor U77210 ( n62566, n823, n42015 );
nand U77211 ( n57363, n62537, n62538 );
nor U77212 ( n62538, n62539, n62540 );
nor U77213 ( n62537, n61296, n47420 );
nor U77214 ( n62540, n754, n76061 );
nand U77215 ( n72680, n72707, n72708 );
or U77216 ( n72707, n72672, n72670 );
nand U77217 ( n72708, n72673, n72709 );
nand U77218 ( n72709, n72670, n72672 );
nand U77219 ( n71089, n1027, n71083 );
not U77220 ( n1027, n71086 );
nand U77221 ( n71629, n72500, n72501 );
nand U77222 ( n72501, n72502, n72503 );
nor U77223 ( n72500, n72504, n72505 );
nor U77224 ( n62653, n62586, n61618 );
nand U77225 ( n71126, n71364, n71365 );
nand U77226 ( n71365, n71321, n1048 );
nor U77227 ( n71364, n71367, n71368 );
nor U77228 ( n71367, n71366, n71369 );
not U77229 ( n1048, n71320 );
nor U77230 ( n71368, n71319, n1040 );
not U77231 ( n1040, n71322 );
and U77232 ( n71490, n71644, n71645 );
nand U77233 ( n71645, n71646, n71647 );
nor U77234 ( n71644, n71648, n71649 );
and U77235 ( n71649, n1052, n71647 );
xor U77236 ( n71319, n71316, n71370 );
xor U77237 ( n71370, n71140, n71315 );
xor U77238 ( n71369, n71320, n71319 );
nand U77239 ( n71942, n1037, n71531 );
nand U77240 ( n72654, n1124, n72503 );
nand U77241 ( n72524, n72735, n72736 );
or U77242 ( n72735, n72719, n72717 );
nand U77243 ( n72736, n72720, n72737 );
nand U77244 ( n72737, n72717, n72719 );
nand U77245 ( n72734, n72733, n72524 );
buf U77246 ( n76391, n75765 );
nand U77247 ( n62280, n538, n61612 );
and U77248 ( n72505, n72649, n72503 );
nand U77249 ( n56372, n62354, n62355 );
nor U77250 ( n62355, n62356, n62357 );
nor U77251 ( n62354, n61599, n46555 );
nor U77252 ( n62356, n764, n76065 );
nor U77253 ( n62369, n757, n62370 );
nor U77254 ( n62370, n62371, n62372 );
nand U77255 ( n62371, n62377, n62378 );
nand U77256 ( n62372, n62373, n62374 );
nand U77257 ( n71026, n71801, n71802 );
nand U77258 ( n71802, n71803, n1047 );
nor U77259 ( n71801, n71804, n71805 );
nor U77260 ( n71805, n71806, n71807 );
and U77261 ( n71804, n71807, n75723 );
nor U77262 ( n75723, n71810, n1047 );
nor U77263 ( n71976, n71977, n1118 );
nor U77264 ( n72257, n72258, n1193 );
nand U77265 ( n72260, n72333, n72334 );
nand U77266 ( n72333, n72248, n72245 );
nand U77267 ( n72334, n72247, n72335 );
or U77268 ( n72335, n72245, n72248 );
nand U77269 ( n71926, n71965, n71966 );
nand U77270 ( n71965, n71913, n71912 );
nand U77271 ( n71966, n71914, n71967 );
or U77272 ( n71967, n71912, n71913 );
not U77273 ( n1154, n72163 );
nor U77274 ( n72253, n72254, n72255 );
nor U77275 ( n72254, n72256, n72257 );
and U77276 ( n72256, n72258, n1193 );
nor U77277 ( n72157, n72158, n72159 );
nor U77278 ( n72158, n72160, n72161 );
nor U77279 ( n72160, n72162, n72163 );
nor U77280 ( n71972, n71973, n71974 );
nor U77281 ( n71973, n71975, n71976 );
and U77282 ( n71975, n71977, n1118 );
and U77283 ( n71809, n71810, n71811 );
and U77284 ( n71794, n71915, n71916 );
nand U77285 ( n71916, n71917, n1089 );
nor U77286 ( n71915, n71918, n71919 );
nor U77287 ( n71918, n1088, n71925 );
and U77288 ( n71799, n71831, n71832 );
nand U77289 ( n71832, n71686, n71691 );
nor U77290 ( n71831, n71682, n71688 );
nand U77291 ( n71979, n72113, n72114 );
or U77292 ( n72113, n71982, n71985 );
nand U77293 ( n72114, n71984, n72115 );
nand U77294 ( n72115, n71985, n71982 );
nand U77295 ( n71691, n71833, n71834 );
nand U77296 ( n71833, n71794, n71795 );
nand U77297 ( n71834, n71796, n71835 );
or U77298 ( n71835, n71795, n71794 );
nand U77299 ( n62308, n62290, n62398 );
nand U77300 ( n62398, n62254, n62253 );
nand U77301 ( n71551, n72397, n72398 );
nand U77302 ( n72397, n72381, n72380 );
nand U77303 ( n72398, n72382, n72399 );
or U77304 ( n72399, n72380, n72381 );
nand U77305 ( n72396, n72395, n71551 );
nor U77306 ( n39113, n39114, n39115 );
nand U77307 ( n39114, n39120, n39121 );
nand U77308 ( n39115, n39116, n39117 );
nor U77309 ( n39121, n39122, n39123 );
nand U77310 ( n62281, n538, n61613 );
nand U77311 ( n46553, n46554, n45758 );
nand U77312 ( n46554, n76858, n46555 );
nand U77313 ( n38995, n38996, n38973 );
nand U77314 ( n38996, n2125, n38999 );
nand U77315 ( n38999, n1875, n38948 );
xor U77316 ( n45482, n45483, n45484 );
and U77317 ( n62586, n42014, n62665 );
nand U77318 ( n39188, n39189, n39190 );
nand U77319 ( n39189, n39192, n39161 );
nand U77320 ( n39190, n39191, n39161 );
nor U77321 ( n39192, n39193, n38956 );
xnor U77322 ( n72644, n72670, n72671 );
xnor U77323 ( n72671, n72672, n72673 );
nand U77324 ( n72377, n72418, n72419 );
or U77325 ( n72418, n72363, n72366 );
nand U77326 ( n72419, n72420, n72365 );
nand U77327 ( n72420, n72366, n72363 );
nor U77328 ( n72643, n72646, n1182 );
not U77329 ( n1144, n72469 );
nor U77330 ( n72463, n72464, n72465 );
nor U77331 ( n72464, n72466, n72467 );
nor U77332 ( n72466, n72468, n72469 );
nand U77333 ( n72279, n72306, n72307 );
or U77334 ( n72306, n72270, n72272 );
nand U77335 ( n72307, n72308, n72271 );
nand U77336 ( n72308, n72272, n72270 );
xor U77337 ( n38151, n38834, n38770 );
xnor U77338 ( n71374, n71485, n71547 );
xnor U77339 ( n71547, n71483, n71484 );
nand U77340 ( n72513, n1127, n71578 );
and U77341 ( n39221, n39173, n75724 );
or U77342 ( n75724, n37402, n2112 );
nand U77343 ( n71591, n72535, n72536 );
or U77344 ( n72535, n72540, n72539 );
nand U77345 ( n72536, n72537, n72538 );
nand U77346 ( n72538, n72539, n72540 );
nand U77347 ( n72534, n72533, n71591 );
not U77348 ( n2032, n40325 );
nor U77349 ( n62316, n62319, n62320 );
nor U77350 ( n62319, n62308, n62322 );
nor U77351 ( n62320, n542, n62321 );
nand U77352 ( n62322, n62289, n41937 );
nor U77353 ( n71806, n71808, n71809 );
nor U77354 ( n71808, n71810, n71811 );
nand U77355 ( n71388, n71632, n71633 );
or U77356 ( n71632, n71637, n71636 );
nand U77357 ( n71633, n71634, n71635 );
nand U77358 ( n71634, n71636, n71637 );
and U77359 ( n71485, n71554, n71555 );
nand U77360 ( n71555, n71389, n1093 );
nor U77361 ( n71554, n71556, n71557 );
not U77362 ( n1093, n71387 );
nor U77363 ( n39236, n2109, n39238 );
nor U77364 ( n39238, n39239, n39240 );
nand U77365 ( n39239, n39246, n39247 );
nand U77366 ( n39240, n39241, n39242 );
nor U77367 ( n62386, n62388, n62389 );
and U77368 ( n62389, n62351, n835 );
nor U77369 ( n62388, n61624, n62308 );
xnor U77370 ( n72091, n72269, n72270 );
xnor U77371 ( n72269, n72271, n72272 );
nand U77372 ( n72175, n72194, n72195 );
nand U77373 ( n72195, n72091, n72088 );
nor U77374 ( n72194, n72090, n72084 );
nand U77375 ( n72406, n72557, n72558 );
or U77376 ( n72557, n72414, n72417 );
nand U77377 ( n72558, n72559, n72416 );
nand U77378 ( n72559, n72417, n72414 );
nor U77379 ( n72601, n72602, n72603 );
nor U77380 ( n72602, n72604, n72605 );
nor U77381 ( n72604, n72606, n72607 );
and U77382 ( n72605, n72606, n72607 );
nand U77383 ( n72410, n72411, n72406 );
nor U77384 ( n72086, n72087, n72088 );
nor U77385 ( n72087, n72089, n72090 );
nor U77386 ( n72089, n1074, n72091 );
nand U77387 ( n71952, n72079, n72080 );
nand U77388 ( n72079, n72054, n72056 );
nand U77389 ( n72080, n72057, n72081 );
or U77390 ( n72081, n72056, n72054 );
and U77391 ( n72057, n72082, n72083 );
nand U77392 ( n72083, n72084, n1084 );
nor U77393 ( n72082, n72085, n72086 );
nor U77394 ( n72085, n1084, n72092 );
xor U77395 ( n72208, n72363, n72364 );
xor U77396 ( n72364, n72365, n72366 );
xor U77397 ( n72048, n72169, n72170 );
xor U77398 ( n72169, n72171, n72172 );
nor U77399 ( n72207, n72210, n1113 );
buf U77400 ( n76460, n75766 );
nand U77401 ( n72052, n72096, n72097 );
nand U77402 ( n72096, n72038, n72040 );
nand U77403 ( n72097, n72041, n72098 );
or U77404 ( n72098, n72040, n72038 );
nand U77405 ( n71829, n71960, n71961 );
nand U77406 ( n71960, n71927, n71930 );
nand U77407 ( n71961, n71929, n71962 );
or U77408 ( n71962, n71930, n71927 );
nor U77409 ( n72355, n72356, n1190 );
nor U77410 ( n71970, n71977, n1117 );
nand U77411 ( n72040, n72111, n72112 );
nand U77412 ( n72112, n71974, n71979 );
nor U77413 ( n72111, n71970, n71976 );
not U77414 ( n1117, n71974 );
nand U77415 ( n72358, n72444, n72445 );
nand U77416 ( n72444, n72346, n72343 );
nand U77417 ( n72445, n72345, n72446 );
or U77418 ( n72446, n72343, n72346 );
nor U77419 ( n72220, n72221, n72222 );
nor U77420 ( n72221, n72223, n72224 );
nor U77421 ( n72223, n72225, n72226 );
not U77422 ( n1152, n72226 );
nor U77423 ( n71823, n71824, n71825 );
nor U77424 ( n71824, n71826, n71827 );
nor U77425 ( n71826, n71828, n71829 );
nor U77426 ( n72351, n72352, n72353 );
nor U77427 ( n72352, n72354, n72355 );
and U77428 ( n72354, n72356, n1190 );
and U77429 ( n71827, n71828, n71829 );
xnor U77430 ( n72590, n72631, n72632 );
xnor U77431 ( n72632, n72633, n72634 );
nor U77432 ( n72589, n72592, n1183 );
not U77433 ( n1047, n71811 );
and U77434 ( n62393, n62351, n824 );
nand U77435 ( n72496, n72610, n72611 );
nand U77436 ( n72611, n72603, n72607 );
nor U77437 ( n72610, n72605, n72599 );
nand U77438 ( n71564, n72492, n72493 );
nand U77439 ( n72492, n72497, n72496 );
nand U77440 ( n72493, n72494, n72495 );
or U77441 ( n72495, n72496, n72497 );
nand U77442 ( n72491, n72490, n71564 );
nand U77443 ( n71155, n71480, n71481 );
nand U77444 ( n71480, n71485, n71484 );
nand U77445 ( n71481, n71482, n71483 );
or U77446 ( n71482, n71484, n71485 );
nand U77447 ( n71316, n71378, n71379 );
or U77448 ( n71379, n71154, n71155 );
nor U77449 ( n71378, n71381, n71382 );
nor U77450 ( n71382, n71156, n71153 );
and U77451 ( n71321, n71366, n71319 );
nand U77452 ( n62326, n62327, n62306 );
nand U77453 ( n62327, n758, n62330 );
nand U77454 ( n62330, n542, n62289 );
or U77455 ( n71830, n71828, n1064 );
nand U77456 ( n72088, n72196, n72197 );
nand U77457 ( n72196, n72170, n72171 );
nand U77458 ( n72197, n72172, n72198 );
or U77459 ( n72198, n72171, n72170 );
and U77460 ( n72084, n1074, n72088 );
not U77461 ( n1143, n72607 );
or U77462 ( n72608, n72606, n1143 );
xor U77463 ( n71908, n71982, n71983 );
xor U77464 ( n71983, n71984, n71985 );
nand U77465 ( n71795, n71836, n71837 );
nand U77466 ( n71837, n71787, n71792 );
nor U77467 ( n71836, n71783, n71789 );
nand U77468 ( n71792, n71838, n71839 );
nand U77469 ( n71838, n71778, n71779 );
nand U77470 ( n71839, n71780, n71840 );
or U77471 ( n71840, n71779, n71778 );
nor U77472 ( n71903, n71904, n71905 );
nor U77473 ( n71904, n71906, n71907 );
nor U77474 ( n71906, n1103, n71908 );
and U77475 ( n71778, n71899, n71900 );
nand U77476 ( n71900, n71901, n1119 );
nor U77477 ( n71899, n71902, n71903 );
nor U77478 ( n71902, n1119, n71909 );
nand U77479 ( n72283, n72284, n72279 );
or U77480 ( n62374, n62351, n62272 );
xnor U77481 ( n71787, n71911, n71912 );
xnor U77482 ( n71911, n71913, n71914 );
not U77483 ( n1115, n72110 );
and U77484 ( n72041, n72099, n72100 );
nand U77485 ( n72100, n72101, n1115 );
nor U77486 ( n72099, n72102, n72103 );
nor U77487 ( n72102, n1114, n72109 );
and U77488 ( n72599, n72606, n72603 );
nand U77489 ( n39103, n2038, n39104 );
nand U77490 ( n71912, n71980, n71981 );
nand U77491 ( n71981, n71908, n71905 );
nor U77492 ( n71980, n71901, n71907 );
and U77493 ( n71580, n72508, n71578 );
nand U77494 ( n61450, n61587, n61588 );
nand U77495 ( n61588, n61589, n61590 );
nand U77496 ( n61449, n61450, n61412 );
nand U77497 ( n61589, n62249, n62250 );
nand U77498 ( n62250, n62251, n62252 );
and U77499 ( n62251, n62253, n62254 );
nand U77500 ( n72684, n72685, n72680 );
or U77501 ( n71120, n71126, n71125 );
xnor U77502 ( n71825, n72054, n72055 );
xnor U77503 ( n72055, n72056, n72057 );
and U77504 ( n71821, n71828, n71825 );
xnor U77505 ( n71921, n72038, n72039 );
xnor U77506 ( n72039, n72040, n72041 );
nand U77507 ( n71930, n71963, n71964 );
nand U77508 ( n71964, n71921, n71926 );
nor U77509 ( n71963, n71917, n71923 );
xnor U77510 ( n71686, n71927, n71928 );
xnor U77511 ( n71928, n71929, n71930 );
nand U77512 ( n71991, n72137, n72138 );
nand U77513 ( n72138, n72139, n1195 );
nor U77514 ( n72137, n72140, n72141 );
nor U77515 ( n72140, n1194, n72147 );
nand U77516 ( n72148, n72235, n72236 );
nand U77517 ( n72235, n72136, n72133 );
nand U77518 ( n72236, n72135, n72237 );
or U77519 ( n72237, n72133, n72136 );
not U77520 ( n1157, n72036 );
and U77521 ( n72152, n72233, n72234 );
nand U77522 ( n72234, n72143, n72148 );
nor U77523 ( n72233, n72139, n72145 );
and U77524 ( n71985, n72116, n72117 );
nand U77525 ( n72117, n72032, n72036 );
nor U77526 ( n72116, n72028, n72034 );
nand U77527 ( n72587, n72621, n72622 );
or U77528 ( n72621, n72579, n72577 );
nand U77529 ( n72622, n72580, n72623 );
nand U77530 ( n72623, n72577, n72579 );
nand U77531 ( n71118, n71125, n71126 );
xor U77532 ( n72143, n72245, n72246 );
xor U77533 ( n72246, n72247, n72248 );
xor U77534 ( n38167, n2135, n38837 );
nand U77535 ( n72171, n72211, n72212 );
nand U77536 ( n72212, n72105, n72110 );
nor U77537 ( n72211, n72101, n72107 );
nor U77538 ( n72030, n72031, n72032 );
nor U77539 ( n72031, n72033, n72034 );
nor U77540 ( n72033, n72035, n72036 );
and U77541 ( n71901, n1103, n71905 );
nor U77542 ( n62435, n752, n62436 );
not U77543 ( n752, n41920 );
nor U77544 ( n62436, n62437, n62438 );
nand U77545 ( n62437, n62443, n62444 );
nand U77546 ( n56888, n62421, n62422 );
nor U77547 ( n62422, n62423, n62424 );
nor U77548 ( n62421, n61296, n46942 );
nor U77549 ( n62424, n759, n76064 );
nand U77550 ( n62438, n62439, n62440 );
or U77551 ( n62440, n62395, n62272 );
nor U77552 ( n62439, n62441, n62442 );
nor U77553 ( n62441, n540, n61624 );
not U77554 ( n1943, n37585 );
nand U77555 ( n72164, n1129, n72163 );
xnor U77556 ( n71387, n71479, n71560 );
xnor U77557 ( n71560, n71477, n71478 );
and U77558 ( n71032, n71680, n71681 );
nand U77559 ( n71681, n71682, n1067 );
nor U77560 ( n71680, n71683, n71684 );
nor U77561 ( n71683, n1065, n71690 );
and U77562 ( n71027, n71674, n71675 );
nand U77563 ( n71674, n71041, n71043 );
nand U77564 ( n71675, n71044, n71676 );
or U77565 ( n71676, n71043, n71041 );
nand U77566 ( n71129, n71317, n71318 );
nand U77567 ( n71318, n71319, n71320 );
nor U77568 ( n71317, n71321, n71322 );
nand U77569 ( n38179, n38972, n38973 );
nand U77570 ( n38972, n2125, n38974 );
or U77571 ( n38974, n38975, n2127 );
xor U77572 ( n71156, n71168, n71384 );
xor U77573 ( n71384, n71163, n71167 );
nand U77574 ( n71163, n71385, n71386 );
nand U77575 ( n71386, n71387, n71388 );
nor U77576 ( n71385, n71389, n1077 );
not U77577 ( n1077, n71390 );
nand U77578 ( n72641, n72660, n72661 );
or U77579 ( n72660, n72633, n72631 );
nand U77580 ( n72661, n72634, n72662 );
nand U77581 ( n72662, n72631, n72633 );
nand U77582 ( n72645, n72646, n72641 );
nor U77583 ( n39193, n2112, n39194 );
nor U77584 ( n62556, n62465, n62586 );
nor U77585 ( n62554, n62556, n61618 );
xor U77586 ( n72105, n72265, n72266 );
xor U77587 ( n72266, n72267, n72268 );
and U77588 ( n72267, n72326, n72327 );
nand U77589 ( n72327, n72222, n72226 );
nor U77590 ( n72326, n72218, n72224 );
nand U77591 ( n62580, n62581, n62582 );
nand U77592 ( n62581, n62584, n62555 );
nand U77593 ( n62582, n62583, n62555 );
nor U77594 ( n62584, n62585, n62272 );
nor U77595 ( n39175, n38872, n39134 );
not U77596 ( n1155, n72032 );
xor U77597 ( n72255, n72343, n72344 );
xor U77598 ( n72344, n72345, n72346 );
xor U77599 ( n38199, n38975, n2124 );
nand U77600 ( n62306, n62328, n62329 );
nor U77601 ( n62328, n763, n760 );
nand U77602 ( n62329, n62308, n62325 );
nand U77603 ( n39242, n39194, n2038 );
nand U77604 ( n57455, n62629, n62630 );
nor U77605 ( n62630, n62631, n62632 );
nor U77606 ( n62629, n61599, n47964 );
nor U77607 ( n62631, n750, n76064 );
and U77608 ( n62643, n62567, n75725 );
or U77609 ( n75725, n747, n62465 );
and U77610 ( n72167, n72228, n72229 );
nand U77611 ( n72229, n72159, n72163 );
nor U77612 ( n72228, n72155, n72161 );
nand U77613 ( n72470, n1125, n72465 );
nand U77614 ( n72365, n72421, n72422 );
nand U77615 ( n72422, n72320, n72324 );
nor U77616 ( n72421, n72322, n72316 );
and U77617 ( n72316, n72323, n72320 );
and U77618 ( n39177, n75726, n75727 );
nand U77619 ( n75726, n39137, n38861 );
nand U77620 ( n75727, n39134, n2047 );
nor U77621 ( n72251, n72258, n1192 );
not U77622 ( n1165, n72733 );
nand U77623 ( n47962, n47963, n45758 );
nand U77624 ( n47963, n76858, n47964 );
nand U77625 ( n71956, n71957, n71952 );
nand U77626 ( n71402, n71626, n71627 );
or U77627 ( n71626, n71631, n71630 );
nand U77628 ( n71627, n71628, n71629 );
nand U77629 ( n71628, n71630, n71631 );
not U77630 ( n1153, n72159 );
nand U77631 ( n71978, n71977, n71979 );
not U77632 ( n674, n42077 );
nand U77633 ( n72259, n72258, n72260 );
nor U77634 ( n64811, n674, n64813 );
nor U77635 ( n64813, n41550, n42082 );
nand U77636 ( n38268, n39277, n39278 );
nor U77637 ( n39278, n39279, n39280 );
nor U77638 ( n39277, n39304, n39305 );
nand U77639 ( n39280, n39281, n39282 );
nor U77640 ( n39304, n2103, n39306 );
nor U77641 ( n39306, n39307, n39308 );
nand U77642 ( n39307, n39313, n39314 );
nand U77643 ( n39308, n39309, n39310 );
xor U77644 ( n72373, n72414, n72415 );
xor U77645 ( n72415, n72416, n72417 );
nand U77646 ( n72416, n72560, n72561 );
nand U77647 ( n72561, n72469, n72465 );
nor U77648 ( n72560, n72467, n72461 );
not U77649 ( n1142, n72603 );
nor U77650 ( n62658, n744, n62660 );
nor U77651 ( n62660, n62661, n62662 );
nand U77652 ( n62661, n62668, n62669 );
nand U77653 ( n62662, n62663, n62664 );
not U77654 ( n1883, n39183 );
nand U77655 ( n71178, n71474, n71475 );
nand U77656 ( n71474, n71479, n71478 );
nand U77657 ( n71475, n71476, n71477 );
or U77658 ( n71476, n71478, n71479 );
nand U77659 ( n71168, n71391, n71392 );
or U77660 ( n71392, n71177, n71178 );
nor U77661 ( n71391, n71394, n71395 );
nor U77662 ( n71395, n71179, n71176 );
nor U77663 ( n72318, n72319, n72320 );
nor U77664 ( n72319, n72321, n72322 );
nor U77665 ( n72321, n72323, n72324 );
nand U77666 ( n72440, n72567, n72568 );
nand U77667 ( n72567, n72458, n72455 );
nand U77668 ( n72568, n72457, n72569 );
or U77669 ( n72569, n72455, n72458 );
nor U77670 ( n36605, n1988, n36606 );
not U77671 ( n1988, n36608 );
nand U77672 ( n36606, n36607, n36571 );
nand U77673 ( n36607, n1844, n36570 );
not U77674 ( n1844, n36569 );
nor U77675 ( n36604, n36608, n36609 );
nand U77676 ( n36609, n36610, n36570 );
and U77677 ( n72322, n72323, n72324 );
nor U77678 ( n62452, n62454, n62455 );
and U77679 ( n62455, n62395, n835 );
nor U77680 ( n62454, n61624, n62254 );
xor U77681 ( n72353, n72455, n72456 );
xor U77682 ( n72456, n72457, n72458 );
nor U77683 ( n72349, n72356, n1187 );
not U77684 ( n1150, n72222 );
nand U77685 ( n72205, n72311, n72312 );
or U77686 ( n72311, n72265, n72267 );
nand U77687 ( n72312, n72268, n72313 );
nand U77688 ( n72313, n72267, n72265 );
nor U77689 ( n39170, n2039, n39137 );
not U77690 ( n1167, n72685 );
nor U77691 ( n71571, n71401, n71404 );
xor U77692 ( n71179, n71191, n71398 );
xor U77693 ( n71398, n71186, n71190 );
nand U77694 ( n71186, n71399, n71400 );
nand U77695 ( n71400, n71401, n71402 );
nor U77696 ( n71399, n71403, n1104 );
not U77697 ( n1104, n71404 );
nand U77698 ( n72227, n1128, n72226 );
nand U77699 ( n72357, n72356, n72358 );
not U77700 ( n1149, n72324 );
or U77701 ( n72325, n72323, n1149 );
nor U77702 ( n40998, n599, n40999 );
not U77703 ( n599, n41001 );
nand U77704 ( n40999, n41000, n40966 );
nand U77705 ( n41000, n518, n40965 );
not U77706 ( n518, n40964 );
and U77707 ( n62459, n62395, n824 );
and U77708 ( n62458, n62395, n825 );
nor U77709 ( n40997, n41001, n41002 );
nand U77710 ( n41002, n41003, n40965 );
xor U77711 ( n71401, n71473, n71573 );
xor U77712 ( n71573, n71471, n71472 );
nand U77713 ( n71473, n71581, n71582 );
nand U77714 ( n71582, n71418, n1148 );
nor U77715 ( n71581, n71584, n71585 );
nor U77716 ( n71584, n71583, n71586 );
nor U77717 ( n71585, n71416, n1135 );
not U77718 ( n1135, n71419 );
not U77719 ( n1148, n71417 );
nand U77720 ( n71471, n71575, n71576 );
nand U77721 ( n71576, n71577, n71578 );
nor U77722 ( n71575, n71579, n71580 );
and U77723 ( n72461, n72468, n72465 );
xnor U77724 ( n45471, n45473, n45474 );
not U77725 ( n535, n62760 );
nand U77726 ( n62757, n62969, n62970 );
nand U77727 ( n62969, n535, n822 );
nand U77728 ( n62970, n535, n61612 );
nand U77729 ( n57498, n62730, n62731 );
nor U77730 ( n62731, n62732, n62733 );
nor U77731 ( n62730, n61296, n48079 );
nor U77732 ( n62733, n745, n76063 );
nor U77733 ( n62751, n62753, n62754 );
nor U77734 ( n62754, n559, n61618 );
nor U77735 ( n62753, n734, n62755 );
nor U77736 ( n62755, n62756, n62757 );
not U77737 ( n1872, n39186 );
not U77738 ( n1174, n72533 );
nand U77739 ( n39178, n2005, n39134 );
nor U77740 ( n72006, n72007, n1198 );
not U77741 ( n1198, n72009 );
and U77742 ( n71994, n72121, n72122 );
nand U77743 ( n72122, n72004, n72009 );
nor U77744 ( n72121, n72000, n72006 );
xor U77745 ( n72004, n72133, n72134 );
xor U77746 ( n72134, n72135, n72136 );
nor U77747 ( n72000, n72007, n1197 );
nand U77748 ( n71152, n71153, n71154 );
nand U77749 ( n71130, n71131, n71132 );
nand U77750 ( n71131, n71141, n71142 );
nand U77751 ( n71132, n71133, n71134 );
nor U77752 ( n71141, n71314, n71139 );
and U77753 ( n39898, n39943, n39891 );
not U77754 ( n1145, n72320 );
nand U77755 ( n71779, n71841, n71842 );
nand U77756 ( n71842, n71771, n71776 );
nor U77757 ( n71841, n71767, n71773 );
not U77758 ( n1120, n71771 );
nor U77759 ( n62296, n61443, n46221 );
nand U77760 ( n72209, n72210, n72205 );
and U77761 ( n71030, n71692, n71693 );
nand U77762 ( n71692, n71037, n71039 );
nand U77763 ( n71693, n71040, n71694 );
or U77764 ( n71694, n71039, n71037 );
and U77765 ( n71034, n71781, n71782 );
nand U77766 ( n71782, n71783, n1092 );
nor U77767 ( n71781, n71784, n71785 );
nor U77768 ( n71784, n1090, n71791 );
nand U77769 ( n71039, n71695, n71696 );
nand U77770 ( n71695, n71034, n71035 );
nand U77771 ( n71696, n71036, n71697 );
or U77772 ( n71697, n71035, n71034 );
and U77773 ( n71139, n71316, n71315 );
or U77774 ( n39310, n39127, n38956 );
xnor U77775 ( n72436, n72577, n72578 );
xnor U77776 ( n72578, n72579, n72580 );
nand U77777 ( n41489, n41603, n41604 );
nor U77778 ( n41603, n41879, n41880 );
nor U77779 ( n41604, n41605, n41606 );
nor U77780 ( n41880, n41881, n41882 );
nor U77781 ( n41621, n41625, n41626 );
nor U77782 ( n41626, n41627, n41628 );
nor U77783 ( n41625, n41629, n41630 );
nand U77784 ( n41630, n41631, n41632 );
nor U77785 ( n41675, n41676, n41677 );
nand U77786 ( n41677, n41678, n41679 );
nand U77787 ( n41676, n41686, n41687 );
nor U77788 ( n41678, n41680, n41681 );
nand U77789 ( n41618, n41619, n41620 );
nand U77790 ( n41619, n41840, n41841 );
nand U77791 ( n41620, n41621, n41622 );
nand U77792 ( n41622, n41623, n41624 );
nor U77793 ( n41717, n41718, n41719 );
nor U77794 ( n41718, n41738, n41739 );
nor U77795 ( n41719, n41720, n41721 );
nand U77796 ( n41739, n41726, n642 );
nor U77797 ( n41610, n41611, n41612 );
and U77798 ( n41611, n41847, n41846 );
nand U77799 ( n41612, n41613, n41614 );
nand U77800 ( n41613, n41842, n41843 );
nand U77801 ( n41614, n41615, n41616 );
nor U77802 ( n41615, n41844, n41845 );
nor U77803 ( n41616, n41617, n41618 );
nor U77804 ( n41844, n41623, n41624 );
and U77805 ( n41629, n41628, n41627 );
nor U77806 ( n39222, n39223, n37325 );
nor U77807 ( n39223, n39224, n39225 );
nor U77808 ( n39224, n38872, n39183 );
nand U77809 ( n39225, n39226, n39227 );
nand U77810 ( n39226, n1883, n2047 );
not U77811 ( n1158, n71856 );
not U77812 ( n1122, n71776 );
nor U77813 ( n71850, n71851, n71852 );
nor U77814 ( n71851, n71853, n71854 );
nor U77815 ( n71853, n71855, n71856 );
nor U77816 ( n62585, n62465, n62586 );
xor U77817 ( n71586, n71417, n71416 );
nand U77818 ( n71191, n71405, n71406 );
or U77819 ( n71406, n71200, n71201 );
nor U77820 ( n71405, n71408, n71409 );
nor U77821 ( n71409, n71202, n71199 );
nand U77822 ( n71201, n71468, n71469 );
or U77823 ( n71468, n71473, n71472 );
nand U77824 ( n71469, n71470, n71471 );
nand U77825 ( n71470, n71472, n71473 );
nand U77826 ( n62453, n837, n62395 );
and U77827 ( n71898, n71989, n71990 );
nand U77828 ( n71990, n71856, n71852 );
nor U77829 ( n71989, n71848, n71854 );
nor U77830 ( n71138, n71315, n71316 );
xor U77831 ( n71202, n71216, n71412 );
xor U77832 ( n71412, n71211, n71215 );
nand U77833 ( n71211, n71414, n71415 );
nand U77834 ( n71415, n71416, n71417 );
nor U77835 ( n71414, n71418, n71419 );
nand U77836 ( n72591, n72592, n72587 );
nand U77837 ( n41488, n41489, n76925 );
nand U77838 ( n72037, n1130, n72036 );
nor U77839 ( n39279, n39296, n39297 );
nor U77840 ( n39297, n2108, n2105 );
nor U77841 ( n39296, n39298, n39299 );
nand U77842 ( n39298, n39302, n39303 );
nand U77843 ( n39299, n39300, n39301 );
nand U77844 ( n39300, n2038, n39127 );
nand U77845 ( n39301, n2043, n39127 );
nor U77846 ( n62764, n739, n62766 );
nor U77847 ( n62766, n62767, n62768 );
nand U77848 ( n62767, n62773, n62774 );
nand U77849 ( n62768, n62769, n62770 );
nand U77850 ( n39303, n2045, n39127 );
nor U77851 ( n62240, n61443, n45999 );
not U77852 ( n642, n41721 );
nand U77853 ( n39302, n2044, n39127 );
nand U77854 ( n41581, n62463, n62464 );
nand U77855 ( n62464, n750, n76386 );
nor U77856 ( n62463, n62465, n742 );
not U77857 ( n742, n62466 );
nand U77858 ( n62466, n743, n76385 );
nand U77859 ( n39227, n1872, n38861 );
xor U77860 ( n38212, n38905, n2118 );
and U77861 ( n39078, n38212, n2033 );
not U77862 ( n1159, n71716 );
nor U77863 ( n72002, n72003, n72004 );
nor U77864 ( n72003, n72005, n72006 );
and U77865 ( n72005, n72007, n1198 );
and U77866 ( n71762, n71858, n71859 );
nand U77867 ( n71859, n71716, n71720 );
nor U77868 ( n71858, n71712, n71718 );
not U77869 ( n670, n41550 );
nor U77870 ( n37530, n2132, n37533 );
nor U77871 ( n37533, n37534, n2129 );
nor U77872 ( n37534, n2120, n37536 );
nand U77873 ( n37536, n37460, n37537 );
nand U77874 ( n37121, n37305, n37306 );
nand U77875 ( n37306, n2032, n37307 );
nand U77876 ( n37305, n37308, n2038 );
nor U77877 ( n37570, n37575, n37576 );
nand U77878 ( n37576, n37577, n37578 );
nand U77879 ( n37575, n37467, n37580 );
nand U77880 ( n37578, n1943, n37443 );
and U77881 ( n37308, n37514, n37515 );
nor U77882 ( n37515, n37516, n37517 );
nor U77883 ( n37514, n37523, n37524 );
nand U77884 ( n37517, n37476, n37518 );
nand U77885 ( n37589, n37590, n37591 );
nor U77886 ( n37590, n37266, n37274 );
nand U77887 ( n37580, n37581, n37582 );
nor U77888 ( n37582, n1934, n1939 );
nor U77889 ( n37581, n37584, n37585 );
nor U77890 ( n37584, n1920, n37586 );
nand U77891 ( n37564, n37565, n37491 );
nand U77892 ( n37565, n37566, n1962 );
not U77893 ( n1962, n37488 );
nor U77894 ( n37566, n37570, n37571 );
nand U77895 ( n36563, n36568, n36569 );
nand U77896 ( n36568, n36570, n36571 );
nand U77897 ( n41528, n737, n76386 );
xor U77898 ( n71037, n71793, n71794 );
xor U77899 ( n71793, n71795, n71796 );
nand U77900 ( n40958, n40963, n40964 );
nand U77901 ( n40963, n40965, n40966 );
nor U77902 ( n37516, n2190, n37522 );
not U77903 ( n1200, n71874 );
not U77904 ( n1160, n71720 );
and U77905 ( n71759, n71863, n71864 );
nand U77906 ( n71864, n71865, n1200 );
nor U77907 ( n71863, n71866, n71867 );
nor U77908 ( n71866, n1199, n71873 );
xnor U77909 ( MUL_1411_U439, n71045, n71046 );
xnor U77910 ( n71046, n71047, n71048 );
nor U77911 ( n39313, n39317, n39318 );
nor U77912 ( n39318, n2002, n39292 );
nor U77913 ( n39317, n39323, n39294 );
and U77914 ( n39323, n39403, n39404 );
nand U77915 ( n39403, n2005, n39369 );
nand U77916 ( n39404, n2047, n39369 );
nand U77917 ( n65342, n65344, n65345 );
nand U77918 ( n65345, n65346, n65341 );
nor U77919 ( n65344, n65347, n65348 );
and U77920 ( n71848, n71855, n71852 );
and U77921 ( n40824, n76386, n41264 );
nand U77922 ( n41246, n41287, n41288 );
nand U77923 ( n41287, n40908, n40907 );
nand U77924 ( n41288, n608, n40905 );
not U77925 ( n1168, n72646 );
nor U77926 ( n62569, n61624, n62473 );
xor U77927 ( n38230, n39137, n2114 );
nand U77928 ( n71433, n71614, n71615 );
or U77929 ( n71614, n71619, n71618 );
nand U77930 ( n71615, n71616, n71617 );
nand U77931 ( n71617, n71618, n71619 );
and U77932 ( n71418, n71583, n71416 );
xnor U77933 ( n71432, n71460, n71600 );
xnor U77934 ( n71600, n71461, n71458 );
nor U77935 ( n62951, n62965, n41932 );
nor U77936 ( n62965, n62966, n62967 );
nand U77937 ( n62966, n62973, n62974 );
nand U77938 ( n62967, n62968, n534 );
nand U77939 ( n57589, n62935, n62936 );
nor U77940 ( n62936, n62937, n62938 );
nor U77941 ( n62935, n62948, n48337 );
and U77942 ( n62937, n48336, n76077 );
and U77943 ( n62783, n62957, n62958 );
nand U77944 ( n62957, n822, n62760 );
nand U77945 ( n62958, n61612, n62760 );
nor U77946 ( n62773, n62777, n62778 );
nor U77947 ( n62778, n820, n62684 );
nor U77948 ( n62777, n62783, n62686 );
or U77949 ( n62770, n62462, n62272 );
nand U77950 ( n48333, n48334, n48335 );
nand U77951 ( n48335, n568, n48336 );
nand U77952 ( n48334, n76857, n48337 );
and U77953 ( n39737, n39744, n39792 );
nand U77954 ( n39286, n39415, n39416 );
nand U77955 ( n39415, n1887, n2005 );
nand U77956 ( n39416, n1887, n2047 );
nor U77957 ( n39398, n2048, n39399 );
nor U77958 ( n39399, n39400, n39401 );
nand U77959 ( n39400, n39407, n39408 );
nand U77960 ( n39401, n39402, n39323 );
nand U77961 ( n38661, n39381, n39382 );
nor U77962 ( n39382, n39383, n39384 );
nor U77963 ( n39381, n39394, n38300 );
nand U77964 ( n39384, n39385, n39386 );
not U77965 ( n1169, n72592 );
nand U77966 ( n71160, n71167, n71168 );
nand U77967 ( n71157, n71164, n71165 );
nand U77968 ( n71165, n71162, n71166 );
nand U77969 ( n71166, n71160, n71163 );
nand U77970 ( n38284, n39351, n39352 );
nor U77971 ( n39351, n39371, n39372 );
nor U77972 ( n39352, n39353, n39354 );
nand U77973 ( n39371, n39375, n39376 );
nor U77974 ( n39366, n39370, n39347 );
nor U77975 ( n39370, n2049, n1887 );
nand U77976 ( n39353, n39363, n39364 );
nand U77977 ( n39363, n39365, n2005 );
nand U77978 ( n39364, n39365, n2047 );
nor U77979 ( n39365, n39366, n39367 );
nand U77980 ( n38296, n38297, n38298 );
nand U77981 ( n38298, n76819, n38299 );
nand U77982 ( n38297, n76812, n38300 );
nand U77983 ( n47602, n44985, n47683 );
nand U77984 ( n47480, n7610, n47533 );
nand U77985 ( n47297, n7584, n47333 );
not U77986 ( n7584, n47432 );
nand U77987 ( n47432, n7597, n47479 );
not U77988 ( n7597, n47480 );
nand U77989 ( n47281, n7573, n47288 );
not U77990 ( n7573, n47297 );
nor U77991 ( n47863, n7803, n7797 );
nand U77992 ( n47382, n47856, n7810 );
nand U77993 ( n47392, n47863, n7810 );
nand U77994 ( n47385, n47856, n7808 );
nand U77995 ( n47395, n47863, n7808 );
nand U77996 ( n62750, n835, n62462 );
nor U77997 ( n39411, n39412, n39413 );
nand U77998 ( n39412, n39423, n39424 );
nand U77999 ( n39413, n39414, n1882 );
nand U78000 ( n39424, n1869, n38861 );
nor U78001 ( n71598, n71432, n71435 );
or U78002 ( n71162, n71168, n71167 );
nor U78003 ( n62842, n62846, n62847 );
nor U78004 ( n62846, n728, n535 );
nand U78005 ( n62838, n62839, n62840 );
nand U78006 ( n62839, n825, n62848 );
nand U78007 ( n62840, n62841, n61613 );
nor U78008 ( n62841, n62842, n62843 );
nand U78009 ( n48210, n62835, n62836 );
nor U78010 ( n62835, n62859, n62860 );
nor U78011 ( n62836, n62837, n62838 );
nand U78012 ( n62859, n62863, n62864 );
nand U78013 ( n62752, n824, n62462 );
nand U78014 ( n71216, n71420, n71421 );
nand U78015 ( n71421, n71222, n1163 );
nor U78016 ( n71420, n71424, n71425 );
nor U78017 ( n71425, n71423, n71221 );
nor U78018 ( n71424, n71426, n71427 );
xor U78019 ( n71427, n71423, n71422 );
nand U78020 ( n71234, n71430, n71431 );
nand U78021 ( n71431, n71432, n71433 );
nor U78022 ( n71430, n71434, n1175 );
not U78023 ( n1175, n71435 );
nand U78024 ( n71857, n1132, n71852 );
nor U78025 ( n62423, n61443, n46938 );
not U78026 ( n1869, n39291 );
nor U78027 ( n39358, n39361, n39347 );
nor U78028 ( n39361, n2049, n1869 );
nand U78029 ( n39354, n39355, n39356 );
nand U78030 ( n39355, n2045, n39362 );
nand U78031 ( n39356, n39357, n38861 );
nor U78032 ( n39357, n39358, n39359 );
nor U78033 ( n71173, n71174, n71175 );
and U78034 ( n71174, n71178, n71179 );
nand U78035 ( n71175, n71176, n71177 );
not U78036 ( n1069, n71164 );
nand U78037 ( n47360, n47839, n7810 );
nor U78038 ( n72439, n1223, n1173 );
nand U78039 ( n47363, n47839, n7808 );
nand U78040 ( n39281, n38262, n38861 );
and U78041 ( n62571, n75728, n75729 );
nand U78042 ( n75728, n62473, n61613 );
nand U78043 ( n75729, n62473, n61612 );
not U78044 ( n1974, n37492 );
xor U78045 ( n39362, n37344, n39316 );
nand U78046 ( n26622, n24311, n26703 );
nand U78047 ( n59764, n57434, n59845 );
nand U78048 ( n68623, n65893, n68704 );
nand U78049 ( n68501, n5823, n68554 );
nand U78050 ( n68328, n5797, n68365 );
not U78051 ( n5797, n68453 );
nand U78052 ( n26500, n4054, n26553 );
nand U78053 ( n59639, n6687, n59695 );
nand U78054 ( n26327, n4033, n26364 );
not U78055 ( n4033, n26452 );
nand U78056 ( n59466, n6665, n59503 );
not U78057 ( n6665, n59591 );
nand U78058 ( n68453, n5809, n68500 );
not U78059 ( n5809, n68501 );
nand U78060 ( n26452, n4043, n26499 );
not U78061 ( n4043, n26500 );
nand U78062 ( n59591, n6675, n59638 );
not U78063 ( n6675, n59639 );
nand U78064 ( n68312, n5785, n68319 );
not U78065 ( n5785, n68328 );
nand U78066 ( n26311, n4024, n26318 );
not U78067 ( n4024, n26327 );
nand U78068 ( n59450, n6657, n59457 );
not U78069 ( n6657, n59466 );
nand U78070 ( n39376, n2044, n39362 );
nor U78071 ( n68883, n6015, n6009 );
nor U78072 ( n26884, n4238, n4232 );
nor U78073 ( n60024, n6870, n6864 );
nand U78074 ( n71758, n71875, n71876 );
nand U78075 ( n71876, n71751, n71756 );
nor U78076 ( n71875, n71747, n71753 );
not U78077 ( n1203, n71756 );
nand U78078 ( n68414, n68876, n6023 );
nand U78079 ( n26413, n26877, n4245 );
nand U78080 ( n59552, n60017, n6878 );
nand U78081 ( n68424, n68883, n6023 );
nand U78082 ( n26423, n26884, n4245 );
nand U78083 ( n59562, n60024, n6878 );
nand U78084 ( n68417, n68876, n6020 );
nand U78085 ( n26416, n26877, n4243 );
nand U78086 ( n59555, n60017, n6875 );
and U78087 ( n71891, n72010, n72011 );
nand U78088 ( n72011, n71869, n71874 );
nor U78089 ( n72010, n71865, n71871 );
nand U78090 ( n68427, n68883, n6020 );
nand U78091 ( n26426, n26884, n4243 );
nand U78092 ( n59565, n60024, n6875 );
nand U78093 ( n39375, n2043, n39362 );
not U78094 ( n1199, n71869 );
or U78095 ( n39556, n37491, n37500 );
nor U78096 ( n62852, n62855, n62856 );
nor U78097 ( n62855, n62760, n62847 );
nor U78098 ( n62856, n535, n62845 );
nand U78099 ( n71299, n71456, n71457 );
or U78100 ( n71456, n71461, n71460 );
nand U78101 ( n71457, n71458, n71459 );
nand U78102 ( n71459, n71460, n71461 );
nor U78103 ( n71439, n71438, n71441 );
xor U78104 ( n71441, n71299, n71298 );
nand U78105 ( n47370, n47846, n7810 );
nand U78106 ( n68392, n68859, n6023 );
nand U78107 ( n26391, n26860, n4245 );
nand U78108 ( n59530, n60000, n6878 );
nand U78109 ( n47373, n47846, n7808 );
nand U78110 ( n68395, n68859, n6020 );
nand U78111 ( n26394, n26860, n4243 );
nand U78112 ( n59533, n60000, n6875 );
nand U78113 ( n48075, n62761, n62762 );
and U78114 ( n62761, n739, n62763 );
nand U78115 ( n62762, n535, n62684 );
nand U78116 ( n62763, n62684, n62686 );
nand U78117 ( n71221, n71426, n71422 );
nand U78118 ( n72008, n72007, n72009 );
nor U78119 ( n39290, n39291, n2058 );
nor U78120 ( n36715, n36716, n36717 );
nand U78121 ( n36717, n36718, n36719 );
nand U78122 ( n36719, n1845, n1963 );
nand U78123 ( n36530, n36724, n36725 );
nand U78124 ( n36725, n36726, n36727 );
nor U78125 ( n39367, n39368, n39349 );
nor U78126 ( n39368, n2057, n39369 );
nand U78127 ( n41100, n40929, n41418 );
nor U78128 ( n41419, n41107, n41420 );
nor U78129 ( n41420, n41100, n41108 );
nor U78130 ( n39359, n39360, n39349 );
nor U78131 ( n39360, n2057, n39291 );
nand U78132 ( n39658, n37491, n39674 );
nor U78133 ( n39657, n39594, n38956 );
nor U78134 ( n39601, n37500, n39602 );
nor U78135 ( n39602, n39603, n39604 );
nor U78136 ( n39603, n2034, n37492 );
nand U78137 ( n38670, n39564, n39565 );
nor U78138 ( n39565, n39566, n39567 );
nor U78139 ( n39564, n39582, n38354 );
nand U78140 ( n39567, n39568, n39569 );
nand U78141 ( n39597, n39598, n39599 );
nand U78142 ( n39599, n1865, n38861 );
nor U78143 ( n39598, n39600, n39601 );
nor U78144 ( n39600, n39605, n39488 );
and U78145 ( n39414, n75730, n75731 );
nand U78146 ( n75730, n39378, n2043 );
nand U78147 ( n75731, n39378, n2038 );
nor U78148 ( n62843, n62844, n62845 );
nor U78149 ( n62844, n732, n62760 );
and U78150 ( n39423, n75732, n75733 );
nand U78151 ( n75732, n39378, n2045 );
nand U78152 ( n75733, n39378, n2044 );
nor U78153 ( n41289, n608, n40905 );
nand U78154 ( n62974, n535, n61613 );
not U78155 ( n1202, n71751 );
nor U78156 ( n71440, n71298, n71301 );
xor U78157 ( n38247, n39186, n2109 );
nand U78158 ( n40829, n76386, n76844 );
not U78159 ( n608, n40906 );
nand U78160 ( n68402, n68866, n6023 );
nand U78161 ( n26401, n26867, n4245 );
nand U78162 ( n59540, n60007, n6878 );
nor U78163 ( n37403, n37271, n37266 );
not U78164 ( n1162, n71423 );
nand U78165 ( n68405, n68866, n6020 );
nand U78166 ( n26404, n26867, n4243 );
nand U78167 ( n59543, n60007, n6875 );
nand U78168 ( n40928, n41108, n41109 );
or U78169 ( n41109, n41110, n41111 );
nor U78170 ( n41099, n41100, n41101 );
nand U78171 ( n41101, n41102, n41103 );
nand U78172 ( n41103, n519, n588 );
nor U78173 ( n62953, n62954, n62955 );
nand U78174 ( n62954, n62961, n62962 );
nand U78175 ( n62955, n62956, n62783 );
nand U78176 ( n62962, n61613, n62760 );
nor U78177 ( n62644, n62645, n41918 );
nor U78178 ( n62645, n62646, n62647 );
nor U78179 ( n62646, n61624, n62577 );
nand U78180 ( n62647, n62648, n62649 );
nand U78181 ( n62649, n537, n61613 );
nand U78182 ( n62648, n537, n61612 );
not U78183 ( n1920, n37592 );
xor U78184 ( n71070, n71777, n71778 );
xor U78185 ( n71777, n71779, n71780 );
nand U78186 ( n71035, n71698, n71699 );
nand U78187 ( n71698, n71070, n71073 );
nand U78188 ( n71699, n71072, n71700 );
or U78189 ( n71700, n71073, n71070 );
nand U78190 ( n36716, n37051, n36531 );
nor U78191 ( n37052, n36723, n37053 );
nor U78192 ( n37053, n36716, n36724 );
nand U78193 ( n39408, n38861, n39291 );
nand U78194 ( n64381, n64383, n64384 );
nand U78195 ( n64384, n64385, n64380 );
nor U78196 ( n64383, n64386, n64387 );
nor U78197 ( n39456, n1992, n39457 );
nor U78198 ( n39457, n39458, n39459 );
nand U78199 ( n39458, n39464, n39465 );
nand U78200 ( n39459, n39460, n39461 );
nand U78201 ( n38664, n39435, n39436 );
nor U78202 ( n39436, n39437, n39438 );
nor U78203 ( n39435, n39452, n38322 );
nand U78204 ( n39438, n39439, n39440 );
not U78205 ( n1124, n72649 );
nand U78206 ( n71505, n71765, n71766 );
nand U78207 ( n71766, n71767, n1122 );
nor U78208 ( n71765, n71768, n71769 );
nor U78209 ( n71768, n1120, n71775 );
nand U78210 ( n71073, n71701, n71702 );
or U78211 ( n71701, n71505, n71507 );
nand U78212 ( n71702, n71506, n71703 );
nand U78213 ( n71703, n71507, n71505 );
nand U78214 ( n48074, n62758, n62759 );
nor U78215 ( n62758, n739, n734 );
nand U78216 ( n62759, n727, n62760 );
and U78217 ( n39594, n37491, n39674 );
not U78218 ( n1163, n71422 );
and U78219 ( n39464, n75734, n75735 );
nand U78220 ( n75734, n39426, n38861 );
nand U78221 ( n75735, n39419, n2047 );
xor U78222 ( n62848, n41933, n62776 );
nand U78223 ( n62864, n824, n62848 );
nand U78224 ( n62863, n835, n62848 );
and U78225 ( n71300, n71438, n71298 );
nor U78226 ( n39473, n39475, n39476 );
and U78227 ( n39476, n39430, n2043 );
nor U78228 ( n39475, n38872, n39419 );
nor U78229 ( n39470, n39471, n39472 );
nand U78230 ( n39471, n39477, n39478 );
nand U78231 ( n39472, n39473, n39474 );
nor U78232 ( n39478, n39479, n39480 );
nor U78233 ( n62732, n61443, n62741 );
and U78234 ( n62968, n75736, n75737 );
nand U78235 ( n75736, n62866, n835 );
nand U78236 ( n75737, n62866, n837 );
not U78237 ( n7493, n46441 );
not U78238 ( n5707, n67505 );
not U78239 ( n3949, n25500 );
not U78240 ( n6582, n58637 );
or U78241 ( n71185, n71191, n71190 );
not U78242 ( n697, n41540 );
and U78243 ( n64032, n41540, n64226 );
nand U78244 ( n57728, n63980, n63981 );
nor U78245 ( n63981, n63982, n63983 );
nor U78246 ( n63980, n63993, n48685 );
and U78247 ( n63982, n48684, n76078 );
nand U78248 ( n63996, n64005, n64006 );
nand U78249 ( n64005, n64017, n41924 );
nand U78250 ( n64006, n702, n64007 );
nand U78251 ( n64017, n64018, n64019 );
nand U78252 ( n64007, n64008, n64009 );
nor U78253 ( n64008, n64015, n64016 );
nor U78254 ( n64009, n64010, n64011 );
nor U78255 ( n64015, n832, n63306 );
nor U78256 ( n62539, n61443, n47416 );
nand U78257 ( n71183, n71190, n71191 );
nor U78258 ( n64214, n64032, n62272 );
nor U78259 ( n64210, n64032, n61618 );
nand U78260 ( n64212, n41540, n64226 );
nor U78261 ( n62822, n61443, n48209 );
nand U78262 ( n48209, n62829, n62830 );
nand U78263 ( n62830, n733, n62831 );
nand U78264 ( n62829, n725, n62833 );
nand U78265 ( n62831, n62760, n62832 );
and U78266 ( n62973, n75738, n75739 );
nand U78267 ( n75738, n62866, n825 );
nand U78268 ( n75739, n62866, n824 );
nand U78269 ( n57634, n63255, n63256 );
nor U78270 ( n63256, n63257, n63258 );
nor U78271 ( n63255, n63270, n48458 );
nor U78272 ( n63257, n730, n76061 );
nor U78273 ( n63273, n63288, n41925 );
nor U78274 ( n63288, n63289, n63290 );
nand U78275 ( n63289, n63295, n63296 );
nand U78276 ( n63290, n63291, n63292 );
nor U78277 ( n63291, n63293, n63294 );
and U78278 ( n63294, n62979, n835 );
nor U78279 ( n63293, n61624, n62677 );
nor U78280 ( n63295, n63301, n63302 );
nor U78281 ( n63301, n833, n62677 );
nor U78282 ( n63302, n832, n62677 );
nand U78283 ( n48681, n48682, n48683 );
nand U78284 ( n48683, n568, n48684 );
nand U78285 ( n48682, n76857, n48685 );
nand U78286 ( n36524, n36529, n36530 );
nand U78287 ( n36529, n1963, n36531 );
and U78288 ( n39480, n39430, n2044 );
and U78289 ( n39479, n39430, n2045 );
not U78290 ( n1127, n72508 );
xor U78291 ( n71187, n71192, n71193 );
xor U78292 ( n71192, n71203, n71204 );
xor U78293 ( n71193, n71194, n71195 );
nor U78294 ( n71204, n1232, n1079 );
nor U78295 ( n71194, n71197, n71198 );
and U78296 ( n71197, n71201, n71202 );
nand U78297 ( n71198, n71199, n71200 );
nand U78298 ( n41529, n754, n76385 );
or U78299 ( n39461, n39430, n38956 );
nand U78300 ( n40922, n40927, n40928 );
nand U78301 ( n40927, n588, n40929 );
nor U78302 ( n63275, n63276, n63277 );
nand U78303 ( n63276, n63282, n63283 );
nand U78304 ( n63277, n63278, n63279 );
nor U78305 ( n63283, n63284, n63285 );
and U78306 ( n63282, n75740, n75741 );
nand U78307 ( n75740, n62677, n61613 );
nand U78308 ( n75741, n62677, n61612 );
nand U78309 ( n38276, n39343, n39344 );
nand U78310 ( n39344, n2055, n39345 );
nand U78311 ( n39343, n2050, n39348 );
not U78312 ( n2055, n39347 );
or U78313 ( n39348, n39291, n2057 );
nand U78314 ( n38338, n39526, n39527 );
nor U78315 ( n39526, n39545, n39546 );
nor U78316 ( n39527, n39528, n39529 );
nand U78317 ( n39545, n39549, n39550 );
nor U78318 ( n39541, n39544, n1978 );
nor U78319 ( n39544, n1979, n1880 );
not U78320 ( n1880, n39488 );
nand U78321 ( n38667, n39506, n39507 );
nor U78322 ( n39507, n39508, n39509 );
nor U78323 ( n39506, n39525, n38338 );
nand U78324 ( n39509, n39510, n39511 );
nand U78325 ( n39528, n39538, n39539 );
nand U78326 ( n39538, n39540, n2005 );
nand U78327 ( n39539, n39540, n2047 );
nor U78328 ( n39540, n39541, n39542 );
nand U78329 ( n39345, n39291, n39346 );
not U78330 ( n1865, n39490 );
nand U78331 ( n39529, n39530, n39531 );
nand U78332 ( n39530, n39537, n2045 );
nand U78333 ( n39531, n39532, n38861 );
nor U78334 ( n39532, n39533, n39534 );
nand U78335 ( n38334, n38335, n38336 );
nand U78336 ( n38336, n76820, n38337 );
nand U78337 ( n38335, n76812, n38338 );
nor U78338 ( n63284, n61618, n62979 );
and U78339 ( n71507, n71704, n71705 );
or U78340 ( n71704, n71066, n71069 );
nand U78341 ( n71705, n71068, n71706 );
nand U78342 ( n71706, n71069, n71066 );
nand U78343 ( n62686, n62832, n62779 );
nor U78344 ( n39591, n37500, n39594 );
nor U78345 ( n71596, n1173, n1227 );
nor U78346 ( n39542, n39543, n39524 );
nor U78347 ( n39543, n39495, n39488 );
nand U78348 ( n39616, n39617, n39618 );
nand U78349 ( n39617, n39620, n39590 );
nand U78350 ( n39618, n39619, n39590 );
nor U78351 ( n39620, n39591, n38956 );
xor U78352 ( n48328, n62760, n724 );
and U78353 ( n39646, n39604, n75742 );
or U78354 ( n75742, n1974, n37500 );
nand U78355 ( n38673, n39630, n39631 );
nor U78356 ( n39631, n39632, n39633 );
nor U78357 ( n39630, n39643, n38370 );
nor U78358 ( n39632, n2175, n38604 );
nand U78359 ( n38366, n38367, n38368 );
nand U78360 ( n38368, n76820, n38369 );
nand U78361 ( n38367, n76812, n38370 );
xor U78362 ( n38291, n39291, n2048 );
and U78363 ( n39383, n38291, n2033 );
and U78364 ( n62676, n62678, n727 );
and U78365 ( n62678, n62679, n62680 );
nor U78366 ( n39659, n1973, n39661 );
nor U78367 ( n39661, n39662, n39663 );
nand U78368 ( n39662, n39672, n39673 );
nand U78369 ( n39663, n39664, n39665 );
nor U78370 ( n39534, n39535, n39524 );
nor U78371 ( n39535, n39495, n39490 );
nand U78372 ( n41635, n76386, n76380 );
not U78373 ( n533, n63306 );
nor U78374 ( n63685, n63689, n63690 );
nor U78375 ( n63689, n63691, n63668 );
nor U78376 ( n63691, n704, n533 );
not U78377 ( n704, n63307 );
nand U78378 ( n57678, n63655, n63656 );
nor U78379 ( n63656, n63657, n63658 );
nor U78380 ( n63655, n63678, n48575 );
nor U78381 ( n63657, n720, n76060 );
nand U78382 ( n63682, n63683, n63684 );
nand U78383 ( n63683, n825, n63686 );
nand U78384 ( n63684, n63685, n61613 );
nand U78385 ( n48575, n63679, n63680 );
nor U78386 ( n63679, n63697, n63698 );
nor U78387 ( n63680, n63681, n63682 );
nand U78388 ( n63697, n63701, n63702 );
nand U78389 ( n63681, n63687, n63688 );
nand U78390 ( n63687, n63692, n822 );
nand U78391 ( n63688, n63685, n61612 );
nor U78392 ( n63692, n63693, n63690 );
and U78393 ( n63296, n75743, n75744 );
nand U78394 ( n75743, n62979, n825 );
nand U78395 ( n75744, n62979, n824 );
not U78396 ( n1125, n72468 );
not U78397 ( n76378, n76381 );
nor U78398 ( n63690, n63694, n63670 );
nor U78399 ( n63694, n709, n63306 );
or U78400 ( n63279, n62979, n62272 );
xor U78401 ( MUL_1411_U440, n71041, n71042 );
xor U78402 ( n71042, n71043, n71044 );
not U78403 ( n1129, n72162 );
not U78404 ( n76379, n76381 );
nor U78405 ( n71438, n1173, n1225 );
nand U78406 ( n41521, n759, n76385 );
nand U78407 ( n41632, n76386, n76010 );
nor U78408 ( n64011, n833, n63306 );
nand U78409 ( n37443, n37442, n37579 );
not U78410 ( n1965, n37573 );
nor U78411 ( n37467, n1958, n1965 );
not U78412 ( n1958, n37574 );
nor U78413 ( n64016, n61624, n63306 );
nor U78414 ( n71714, n71715, n71716 );
nor U78415 ( n71715, n71717, n71718 );
nor U78416 ( n71717, n71719, n71720 );
not U78417 ( n1128, n72225 );
nand U78418 ( n63292, n837, n62979 );
nand U78419 ( n57998, n64187, n64188 );
nor U78420 ( n64188, n64189, n64190 );
nor U78421 ( n64187, n64202, n48803 );
nor U78422 ( n64189, n707, n76063 );
nor U78423 ( n39593, n37500, n39594 );
and U78424 ( n39487, n39491, n39492 );
nand U78425 ( n39608, n37100, n39488 );
xor U78426 ( n71248, n71288, n71289 );
nor U78427 ( n71289, n71290, n71291 );
nand U78428 ( n71288, n71296, n71297 );
nor U78429 ( n71291, n71292, n71293 );
nor U78430 ( n71296, n71300, n1177 );
not U78431 ( n1177, n71301 );
nand U78432 ( n71223, n71225, n71226 );
nand U78433 ( n71226, n71227, n71228 );
nand U78434 ( n71225, n71235, n71236 );
nor U78435 ( n71227, n71231, n71232 );
xnor U78436 ( n71236, n71230, n71229 );
not U78437 ( n637, n42087 );
nor U78438 ( n41551, n41552, n41553 );
nor U78439 ( n41552, n668, n41554 );
nor U78440 ( n41554, n41555, n41556 );
nor U78441 ( n41555, n41570, n41571 );
nand U78442 ( n41505, n41512, n41513 );
nand U78443 ( n41512, n779, n76385 );
nand U78444 ( n41513, n41514, n41515 );
nor U78445 ( n41514, n41597, n770 );
nand U78446 ( n41523, n41524, n41525 );
nor U78447 ( n41524, n41580, n41581 );
nor U78448 ( n41525, n41526, n41527 );
nor U78449 ( n41580, n41582, n41530 );
nand U78450 ( n41561, n41563, n41564 );
nand U78451 ( n41564, n41565, n634 );
nor U78452 ( n41565, n653, n41567 );
not U78453 ( n634, n41566 );
nand U78454 ( n41545, n41547, n41548 );
nor U78455 ( n41548, n688, n683 );
nor U78456 ( n41547, n41549, n41550 );
nor U78457 ( n41549, n674, n41551 );
nor U78458 ( n64224, n64227, n64228 );
nor U78459 ( n64227, n532, n64229 );
nor U78460 ( n64228, n61618, n64212 );
nor U78461 ( n64229, n61613, n41469 );
nor U78462 ( n63693, n63696, n63668 );
and U78463 ( n63696, n63307, n63306 );
nor U78464 ( n64004, n699, n64032 );
nand U78465 ( n64027, n64028, n64029 );
nand U78466 ( n64028, n64031, n64001 );
nand U78467 ( n64029, n64030, n64001 );
nor U78468 ( n64031, n64004, n62272 );
nand U78469 ( n63997, n63998, n63999 );
nand U78470 ( n63999, n64000, n64001 );
nand U78471 ( n63998, n64003, n64001 );
nor U78472 ( n64000, n64002, n61618 );
nand U78473 ( n39550, n39537, n2044 );
nand U78474 ( n38386, n39704, n39705 );
nor U78475 ( n39705, n39706, n39707 );
nor U78476 ( n39704, n39719, n39720 );
nor U78477 ( n39707, n39708, n37373 );
nor U78478 ( n39719, n1968, n39721 );
nor U78479 ( n39721, n39722, n39723 );
nand U78480 ( n39722, n39728, n39729 );
nand U78481 ( n39723, n39724, n39725 );
nand U78482 ( n38676, n39686, n39687 );
nor U78483 ( n39687, n39688, n39689 );
nor U78484 ( n39686, n39703, n38386 );
nor U78485 ( n39688, n2174, n38604 );
nand U78486 ( n39673, n39594, n2044 );
nand U78487 ( n39549, n39537, n2043 );
nor U78488 ( n64002, n699, n64032 );
nand U78489 ( n33867, n31607, n33948 );
nand U78490 ( n33745, n3224, n33798 );
nand U78491 ( n33572, n3198, n33609 );
not U78492 ( n3198, n33697 );
nand U78493 ( n33697, n3210, n33744 );
not U78494 ( n3210, n33745 );
nand U78495 ( n33556, n3187, n33563 );
not U78496 ( n3187, n33572 );
nand U78497 ( n39607, n38861, n39490 );
nor U78498 ( n34129, n3400, n3394 );
nand U78499 ( n33658, n34122, n3408 );
nand U78500 ( n33668, n34129, n3408 );
nand U78501 ( n33661, n34122, n3405 );
nand U78502 ( n33671, n34129, n3405 );
nand U78503 ( n41854, n41865, n777 );
nor U78504 ( n41865, n41867, n41868 );
not U78505 ( n777, n41866 );
nor U78506 ( n41867, n41871, n41872 );
nand U78507 ( n41866, n41890, n41891 );
nor U78508 ( n41891, n41892, n41893 );
nor U78509 ( n41890, n41896, n41882 );
and U78510 ( n41892, n41886, n41885 );
xor U78511 ( n48453, n62677, n718 );
nand U78512 ( n63258, n63259, n63260 );
nand U78513 ( n63260, n48452, n76078 );
nand U78514 ( n63259, n48453, n827 );
xor U78515 ( n71228, n71229, n71230 );
xor U78516 ( n38314, n39426, n1992 );
and U78517 ( n39437, n38314, n2033 );
not U78518 ( n1130, n72035 );
nor U78519 ( n41896, n41899, n41900 );
or U78520 ( n71210, n71216, n71215 );
and U78521 ( n62249, n62288, n62289 );
and U78522 ( n62288, n62290, n62291 );
nand U78523 ( n33636, n34105, n3408 );
nand U78524 ( n33639, n34105, n3405 );
and U78525 ( n41893, n41888, n41887 );
nand U78526 ( n71208, n71215, n71216 );
nor U78527 ( n71235, n71304, n71233 );
nor U78528 ( n71304, n1170, n71232 );
not U78529 ( n1170, n71234 );
nand U78530 ( n71220, n71221, n1137 );
not U78531 ( n1137, n71222 );
nand U78532 ( n64223, n64032, n835 );
nor U78533 ( n41579, n42092, n41567 );
nand U78534 ( n64225, n64032, n824 );
and U78535 ( n71509, n71722, n71723 );
nand U78536 ( n71722, n71062, n71064 );
nand U78537 ( n71723, n71065, n71724 );
or U78538 ( n71724, n71064, n71062 );
nand U78539 ( n33646, n34112, n3408 );
nor U78540 ( n42031, n42032, n42026 );
nor U78541 ( n42032, n42033, n42034 );
nor U78542 ( n42033, n42050, n42051 );
nor U78543 ( n42034, n747, n42035 );
nor U78544 ( n42035, n42036, n42037 );
nand U78545 ( n42036, n42046, n42047 );
nand U78546 ( n42037, n42038, n740 );
nand U78547 ( n42047, n42048, n694 );
nand U78548 ( n41517, n764, n76385 );
nand U78549 ( n33649, n34112, n3405 );
not U78550 ( n532, n64024 );
nor U78551 ( n39647, n39648, n37374 );
nor U78552 ( n39648, n39649, n39650 );
nor U78553 ( n39650, n2039, n39614 );
nor U78554 ( n39649, n2002, n39611 );
nand U78555 ( n39665, n38861, n39614 );
nand U78556 ( n71512, n71745, n71746 );
nand U78557 ( n71746, n71747, n1203 );
nor U78558 ( n71745, n71748, n71749 );
nor U78559 ( n71748, n1202, n71755 );
nor U78560 ( n41617, n41842, n41843 );
nand U78561 ( n38310, n38311, n38312 );
nand U78562 ( n38312, n76447, n2892 );
nand U78563 ( n38311, n38314, n76442 );
nor U78564 ( n41845, n41846, n41847 );
nor U78565 ( n64362, n64364, n64365 );
and U78566 ( n64364, n64232, n61439 );
nor U78567 ( n64365, n61618, n63706 );
nor U78568 ( n64356, n693, n64357 );
nor U78569 ( n64357, n64358, n64359 );
nand U78570 ( n64359, n64360, n64361 );
nand U78571 ( n64358, n64362, n64363 );
nand U78572 ( n58227, n64335, n64336 );
nor U78573 ( n64336, n64337, n64338 );
nor U78574 ( n64335, n64352, n48920 );
nor U78575 ( n64337, n700, n76060 );
nand U78576 ( n38329, n39519, n39520 );
nand U78577 ( n39520, n39521, n39522 );
nand U78578 ( n39519, n1980, n39523 );
nand U78579 ( n39522, n39490, n39491 );
or U78580 ( n39523, n39490, n39495 );
nor U78581 ( n71231, n71233, n71234 );
and U78582 ( n39728, n75745, n75746 );
nand U78583 ( n75745, n37100, n39678 );
nand U78584 ( n75746, n39668, n38861 );
nand U78585 ( n64019, n822, n63306 );
nand U78586 ( n41570, n41575, n41576 );
nor U78587 ( n41576, n637, n657 );
and U78588 ( n41575, n41563, n41568 );
nor U78589 ( n41605, n41864, n41854 );
nor U78590 ( n41864, n41873, n41874 );
and U78591 ( n41874, n41872, n41871 );
nor U78592 ( n41873, n41860, n41861 );
nand U78593 ( n71297, n71298, n71299 );
and U78594 ( n62467, n42015, n42014 );
nand U78595 ( n40842, n41213, n41214 );
nand U78596 ( n41213, n41215, n41216 );
nand U78597 ( n41214, n40945, n40942 );
buf U78598 ( n76010, n76382 );
or U78599 ( n39725, n39554, n38956 );
nand U78600 ( n71721, n1133, n71720 );
xor U78601 ( n63686, n63300, n712 );
nor U78602 ( n37254, n2167, n76801 );
nand U78603 ( n63702, n824, n63686 );
nand U78604 ( n48445, n48450, n48451 );
nand U78605 ( n48451, n48452, n568 );
nand U78606 ( n48450, n48453, n45754 );
nand U78607 ( n63701, n835, n63686 );
not U78608 ( n553, n66441 );
nor U78609 ( n41868, n41869, n41870 );
and U78610 ( n48567, n63665, n63666 );
nand U78611 ( n63666, n708, n63667 );
nand U78612 ( n63665, n703, n63669 );
not U78613 ( n708, n63668 );
or U78614 ( n63669, n63306, n709 );
nor U78615 ( n41597, n76385, n775 );
nand U78616 ( n41980, n41993, n41994 );
nand U78617 ( n41993, n42012, n42013 );
nand U78618 ( n41994, n41995, n41996 );
nor U78619 ( n42013, n738, n41585 );
not U78620 ( n769, n42026 );
not U78621 ( n633, n41987 );
not U78622 ( n1207, n71258 );
xnor U78623 ( n41216, n593, n41222 );
nor U78624 ( n41222, n41223, n40824 );
nor U78625 ( n41223, n764, n40825 );
nand U78626 ( n63667, n63306, n63307 );
not U78627 ( n592, n40965 );
nand U78628 ( n39714, n39715, n39716 );
nand U78629 ( n39715, n2038, n39554 );
nand U78630 ( n39716, n2043, n39554 );
nand U78631 ( n39718, n2045, n39554 );
xnor U78632 ( n38346, n39490, n39581 );
nor U78633 ( n64513, n64385, n64379 );
nand U78634 ( n58435, n64488, n64489 );
nor U78635 ( n64489, n64490, n64491 );
nor U78636 ( n64488, n64501, n49035 );
and U78637 ( n64490, n49034, n76081 );
nor U78638 ( n64516, n64386, n64517 );
nor U78639 ( n64517, n64387, n530 );
and U78640 ( n49026, n64509, n64510 );
nand U78641 ( n64510, n64511, n64512 );
nand U78642 ( n64509, n64516, n64380 );
nor U78643 ( n64511, n64387, n64515 );
nand U78644 ( n39717, n2044, n39554 );
not U78645 ( n595, n40841 );
nor U78646 ( n64366, n64367, n64368 );
nand U78647 ( n64368, n64369, n64370 );
nand U78648 ( n64367, n64371, n64372 );
nand U78649 ( n64369, n837, n63706 );
nor U78650 ( n64371, n64373, n64374 );
nor U78651 ( n64373, n819, n64232 );
and U78652 ( n64374, n63706, n825 );
nand U78653 ( n49031, n49032, n49033 );
nand U78654 ( n49033, n568, n49034 );
nand U78655 ( n49032, n76857, n49035 );
nand U78656 ( n38679, n39759, n39760 );
nor U78657 ( n39760, n39761, n39762 );
nor U78658 ( n39759, n39774, n38401 );
nand U78659 ( n39762, n39763, n39764 );
nand U78660 ( n39777, n39782, n39783 );
nand U78661 ( n39782, n2045, n39781 );
nand U78662 ( n39783, n39784, n39785 );
nand U78663 ( n39785, n39786, n39787 );
nor U78664 ( n39784, n2002, n39789 );
nor U78665 ( n39789, n39790, n39791 );
and U78666 ( n39790, n39792, n39788 );
not U78667 ( n657, n41569 );
nand U78668 ( n38397, n38398, n38399 );
nand U78669 ( n38399, n76820, n38400 );
nand U78670 ( n38398, n76812, n38401 );
not U78671 ( n3105, n32740 );
xor U78672 ( n48676, n63306, n702 );
and U78673 ( n41522, n42102, n75747 );
or U78674 ( n75747, n750, n76385 );
nor U78675 ( n42027, n42063, n42026 );
nor U78676 ( n42063, n42069, n42070 );
nand U78677 ( n42069, n41521, n41517 );
nand U78678 ( n42070, n42071, n42072 );
nand U78679 ( n42071, n41985, n41566 );
or U78680 ( n64360, n63706, n62272 );
nand U78681 ( n38342, n38343, n38344 );
nand U78682 ( n38344, n76447, n2889 );
nand U78683 ( n38343, n1867, n76443 );
not U78684 ( n1867, n38346 );
nor U78685 ( n37246, n2168, n76801 );
not U78686 ( n1132, n71855 );
nor U78687 ( n41879, n41889, n41866 );
nor U78688 ( n41889, n41901, n41902 );
and U78689 ( n41901, n41870, n41869 );
and U78690 ( n41902, n41900, n41899 );
nor U78691 ( n40846, n40945, n40942 );
not U78692 ( n1864, n39803 );
nand U78693 ( n39794, n39795, n39796 );
nand U78694 ( n39796, n2038, n39781 );
nand U78695 ( n39795, n1863, n38861 );
nand U78696 ( n39773, n39799, n39800 );
nand U78697 ( n39799, n1960, n39802 );
nand U78698 ( n39800, n39786, n39801 );
not U78699 ( n1960, n39791 );
nor U78700 ( n41504, n76385, n779 );
buf U78701 ( n76011, n76382 );
not U78702 ( n76380, n76381 );
not U78703 ( n1984, n36570 );
nor U78704 ( n40847, n41215, n41216 );
nand U78705 ( n41855, n41856, n41857 );
nand U78706 ( n41856, n41860, n41861 );
or U78707 ( n41857, n41841, n41840 );
nand U78708 ( n64370, n835, n63706 );
not U78709 ( n2058, n39292 );
nor U78710 ( n42012, n42017, n42018 );
nand U78711 ( n42018, n769, n42019 );
nand U78712 ( n42019, n42020, n42021 );
nand U78713 ( n42021, n719, n41586 );
nand U78714 ( n64372, n824, n63706 );
nand U78715 ( n42072, n42073, n42074 );
nor U78716 ( n42074, n42075, n42076 );
nand U78717 ( n42076, n41543, n42077 );
nor U78718 ( n42075, n42078, n41553 );
xor U78719 ( n38364, n39614, n1973 );
nand U78720 ( n39633, n39634, n39635 );
nand U78721 ( n39634, n76797, n38369 );
nand U78722 ( n39635, n2033, n38364 );
nand U78723 ( n39802, n39803, n39792 );
not U78724 ( n1892, n38833 );
not U78725 ( n610, n41019 );
not U78726 ( n2112, n37542 );
nor U78727 ( n41881, n41883, n41884 );
nor U78728 ( n41883, n41887, n41888 );
nor U78729 ( n41884, n41885, n41886 );
nand U78730 ( n38682, n39815, n39816 );
nor U78731 ( n39816, n39817, n39818 );
nor U78732 ( n39815, n39830, n38417 );
nand U78733 ( n39818, n39819, n39820 );
nor U78734 ( n38106, n38109, n38110 );
not U78735 ( n2052, n39294 );
nor U78736 ( n39833, n2002, n39837 );
xor U78737 ( n39837, n39829, n39788 );
nand U78738 ( n58782, n64776, n64777 );
nor U78739 ( n64777, n64778, n64779 );
nor U78740 ( n64776, n64792, n49145 );
nor U78741 ( n64778, n689, n76059 );
xor U78742 ( n39781, n37356, n39731 );
nand U78743 ( n39778, n39779, n39780 );
nand U78744 ( n39779, n2043, n39781 );
nand U78745 ( n39780, n2044, n39781 );
xor U78746 ( n45442, n45443, n45444 );
and U78747 ( n71515, n71728, n71729 );
nand U78748 ( n71728, n71058, n71061 );
nand U78749 ( n71729, n71060, n71730 );
or U78750 ( n71730, n71061, n71058 );
not U78751 ( n734, n62684 );
nor U78752 ( n64205, n64024, n64215 );
nand U78753 ( n64215, n698, n64216 );
nand U78754 ( n41920, n62253, n62290 );
nand U78755 ( n41599, n41909, n41910 );
nor U78756 ( n41909, n41940, n41941 );
nor U78757 ( n41910, n41911, n41912 );
nand U78758 ( n41940, n41953, n41954 );
nand U78759 ( n41912, n41913, n41914 );
nor U78760 ( n41913, n41921, n41922 );
nor U78761 ( n41914, n41915, n41916 );
nand U78762 ( n41922, n41923, n41924 );
nor U78763 ( n37242, n2169, n76801 );
nand U78764 ( n41936, n62325, n62289 );
nand U78765 ( n41911, n41927, n41928 );
nor U78766 ( n41928, n41929, n41930 );
nor U78767 ( n41927, n41934, n41935 );
nand U78768 ( n41930, n41931, n41932 );
nand U78769 ( n41926, n61590, n61587 );
nand U78770 ( n41921, n41925, n41926 );
not U78771 ( n1133, n71719 );
nor U78772 ( n64797, n64798, n64799 );
nor U78773 ( n64798, n64800, n64525 );
nor U78774 ( n64799, n819, n64513 );
nand U78775 ( n37454, n37554, n37593 );
nand U78776 ( n41937, n62331, n62291 );
xor U78777 ( n48798, n64024, n698 );
nand U78778 ( n64190, n64191, n64192 );
nand U78779 ( n64192, n48797, n76075 );
nand U78780 ( n64191, n48798, n827 );
nor U78781 ( n40817, n600, n40707 );
not U78782 ( n600, n40832 );
nand U78783 ( n41918, n62578, n62575 );
nand U78784 ( n41933, n62779, n62782 );
nand U78785 ( n41917, n62679, n62681 );
nor U78786 ( n62851, n61624, n62853 );
nand U78787 ( n62853, n62857, n62858 );
nand U78788 ( n62857, n732, n725 );
nand U78789 ( n62858, n728, n733 );
not U78790 ( n733, n62847 );
not U78791 ( n2105, n37546 );
not U78792 ( n1985, n37498 );
xor U78793 ( n40901, n40907, n40908 );
nand U78794 ( n41919, n62474, n62471 );
nor U78795 ( n65823, n65346, n65340 );
nand U78796 ( n49381, n65810, n65811 );
nor U78797 ( n65811, n65812, n65813 );
nor U78798 ( n65810, n65817, n65818 );
nor U78799 ( n65812, n65354, n65815 );
nand U78800 ( n65801, n65819, n65820 );
nand U78801 ( n65820, n65821, n65822 );
nand U78802 ( n65819, n65825, n65341 );
nor U78803 ( n65821, n41939, n65348 );
nand U78804 ( n59661, n65795, n65796 );
nor U78805 ( n65796, n65797, n65798 );
nor U78806 ( n65795, n65809, n49381 );
and U78807 ( n65797, n49380, n76080 );
nor U78808 ( n65825, n65347, n65826 );
nor U78809 ( n65826, n65348, n529 );
not U78810 ( n668, n42082 );
nor U78811 ( n40819, n612, n40832 );
not U78812 ( n612, n40707 );
nand U78813 ( n38685, n39860, n39861 );
nor U78814 ( n39861, n39862, n39863 );
nor U78815 ( n39860, n39874, n38433 );
nor U78816 ( n39862, n2170, n38604 );
nand U78817 ( n39878, n39879, n39880 );
nand U78818 ( n39880, n39881, n39742 );
nand U78819 ( n39879, n1952, n39882 );
nor U78820 ( n39881, n2002, n1952 );
nand U78821 ( n38692, n39916, n39917 );
nor U78822 ( n39917, n39918, n39919 );
nor U78823 ( n39916, n39932, n38449 );
nand U78824 ( n39919, n39920, n39921 );
nand U78825 ( n39930, n39944, n39898 );
nor U78826 ( n39944, n1949, n39945 );
nor U78827 ( n39945, n1942, n39942 );
nand U78828 ( n49377, n49378, n49379 );
nand U78829 ( n49379, n568, n49380 );
nand U78830 ( n49378, n76857, n49381 );
xor U78831 ( n64518, n687, n64376 );
nand U78832 ( n64521, n64522, n64523 );
nand U78833 ( n64522, n837, n64518 );
nand U78834 ( n64523, n835, n64518 );
nand U78835 ( n65336, n65354, n61410 );
and U78836 ( n65334, n75748, n65336 );
or U78837 ( n75748, n823, n42077 );
nor U78838 ( n65330, n65331, n41931 );
nor U78839 ( n65331, n65332, n65333 );
nor U78840 ( n65333, n819, n64804 );
nor U78841 ( n65332, n669, n65334 );
nand U78842 ( n59154, n65309, n65310 );
nor U78843 ( n65310, n65311, n65312 );
nor U78844 ( n65309, n65326, n49268 );
nor U78845 ( n65311, n684, n76065 );
xor U78846 ( MUL_1411_U441, n71037, n71038 );
xor U78847 ( n71038, n71039, n71040 );
not U78848 ( n1890, n39031 );
nor U78849 ( n62315, n61624, n62317 );
or U78850 ( n62317, n75749, n75750 );
nor U78851 ( n75749, n62325, n763 );
nor U78852 ( n75750, n41517, n759 );
nand U78853 ( n62845, n727, n62782 );
xnor U78854 ( n38409, n39829, n1864 );
not U78855 ( n1095, n72411 );
nor U78856 ( n37234, n2170, n76801 );
nor U78857 ( n36274, n36275, n36276 );
nand U78858 ( n36275, n36280, n36281 );
nand U78859 ( n36276, n36277, n36278 );
nand U78860 ( n36278, n1847, n36279 );
not U78861 ( n1847, n36813 );
xor U78862 ( n49137, n530, n64784 );
nand U78863 ( n64779, n64780, n64781 );
nand U78864 ( n64781, n49140, n76079 );
nand U78865 ( n64780, n49137, n827 );
and U78866 ( n40827, n75751, n40829 );
or U78867 ( n75751, n775, n40830 );
not U78868 ( n1097, n72490 );
nor U78869 ( n72376, n1100, n1234 );
nand U78870 ( n48790, n48795, n48796 );
nand U78871 ( n48796, n48797, n568 );
nand U78872 ( n48795, n48798, n45754 );
xnor U78873 ( n38427, n37337, n39739 );
and U78874 ( n39877, n38861, n38427 );
nand U78875 ( n38405, n38406, n38407 );
nand U78876 ( n38407, n76447, n2915 );
nand U78877 ( n38406, n1862, n76443 );
not U78878 ( n1862, n38409 );
nand U78879 ( n39931, n39940, n39941 );
nor U78880 ( n39940, n1945, n1942 );
nand U78881 ( n39941, n39942, n39943 );
nand U78882 ( n39886, n39908, n38792 );
nand U78883 ( n42051, n42093, n42002 );
nor U78884 ( n42093, n685, n42006 );
xor U78885 ( n48915, n64232, n693 );
nor U78886 ( n40678, n40679, n40680 );
nand U78887 ( n40679, n40684, n40685 );
nand U78888 ( n40680, n40681, n40682 );
nand U78889 ( n40682, n520, n40683 );
not U78890 ( n520, n41194 );
nor U78891 ( n65936, n65942, n665 );
nor U78892 ( n65942, n65943, n65944 );
and U78893 ( n65943, n61410, n64809 );
nor U78894 ( n65944, n819, n529 );
nand U78895 ( n60122, n65918, n65919 );
nor U78896 ( n65919, n65920, n65921 );
nor U78897 ( n65918, n65933, n49577 );
nand U78898 ( n65921, n65922, n65923 );
nand U78899 ( n62321, n62252, n62291 );
not U78900 ( n760, n62289 );
not U78901 ( n555, n64525 );
nand U78902 ( n14293, n11304, n14412 );
nand U78903 ( n14140, n4957, n14207 );
nand U78904 ( n13927, n4930, n13964 );
not U78905 ( n4930, n14080 );
nand U78906 ( n14080, n4943, n14139 );
not U78907 ( n4943, n14140 );
nand U78908 ( n13907, n4921, n13915 );
not U78909 ( n4921, n13927 );
nand U78910 ( n12218, n4914, n12660 );
nand U78911 ( n14037, n14619, n5153 );
nand U78912 ( n14033, n14619, n5155 );
not U78913 ( n7595, n47533 );
nor U78914 ( n14628, n5148, n5142 );
nand U78915 ( n36502, n36895, n36510 );
xor U78916 ( n11662, n11663, n11664 );
nor U78917 ( n36896, n36701, n36898 );
nor U78918 ( n36898, n36502, n36698 );
nand U78919 ( n14049, n14628, n5153 );
nand U78920 ( n14045, n14628, n5155 );
xnor U78921 ( n38459, n39942, n37355 );
nand U78922 ( n38465, n39974, n39975 );
nor U78923 ( n39975, n39976, n39977 );
nor U78924 ( n39974, n39983, n39984 );
nor U78925 ( n39977, n39848, n39978 );
nand U78926 ( n38695, n39959, n39960 );
nor U78927 ( n39960, n39961, n39962 );
nor U78928 ( n39959, n39973, n38465 );
nor U78929 ( n39961, n2168, n38604 );
nor U78930 ( n65939, n65940, n65941 );
nor U78931 ( n65940, n823, n64809 );
nor U78932 ( n65941, n819, n65823 );
nand U78933 ( n41585, n42014, n42015 );
nand U78934 ( n41530, n41583, n41584 );
nor U78935 ( n41583, n738, n41587 );
nor U78936 ( n41584, n735, n41585 );
nor U78937 ( n41587, n729, n41588 );
xor U78938 ( n47690, n44985, n47683 );
not U78939 ( n5808, n68554 );
not U78940 ( n6674, n59695 );
not U78941 ( n4042, n26553 );
not U78942 ( n715, n41809 );
nand U78943 ( n49133, n49134, n49135 );
nand U78944 ( n49135, n76335, n1798 );
nand U78945 ( n49134, n49137, n45754 );
nand U78946 ( n38437, n38438, n38439 );
nand U78947 ( n38439, n76446, n2913 );
nand U78948 ( n38438, n1860, n76443 );
not U78949 ( n1860, n38441 );
xor U78950 ( n68711, n65893, n68704 );
xor U78951 ( n26710, n24311, n26703 );
xor U78952 ( n59852, n57434, n59845 );
not U78953 ( n738, n42016 );
not U78954 ( n2100, n37557 );
not U78955 ( n2020, n36897 );
nand U78956 ( n14009, n14598, n5153 );
nand U78957 ( n14005, n14598, n5155 );
nor U78958 ( n37230, n2172, n76801 );
nand U78959 ( n14022, n14607, n5153 );
xor U78960 ( n45432, n45433, n45434 );
and U78961 ( n62252, n62325, n62331 );
nand U78962 ( n14018, n14607, n5155 );
nand U78963 ( n36810, n36816, n36813 );
nand U78964 ( n36816, n36279, n36281 );
nor U78965 ( n48080, n549, n76385 );
nor U78966 ( n39946, n39948, n39886 );
nor U78967 ( n39948, n1944, n1948 );
nor U78968 ( n65329, n819, n65337 );
nand U78969 ( n65337, n64804, n41931 );
nand U78970 ( n41541, n41543, n41544 );
nand U78971 ( n62824, n48204, n76079 );
nor U78972 ( n65920, n61443, n49569 );
not U78973 ( n1102, n72210 );
nand U78974 ( n38485, n40008, n40009 );
nor U78975 ( n40009, n40010, n40011 );
nor U78976 ( n40008, n40019, n40020 );
nor U78977 ( n40011, n39982, n40012 );
nand U78978 ( n38698, n39993, n39994 );
nor U78979 ( n39994, n39995, n39996 );
nor U78980 ( n39993, n40007, n38485 );
nor U78981 ( n39995, n2167, n38604 );
and U78982 ( n40019, n38819, n38479 );
nand U78983 ( n41191, n41197, n41194 );
nand U78984 ( n41197, n40683, n40685 );
nor U78985 ( n39936, n39908, n39937 );
nand U78986 ( n39937, n38792, n39938 );
nor U78987 ( n65813, n65814, n65336 );
nor U78988 ( n65814, n674, n669 );
and U78989 ( n61599, n76080, n48080 );
nor U78990 ( n37222, n2173, n76802 );
nand U78991 ( n39331, n38279, n76797 );
not U78992 ( n747, n42015 );
xor U78993 ( MUL_1411_U7, n71033, n71034 );
xor U78994 ( n71033, n71035, n71036 );
xnor U78995 ( n49263, n64804, n41931 );
not U78996 ( n770, n42067 );
nor U78997 ( n71569, n1232, n1100 );
nand U78998 ( n39996, n39997, n39998 );
nand U78999 ( n39997, n76798, n38480 );
nand U79000 ( n39998, n2033, n38479 );
nor U79001 ( n41589, n42098, n719 );
and U79002 ( n40057, n40052, n75752 );
and U79003 ( n75752, n40053, n38819 );
nand U79004 ( n38701, n40039, n40040 );
nor U79005 ( n40040, n40041, n40042 );
nor U79006 ( n40039, n40054, n38501 );
nand U79007 ( n40042, n40043, n40044 );
not U79008 ( n7583, n47479 );
nor U79009 ( n41518, n762, n765 );
not U79010 ( n762, n42100 );
not U79011 ( n765, n62273 );
nor U79012 ( n41588, n722, n41589 );
not U79013 ( n722, n41590 );
nand U79014 ( n38497, n38498, n38499 );
nand U79015 ( n38499, n76819, n38500 );
nand U79016 ( n38498, n76812, n38501 );
nand U79017 ( n48198, n48203, n45752 );
nand U79018 ( n48203, n48204, n568 );
nand U79019 ( n39386, n76798, n38299 );
nand U79020 ( n37382, n37434, n37462 );
nor U79021 ( n37462, n37403, n37408 );
nor U79022 ( n37468, n37489, n37490 );
nand U79023 ( n37489, n37491, n37492 );
nand U79024 ( n37427, n37428, n37429 );
nor U79025 ( n37429, n37430, n37431 );
nor U79026 ( n37428, n37458, n37459 );
nor U79027 ( n37430, n37447, n37448 );
nand U79028 ( n42024, n41590, n41586 );
nand U79029 ( n60232, n65996, n65997 );
nor U79030 ( n65997, n65998, n65999 );
nor U79031 ( n65996, n66013, n54623 );
nor U79032 ( n65998, n667, n76064 );
and U79033 ( n66017, n61439, n54618 );
not U79034 ( n5795, n68500 );
not U79035 ( n6664, n59638 );
not U79036 ( n4032, n26499 );
not U79037 ( n3147, n33026 );
nand U79038 ( n38278, n38279, n76818 );
xor U79039 ( n11649, n11650, n11652 );
nor U79040 ( n61586, n774, n61429 );
not U79041 ( n774, n61412 );
nor U79042 ( n37218, n2174, n76802 );
xor U79043 ( n38509, n40028, n37368 );
nand U79044 ( n38704, n40081, n40082 );
nor U79045 ( n40082, n40083, n40084 );
nor U79046 ( n40081, n40098, n38517 );
nand U79047 ( n40084, n40085, n40086 );
not U79048 ( n2120, n37596 );
nand U79049 ( n37455, n37406, n37508 );
nand U79050 ( n37508, n37402, n37502 );
nand U79051 ( n42059, n42089, n42090 );
nor U79052 ( n42090, n674, n657 );
nor U79053 ( n42089, n678, n42083 );
not U79054 ( n678, n41543 );
nand U79055 ( n42055, n645, n42056 );
nor U79056 ( n71407, n1230, n1100 );
or U79057 ( n37311, n37103, n37307 );
nand U79058 ( n39511, n76797, n38337 );
nand U79059 ( n38492, n40052, n40053 );
nand U79060 ( n38472, n38477, n38478 );
nand U79061 ( n38477, n76819, n38480 );
nand U79062 ( n38478, n38479, n76443 );
nand U79063 ( n54638, n66100, n66101 );
nor U79064 ( n66101, n66102, n66103 );
nor U79065 ( n66100, n66110, n66111 );
nor U79066 ( n66103, n66104, n66029 );
nor U79067 ( n66110, n819, n66091 );
nand U79068 ( n60344, n66085, n66086 );
nor U79069 ( n66086, n66087, n66088 );
nor U79070 ( n66085, n66099, n54638 );
and U79071 ( n66087, n54637, n76079 );
nand U79072 ( n37444, n37446, n37266 );
nor U79073 ( n37446, n1932, n37443 );
nand U79074 ( n54634, n54635, n54636 );
nand U79075 ( n54636, n568, n54637 );
nand U79076 ( n54635, n76857, n54638 );
not U79077 ( n2115, n37594 );
not U79078 ( n1932, n37263 );
and U79079 ( n38900, n38945, n38946 );
nand U79080 ( n38946, n38903, n38947 );
nand U79081 ( n38947, n38948, n38949 );
not U79082 ( n649, n42056 );
nor U79083 ( n40118, n1927, n40120 );
not U79084 ( n692, n41546 );
nor U79085 ( n37210, n2175, n76802 );
nand U79086 ( n37448, n2110, n37449 );
nand U79087 ( n37449, n37450, n37451 );
not U79088 ( n2110, n37455 );
nand U79089 ( n37451, n37452, n1983 );
nand U79090 ( n45752, n569, n76385 );
nand U79091 ( n37378, n37379, n37380 );
nand U79092 ( n37379, n37385, n37386 );
nand U79093 ( n37380, n37381, n1924 );
nand U79094 ( n37386, n37387, n37388 );
nand U79095 ( n40122, n40120, n37271 );
nand U79096 ( n66029, n66035, n61410 );
not U79097 ( n527, n66091 );
nand U79098 ( n42083, n41560, n42082 );
not U79099 ( n7572, n47333 );
nor U79100 ( n41996, n41997, n41998 );
nand U79101 ( n41998, n41999, n42000 );
nand U79102 ( n41997, n42002, n644 );
nor U79103 ( n41999, n629, n685 );
nand U79104 ( n49640, n7439, n283 );
nand U79105 ( n37405, n37406, n1957 );
not U79106 ( n1957, n37407 );
nand U79107 ( n37392, n37393, n37394 );
nor U79108 ( n37394, n37395, n37396 );
nor U79109 ( n37393, n37404, n37405 );
nand U79110 ( n37396, n37397, n37398 );
nor U79111 ( n40148, n2034, n40158 );
nor U79112 ( n40158, n40159, n40160 );
nor U79113 ( n40159, n40120, n40161 );
nor U79114 ( n40160, n37369, n1894 );
nand U79115 ( n38707, n40132, n40133 );
nor U79116 ( n40133, n40134, n40135 );
nor U79117 ( n40132, n40145, n38533 );
nand U79118 ( n40135, n40136, n40137 );
not U79119 ( n1894, n40120 );
nand U79120 ( n41950, n712, n41952 );
nand U79121 ( n40703, n76386, n578 );
nand U79122 ( n37423, n37473, n37474 );
nand U79123 ( n37474, n37475, n37476 );
nand U79124 ( n37473, n37415, n37481 );
nand U79125 ( n37475, n37477, n37478 );
nand U79126 ( n37481, n37482, n37483 );
and U79127 ( n37482, n37502, n37503 );
nor U79128 ( n37483, n37484, n37485 );
nor U79129 ( n37484, n37493, n37490 );
nand U79130 ( n38529, n38530, n38531 );
nand U79131 ( n38531, n76819, n38532 );
nand U79132 ( n38530, n76812, n38533 );
not U79133 ( n735, n41586 );
not U79134 ( n5784, n68365 );
not U79135 ( n6655, n59503 );
not U79136 ( n4023, n26364 );
nor U79137 ( n66031, n66033, n66034 );
nand U79138 ( n66033, n41569, n41949 );
nand U79139 ( n66034, n65949, n61410 );
nor U79140 ( n40065, n40067, n40017 );
nor U79141 ( n40067, n1934, n1932 );
not U79142 ( n3209, n33798 );
not U79143 ( n827, n61443 );
not U79144 ( n570, n45363 );
xor U79145 ( n33955, n31607, n33948 );
or U79146 ( n75753, n41477, n45363 );
nand U79147 ( n49372, n76335, n1795 );
nand U79148 ( n54642, n54643, n54644 );
nand U79149 ( n54643, n54646, n45754 );
nand U79150 ( n54644, n76335, n1802 );
nand U79151 ( n48909, n76335, n1800 );
nand U79152 ( n48447, n76335, n1775 );
nand U79153 ( n54615, n54618, n45754 );
nand U79154 ( n48677, n76335, n1773 );
nor U79155 ( n71224, n1229, n1100 );
xor U79156 ( n49644, n49646, n49647 );
not U79157 ( n2132, n37433 );
or U79158 ( n37404, n37408, n37383 );
and U79159 ( n66286, n66281, n75754 );
and U79160 ( n75754, n66282, n61439 );
nand U79161 ( n66282, n66290, n647 );
nor U79162 ( n66290, n640, n66292 );
nor U79163 ( n66292, n638, n66293 );
nand U79164 ( n60564, n66268, n66269 );
nor U79165 ( n66269, n66270, n66271 );
nor U79166 ( n66268, n66283, n54678 );
nand U79167 ( n66271, n66272, n66273 );
nor U79168 ( n66293, n66208, n66362 );
and U79169 ( n66362, n66363, n66206 );
nand U79170 ( n54674, n54675, n54676 );
nand U79171 ( n54676, n568, n54677 );
nand U79172 ( n54675, n76857, n54678 );
not U79173 ( n7563, n47288 );
nand U79174 ( n39764, n76797, n38400 );
not U79175 ( n1072, n72395 );
nand U79176 ( n38524, n40150, n40151 );
nand U79177 ( n40151, n40152, n40153 );
nand U79178 ( n40150, n40155, n40156 );
nor U79179 ( n40152, n40107, n37369 );
not U79180 ( n2137, n37389 );
not U79181 ( n5775, n68319 );
not U79182 ( n6649, n59457 );
not U79183 ( n4017, n26318 );
nor U79184 ( n41507, n42061, n42062 );
not U79185 ( n1944, n37466 );
nand U79186 ( n60461, n66171, n66172 );
nor U79187 ( n66172, n66173, n66174 );
nor U79188 ( n66171, n66188, n54654 );
nor U79189 ( n66173, n654, n76063 );
and U79190 ( n66192, n61439, n54646 );
nand U79191 ( n54915, n76858, n41311 );
nor U79192 ( n36371, n1915, n36372 );
not U79193 ( n1915, n36376 );
nand U79194 ( n36372, n36373, n36374 );
nand U79195 ( n36373, n1848, n36375 );
not U79196 ( n1848, n36778 );
nand U79197 ( n42054, n669, n41543 );
not U79198 ( n1073, n72284 );
nor U79199 ( n36370, n36376, n36377 );
nand U79200 ( n36377, n36378, n36375 );
nand U79201 ( n60669, n66341, n66342 );
nor U79202 ( n66342, n66343, n66344 );
nor U79203 ( n66341, n66357, n54762 );
nand U79204 ( n66344, n66345, n66346 );
nor U79205 ( n37206, n2177, n76802 );
and U79206 ( n33176, n76022, n33160 );
nor U79207 ( n72051, n1238, n1079 );
nor U79208 ( n37415, n37455, n37413 );
nor U79209 ( n40774, n594, n40775 );
not U79210 ( n594, n40779 );
nand U79211 ( n40775, n40776, n40777 );
nand U79212 ( n40776, n522, n40778 );
not U79213 ( n522, n41161 );
not U79214 ( n778, n41952 );
nand U79215 ( n61440, n61445, n61446 );
nand U79216 ( n61446, n61429, n41952 );
nand U79217 ( n61445, n774, n778 );
nand U79218 ( n39820, n76797, n38412 );
nor U79219 ( n40773, n40779, n40780 );
nand U79220 ( n40780, n40781, n40778 );
nand U79221 ( n38505, n38506, n38507 );
nand U79222 ( n38507, n76446, n2919 );
nand U79223 ( n38506, n38509, n76444 );
nand U79224 ( n49571, n49572, n568 );
nand U79225 ( n49139, n49140, n568 );
nand U79226 ( n40153, n40154, n40113 );
not U79227 ( n4942, n14207 );
nor U79228 ( n66270, n61443, n54669 );
nand U79229 ( n54669, n66281, n66282 );
xor U79230 ( MUL_1411_U385, n71070, n71071 );
xor U79231 ( n71071, n71072, n71073 );
nand U79232 ( n54919, n54920, n54921 );
nand U79233 ( n54920, n76857, n54924 );
nand U79234 ( n54921, n568, n54922 );
nand U79235 ( n54817, n54818, n54819 );
nand U79236 ( n54818, n76857, n54821 );
nand U79237 ( n54819, n568, n54820 );
nand U79238 ( n66213, n66219, n61410 );
xor U79239 ( n14392, n11304, n14412 );
nor U79240 ( n71558, n1223, n1079 );
not U79241 ( n685, n41544 );
or U79242 ( n61451, n41952, n61429 );
nor U79243 ( n37198, n2178, n76802 );
nand U79244 ( n16667, n4795, n31 );
nand U79245 ( n36438, n2017, n36840 );
not U79246 ( n2017, n36549 );
nand U79247 ( n36437, n36438, n36439 );
nor U79248 ( n66215, n66217, n66218 );
nand U79249 ( n66217, n41958, n42092 );
nand U79250 ( n66218, n66109, n61410 );
xor U79251 ( n38540, n40154, n37336 );
nand U79252 ( n38710, n40170, n40171 );
nor U79253 ( n40171, n40172, n40173 );
nor U79254 ( n40170, n40186, n38548 );
nor U79255 ( n40172, n2162, n38604 );
nand U79256 ( n36436, n2014, n36549 );
nor U79257 ( n41953, n41960, n41961 );
nand U79258 ( n41960, n41962, n41963 );
nand U79259 ( n41961, n687, n523 );
nor U79260 ( n39581, n39495, n1979 );
not U79261 ( n1979, n39491 );
nand U79262 ( n37327, n1977, n37331 );
nand U79263 ( n37319, n37320, n37321 );
nor U79264 ( n37321, n37322, n37323 );
nor U79265 ( n37320, n37327, n37328 );
nand U79266 ( n37322, n37325, n37326 );
nand U79267 ( n49611, n7439, n277 );
not U79268 ( n665, n65938 );
not U79269 ( n687, n64515 );
not U79270 ( n682, n64784 );
nor U79271 ( n41954, n41955, n41956 );
nand U79272 ( n41956, n41957, n41958 );
nand U79273 ( n41955, n682, n41959 );
not U79274 ( n3197, n33744 );
nand U79275 ( n38411, n76819, n38412 );
xnor U79276 ( n16672, n16674, n16675 );
nor U79277 ( n66296, n66298, n66213 );
nor U79278 ( n66298, n643, n645 );
nor U79279 ( n37336, n40107, n1918 );
not U79280 ( n1918, n40113 );
nand U79281 ( n37318, n37332, n37333 );
nor U79282 ( n37332, n37339, n37340 );
nor U79283 ( n37333, n37334, n37335 );
nand U79284 ( n37339, n37343, n37344 );
nor U79285 ( n66343, n61443, n54754 );
nand U79286 ( n61409, n42061, n61410 );
or U79287 ( n41934, n41938, n41939 );
nand U79288 ( n41931, n64805, n677 );
not U79289 ( n677, n64385 );
nand U79290 ( n37371, n1852, n37372 );
nand U79291 ( n37345, n37363, n37364 );
nor U79292 ( n37364, n37365, n37366 );
nor U79293 ( n37363, n37370, n37371 );
nand U79294 ( n37366, n37367, n37368 );
nor U79295 ( n66287, n66219, n66288 );
nand U79296 ( n66288, n647, n61410 );
nand U79297 ( n36775, n36781, n36778 );
nand U79298 ( n36781, n36375, n36374 );
nand U79299 ( n39921, n76798, n38444 );
not U79300 ( n1850, n37302 );
not U79301 ( n1945, n39938 );
not U79302 ( n1955, n39829 );
or U79303 ( n37365, n1955, n37369 );
nand U79304 ( n41949, n65946, n659 );
not U79305 ( n659, n65346 );
not U79306 ( n2014, n36840 );
xor U79307 ( n38555, n40112, n37329 );
nand U79308 ( n38713, n40209, n40210 );
nor U79309 ( n40210, n40211, n40212 );
nor U79310 ( n40209, n40221, n38563 );
nand U79311 ( n40212, n40213, n40214 );
nand U79312 ( n41959, n632, n66206 );
not U79313 ( n632, n66208 );
nand U79314 ( n41158, n41164, n41161 );
nand U79315 ( n41164, n40778, n40777 );
not U79316 ( n638, n66201 );
nor U79317 ( n41938, n640, n638 );
nand U79318 ( n38559, n38560, n38561 );
nand U79319 ( n38561, n76819, n38562 );
nand U79320 ( n38560, n76812, n38563 );
xnor U79321 ( n54813, n66363, n630 );
nand U79322 ( n60768, n66418, n66419 );
nor U79323 ( n66419, n66420, n66421 );
nor U79324 ( n66418, n66430, n54821 );
nand U79325 ( n66421, n66422, n66423 );
nand U79326 ( n39349, n2052, n39321 );
nor U79327 ( n71393, n1224, n1079 );
nor U79328 ( n37459, n2134, n37460 );
not U79329 ( n2142, n38834 );
nand U79330 ( n37323, n2142, n37324 );
not U79331 ( n1978, n39521 );
nand U79332 ( n37328, n37329, n37330 );
nand U79333 ( n65923, n49572, n76077 );
or U79334 ( n37388, n37389, n37390 );
not U79335 ( n2012, n36838 );
nand U79336 ( n37334, n37337, n37338 );
nor U79337 ( n37194, n2179, n76802 );
nor U79338 ( n66737, n625, n66744 );
not U79339 ( n625, n41923 );
nor U79340 ( n66744, n66745, n66746 );
nor U79341 ( n66746, n823, n66441 );
not U79342 ( n524, n66205 );
nand U79343 ( n60875, n66719, n66720 );
nor U79344 ( n66720, n66721, n66722 );
nor U79345 ( n66719, n66734, n54876 );
nand U79346 ( n66722, n66723, n66724 );
nand U79347 ( n39293, n39292, n39294 );
not U79348 ( n810, n61175 );
not U79349 ( n2021, n36841 );
not U79350 ( n4887, n13249 );
nand U79351 ( n37370, n37373, n37374 );
nor U79352 ( n40277, n2002, n40275 );
nor U79353 ( n40267, n1907, n40276 );
not U79354 ( n1907, n37330 );
nor U79355 ( n40276, n40277, n40278 );
nor U79356 ( n40278, n2034, n40273 );
nand U79357 ( n38716, n40249, n40250 );
nor U79358 ( n40250, n40251, n40252 );
nor U79359 ( n40249, n40264, n38578 );
nor U79360 ( n40251, n2159, n38604 );
not U79361 ( n629, n42001 );
not U79362 ( n2103, n37324 );
nand U79363 ( n40237, n1905, n37411 );
not U79364 ( n4929, n14139 );
nor U79365 ( n38983, n38872, n38985 );
not U79366 ( n2130, n37343 );
not U79367 ( n2049, n39346 );
nand U79368 ( n38443, n76819, n38444 );
nand U79369 ( n41951, n652, n647 );
nor U79370 ( n37186, n2180, n76803 );
nand U79371 ( n38989, n38903, n38945 );
nor U79372 ( n36839, n2013, n36439 );
nand U79373 ( n37340, n37341, n37342 );
xor U79374 ( n54868, n41923, n66205 );
not U79375 ( n3185, n33609 );
xor U79376 ( n38570, n37330, n40275 );
and U79377 ( n40280, n38861, n38570 );
nor U79378 ( n40161, n1922, n1927 );
nor U79379 ( n66437, n66438, n66439 );
nor U79380 ( n66438, n41959, n41573 );
nor U79381 ( n66439, n630, n66371 );
nand U79382 ( n36475, n36482, n36483 );
nand U79383 ( n36483, n36480, n36484 );
nand U79384 ( n36484, n2040, n36478 );
xnor U79385 ( MUL_1411_U14, n71504, n71505 );
xnor U79386 ( n71504, n71506, n71507 );
not U79387 ( n728, n62832 );
nand U79388 ( n40235, n37329, n37411 );
nand U79389 ( n40044, n76798, n38500 );
nand U79390 ( n40119, n37368, n37271 );
not U79391 ( n587, n42201 );
nand U79392 ( n42198, n42294, n45202 );
nand U79393 ( n16630, n4795, n26 );
nor U79394 ( n66420, n61443, n54813 );
nor U79395 ( n61174, n61175, n76074 );
not U79396 ( n1963, n36723 );
not U79397 ( n2127, n38948 );
nor U79398 ( n40156, n40103, n1918 );
not U79399 ( n2018, n36701 );
not U79400 ( n702, n41924 );
nand U79401 ( n37138, n37291, n37292 );
nor U79402 ( n38921, n2134, n2135 );
not U79403 ( n2135, n37331 );
nand U79404 ( n36836, n2012, n36435 );
nor U79405 ( n39161, n2114, n37402 );
not U79406 ( n2114, n37326 );
nor U79407 ( n37132, n2192, n37134 );
not U79408 ( n2144, n37387 );
and U79409 ( n36683, n36684, n76830 );
not U79410 ( n588, n41107 );
not U79411 ( n1952, n37337 );
not U79412 ( n3177, n33563 );
not U79413 ( n574, n42193 );
nand U79414 ( n49583, n7439, n270 );
nor U79415 ( n40274, n2002, n37330 );
not U79416 ( n2079, n37694 );
nand U79417 ( n38039, n38098, n38099 );
nand U79418 ( n38098, n37117, n37745 );
nand U79419 ( n38099, n2087, n37745 );
xor U79420 ( n54914, n41962, n66752 );
nand U79421 ( n60973, n66993, n66994 );
nor U79422 ( n66994, n66995, n66996 );
nor U79423 ( n66993, n67005, n54924 );
nand U79424 ( n66996, n66997, n66998 );
xnor U79425 ( n38585, n37372, n40282 );
not U79426 ( n2028, n38109 );
buf U79427 ( n76813, n2030 );
nor U79428 ( n66721, n61443, n54868 );
or U79429 ( n65815, n823, n41939 );
not U79430 ( n4920, n13964 );
not U79431 ( n1973, n37374 );
nor U79432 ( n37182, n2182, n76803 );
or U79433 ( n37144, n37149, n37148 );
nand U79434 ( n38807, n37390, n38792 );
and U79435 ( n37523, n37528, n37390 );
nand U79436 ( n40137, n76798, n38532 );
not U79437 ( n575, n42194 );
nor U79438 ( n66743, n820, n41923 );
nand U79439 ( n40012, n38792, n37352 );
nand U79440 ( n66273, n76075, n54677 );
not U79441 ( n2048, n37338 );
nor U79442 ( n66104, n657, n653 );
not U79443 ( n724, n41932 );
not U79444 ( n1968, n37373 );
not U79445 ( n698, n41957 );
nor U79446 ( n45748, n76059, n45363 );
not U79447 ( n2124, n37342 );
xor U79448 ( n49588, n49589, n49590 );
nand U79449 ( n39978, n38792, n37355 );
not U79450 ( n2118, n37341 );
not U79451 ( n718, n41925 );
not U79452 ( n1980, n39524 );
not U79453 ( n1992, n37367 );
and U79454 ( n13434, n76603, n13414 );
buf U79455 ( n76798, n2070 );
nand U79456 ( n37690, n37779, n38039 );
nand U79457 ( n47674, n47532, n47681 );
nand U79458 ( n47681, n7610, n47682 );
not U79459 ( n693, n41963 );
not U79460 ( n2109, n37325 );
not U79461 ( n4913, n13915 );
not U79462 ( n703, n63670 );
not U79463 ( n2077, n37689 );
nand U79464 ( n40214, n76798, n38562 );
nor U79465 ( n67215, n61443, n523 );
nand U79466 ( n61070, n67212, n67213 );
nor U79467 ( n67212, n67218, n54995 );
nor U79468 ( n67213, n67214, n67215 );
nor U79469 ( n67218, n623, n76062 );
nor U79470 ( n66995, n54914, n61443 );
nand U79471 ( n66423, n76074, n54820 );
nor U79472 ( n71543, n1235, n1057 );
nand U79473 ( n47532, n7609, n47684 );
nand U79474 ( n47684, n47682, n44985 );
not U79475 ( n1053, n71957 );
xor U79476 ( n47679, n44985, n47682 );
not U79477 ( n7609, n47683 );
xor U79478 ( n47525, n47532, n47533 );
xor U79479 ( MUL_1411_U386, n71066, n71067 );
xor U79480 ( n71067, n71068, n71069 );
nand U79481 ( n33939, n33797, n33946 );
nand U79482 ( n33946, n3224, n33947 );
nand U79483 ( n16594, n4795, n21 );
nand U79484 ( n68695, n68553, n68702 );
nand U79485 ( n68702, n5823, n68703 );
nand U79486 ( n26694, n26552, n26701 );
nand U79487 ( n26701, n4054, n26702 );
nand U79488 ( n59836, n59694, n59843 );
nand U79489 ( n59843, n6687, n59844 );
nand U79490 ( n66998, n76081, n54922 );
nor U79491 ( n71380, n1234, n1057 );
nand U79492 ( n33797, n3223, n33949 );
nand U79493 ( n33949, n33947, n31607 );
nand U79494 ( n47482, n7592, n47540 );
nand U79495 ( n26552, n4053, n26704 );
nand U79496 ( n26704, n26702, n24311 );
nand U79497 ( n59694, n6685, n59846 );
nand U79498 ( n59846, n59844, n57434 );
nand U79499 ( n68553, n5822, n68705 );
nand U79500 ( n68705, n68703, n65893 );
nor U79501 ( n37098, n2044, n2045 );
not U79502 ( n2004, n36843 );
buf U79503 ( n76804, n76800 );
buf U79504 ( n76800, n2065 );
xor U79505 ( n33944, n31607, n33947 );
xor U79506 ( n68700, n65893, n68703 );
xor U79507 ( n26699, n24311, n26702 );
xor U79508 ( n59841, n57434, n59844 );
not U79509 ( n3223, n33948 );
nor U79510 ( n37164, n2185, n76803 );
not U79511 ( n5822, n68704 );
not U79512 ( n6685, n59845 );
not U79513 ( n4053, n26703 );
not U79514 ( n2087, n37108 );
xor U79515 ( n33790, n33797, n33798 );
xor U79516 ( n68546, n68553, n68554 );
xor U79517 ( n26545, n26552, n26553 );
xor U79518 ( n59687, n59694, n59695 );
nand U79519 ( n49537, n7439, n264 );
nand U79520 ( n14400, n14205, n14409 );
nand U79521 ( n14409, n4957, n14410 );
nand U79522 ( n47443, n47532, n47533 );
nand U79523 ( n14205, n4955, n14413 );
nand U79524 ( n14413, n14410, n11304 );
nand U79525 ( n33747, n3205, n33805 );
xor U79526 ( n47618, n47602, n47533 );
xor U79527 ( n47337, n47332, n47333 );
nand U79528 ( n68503, n5804, n68561 );
nand U79529 ( n26502, n4038, n26560 );
nand U79530 ( n59641, n6670, n59702 );
not U79531 ( n2080, n37745 );
xor U79532 ( n14407, n11304, n14410 );
not U79533 ( n4955, n14412 );
xor U79534 ( n14197, n14205, n14207 );
nand U79535 ( n33708, n33797, n33798 );
nand U79536 ( n26463, n26552, n26553 );
nand U79537 ( n59602, n59694, n59695 );
nand U79538 ( n68464, n68553, n68554 );
not U79539 ( n579, n41445 );
not U79540 ( n1037, n71937 );
nand U79541 ( n14143, n4938, n14215 );
xor U79542 ( n47350, n47432, n47333 );
xor U79543 ( n33613, n33608, n33609 );
xor U79544 ( n68369, n68364, n68365 );
xor U79545 ( n26368, n26363, n26364 );
xor U79546 ( n59507, n59502, n59503 );
nand U79547 ( n40884, n579, n41476 );
nand U79548 ( n41476, n41477, n41478 );
nand U79549 ( n41478, n41311, n41443 );
nor U79550 ( n37153, n2188, n76803 );
nand U79551 ( n16557, n4795, n16 );
xor U79552 ( n33883, n33867, n33798 );
xor U79553 ( n68639, n68623, n68554 );
xor U79554 ( n26638, n26622, n26553 );
xor U79555 ( n59780, n59764, n59695 );
nand U79556 ( n14094, n14205, n14207 );
or U79557 ( n36488, n36292, n76039 );
nand U79558 ( n49508, n7439, n258 );
not U79559 ( n76255, n76256 );
xor U79560 ( n14313, n14293, n14207 );
xor U79561 ( n33626, n33697, n33609 );
xor U79562 ( n13969, n13963, n13964 );
xor U79563 ( n68382, n68453, n68365 );
xor U79564 ( n26381, n26452, n26364 );
xor U79565 ( n59520, n59591, n59503 );
nand U79566 ( n36801, n2892, n36292 );
nand U79567 ( n36576, n2889, n36292 );
nand U79568 ( n36326, n2918, n36292 );
nand U79569 ( n36536, n2915, n36292 );
nand U79570 ( n36359, n2913, n36292 );
nand U79571 ( n36466, n2910, n36292 );
nand U79572 ( n36821, n2919, n36292 );
and U79573 ( n47240, n47332, n47333 );
nor U79574 ( n37149, n2189, n76804 );
not U79575 ( n76425, n76426 );
xor U79576 ( n13993, n14080, n13964 );
xor U79577 ( MUL_1411_U387, n71062, n71063 );
xor U79578 ( n71063, n71064, n71065 );
nand U79579 ( n49475, n7439, n252 );
buf U79580 ( n76814, n2030 );
and U79581 ( n33516, n33608, n33609 );
and U79582 ( n26270, n26363, n26364 );
and U79583 ( n59409, n59502, n59503 );
and U79584 ( n68271, n68364, n68365 );
xnor U79585 ( n47245, n47287, n7530 );
nand U79586 ( n47287, n47240, n47288 );
nand U79587 ( n16520, n4795, n11 );
buf U79588 ( n75996, n76257 );
buf U79589 ( n75994, n76257 );
buf U79590 ( n75995, n76257 );
nand U79591 ( n26904, n26918, n23826 );
nand U79592 ( n60044, n60058, n56950 );
nand U79593 ( n28485, n28726, n28727 );
nor U79594 ( n28726, n26903, n28336 );
nor U79595 ( n28727, n3978, n26904 );
nand U79596 ( n61790, n62031, n62032 );
nor U79597 ( n62031, n60043, n61558 );
nor U79598 ( n62032, n6610, n60044 );
and U79599 ( n75755, n56380, n6610 );
and U79600 ( n75756, n23256, n3978 );
nand U79601 ( n68903, n68917, n65424 );
nand U79602 ( n70390, n70631, n70632 );
nor U79603 ( n70631, n68902, n70274 );
nor U79604 ( n70632, n5735, n68903 );
and U79605 ( n75757, n64736, n5735 );
nand U79606 ( n34149, n34163, n31170 );
nand U79607 ( n35664, n35905, n35906 );
nor U79608 ( n35905, n34148, n35546 );
nor U79609 ( n35906, n3134, n34149 );
and U79610 ( n75758, n30577, n3134 );
not U79611 ( n4059, n24601 );
not U79612 ( n6692, n57733 );
not U79613 ( n5830, n66409 );
not U79614 ( n3232, n31817 );
not U79615 ( n3978, n23077 );
not U79616 ( n6610, n56198 );
not U79617 ( n5735, n64567 );
not U79618 ( n3134, n30408 );
not U79619 ( n6699, n61512 );
not U79620 ( n4067, n28290 );
not U79621 ( n5842, n70246 );
not U79622 ( n3242, n35518 );
not U79623 ( n2062, n36492 );
not U79624 ( n825, n61618 );
not U79625 ( n585, n41229 );
nor U79626 ( n41467, n824, n825 );
and U79627 ( n13857, n13963, n13964 );
xnor U79628 ( n33521, n33562, n3143 );
nand U79629 ( n33562, n33516, n33563 );
xnor U79630 ( n68276, n68318, n5744 );
nand U79631 ( n68318, n68271, n68319 );
xnor U79632 ( n26275, n26317, n3987 );
nand U79633 ( n26317, n26270, n26318 );
xnor U79634 ( n59414, n59456, n6619 );
nand U79635 ( n59456, n59409, n59457 );
buf U79636 ( n76017, n76427 );
buf U79637 ( n76016, n76427 );
buf U79638 ( n76015, n76427 );
buf U79639 ( n76744, n76740 );
nand U79640 ( n28481, n28648, n28649 );
nor U79641 ( n28648, n23826, n26918 );
nor U79642 ( n28649, n26903, n28650 );
nand U79643 ( n28650, n28336, n23077 );
nand U79644 ( n61786, n61953, n61954 );
nor U79645 ( n61953, n56950, n60058 );
nor U79646 ( n61954, n60043, n61955 );
nand U79647 ( n61955, n61558, n56198 );
nor U79648 ( n28565, n28481, n26905 );
nor U79649 ( n61870, n61786, n60045 );
nand U79650 ( n70386, n70553, n70554 );
nor U79651 ( n70553, n65424, n68917 );
nor U79652 ( n70554, n68902, n70555 );
nand U79653 ( n70555, n70274, n64567 );
nor U79654 ( n70470, n70386, n68904 );
nand U79655 ( n35660, n35827, n35828 );
nor U79656 ( n35827, n31170, n34163 );
nor U79657 ( n35828, n34148, n35829 );
nand U79658 ( n35829, n35546, n30408 );
nor U79659 ( n35744, n35660, n34150 );
buf U79660 ( n76742, n76740 );
buf U79661 ( n76439, n76437 );
buf U79662 ( n76438, n76437 );
buf U79663 ( n76677, n76673 );
nand U79664 ( n16479, n4795, n6 );
buf U79665 ( n76675, n76673 );
buf U79666 ( n76442, n76441 );
buf U79667 ( n76443, n76441 );
buf U79668 ( n76446, n76445 );
buf U79669 ( n76440, n76437 );
buf U79670 ( n76447, n76445 );
buf U79671 ( n76444, n76441 );
nand U79672 ( n38474, n76446, n2910 );
nand U79673 ( n38375, n76447, n2918 );
buf U79674 ( n76448, n76445 );
nand U79675 ( n29177, n3232, n35518 );
nand U79676 ( n32586, n76774, n3387 );
not U79677 ( n7618, n45509 );
nand U79678 ( n21864, n4059, n28290 );
nand U79679 ( n62899, n5830, n70246 );
nand U79680 ( n54955, n6692, n61512 );
nand U79681 ( n42390, n7618, n49449 );
nand U79682 ( n67351, n76708, n6002 );
nand U79683 ( n46290, n76660, n7789 );
nand U79684 ( n25344, n76754, n4224 );
nand U79685 ( n58483, n76687, n6857 );
not U79686 ( n4047, n26905 );
not U79687 ( n6679, n60045 );
not U79688 ( n5815, n68904 );
not U79689 ( n3217, n34150 );
nand U79690 ( n24316, n4009, n26918 );
nand U79691 ( n57439, n6642, n60058 );
not U79692 ( n4009, n23826 );
not U79693 ( n6642, n56950 );
nand U79694 ( n65898, n5768, n68917 );
not U79695 ( n5768, n65424 );
nand U79696 ( n31612, n3169, n34163 );
not U79697 ( n3169, n31170 );
not U79698 ( n7520, n43725 );
not U79699 ( n4035, n28336 );
not U79700 ( n6668, n61558 );
not U79701 ( n5802, n70274 );
not U79702 ( n3203, n35546 );
not U79703 ( n2027, n36489 );
not U79704 ( n7603, n47884 );
not U79705 ( n4964, n11733 );
nand U79706 ( n8304, n4964, n16448 );
nand U79707 ( n12677, n76727, n5134 );
not U79708 ( n7589, n49545 );
not U79709 ( n4782, n12150 );
not U79710 ( n3045, n32252 );
not U79711 ( n5647, n66891 );
not U79712 ( n3044, n32317 );
not U79713 ( n7422, n45940 );
not U79714 ( n3889, n25015 );
not U79715 ( n6522, n58150 );
not U79716 ( n5645, n66956 );
not U79717 ( n7420, n46016 );
not U79718 ( n3888, n25080 );
not U79719 ( n6520, n58215 );
not U79720 ( n4875, n9804 );
not U79721 ( n4949, n14654 );
buf U79722 ( n76409, n75777 );
nand U79723 ( n22756, n24601, n28290 );
nand U79724 ( n55870, n57733, n61512 );
nand U79725 ( n64094, n66409, n70246 );
nand U79726 ( n30077, n31817, n35518 );
nor U79727 ( n41473, n835, n837 );
and U79728 ( n41470, n41472, n41473 );
nand U79729 ( n47883, n47897, n44495 );
not U79730 ( n4935, n16567 );
buf U79731 ( n76743, n76740 );
not U79732 ( n4778, n12253 );
not U79733 ( n4777, n12334 );
xnor U79734 ( n13863, n13914, n4885 );
nand U79735 ( n13914, n13857, n13915 );
not U79736 ( n3192, n34148 );
not U79737 ( n5790, n68902 );
not U79738 ( n6659, n60043 );
not U79739 ( n7578, n47882 );
not U79740 ( n4027, n26903 );
nor U79741 ( n39605, n2047, n2005 );
nor U79742 ( n36947, n2175, n76454 );
nor U79743 ( n36540, n2188, n76455 );
nor U79744 ( n36495, n2183, n76455 );
nor U79745 ( n36658, n2168, n76454 );
nor U79746 ( n36687, n2182, n76454 );
nor U79747 ( n36389, n2180, n76455 );
nor U79748 ( n36754, n2170, n76454 );
nor U79749 ( n36453, n2167, n76455 );
nor U79750 ( n36406, n2192, n76455 );
nor U79751 ( n36709, n2173, n76454 );
nor U79752 ( n36519, n2172, n76455 );
nor U79753 ( n36825, n2189, n76454 );
nor U79754 ( n36640, n2162, n76454 );
nor U79755 ( n36365, n2160, n76455 );
buf U79756 ( n76676, n76673 );
nor U79757 ( n36805, n2164, n76454 );
nor U79758 ( n36621, n2187, n76455 );
nor U79759 ( n36599, n2178, n76455 );
nor U79760 ( n36788, n2179, n76454 );
nor U79761 ( n36580, n2163, n76455 );
nor U79762 ( n36738, n2184, n76454 );
nor U79763 ( n36558, n2177, n76455 );
nand U79764 ( n14653, n14670, n10697 );
not U79765 ( n837, n62272 );
nor U79766 ( n36346, n2169, n76456 );
nor U79767 ( n36330, n2185, n76456 );
nor U79768 ( n36313, n2174, n76456 );
nor U79769 ( n36296, n2190, n76456 );
nor U79770 ( n36268, n2165, n76456 );
not U79771 ( n4925, n14652 );
nor U79772 ( n32562, n76776, n76480 );
buf U79773 ( n76776, n3062 );
nor U79774 ( n67327, n76710, n76202 );
nor U79775 ( n25320, n76758, n76526 );
nor U79776 ( n58459, n76691, n76268 );
buf U79777 ( n76758, n3905 );
buf U79778 ( n76691, n6538 );
buf U79779 ( n76710, n5663 );
and U79780 ( n37101, n37103, n37104 );
nor U79781 ( n46266, n76662, n76346 );
buf U79782 ( n76662, n7437 );
nor U79783 ( n40329, n2157, n38604 );
nor U79784 ( n62834, n743, n76062 );
not U79785 ( n7530, n46277 );
or U79786 ( n40881, n40696, n76041 );
nor U79787 ( n12638, n76729, n76607 );
buf U79788 ( n76729, n4793 );
nand U79789 ( n40714, n41067, n41308 );
nand U79790 ( n41308, n41309, n76925 );
nand U79791 ( n41309, n603, n41310 );
nand U79792 ( n41310, n41311, n617 );
nand U79793 ( n41182, n1775, n40696 );
nand U79794 ( n40971, n1773, n40696 );
nand U79795 ( n40731, n1800, n40696 );
nand U79796 ( n40934, n1798, n40696 );
nand U79797 ( n40764, n1795, n40696 );
nand U79798 ( n40868, n1793, n40696 );
nand U79799 ( n41202, n1802, n40696 );
nor U79800 ( n41063, n623, n76111 );
nor U79801 ( n41186, n654, n76106 );
nor U79802 ( n40718, n700, n76107 );
nor U79803 ( n41014, n750, n40708 );
nor U79804 ( n41153, n623, n40708 );
nor U79805 ( n41122, n743, n40708 );
nor U79806 ( n40891, n737, n40708 );
nor U79807 ( n41137, n684, n76109 );
nor U79808 ( n40855, n667, n76113 );
buf U79809 ( n76113, n40691 );
nor U79810 ( n40735, n745, n40708 );
nor U79811 ( n40792, n737, n76114 );
buf U79812 ( n76114, n40691 );
nor U79813 ( n36770, n2157, n36489 );
not U79814 ( n584, n40708 );
not U79815 ( n617, n41443 );
nand U79816 ( n41469, n832, n61624 );
nor U79817 ( n40872, n624, n40708 );
nor U79818 ( n40751, n679, n76106 );
nor U79819 ( n40700, n764, n40708 );
nor U79820 ( n40938, n754, n40708 );
nor U79821 ( n41078, n730, n40708 );
nor U79822 ( n41315, n707, n76105 );
nor U79823 ( n41169, n730, n76107 );
nor U79824 ( n40975, n650, n76111 );
nor U79825 ( n41027, n648, n76109 );
buf U79826 ( n76638, n75775 );
nor U79827 ( n40809, n768, n40708 );
nor U79828 ( n41045, n672, n76112 );
not U79829 ( n3143, n32573 );
nor U79830 ( n40917, n689, n76113 );
nor U79831 ( n40992, n720, n76110 );
nor U79832 ( n41093, n695, n76110 );
nor U79833 ( n40768, n639, n76105 );
nand U79834 ( n41067, n41447, n617 );
not U79835 ( n5744, n67338 );
not U79836 ( n6619, n58470 );
not U79837 ( n3987, n25331 );
nor U79838 ( n40953, n714, n76112 );
nor U79839 ( n40672, n660, n76108 );
buf U79840 ( n76777, n3062 );
nor U79841 ( n36470, n2155, n36489 );
nor U79842 ( n41064, n41065, n41066 );
nand U79843 ( n41065, n41068, n76925 );
nand U79844 ( n41066, n603, n41067 );
nand U79845 ( n41068, n41475, n41311 );
nor U79846 ( n41475, n41443, n41445 );
buf U79847 ( n76759, n3905 );
buf U79848 ( n76711, n5663 );
buf U79849 ( n76692, n6538 );
buf U79850 ( n76663, n7437 );
nand U79851 ( n36681, n37107, n76409 );
nor U79852 ( n37107, n2090, n37108 );
nor U79853 ( n28569, n26905, n28336 );
nor U79854 ( n61874, n60045, n61558 );
nor U79855 ( n28568, n4009, n26918 );
nor U79856 ( n61873, n6642, n60058 );
nor U79857 ( n70474, n68904, n70274 );
nor U79858 ( n35748, n34150, n35546 );
nor U79859 ( n70473, n5768, n68917 );
nor U79860 ( n35747, n3169, n34163 );
buf U79861 ( n76730, n4793 );
nand U79862 ( n35767, n35768, n35769 );
nand U79863 ( n35769, n35770, n34148 );
nand U79864 ( n35768, n3217, n35772 );
nand U79865 ( n35770, n35771, n34149 );
nand U79866 ( n28588, n28589, n28590 );
nand U79867 ( n28590, n28591, n26903 );
nand U79868 ( n28589, n4047, n28593 );
nand U79869 ( n28591, n28592, n26904 );
nand U79870 ( n70493, n70494, n70495 );
nand U79871 ( n70495, n70496, n68902 );
nand U79872 ( n70494, n5815, n70498 );
nand U79873 ( n70496, n70497, n68903 );
nand U79874 ( n61893, n61894, n61895 );
nand U79875 ( n61895, n61896, n60043 );
nand U79876 ( n61894, n6679, n61898 );
nand U79877 ( n61896, n61897, n60044 );
nand U79878 ( n35772, n35773, n35774 );
nor U79879 ( n35774, n35775, n35776 );
nor U79880 ( n35773, n35779, n35780 );
nand U79881 ( n35776, n35777, n30408 );
nand U79882 ( n28593, n28594, n28595 );
nor U79883 ( n28595, n28596, n28597 );
nor U79884 ( n28594, n28600, n28601 );
nand U79885 ( n28597, n28598, n23077 );
nand U79886 ( n70498, n70499, n70500 );
nor U79887 ( n70500, n70501, n70502 );
nor U79888 ( n70499, n70505, n70506 );
nand U79889 ( n70502, n70503, n64567 );
nand U79890 ( n61898, n61899, n61900 );
nor U79891 ( n61900, n61901, n61902 );
nor U79892 ( n61899, n61905, n61906 );
nand U79893 ( n61902, n61903, n56198 );
nand U79894 ( n54265, n54266, n54267 );
nand U79895 ( n54267, n54268, n47882 );
nand U79896 ( n54266, n7603, n54270 );
nand U79897 ( n54268, n54269, n47883 );
nand U79898 ( n54270, n54271, n54272 );
nor U79899 ( n54272, n54273, n54274 );
nor U79900 ( n54271, n54277, n54278 );
nand U79901 ( n54274, n54275, n43725 );
buf U79902 ( n76785, n3040 );
buf U79903 ( n76671, n7417 );
buf U79904 ( n76767, n3884 );
buf U79905 ( n76719, n5642 );
buf U79906 ( n76700, n6517 );
buf U79907 ( n76784, n3040 );
buf U79908 ( n76766, n3884 );
buf U79909 ( n76670, n7417 );
buf U79910 ( n76718, n5642 );
buf U79911 ( n76699, n6517 );
not U79912 ( n7629, n49449 );
xor U79913 ( MUL_1411_U388, n71058, n71059 );
xor U79914 ( n71059, n71060, n71061 );
buf U79915 ( n76786, n3040 );
buf U79916 ( n76768, n3884 );
buf U79917 ( n76701, n6517 );
buf U79918 ( n76672, n7417 );
buf U79919 ( n76720, n5642 );
nor U79920 ( n54213, n7509, n7803 );
nor U79921 ( n35715, n3123, n3400 );
nor U79922 ( n28536, n3965, n4238 );
nor U79923 ( n70441, n5723, n6015 );
nor U79924 ( n61841, n6598, n6870 );
buf U79925 ( n76738, n4773 );
not U79926 ( n583, n40691 );
buf U79927 ( n76737, n4773 );
not U79928 ( n4975, n16448 );
nor U79929 ( n12833, n21341, n21179 );
nand U79930 ( n21341, n14654, n4967 );
nand U79931 ( n9420, n4975, n11733 );
nor U79932 ( n46405, n54324, n54162 );
nand U79933 ( n54324, n47884, n7620 );
nand U79934 ( n43363, n7629, n45509 );
nand U79935 ( n21273, n21274, n21275 );
nand U79936 ( n21275, n21276, n14652 );
nand U79937 ( n21274, n4949, n21278 );
nand U79938 ( n21276, n21277, n14653 );
nand U79939 ( n21278, n21279, n21280 );
nor U79940 ( n21280, n21281, n21282 );
nor U79941 ( n21279, n21285, n21286 );
nand U79942 ( n21282, n21283, n9804 );
buf U79943 ( n76739, n4773 );
not U79944 ( n4885, n12660 );
buf U79945 ( n76401, n75776 );
not U79946 ( n3042, n32553 );
not U79947 ( n3885, n25311 );
not U79948 ( n7418, n46257 );
not U79949 ( n5643, n67209 );
not U79950 ( n6518, n58450 );
nor U79951 ( n35775, n3232, n35546 );
nor U79952 ( n28596, n4059, n28336 );
nor U79953 ( n70501, n5830, n70274 );
nor U79954 ( n61901, n6692, n61558 );
nor U79955 ( n54273, n7618, n49545 );
nand U79956 ( n44990, n7554, n47897 );
not U79957 ( n7554, n44495 );
not U79958 ( n3075, n30405 );
not U79959 ( n5677, n64564 );
not U79960 ( n7462, n43722 );
not U79961 ( n4818, n9800 );
not U79962 ( n3919, n23074 );
not U79963 ( n6552, n56195 );
nor U79964 ( n21294, n4864, n5148 );
nand U79965 ( n11310, n4905, n14670 );
not U79966 ( n4905, n10697 );
not U79967 ( n4774, n12627 );
buf U79968 ( n76111, n76104 );
buf U79969 ( n76107, n76103 );
buf U79970 ( n76106, n76103 );
buf U79971 ( n76110, n76104 );
buf U79972 ( n76109, n76104 );
buf U79973 ( n76105, n76103 );
buf U79974 ( n76112, n76104 );
buf U79975 ( n76108, n76103 );
nand U79976 ( n21175, n21342, n21343 );
nor U79977 ( n21342, n10697, n14670 );
nor U79978 ( n21343, n14652, n21344 );
nand U79979 ( n21344, n16567, n9804 );
nor U79980 ( n21290, n21175, n14654 );
nand U79981 ( n21179, n21420, n21421 );
nor U79982 ( n21420, n14652, n16567 );
nor U79983 ( n21421, n4875, n14653 );
nand U79984 ( n54158, n54325, n54326 );
nor U79985 ( n54325, n44495, n47897 );
nor U79986 ( n54326, n47882, n54327 );
nand U79987 ( n54327, n49545, n43725 );
nor U79988 ( n54242, n54158, n47884 );
nand U79989 ( n54162, n54403, n54404 );
nor U79990 ( n54403, n47882, n49545 );
nor U79991 ( n54404, n7520, n47883 );
nand U79992 ( n35777, n35778, n3169 );
nor U79993 ( n35778, n34148, n35518 );
nand U79994 ( n28598, n28599, n4009 );
nor U79995 ( n28599, n26903, n28290 );
nand U79996 ( n70503, n70504, n5768 );
nor U79997 ( n70504, n68902, n70246 );
nand U79998 ( n61903, n61904, n6642 );
nor U79999 ( n61904, n60043, n61512 );
nand U80000 ( n54275, n54276, n7554 );
nor U80001 ( n54276, n47882, n49449 );
buf U80002 ( n76059, n54990 );
nor U80003 ( n21281, n4964, n16567 );
nor U80004 ( n67469, n70552, n70390 );
nand U80005 ( n70552, n68904, n5833 );
nor U80006 ( n32704, n35826, n35664 );
nand U80007 ( n35826, n34150, n3234 );
nor U80008 ( n25464, n28647, n28485 );
nand U80009 ( n28647, n26905, n4062 );
nor U80010 ( n58601, n61952, n61790 );
nand U80011 ( n61952, n60045, n6694 );
nand U80012 ( n30090, n3242, n31817 );
nand U80013 ( n22769, n4067, n24601 );
nand U80014 ( n64107, n5842, n66409 );
nand U80015 ( n55883, n6699, n57733 );
not U80016 ( n822, n61624 );
nor U80017 ( n28613, n28616, n26905 );
nor U80018 ( n28616, n28617, n28618 );
nand U80019 ( n28617, n28622, n28623 );
nand U80020 ( n28618, n28619, n28620 );
nor U80021 ( n61918, n61921, n60045 );
nor U80022 ( n61921, n61922, n61923 );
nand U80023 ( n61922, n61927, n61928 );
nand U80024 ( n61923, n61924, n61925 );
nor U80025 ( n35792, n35795, n34150 );
nor U80026 ( n35795, n35796, n35797 );
nand U80027 ( n35796, n35801, n35802 );
nand U80028 ( n35797, n35798, n35799 );
nor U80029 ( n70518, n70521, n68904 );
nor U80030 ( n70521, n70522, n70523 );
nand U80031 ( n70522, n70527, n70528 );
nand U80032 ( n70523, n70524, n70525 );
buf U80033 ( n76894, n215 );
buf U80034 ( n76903, n182 );
buf U80035 ( n76877, n453 );
buf U80036 ( n76868, n487 );
nand U80037 ( n12678, n5132, n12679 );
buf U80038 ( n76376, n76377 );
nand U80039 ( n21283, n21284, n4905 );
nor U80040 ( n21284, n14652, n16448 );
nand U80041 ( n43808, n43889, n7520 );
nand U80042 ( n9908, n9965, n4875 );
buf U80043 ( n76895, n215 );
buf U80044 ( n76869, n487 );
buf U80045 ( n76904, n182 );
buf U80046 ( n76878, n453 );
nand U80047 ( n32587, n3384, n32588 );
buf U80048 ( n76896, n215 );
buf U80049 ( n76870, n487 );
buf U80050 ( n76905, n182 );
buf U80051 ( n76879, n453 );
nand U80052 ( n67352, n5999, n67353 );
nand U80053 ( n25345, n4222, n25346 );
nand U80054 ( n58484, n6854, n58485 );
nor U80055 ( n54246, n47884, n49545 );
not U80056 ( n189, n35678 );
not U80057 ( n152, n28499 );
not U80058 ( n460, n70404 );
not U80059 ( n424, n61804 );
nand U80060 ( n46291, n7787, n46292 );
not U80061 ( n494, n54176 );
nor U80062 ( n54290, n54293, n47884 );
nor U80063 ( n54293, n54294, n54295 );
nand U80064 ( n54294, n54299, n54300 );
nand U80065 ( n54295, n54296, n54297 );
nand U80066 ( n35746, n3229, n30408 );
nand U80067 ( n28567, n4057, n23077 );
nand U80068 ( n70472, n5828, n64567 );
nand U80069 ( n61872, n6689, n56198 );
and U80070 ( n35687, n35742, n35743 );
nand U80071 ( n35743, n35744, n35518 );
nor U80072 ( n35742, n32704, n35745 );
nor U80073 ( n35745, n35739, n35746 );
and U80074 ( n28508, n28563, n28564 );
nand U80075 ( n28564, n28565, n28290 );
nor U80076 ( n28563, n25464, n28566 );
nor U80077 ( n28566, n28560, n28567 );
and U80078 ( n70413, n70468, n70469 );
nand U80079 ( n70469, n70470, n70246 );
nor U80080 ( n70468, n67469, n70471 );
nor U80081 ( n70471, n70465, n70472 );
and U80082 ( n61813, n61868, n61869 );
nand U80083 ( n61869, n61870, n61512 );
nor U80084 ( n61868, n58601, n61871 );
nor U80085 ( n61871, n61865, n61872 );
nand U80086 ( n54244, n7615, n43725 );
and U80087 ( n54185, n54240, n54241 );
nand U80088 ( n54241, n54242, n49449 );
nor U80089 ( n54240, n46405, n54243 );
nor U80090 ( n54243, n54237, n54244 );
nand U80091 ( n35761, n3203, n35762 );
nand U80092 ( n35762, n3242, n30408 );
nand U80093 ( n28582, n4035, n28583 );
nand U80094 ( n28583, n4067, n23077 );
nand U80095 ( n70487, n5802, n70488 );
nand U80096 ( n70488, n5842, n64567 );
nand U80097 ( n61887, n6668, n61888 );
nand U80098 ( n61888, n6699, n56198 );
nand U80099 ( n54259, n7589, n54260 );
nand U80100 ( n54260, n7629, n43725 );
not U80101 ( n223, n21202 );
nor U80102 ( n21307, n21310, n14654 );
nor U80103 ( n21310, n21311, n21312 );
nand U80104 ( n21311, n21316, n21317 );
nand U80105 ( n21312, n21313, n21314 );
not U80106 ( n3183, n34163 );
not U80107 ( n4020, n26918 );
not U80108 ( n5782, n68917 );
not U80109 ( n6653, n60058 );
nand U80110 ( n35771, n3183, n35546 );
nand U80111 ( n28592, n4020, n28336 );
nand U80112 ( n70497, n5782, n70274 );
nand U80113 ( n61897, n6653, n61558 );
not U80114 ( n7569, n47897 );
nand U80115 ( n54269, n7569, n49545 );
nor U80116 ( n21271, n14654, n16567 );
nand U80117 ( n21292, n4962, n9804 );
and U80118 ( n21201, n21288, n21289 );
nand U80119 ( n21289, n21290, n16448 );
nor U80120 ( n21288, n12833, n21291 );
nor U80121 ( n21291, n21239, n21292 );
nand U80122 ( n49444, n7439, n245 );
buf U80123 ( n76863, n502 );
buf U80124 ( n76451, n76452 );
buf U80125 ( n76619, n76620 );
and U80126 ( n35802, n35764, n30408 );
and U80127 ( n28623, n28585, n23077 );
and U80128 ( n70528, n70490, n64567 );
and U80129 ( n61928, n61890, n56198 );
and U80130 ( n54300, n54262, n43725 );
buf U80131 ( n76533, n76534 );
buf U80132 ( n76275, n76276 );
buf U80133 ( n76209, n76210 );
nor U80134 ( n35811, n3387, n35812 );
nor U80135 ( n35812, n76774, n32630 );
nor U80136 ( n28632, n4224, n28633 );
nor U80137 ( n28633, n76754, n25390 );
nor U80138 ( n70537, n6002, n70538 );
nor U80139 ( n70538, n76708, n67395 );
nor U80140 ( n61937, n6857, n61938 );
nor U80141 ( n61938, n76687, n58527 );
nor U80142 ( n54309, n7789, n54310 );
nor U80143 ( n54310, n76660, n46331 );
nand U80144 ( n21266, n4935, n21267 );
nand U80145 ( n21267, n4975, n9804 );
buf U80146 ( n76890, n230 );
nand U80147 ( n43350, n45509, n49449 );
buf U80148 ( n76862, n502 );
not U80149 ( n2005, n38872 );
buf U80150 ( n76353, n76354 );
nand U80151 ( n26907, n4222, n23826 );
nand U80152 ( n60047, n6854, n56950 );
nand U80153 ( n34152, n3384, n31170 );
nand U80154 ( n68906, n5999, n65424 );
nor U80155 ( n21293, n4905, n14670 );
nor U80156 ( n54245, n7554, n47897 );
nand U80157 ( n21986, n21997, n22002 );
nand U80158 ( n29301, n29316, n29321 );
nand U80159 ( n63068, n63079, n63084 );
nand U80160 ( n55096, n55107, n55112 );
buf U80161 ( n76864, n502 );
nand U80162 ( n9404, n11733, n16448 );
buf U80163 ( n76889, n230 );
nor U80164 ( n21326, n5134, n21327 );
nor U80165 ( n21327, n76727, n12732 );
and U80166 ( n21317, n21269, n9804 );
not U80167 ( n4918, n14670 );
nand U80168 ( n21277, n4918, n16567 );
nand U80169 ( n35760, n35546, n34150 );
nand U80170 ( n28581, n28336, n26905 );
nand U80171 ( n70486, n70274, n68904 );
nand U80172 ( n61886, n61558, n60045 );
nand U80173 ( n54258, n49545, n47884 );
nor U80174 ( n28615, n28290, n28485 );
nor U80175 ( n61920, n61512, n61790 );
nor U80176 ( n35794, n35518, n35664 );
nor U80177 ( n70520, n70246, n70390 );
not U80178 ( n3073, n30116 );
not U80179 ( n5674, n64129 );
not U80180 ( n3917, n22791 );
not U80181 ( n6549, n55905 );
not U80182 ( n7459, n43385 );
not U80183 ( n4815, n9448 );
nand U80184 ( n30200, n76024, n3677 );
nand U80185 ( n30223, n76024, n3678 );
nand U80186 ( n30242, n76023, n3679 );
nand U80187 ( n30261, n76023, n3680 );
nand U80188 ( n30280, n76023, n3682 );
nand U80189 ( n30299, n76023, n3683 );
nand U80190 ( n30358, n76024, n3687 );
nand U80191 ( n30162, n76023, n3674 );
nand U80192 ( n30181, n76024, n3675 );
nand U80193 ( n43502, n76008, n8092 );
nand U80194 ( n43521, n76008, n8093 );
nand U80195 ( n43540, n76007, n8094 );
nand U80196 ( n43572, n76007, n8095 );
nand U80197 ( n64266, n75992, n6310 );
nand U80198 ( n64285, n75992, n6312 );
nand U80199 ( n64304, n75991, n6313 );
nand U80200 ( n64323, n75991, n6314 );
nand U80201 ( n64403, n75991, n6315 );
nand U80202 ( n64422, n75991, n6317 );
nand U80203 ( n9553, n76037, n5437 );
nand U80204 ( n9577, n76037, n5438 );
nand U80205 ( n9599, n76036, n5439 );
nand U80206 ( n9647, n76036, n5442 );
nand U80207 ( n9674, n76036, n5443 );
nand U80208 ( n9743, n76037, n5447 );
nand U80209 ( n64477, n75992, n6320 );
nand U80210 ( n43591, n76007, n8097 );
nand U80211 ( n43610, n76007, n8098 );
nand U80212 ( n43679, n76008, n8102 );
nand U80213 ( n9623, n76036, n5440 );
nand U80214 ( n43464, n76007, n8089 );
nand U80215 ( n64175, n75991, n6308 );
nand U80216 ( n22837, n76028, n4568 );
nand U80217 ( n55951, n75999, n7200 );
nand U80218 ( n43483, n76008, n8090 );
nand U80219 ( n64247, n75992, n6309 );
nand U80220 ( n22856, n76029, n4569 );
nand U80221 ( n22877, n76029, n4570 );
nand U80222 ( n22896, n76029, n4572 );
nand U80223 ( n22915, n76028, n4573 );
nand U80224 ( n22934, n76028, n4574 );
nand U80225 ( n22953, n76028, n4575 );
nand U80226 ( n22974, n76028, n4577 );
nand U80227 ( n23029, n76029, n4580 );
nand U80228 ( n9505, n76036, n5434 );
nand U80229 ( n9529, n76037, n5435 );
nand U80230 ( n55973, n76000, n7202 );
nand U80231 ( n55992, n76000, n7203 );
nand U80232 ( n56011, n76000, n7204 );
nand U80233 ( n56030, n75999, n7205 );
nand U80234 ( n56049, n75999, n7207 );
nand U80235 ( n56071, n75999, n7208 );
nand U80236 ( n56090, n75999, n7209 );
nand U80237 ( n56145, n76000, n7213 );
not U80238 ( n504, n42527 );
nor U80239 ( n54292, n49449, n54162 );
buf U80240 ( n76062, n54990 );
nand U80241 ( n30322, n76025, n3684 );
nand U80242 ( n30341, n76025, n3685 );
nand U80243 ( n64441, n75993, n6318 );
nand U80244 ( n9698, n76038, n5444 );
nand U80245 ( n9722, n76038, n5445 );
nand U80246 ( n64460, n75993, n6319 );
nand U80247 ( n43629, n76009, n8099 );
nand U80248 ( n43648, n76009, n8100 );
nand U80249 ( n22993, n76030, n4578 );
nand U80250 ( n23012, n76030, n4579 );
nand U80251 ( n56109, n76001, n7210 );
nand U80252 ( n56128, n76001, n7212 );
not U80253 ( n233, n8448 );
nand U80254 ( n21265, n16567, n14654 );
buf U80255 ( n76797, n2070 );
nor U80256 ( n21309, n16448, n21179 );
nand U80257 ( n64216, n64508, n833 );
nor U80258 ( n64508, n822, n61612 );
not U80259 ( n2073, n38604 );
nand U80260 ( n13650, n76925, n76841 );
and U80261 ( n75759, n13650, n76925 );
nor U80262 ( n26817, n23826, n28336 );
nor U80263 ( n59957, n56950, n61558 );
nor U80264 ( n34062, n31170, n35546 );
nor U80265 ( n68816, n65424, n70274 );
nor U80266 ( n47796, n44495, n49545 );
nor U80267 ( n14544, n10697, n16567 );
not U80268 ( n7924, n42489 );
nand U80269 ( n26906, n4047, n24601 );
nand U80270 ( n60046, n6679, n57733 );
nand U80271 ( n34151, n3217, n31817 );
nand U80272 ( n68905, n5815, n66409 );
nand U80273 ( n76157, n21997, n22002 );
nand U80274 ( n76154, n29316, n29321 );
nand U80275 ( n76082, n63079, n63084 );
nand U80276 ( n76085, n55107, n55112 );
nand U80277 ( n11594, n76619, n11733 );
nand U80278 ( n24530, n76533, n24601 );
nand U80279 ( n66323, n76209, n66409 );
nand U80280 ( n57658, n76275, n57733 );
nand U80281 ( n63789, n5630, n6159 );
nand U80282 ( n63893, n5630, n6157 );
nand U80283 ( n29829, n3029, n3544 );
nand U80284 ( n29937, n3029, n3542 );
nand U80285 ( n22510, n3873, n4382 );
nand U80286 ( n22614, n3873, n4379 );
nand U80287 ( n55623, n6505, n7014 );
nand U80288 ( n55727, n6505, n7012 );
nand U80289 ( n40477, n76920, n76794 );
nand U80290 ( n40471, n76395, n76920 );
nand U80291 ( n45391, n76353, n45509 );
nor U80292 ( n26902, n26904, n26905 );
nor U80293 ( n60042, n60044, n60045 );
nor U80294 ( n34147, n34149, n34150 );
nor U80295 ( n68901, n68903, n68904 );
not U80296 ( n7930, n42809 );
not U80297 ( n784, n54990 );
nand U80298 ( n22036, n4643, n76157 );
nand U80299 ( n55146, n7275, n76085 );
nand U80300 ( n29355, n3749, n76154 );
nand U80301 ( n63118, n6383, n76082 );
nand U80302 ( n32911, n3110, n32851 );
not U80303 ( n3110, n32932 );
nand U80304 ( n67672, n5712, n67616 );
not U80305 ( n5712, n67693 );
nand U80306 ( n25667, n3954, n25611 );
not U80307 ( n3954, n25688 );
nand U80308 ( n58807, n6587, n58748 );
not U80309 ( n6587, n58828 );
nand U80310 ( n13239, n13303, n4829 );
not U80311 ( n4829, n13218 );
not U80312 ( n7934, n42979 );
not U80313 ( n7935, n43033 );
buf U80314 ( n76060, n54990 );
buf U80315 ( n76064, n54990 );
buf U80316 ( n76063, n54990 );
buf U80317 ( n76061, n54990 );
not U80318 ( n175, n21987 );
not U80319 ( n209, n29302 );
not U80320 ( n480, n63069 );
not U80321 ( n447, n55097 );
nand U80322 ( n13095, n4854, n13020 );
not U80323 ( n4854, n13122 );
nand U80324 ( n46625, n7498, n46569 );
not U80325 ( n7498, n46646 );
not U80326 ( n5275, n8764 );
not U80327 ( n7937, n43077 );
not U80328 ( n5629, n63070 );
not U80329 ( n3028, n29303 );
not U80330 ( n3872, n21988 );
not U80331 ( n6504, n55098 );
not U80332 ( n483, n63084 );
not U80333 ( n212, n29321 );
not U80334 ( n178, n22002 );
not U80335 ( n449, n55112 );
buf U80336 ( n76065, n54990 );
not U80337 ( n7938, n43129 );
nand U80338 ( n30427, n30577, n3167 );
nand U80339 ( n64586, n64736, n5765 );
not U80340 ( n6147, n63617 );
not U80341 ( n6148, n63732 );
not U80342 ( n6149, n63776 );
not U80343 ( n6150, n63828 );
not U80344 ( n3532, n29718 );
not U80345 ( n3533, n29772 );
not U80346 ( n3534, n29816 );
not U80347 ( n3535, n29872 );
not U80348 ( n3537, n29932 );
not U80349 ( n4372, n22497 );
not U80350 ( n4369, n22397 );
not U80351 ( n4370, n22451 );
not U80352 ( n4373, n22549 );
not U80353 ( n4374, n22609 );
not U80354 ( n7004, n55610 );
not U80355 ( n7002, n55509 );
not U80356 ( n7003, n55566 );
not U80357 ( n7005, n55662 );
not U80358 ( n7007, n55722 );
nor U80359 ( n13890, n13779, n4855 );
not U80360 ( n6152, n63888 );
nor U80361 ( n47268, n47171, n7500 );
nor U80362 ( n31606, n3237, n76486 );
not U80363 ( n3237, n31607 );
nor U80364 ( n65892, n5837, n76219 );
not U80365 ( n5837, n65893 );
nor U80366 ( n31118, n3246, n76487 );
not U80367 ( n3246, n30254 );
nor U80368 ( n65372, n5847, n76220 );
not U80369 ( n5847, n64316 );
not U80370 ( n5279, n8959 );
not U80371 ( n5280, n9027 );
nand U80372 ( n16442, n4795, n1 );
nor U80373 ( n31065, n3239, n76487 );
not U80374 ( n3239, n30245 );
nor U80375 ( n30852, n3180, n76487 );
not U80376 ( n3180, n30193 );
nor U80377 ( n30895, n3189, n76487 );
not U80378 ( n3189, n30207 );
nor U80379 ( n30937, n3200, n76487 );
not U80380 ( n3200, n30216 );
nor U80381 ( n65054, n5779, n76220 );
not U80382 ( n5779, n64259 );
nor U80383 ( n65097, n5788, n76220 );
not U80384 ( n5788, n64269 );
nor U80385 ( n65139, n5799, n76220 );
not U80386 ( n5799, n64278 );
nor U80387 ( n65182, n5812, n76220 );
not U80388 ( n5812, n64288 );
nor U80389 ( n65224, n5825, n76220 );
not U80390 ( n5825, n64297 );
nor U80391 ( n30980, n3213, n76487 );
not U80392 ( n3213, n30226 );
nor U80393 ( n31022, n3227, n76487 );
not U80394 ( n3227, n30235 );
nor U80395 ( n65267, n5839, n76220 );
not U80396 ( n5839, n64307 );
nor U80397 ( n30417, n30122, n76488 );
nor U80398 ( n64576, n64135, n76221 );
not U80399 ( n7939, n43189 );
nand U80400 ( n9827, n9965, n4903 );
nand U80401 ( n43743, n43889, n7552 );
nand U80402 ( n33137, n33164, n33095 );
nand U80403 ( n67893, n67915, n67851 );
nand U80404 ( n25890, n25912, n25848 );
nand U80405 ( n59028, n59050, n58986 );
nor U80406 ( n31179, n3163, n76487 );
not U80407 ( n3163, n30264 );
nor U80408 ( n31237, n3179, n76487 );
not U80409 ( n3179, n30273 );
nor U80410 ( n31281, n3188, n76487 );
not U80411 ( n3188, n30283 );
nor U80412 ( n31322, n3199, n76487 );
not U80413 ( n3199, n30292 );
nor U80414 ( n31362, n3212, n76486 );
not U80415 ( n3212, n30306 );
nor U80416 ( n65491, n5778, n76220 );
not U80417 ( n5778, n64396 );
nor U80418 ( n65531, n5787, n76220 );
not U80419 ( n5787, n64406 );
nor U80420 ( n65572, n5798, n76220 );
not U80421 ( n5798, n64415 );
nor U80422 ( n65612, n5810, n76219 );
not U80423 ( n5810, n64425 );
nor U80424 ( n65433, n5762, n76220 );
not U80425 ( n5762, n64326 );
nor U80426 ( n31403, n3225, n76486 );
not U80427 ( n3225, n30315 );
nor U80428 ( n31443, n3238, n76486 );
not U80429 ( n3238, n30325 );
nor U80430 ( n31484, n3245, n76486 );
not U80431 ( n3245, n30334 );
nor U80432 ( n65653, n5824, n76219 );
not U80433 ( n5824, n64434 );
nor U80434 ( n65693, n5838, n76219 );
not U80435 ( n5838, n64444 );
nor U80436 ( n65734, n5845, n76219 );
not U80437 ( n5845, n64453 );
nor U80438 ( n11303, n4970, n76630 );
not U80439 ( n4970, n11304 );
nor U80440 ( n44984, n7624, n76360 );
not U80441 ( n7624, n44985 );
nor U80442 ( n10699, n4980, n76631 );
not U80443 ( n4980, n9614 );
nand U80444 ( n14657, n5132, n10697 );
nand U80445 ( n12938, n12990, n12879 );
not U80446 ( n5282, n9082 );
nor U80447 ( n10853, n4915, n76631 );
not U80448 ( n4915, n9638 );
nor U80449 ( n10903, n4922, n76631 );
not U80450 ( n4922, n9654 );
nor U80451 ( n10954, n4932, n76631 );
not U80452 ( n4932, n9665 );
nor U80453 ( n11003, n4944, n76630 );
not U80454 ( n4944, n9678 );
nor U80455 ( n11053, n4958, n76630 );
not U80456 ( n4958, n9689 );
nor U80457 ( n11104, n4972, n76630 );
not U80458 ( n4972, n9702 );
nor U80459 ( n11153, n4979, n76630 );
not U80460 ( n4979, n9713 );
nor U80461 ( n44655, n7574, n76361 );
not U80462 ( n7574, n43594 );
nor U80463 ( n44696, n7585, n76361 );
not U80464 ( n7585, n43603 );
nor U80465 ( n44735, n7598, n76360 );
not U80466 ( n7598, n43613 );
nor U80467 ( n44775, n7612, n76360 );
not U80468 ( n7612, n43622 );
nor U80469 ( n44869, n7633, n76360 );
not U80470 ( n7633, n43641 );
nor U80471 ( n44816, n7625, n76360 );
not U80472 ( n7625, n43632 );
nor U80473 ( n44615, n7565, n76361 );
not U80474 ( n7565, n43584 );
nor U80475 ( n10782, n4900, n76631 );
not U80476 ( n4900, n9627 );
nor U80477 ( n44558, n7548, n76361 );
not U80478 ( n7548, n43575 );
not U80479 ( n482, n63079 );
not U80480 ( n210, n29316 );
not U80481 ( n177, n21997 );
not U80482 ( n448, n55107 );
nor U80483 ( n33181, n33142, n3123 );
nand U80484 ( n13385, n13419, n13333 );
nor U80485 ( n67932, n67898, n5723 );
nor U80486 ( n46885, n46851, n7509 );
nor U80487 ( n25929, n25895, n3965 );
nor U80488 ( n59067, n59033, n6598 );
nand U80489 ( n46846, n46868, n46804 );
nor U80490 ( n13215, n13122, n13218 );
nand U80491 ( n67774, n67827, n5688 );
not U80492 ( n5688, n67757 );
nand U80493 ( n46727, n46780, n7473 );
not U80494 ( n7473, n46710 );
nand U80495 ( n25771, n25824, n3930 );
not U80496 ( n3930, n25752 );
nand U80497 ( n58909, n58962, n6563 );
not U80498 ( n6563, n58892 );
nand U80499 ( n33018, n33071, n3087 );
not U80500 ( n3087, n33001 );
nor U80501 ( n32999, n32932, n33001 );
nor U80502 ( n67755, n67693, n67757 );
nor U80503 ( n25750, n25688, n25752 );
nor U80504 ( n58890, n58828, n58892 );
buf U80505 ( n76066, n61173 );
not U80506 ( n5283, n9147 );
nand U80507 ( n47886, n7787, n44495 );
nor U80508 ( n13440, n13392, n4864 );
nor U80509 ( n46708, n46646, n46710 );
not U80510 ( n508, n42517 );
not U80511 ( n5284, n9222 );
nand U80512 ( n67965, n67969, n67913 );
and U80513 ( n67969, n67915, n67970 );
nand U80514 ( n33210, n33214, n33159 );
and U80515 ( n33214, n33164, n33215 );
nand U80516 ( n25962, n25966, n25910 );
and U80517 ( n25966, n25912, n25967 );
nand U80518 ( n59100, n59104, n59048 );
and U80519 ( n59104, n59050, n59105 );
nand U80520 ( n42577, n8164, n76102 );
not U80521 ( n237, n8435 );
buf U80522 ( n76861, n512 );
buf U80523 ( n76888, n240 );
buf U80524 ( n76859, n512 );
buf U80525 ( n76860, n512 );
buf U80526 ( n76886, n240 );
buf U80527 ( n76887, n240 );
nand U80528 ( n68449, n67159, n76708 );
nand U80529 ( n47428, n46195, n76660 );
nand U80530 ( n26448, n25261, n76754 );
nand U80531 ( n59587, n58397, n76687 );
nand U80532 ( n33693, n32503, n76774 );
nand U80533 ( n14076, n12564, n76727 );
nand U80534 ( n8509, n5510, n76172 );
not U80535 ( n3118, n33448 );
not U80536 ( n5719, n68199 );
not U80537 ( n7505, n47168 );
not U80538 ( n3962, n26198 );
not U80539 ( n6594, n59337 );
nand U80540 ( n13477, n13482, n13413 );
and U80541 ( n13482, n13419, n13483 );
nand U80542 ( n46918, n46922, n46866 );
and U80543 ( n46922, n46868, n46923 );
not U80544 ( n4859, n13775 );
nand U80545 ( n46488, n46517, n46431 );
or U80546 ( n46487, n46488, n46388 );
or U80547 ( n25545, n25546, n25447 );
or U80548 ( n32785, n32786, n32687 );
or U80549 ( n67550, n67551, n67452 );
or U80550 ( n58682, n58683, n58584 );
not U80551 ( n5700, n64120 );
not U80552 ( n6575, n55896 );
not U80553 ( n3943, n22782 );
nand U80554 ( n32604, n32588, n32573 );
not U80555 ( n7393, n42500 );
not U80556 ( n7487, n43376 );
not U80557 ( n4751, n8414 );
nand U80558 ( n67369, n67353, n67338 );
nand U80559 ( n25364, n25346, n25331 );
nand U80560 ( n58501, n58485, n58470 );
nor U80561 ( n9395, n4762, n8448 );
not U80562 ( n4844, n9437 );
nand U80563 ( n12887, n12679, n12660 );
not U80564 ( n5168, n18701 );
not U80565 ( n5178, n14734 );
not U80566 ( n5184, n15613 );
nand U80567 ( n46453, n46292, n46277 );
nand U80568 ( n48719, n7833, n47948 );
not U80569 ( n7833, n48240 );
not U80570 ( n7839, n48722 );
nand U80571 ( n22798, n3919, n23077 );
nand U80572 ( n55912, n6552, n56198 );
not U80573 ( n163, n23162 );
and U80574 ( n23825, n23256, n23077 );
and U80575 ( n23819, n23825, n23826 );
not U80576 ( n435, n56283 );
and U80577 ( n56949, n56380, n56198 );
and U80578 ( n56944, n56949, n56950 );
buf U80579 ( n76071, n61173 );
not U80580 ( n5632, n64078 );
not U80581 ( n3030, n30061 );
not U80582 ( n3874, n22738 );
not U80583 ( n6507, n55854 );
nand U80584 ( n64061, n5632, n6015 );
nand U80585 ( n30044, n3030, n3400 );
nand U80586 ( n22721, n3874, n4238 );
nand U80587 ( n55837, n6507, n6870 );
nand U80588 ( n56217, n56380, n6639 );
nand U80589 ( n23096, n23256, n4007 );
nor U80590 ( n15917, n5178, n15062 );
nand U80591 ( n68011, n68044, n67970 );
nand U80592 ( n46976, n47009, n46923 );
nand U80593 ( n26008, n26041, n25967 );
nand U80594 ( n13534, n13575, n13483 );
nand U80595 ( n59146, n59182, n59105 );
nand U80596 ( n33252, n33285, n33215 );
not U80597 ( n5720, n68098 );
not U80598 ( n3119, n33341 );
not U80599 ( n7507, n47067 );
not U80600 ( n3963, n26095 );
not U80601 ( n6595, n59236 );
nor U80602 ( n15812, n5178, n5205 );
nor U80603 ( n48884, n7833, n7859 );
not U80604 ( n4835, n13632 );
not U80605 ( n4834, n13758 );
not U80606 ( n4833, n13939 );
and U80607 ( n57433, n57434, n437 );
and U80608 ( n24310, n24311, n164 );
and U80609 ( n24109, n22986, n164 );
and U80610 ( n24190, n23005, n164 );
and U80611 ( n23987, n22956, n164 );
and U80612 ( n24028, n22967, n164 );
and U80613 ( n24068, n22977, n164 );
and U80614 ( n57069, n56064, n437 );
and U80615 ( n57109, n56074, n437 );
and U80616 ( n57150, n56083, n437 );
and U80617 ( n57190, n56093, n437 );
and U80618 ( n23947, n22946, n164 );
and U80619 ( n57231, n56102, n437 );
and U80620 ( n57271, n56112, n437 );
and U80621 ( n57312, n56121, n437 );
and U80622 ( n24149, n22996, n164 );
not U80623 ( n5715, n68511 );
not U80624 ( n3114, n33755 );
not U80625 ( n4857, n14153 );
not U80626 ( n7502, n47490 );
not U80627 ( n3958, n26510 );
not U80628 ( n6590, n59649 );
and U80629 ( n23820, n22927, n164 );
and U80630 ( n56945, n56042, n437 );
nand U80631 ( n46430, n46389, n46431 );
not U80632 ( n4860, n13642 );
buf U80633 ( n76769, n3823 );
buf U80634 ( n76770, n3823 );
buf U80635 ( n76067, n61173 );
buf U80636 ( n76068, n61173 );
buf U80637 ( n76069, n61173 );
buf U80638 ( n76771, n3823 );
buf U80639 ( n76070, n61173 );
buf U80640 ( n76721, n5580 );
buf U80641 ( n76702, n6455 );
buf U80642 ( n76722, n5580 );
buf U80643 ( n76703, n6455 );
buf U80644 ( n76704, n6455 );
buf U80645 ( n76723, n5580 );
buf U80646 ( n76072, n61173 );
buf U80647 ( n76073, n61173 );
not U80648 ( n5692, n68185 );
not U80649 ( n7477, n47154 );
not U80650 ( n3934, n26184 );
not U80651 ( n6567, n59323 );
not U80652 ( n3090, n33438 );
buf U80653 ( n76679, n7344 );
buf U80654 ( n76680, n7344 );
not U80655 ( n4268, n26969 );
not U80656 ( n6900, n60109 );
not U80657 ( n4274, n27642 );
not U80658 ( n6907, n60795 );
not U80659 ( n3430, n34214 );
not U80660 ( n6045, n68968 );
not U80661 ( n3437, n34887 );
not U80662 ( n6052, n69629 );
buf U80663 ( n76748, n4712 );
not U80664 ( n7408, n43332 );
buf U80665 ( n76747, n4712 );
buf U80666 ( n76746, n4712 );
buf U80667 ( n76681, n7344 );
nand U80668 ( n43315, n7408, n7803 );
nand U80669 ( n47885, n7603, n45509 );
nand U80670 ( n14655, n4949, n11733 );
nor U80671 ( n27792, n4268, n4292 );
nor U80672 ( n60940, n6900, n6924 );
nor U80673 ( n35033, n3430, n3454 );
nor U80674 ( n69771, n6045, n6069 );
not U80675 ( n4763, n9383 );
nand U80676 ( n9362, n4763, n5148 );
nor U80677 ( n27874, n4268, n27213 );
nor U80678 ( n61021, n6900, n60358 );
nor U80679 ( n69849, n6045, n69208 );
nor U80680 ( n35113, n3430, n34458 );
not U80681 ( n7834, n49158 );
nand U80682 ( n33494, n32664, n33451 );
nand U80683 ( n13829, n12775, n13779 );
nand U80684 ( n68249, n67429, n68202 );
nand U80685 ( n47218, n46365, n47171 );
nand U80686 ( n26248, n25424, n26201 );
nand U80687 ( n59387, n58561, n59340 );
nor U80688 ( n48141, n7859, n48240 );
nor U80689 ( n48882, n7857, n7838 );
not U80690 ( n7838, n48418 );
and U80691 ( n31116, n30577, n30408 );
and U80692 ( n65370, n64736, n64567 );
nand U80693 ( n27052, n28289, n24601 );
nand U80694 ( n27128, n28289, n23077 );
nand U80695 ( n27074, n28289, n28336 );
nand U80696 ( n27085, n28289, n26903 );
nand U80697 ( n27063, n28289, n26905 );
nand U80698 ( n27096, n28289, n26918 );
nand U80699 ( n60240, n61511, n60058 );
nand U80700 ( n60215, n61511, n61558 );
nand U80701 ( n60204, n61511, n60045 );
nand U80702 ( n60226, n61511, n60043 );
nand U80703 ( n60193, n61511, n57733 );
nand U80704 ( n60272, n61511, n56198 );
nand U80705 ( n34340, n35517, n34163 );
nand U80706 ( n34351, n35517, n31170 );
nand U80707 ( n34318, n35517, n35546 );
nand U80708 ( n34307, n35517, n34150 );
nand U80709 ( n69059, n70245, n68904 );
nand U80710 ( n69070, n70245, n70274 );
nand U80711 ( n69103, n70245, n65424 );
nand U80712 ( n69092, n70245, n68917 );
nand U80713 ( n34296, n35517, n31817 );
nand U80714 ( n34372, n35517, n30408 );
nand U80715 ( n34329, n35517, n34148 );
nand U80716 ( n69048, n70245, n66409 );
nand U80717 ( n69124, n70245, n64567 );
nand U80718 ( n69081, n70245, n68902 );
nor U80719 ( n15809, n5202, n5183 );
not U80720 ( n5183, n14728 );
nand U80721 ( n30480, n31116, n31170 );
nand U80722 ( n64639, n65370, n65424 );
nor U80723 ( n14957, n5205, n14734 );
and U80724 ( n10695, n9965, n9804 );
and U80725 ( n44494, n43889, n43725 );
not U80726 ( n3099, n30103 );
nand U80727 ( n14209, n4848, n12574 );
not U80728 ( n4937, n14215 );
nand U80729 ( n60100, n60101, n60102 );
nand U80730 ( n60101, n6512, n60106 );
nand U80731 ( n60102, n60103, n60104 );
nand U80732 ( n60106, n6902, n60107 );
nand U80733 ( n26960, n26961, n26962 );
nand U80734 ( n26961, n3879, n26966 );
nand U80735 ( n26962, n26963, n26964 );
nand U80736 ( n26966, n4269, n26967 );
nand U80737 ( n34205, n34206, n34207 );
nand U80738 ( n34206, n3035, n34211 );
nand U80739 ( n34207, n34208, n34209 );
nand U80740 ( n34211, n3432, n34212 );
nand U80741 ( n68959, n68960, n68961 );
nand U80742 ( n68960, n5637, n68965 );
nand U80743 ( n68961, n68962, n68963 );
nand U80744 ( n68965, n6047, n68966 );
nand U80745 ( n13152, n5218, n12732 );
nand U80746 ( n68556, n5704, n67167 );
nand U80747 ( n47535, n7490, n46203 );
nand U80748 ( n26555, n3947, n25269 );
nand U80749 ( n59697, n6579, n58405 );
not U80750 ( n5803, n68561 );
not U80751 ( n4037, n26560 );
not U80752 ( n6669, n59702 );
not U80753 ( n7590, n47540 );
nand U80754 ( n33800, n3103, n32511 );
not U80755 ( n3204, n33805 );
nand U80756 ( n67850, n67851, n67827 );
nand U80757 ( n33094, n33095, n33071 );
nand U80758 ( n46803, n46804, n46780 );
nand U80759 ( n25847, n25848, n25824 );
nand U80760 ( n58985, n58986, n58962 );
nand U80761 ( n13332, n13333, n13303 );
nand U80762 ( n67615, n67616, n67578 );
nand U80763 ( n32850, n32851, n32813 );
nand U80764 ( n46568, n46569, n46517 );
nand U80765 ( n25610, n25611, n25573 );
nand U80766 ( n13019, n13020, n12990 );
nand U80767 ( n58747, n58748, n58710 );
nand U80768 ( n46663, n7872, n46331 );
nand U80769 ( n67710, n6082, n67395 );
nand U80770 ( n25705, n4304, n25390 );
nand U80771 ( n58845, n6937, n58527 );
nand U80772 ( n32956, n3467, n32630 );
nand U80773 ( n13003, n5217, n12732 );
nor U80774 ( n28163, n27085, n28128 );
nor U80775 ( n61327, n60226, n61283 );
nor U80776 ( n28135, n27052, n28128 );
nor U80777 ( n28194, n27128, n28128 );
nor U80778 ( n28171, n27096, n28128 );
nor U80779 ( n61335, n60240, n61283 );
nor U80780 ( n61303, n60193, n61283 );
nor U80781 ( n61358, n60272, n61283 );
nor U80782 ( n28151, n27074, n28128 );
nor U80783 ( n28143, n27063, n28128 );
nor U80784 ( n61319, n60215, n61283 );
nor U80785 ( n61311, n60204, n61283 );
nand U80786 ( n27039, n28289, n28290 );
nand U80787 ( n60180, n61511, n61512 );
nand U80788 ( n60251, n61511, n56950 );
nand U80789 ( n27107, n28289, n23826 );
nand U80790 ( n49462, n47948, n48240 );
nor U80791 ( n35394, n34329, n35363 );
nor U80792 ( n70126, n69081, n70095 );
nor U80793 ( n35370, n34296, n35363 );
nor U80794 ( n35404, n34340, n35363 );
nor U80795 ( n35412, n34351, n35363 );
nor U80796 ( n35427, n34372, n35363 );
nor U80797 ( n70102, n69048, n70095 );
nor U80798 ( n70142, n69103, n70095 );
nor U80799 ( n70157, n69124, n70095 );
nor U80800 ( n70134, n69092, n70095 );
nor U80801 ( n35386, n34318, n35363 );
nor U80802 ( n35378, n34307, n35363 );
nor U80803 ( n70110, n69059, n70095 );
nor U80804 ( n70118, n69070, n70095 );
nand U80805 ( n34283, n35517, n35518 );
nand U80806 ( n69035, n70245, n70246 );
nor U80807 ( n47881, n47883, n47884 );
nor U80808 ( n14650, n14653, n14654 );
nand U80809 ( n13413, n13392, n12732 );
nand U80810 ( n33159, n33142, n32630 );
nand U80811 ( n46866, n46851, n46331 );
nand U80812 ( n67913, n67898, n67395 );
nand U80813 ( n25910, n25895, n25390 );
nand U80814 ( n59048, n59033, n58527 );
nand U80815 ( n67634, n6080, n67395 );
nand U80816 ( n25629, n4303, n25390 );
nand U80817 ( n58766, n6935, n58527 );
nand U80818 ( n32873, n3465, n32630 );
not U80819 ( n7855, n47935 );
nor U80820 ( n28125, n27039, n28128 );
nor U80821 ( n61343, n60251, n61283 );
nor U80822 ( n61280, n60180, n61283 );
nor U80823 ( n28179, n27107, n28128 );
and U80824 ( n43797, n44494, n44495 );
and U80825 ( n9894, n10695, n10697 );
and U80826 ( n46589, n7870, n46331 );
nand U80827 ( n14307, n4848, n12595 );
nand U80828 ( n68634, n5704, n67184 );
nand U80829 ( n26633, n3947, n25286 );
nand U80830 ( n59775, n6579, n58422 );
nand U80831 ( n47613, n7490, n46232 );
nand U80832 ( n33878, n3103, n32528 );
nor U80833 ( n23086, n22797, n23096 );
nor U80834 ( n56207, n55911, n56217 );
not U80835 ( n4868, n13217 );
nor U80836 ( n27788, n4288, n4273 );
nor U80837 ( n60936, n6920, n6905 );
not U80838 ( n4273, n26964 );
not U80839 ( n6905, n60104 );
nor U80840 ( n35029, n3450, n3435 );
nor U80841 ( n69767, n6065, n6050 );
not U80842 ( n3435, n34209 );
not U80843 ( n6050, n68963 );
not U80844 ( n4870, n12993 );
not U80845 ( n3127, n33000 );
not U80846 ( n5728, n67756 );
not U80847 ( n3970, n25751 );
not U80848 ( n6603, n58891 );
not U80849 ( n7514, n46709 );
not U80850 ( n7515, n46570 );
not U80851 ( n5730, n67617 );
not U80852 ( n3129, n32852 );
not U80853 ( n3973, n25612 );
not U80854 ( n6605, n58749 );
nand U80855 ( n31756, n217, n31817 );
not U80856 ( n217, n31725 );
nor U80857 ( n34370, n3454, n34214 );
nor U80858 ( n69122, n6069, n68968 );
nor U80859 ( n27126, n4292, n26969 );
nor U80860 ( n60270, n6924, n60109 );
nand U80861 ( n12895, n12948, n12949 );
nand U80862 ( n12948, n5215, n9812 );
nand U80863 ( n12949, n5215, n12777 );
nor U80864 ( n47946, n47947, n7832 );
nor U80865 ( n47947, n7833, n47948 );
and U80866 ( n46361, n46352, n43731 );
not U80867 ( n76150, n76143 );
not U80868 ( n76147, n76142 );
not U80869 ( n76148, n76143 );
not U80870 ( n76146, n76142 );
not U80871 ( n76149, n76143 );
not U80872 ( n76152, n76144 );
not U80873 ( n76151, n76144 );
not U80874 ( n76145, n76142 );
not U80875 ( n76153, n76143 );
nand U80876 ( n30123, n3075, n30408 );
nand U80877 ( n43392, n7462, n43725 );
nand U80878 ( n64136, n5677, n64567 );
nand U80879 ( n9457, n4818, n9804 );
nand U80880 ( n44192, n44531, n7810 );
nand U80881 ( n10335, n10742, n5155 );
nand U80882 ( n30832, n31152, n3408 );
nand U80883 ( n65034, n65406, n6023 );
nand U80884 ( n30670, n30745, n30746 );
nand U80885 ( n10134, n10230, n10232 );
nand U80886 ( n64876, n64951, n64952 );
nand U80887 ( n44031, n44108, n44109 );
nand U80888 ( n30581, n30656, n30657 );
nand U80889 ( n10024, n10109, n10110 );
nand U80890 ( n64740, n64862, n64863 );
nand U80891 ( n43940, n44015, n44016 );
nand U80892 ( n30491, n30566, n30567 );
nand U80893 ( n9912, n10011, n10012 );
nand U80894 ( n64650, n64725, n64726 );
nand U80895 ( n43811, n43927, n43928 );
nor U80896 ( n30656, n30670, n30671 );
nor U80897 ( n10109, n10134, n10135 );
nor U80898 ( n64862, n64876, n64877 );
nor U80899 ( n44015, n44031, n44032 );
nor U80900 ( n30566, n30581, n30582 );
nor U80901 ( n10011, n10024, n10025 );
nor U80902 ( n64725, n64740, n64741 );
nor U80903 ( n43927, n43940, n43941 );
nor U80904 ( n30476, n30491, n30492 );
nor U80905 ( n9888, n9912, n9913 );
nor U80906 ( n64635, n64650, n64651 );
nor U80907 ( n43792, n43811, n43812 );
nand U80908 ( n23525, n23860, n4245 );
nand U80909 ( n56647, n56984, n6878 );
nand U80910 ( n23260, n23342, n23343 );
nand U80911 ( n56384, n56466, n56467 );
nand U80912 ( n23167, n23246, n23247 );
nand U80913 ( n56288, n56367, n56368 );
nand U80914 ( n23359, n23435, n23436 );
nand U80915 ( n56483, n56557, n56558 );
nor U80916 ( n23246, n23260, n23261 );
nor U80917 ( n56367, n56384, n56385 );
nor U80918 ( n23145, n23167, n23168 );
nor U80919 ( n56266, n56288, n56289 );
nor U80920 ( n23342, n23359, n23360 );
nor U80921 ( n56466, n56483, n56484 );
nand U80922 ( n44197, n44531, n7808 );
nand U80923 ( n10342, n10742, n5153 );
nand U80924 ( n30837, n31152, n3405 );
nand U80925 ( n65039, n65406, n6020 );
nand U80926 ( n23530, n23860, n4243 );
nand U80927 ( n56652, n56984, n6875 );
not U80928 ( n5200, n15062 );
xor U80929 ( n22804, n23146, n23145 );
xor U80930 ( n55918, n56267, n56266 );
nand U80931 ( n67511, n67559, n67560 );
nand U80932 ( n67559, n6079, n67413 );
nand U80933 ( n67560, n6079, n64573 );
nand U80934 ( n32746, n32794, n32795 );
nand U80935 ( n32794, n3464, n32648 );
nand U80936 ( n32795, n3464, n30414 );
nand U80937 ( n46447, n46496, n46497 );
nand U80938 ( n46496, n7869, n46349 );
nand U80939 ( n46497, n7869, n43731 );
nand U80940 ( n25506, n25554, n25555 );
nand U80941 ( n25554, n4302, n25408 );
nand U80942 ( n25555, n4302, n23083 );
nand U80943 ( n58643, n58691, n58692 );
nand U80944 ( n58691, n6934, n58545 );
nand U80945 ( n58692, n6934, n56204 );
xnor U80946 ( n30129, n30477, n30476 );
xnor U80947 ( n64142, n64636, n64635 );
xnor U80948 ( n43398, n43793, n43792 );
xnor U80949 ( n9464, n9889, n9888 );
and U80950 ( n25420, n25411, n23083 );
and U80951 ( n58557, n58548, n56204 );
and U80952 ( n32660, n32651, n30414 );
and U80953 ( n67425, n67416, n64573 );
nand U80954 ( n14548, n4977, n14482 );
not U80955 ( n4287, n27213 );
not U80956 ( n6919, n60358 );
not U80957 ( n6064, n69208 );
not U80958 ( n3449, n34458 );
xor U80959 ( n22814, n23167, n23168 );
xor U80960 ( n55928, n56288, n56289 );
nand U80961 ( n26820, n4068, n26768 );
nand U80962 ( n59960, n6700, n59908 );
nand U80963 ( n47799, n7630, n47746 );
nand U80964 ( n34065, n3243, n34011 );
nand U80965 ( n68819, n5843, n68767 );
xnor U80966 ( n30139, n30491, n30492 );
xnor U80967 ( n64152, n64650, n64651 );
xnor U80968 ( n43408, n43811, n43812 );
xnor U80969 ( n9477, n9912, n9913 );
not U80970 ( n5179, n15679 );
nor U80971 ( n48138, n48418, n7857 );
nor U80972 ( n14953, n14728, n5202 );
xnor U80973 ( n22822, n23247, n23246 );
xnor U80974 ( n55936, n56368, n56367 );
xnor U80975 ( n30147, n30567, n30566 );
xnor U80976 ( n64160, n64726, n64725 );
xnor U80977 ( n43416, n43928, n43927 );
xnor U80978 ( n9487, n10012, n10011 );
not U80979 ( n4269, n27705 );
not U80980 ( n3432, n34950 );
not U80981 ( n6047, n69690 );
not U80982 ( n6902, n60856 );
nor U80983 ( n54137, n46407, n43356 );
nor U80984 ( n35639, n32706, n30083 );
nor U80985 ( n28460, n25466, n22762 );
nor U80986 ( n21154, n12835, n9412 );
nor U80987 ( n70365, n67471, n64100 );
nor U80988 ( n61765, n58603, n55876 );
xor U80989 ( n22830, n23260, n23261 );
xor U80990 ( n55944, n56384, n56385 );
not U80991 ( n4978, n14410 );
not U80992 ( n7632, n47682 );
not U80993 ( n3244, n33947 );
not U80994 ( n5844, n68703 );
not U80995 ( n6702, n59844 );
not U80996 ( n4069, n26702 );
xnor U80997 ( n30155, n30581, n30582 );
xnor U80998 ( n64168, n64740, n64741 );
xnor U80999 ( n43457, n43940, n43941 );
xnor U81000 ( n9497, n10024, n10025 );
nor U81001 ( n27136, n26964, n4288 );
nor U81002 ( n60280, n60104, n6920 );
nor U81003 ( n34381, n34209, n3450 );
nor U81004 ( n69133, n68963, n6065 );
xor U81005 ( n55957, n56467, n56466 );
xor U81006 ( n22840, n23343, n23342 );
xnor U81007 ( n30165, n30657, n30656 );
xnor U81008 ( n64178, n64863, n64862 );
xnor U81009 ( n43467, n44016, n44015 );
xnor U81010 ( n9509, n10110, n10109 );
not U81011 ( n76496, n76498 );
not U81012 ( n76639, n76641 );
not U81013 ( n76367, n76369 );
not U81014 ( n76549, n76551 );
xnor U81015 ( n55966, n56483, n56484 );
xnor U81016 ( n22849, n23359, n23360 );
not U81017 ( n76229, n76231 );
xnor U81018 ( n30174, n30670, n30671 );
xnor U81019 ( n64240, n64876, n64877 );
xnor U81020 ( n43476, n44031, n44032 );
xnor U81021 ( n9520, n10134, n10135 );
not U81022 ( n76295, n76297 );
xor U81023 ( n22859, n23436, n23435 );
xor U81024 ( n55976, n56558, n56557 );
xnor U81025 ( n30184, n30746, n30745 );
xnor U81026 ( n64250, n64952, n64951 );
xnor U81027 ( n43486, n44109, n44108 );
xnor U81028 ( n9533, n10232, n10230 );
not U81029 ( n76497, n76498 );
not U81030 ( n76640, n76641 );
not U81031 ( n76368, n76369 );
not U81032 ( n76550, n76551 );
nand U81033 ( n48122, n49448, n43725 );
nand U81034 ( n14934, n16447, n9804 );
not U81035 ( n76230, n76231 );
not U81036 ( n76296, n76297 );
nor U81037 ( n16329, n14934, n16237 );
not U81038 ( n7634, n43565 );
not U81039 ( n4945, n9580 );
not U81040 ( n4959, n9590 );
not U81041 ( n4923, n9557 );
not U81042 ( n4916, n9544 );
not U81043 ( n7599, n43524 );
not U81044 ( n7613, n43533 );
not U81045 ( n7567, n43495 );
not U81046 ( n7575, n43505 );
not U81047 ( n7627, n43543 );
not U81048 ( n4973, n9603 );
not U81049 ( n4933, n9568 );
not U81050 ( n7587, n43514 );
nand U81051 ( n14854, n16447, n14654 );
nand U81052 ( n48051, n49448, n47884 );
nand U81053 ( n16158, n5197, n4756 );
nand U81054 ( n49197, n7852, n7400 );
nand U81055 ( n14868, n16447, n16567 );
nand U81056 ( n48062, n49448, n49545 );
nand U81057 ( n16168, n5197, n4755 );
nand U81058 ( n49205, n7852, n7399 );
nand U81059 ( n14840, n16447, n11733 );
nand U81060 ( n48040, n49448, n45509 );
nand U81061 ( n16148, n5197, n4757 );
nand U81062 ( n49189, n7852, n7402 );
nand U81063 ( n48087, n49448, n47882 );
nand U81064 ( n14882, n16447, n14652 );
nand U81065 ( n16178, n5197, n4754 );
nand U81066 ( n49213, n7852, n7398 );
nand U81067 ( n14895, n16447, n14670 );
nand U81068 ( n48098, n49448, n47897 );
nand U81069 ( n16188, n5197, n4753 );
nand U81070 ( n49221, n7852, n7397 );
nand U81071 ( n14824, n16447, n16448 );
nand U81072 ( n48027, n49448, n49449 );
nand U81073 ( n16127, n5197, n4758 );
nand U81074 ( n49177, n7852, n7403 );
nand U81075 ( n14909, n16447, n10697 );
nand U81076 ( n48109, n49448, n44495 );
nand U81077 ( n49229, n7852, n7395 );
nand U81078 ( n16198, n5197, n4752 );
or U81079 ( n48779, n7849, n48784 );
or U81080 ( n15692, n5194, n15698 );
nand U81081 ( n48433, n48140, n7847 );
or U81082 ( n34948, n3447, n34951 );
or U81083 ( n69688, n6062, n69691 );
or U81084 ( n27703, n4284, n27706 );
or U81085 ( n60854, n6917, n60857 );
not U81086 ( n6515, n60090 );
not U81087 ( n3883, n26950 );
not U81088 ( n3039, n34195 );
not U81089 ( n5640, n68949 );
not U81090 ( n7439, n49648 );
not U81091 ( n7443, n49152 );
not U81092 ( n7447, n48769 );
not U81093 ( n4803, n15678 );
not U81094 ( n4805, n15470 );
not U81095 ( n4804, n15577 );
not U81096 ( n4799, n16098 );
not U81097 ( n4800, n15990 );
not U81098 ( n4802, n15892 );
not U81099 ( n7449, n48598 );
not U81100 ( n5195, n18709 );
not U81101 ( n7850, n51665 );
not U81102 ( n7445, n48963 );
not U81103 ( n7448, n48692 );
not U81104 ( n7444, n49058 );
not U81105 ( n7442, n49327 );
nand U81106 ( n60089, n6920, n60090 );
nand U81107 ( n26949, n4288, n26950 );
nand U81108 ( n34194, n3450, n34195 );
nand U81109 ( n68948, n6065, n68949 );
not U81110 ( n4795, n16677 );
not U81111 ( n4798, n16309 );
not U81112 ( n4797, n16412 );
not U81113 ( n7440, n49420 );
not U81114 ( n7415, n47930 );
not U81115 ( n4772, n14710 );
not U81116 ( n7354, n42409 );
not U81117 ( n3833, n21883 );
not U81118 ( n4720, n8328 );
not U81119 ( n6465, n54974 );
not U81120 ( n2989, n29200 );
not U81121 ( n5590, n62918 );
xor U81122 ( n50018, n50080, n50009 );
xor U81123 ( n50080, n50010, n1452 );
xor U81124 ( n49742, n50088, n49756 );
xor U81125 ( n50088, n49755, n1507 );
xnor U81126 ( n50070, n50078, n50025 );
xor U81127 ( n50078, n50024, n50022 );
nand U81128 ( n49822, n50190, n50191 );
nand U81129 ( n50190, n50195, n49977 );
nand U81130 ( n50191, n1675, n50192 );
nand U81131 ( n50195, n49974, n49976 );
nand U81132 ( n49780, n50142, n50143 );
nand U81133 ( n50142, n50147, n49981 );
nand U81134 ( n50143, n1609, n50144 );
nand U81135 ( n50147, n49978, n49980 );
nand U81136 ( n49797, n50166, n50167 );
nand U81137 ( n50166, n50171, n49813 );
nand U81138 ( n50167, n1643, n50168 );
nand U81139 ( n50171, n49810, n49812 );
nand U81140 ( n49996, n50118, n50119 );
nand U81141 ( n50118, n50123, n49986 );
nand U81142 ( n50119, n1578, n50120 );
nand U81143 ( n50123, n49983, n49985 );
nand U81144 ( n49844, n50214, n50215 );
nand U81145 ( n50215, n1699, n50216 );
nand U81146 ( n50214, n50219, n49966 );
not U81147 ( n1699, n49966 );
xor U81148 ( n50238, n50239, n50240 );
xor U81149 ( n50192, n50193, n50194 );
xor U81150 ( n50261, n50262, n1745 );
xor U81151 ( n50044, n50045, n1320 );
nand U81152 ( n50240, n50248, n50249 );
nand U81153 ( n50249, n49951, n1738 );
nor U81154 ( n50248, n50251, n50252 );
nor U81155 ( n50251, n1725, n50254 );
nand U81156 ( n50218, n50226, n50227 );
nand U81157 ( n50227, n49961, n1717 );
nor U81158 ( n50226, n50228, n50229 );
nor U81159 ( n50228, n49959, n50231 );
nand U81160 ( n50098, n50106, n50107 );
nand U81161 ( n50107, n49995, n1575 );
nor U81162 ( n50106, n50108, n50109 );
nor U81163 ( n50108, n49993, n50111 );
nand U81164 ( n50146, n50154, n50155 );
nand U81165 ( n50155, n49798, n1639 );
nor U81166 ( n50154, n50157, n50158 );
nor U81167 ( n50157, n49804, n50161 );
nand U81168 ( n50194, n50202, n50203 );
nand U81169 ( n50203, n49843, n1693 );
nor U81170 ( n50202, n50204, n50205 );
nor U81171 ( n50204, n49972, n50207 );
nand U81172 ( n50170, n50178, n50179 );
nand U81173 ( n50179, n49823, n1674 );
nor U81174 ( n50178, n50181, n50182 );
nor U81175 ( n50181, n49829, n50185 );
nand U81176 ( n50122, n50130, n50131 );
nand U81177 ( n50131, n49781, n1607 );
nor U81178 ( n50130, n50133, n50134 );
nor U81179 ( n50133, n49787, n50137 );
nand U81180 ( n50287, n50295, n50296 );
nand U81181 ( n50295, n50300, n49908 );
nand U81182 ( n50296, n1760, n50297 );
xor U81183 ( n50300, n50298, n50299 );
nand U81184 ( n49908, n50301, n50302 );
nand U81185 ( n50302, n50303, n1762 );
not U81186 ( n1762, n50304 );
nor U81187 ( n50205, n50206, n49973 );
xor U81188 ( n50206, n49844, n49972 );
nor U81189 ( n50252, n50253, n49950 );
nor U81190 ( n50253, n49868, n49869 );
nor U81191 ( n50109, n50110, n49994 );
nor U81192 ( n50110, n49768, n49769 );
nand U81193 ( n50270, n50271, n50272 );
nand U81194 ( n50272, n49886, n1755 );
nor U81195 ( n50271, n50274, n50275 );
nor U81196 ( n50274, n1747, n50278 );
nand U81197 ( n50053, n50054, n50055 );
nand U81198 ( n50055, n49714, n1362 );
nor U81199 ( n50054, n50057, n50058 );
nor U81200 ( n50057, n49719, n50061 );
nand U81201 ( n50219, n49963, n49965 );
or U81202 ( n50035, n50069, n50070 );
or U81203 ( n49912, n50287, n50286 );
or U81204 ( n49997, n50098, n50097 );
buf U81205 ( n76653, n8230 );
xor U81206 ( n50068, n50069, n50070 );
or U81207 ( n49953, n50240, n50239 );
xor U81208 ( n50096, n50097, n50098 );
nand U81209 ( n49700, n1320, n50045 );
xor U81210 ( n50285, n50286, n50287 );
nand U81211 ( n49955, n50239, n50240 );
nand U81212 ( n49976, n50193, n50194 );
nand U81213 ( n49999, n50097, n50098 );
nor U81214 ( n49718, n49713, n49719 );
nand U81215 ( n49875, n1745, n50262 );
nor U81216 ( n49803, n49797, n49804 );
nor U81217 ( n49786, n49780, n49787 );
nand U81218 ( n50038, n50070, n50069 );
nor U81219 ( n49828, n49822, n49829 );
or U81220 ( n49974, n50194, n50193 );
nor U81221 ( n49869, n49952, n1725 );
nor U81222 ( n49891, n49885, n1747 );
nor U81223 ( n49769, n49996, n49993 );
nor U81224 ( n49859, n49962, n49959 );
nand U81225 ( n49915, n50287, n50286 );
nand U81226 ( n49877, n1743, n50270 );
not U81227 ( n1743, n50262 );
nor U81228 ( n50536, n50303, n50304 );
nand U81229 ( n49914, n50289, n50290 );
nand U81230 ( n50289, n50294, n50293 );
nand U81231 ( n50290, n50291, n50292 );
or U81232 ( n50291, n50293, n50294 );
nand U81233 ( n49702, n1315, n50053 );
not U81234 ( n1315, n50045 );
and U81235 ( n49675, n49684, n49685 );
nand U81236 ( n49684, n49690, n49691 );
nand U81237 ( n49685, n1245, n49686 );
nand U81238 ( n49691, n49689, n49692 );
not U81239 ( n1245, n49690 );
nand U81240 ( n49686, n49687, n49688 );
nand U81241 ( n49688, n1278, n49689 );
nand U81242 ( n49692, n49687, n49693 );
xor U81243 ( n50519, n50527, n50294 );
xnor U81244 ( n50527, n50293, n50292 );
nand U81245 ( n50281, n50519, n50518 );
not U81246 ( n1758, n50790 );
nand U81247 ( n50282, n50521, n50522 );
nand U81248 ( n50521, n50525, n50526 );
nand U81249 ( n50522, n50523, n50524 );
or U81250 ( n50524, n50525, n50526 );
or U81251 ( n50279, n50518, n50519 );
nand U81252 ( n50111, n49996, n49994 );
xor U81253 ( n16787, n17143, n16801 );
xor U81254 ( n17143, n16800, n2629 );
xor U81255 ( n17057, n16787, n17136 );
xnor U81256 ( n17136, n16788, n16789 );
not U81257 ( n82, n15368 );
nand U81258 ( n16930, n17337, n17338 );
nand U81259 ( n17338, n2872, n17339 );
nand U81260 ( n17337, n17342, n16960 );
not U81261 ( n2872, n16960 );
nand U81262 ( n16867, n17244, n17245 );
nand U81263 ( n17244, n17249, n17023 );
nand U81264 ( n17245, n2794, n17246 );
nand U81265 ( n17249, n17020, n17022 );
nand U81266 ( n16825, n17196, n17197 );
nand U81267 ( n17196, n17201, n17027 );
nand U81268 ( n17197, n2730, n17198 );
nand U81269 ( n17201, n17024, n17026 );
nand U81270 ( n16842, n17220, n17221 );
nand U81271 ( n17220, n17225, n16858 );
nand U81272 ( n17221, n2764, n17222 );
nand U81273 ( n17225, n16855, n16857 );
nand U81274 ( n17042, n17172, n17173 );
nand U81275 ( n17172, n17177, n17032 );
nand U81276 ( n17173, n2699, n17174 );
nand U81277 ( n17177, n17029, n17031 );
xnor U81278 ( n17123, n17071, n17124 );
xor U81279 ( n17124, n17068, n17070 );
nand U81280 ( n16889, n17268, n17269 );
nand U81281 ( n17269, n2815, n17270 );
nand U81282 ( n17268, n17273, n17011 );
not U81283 ( n2815, n17011 );
xor U81284 ( n17292, n17293, n17294 );
xor U81285 ( n17315, n17316, n2863 );
xor U81286 ( n17090, n17091, n2438 );
xor U81287 ( n17114, n17115, n2514 );
nand U81288 ( n17294, n17302, n17303 );
nand U81289 ( n17303, n16996, n2855 );
nor U81290 ( n17302, n17305, n17306 );
nor U81291 ( n17305, n2844, n17308 );
nand U81292 ( n17272, n17280, n17281 );
nand U81293 ( n17281, n17006, n2834 );
nor U81294 ( n17280, n17282, n17283 );
nor U81295 ( n17282, n17004, n17285 );
nand U81296 ( n17152, n17160, n17161 );
nand U81297 ( n17161, n17041, n2697 );
nor U81298 ( n17160, n17162, n17163 );
nor U81299 ( n17162, n17039, n17165 );
nand U81300 ( n17200, n17208, n17209 );
nand U81301 ( n17209, n16843, n2763 );
nor U81302 ( n17208, n17211, n17212 );
nor U81303 ( n17211, n16849, n17215 );
nand U81304 ( n17248, n17256, n17257 );
nand U81305 ( n17257, n16888, n2812 );
nor U81306 ( n17256, n17258, n17259 );
nor U81307 ( n17258, n17018, n17261 );
nand U81308 ( n17224, n17232, n17233 );
nand U81309 ( n17233, n16868, n2793 );
nor U81310 ( n17232, n17235, n17236 );
nor U81311 ( n17235, n16874, n17239 );
nand U81312 ( n17176, n17184, n17185 );
nand U81313 ( n17185, n16826, n2728 );
nor U81314 ( n17184, n17187, n17188 );
nor U81315 ( n17187, n16832, n17191 );
nand U81316 ( n17341, n17349, n17350 );
nand U81317 ( n17349, n17354, n16953 );
nand U81318 ( n17350, n2877, n17351 );
xor U81319 ( n17354, n17353, n17352 );
nand U81320 ( n16953, n17355, n17356 );
nand U81321 ( n17356, n17357, n2878 );
not U81322 ( n2878, n17358 );
nor U81323 ( n17259, n17260, n17019 );
xor U81324 ( n17260, n16889, n17018 );
nor U81325 ( n17306, n17307, n16995 );
nor U81326 ( n17307, n16913, n16914 );
nor U81327 ( n17163, n17164, n17040 );
nor U81328 ( n17164, n16813, n16814 );
nand U81329 ( n17324, n17325, n17326 );
nand U81330 ( n17326, n16931, n2870 );
nor U81331 ( n17325, n17328, n17329 );
nor U81332 ( n17328, n16936, n17332 );
nand U81333 ( n17099, n17100, n17101 );
nand U81334 ( n17101, n16758, n2478 );
nor U81335 ( n17100, n17103, n17104 );
nor U81336 ( n17103, n16763, n17107 );
nand U81337 ( n17273, n17008, n17010 );
nand U81338 ( n17342, n16958, n16961 );
or U81339 ( n17043, n17152, n17151 );
buf U81340 ( n76654, n8224 );
xor U81341 ( n17150, n17151, n17152 );
or U81342 ( n16998, n17294, n17293 );
nand U81343 ( n16744, n2438, n17091 );
nand U81344 ( n17000, n17293, n17294 );
nand U81345 ( n17081, n17115, n2514 );
nand U81346 ( n17045, n17151, n17152 );
nand U81347 ( n14846, n49635, n49636 );
nor U81348 ( n49636, n49637, n49638 );
nor U81349 ( n49635, n49656, n49657 );
nand U81350 ( n49638, n49639, n49640 );
nand U81351 ( n16920, n2863, n17316 );
nor U81352 ( n16848, n16842, n16849 );
nor U81353 ( n16831, n16825, n16832 );
nor U81354 ( n16873, n16867, n16874 );
nor U81355 ( n16914, n16997, n2844 );
nor U81356 ( n16935, n16930, n16936 );
nor U81357 ( n16814, n17042, n17039 );
nor U81358 ( n16904, n17007, n17004 );
nor U81359 ( n16762, n16757, n16763 );
nand U81360 ( n16922, n2859, n17324 );
not U81361 ( n2859, n17316 );
nand U81362 ( n16960, n17343, n17344 );
nand U81363 ( n17343, n17348, n17347 );
nand U81364 ( n17344, n17345, n17346 );
or U81365 ( n17345, n17347, n17348 );
nor U81366 ( n17577, n17357, n17358 );
nand U81367 ( n16746, n2433, n17099 );
not U81368 ( n2433, n17091 );
nand U81369 ( n17084, n17123, n2512 );
not U81370 ( n2512, n17115 );
xor U81371 ( n50517, n50518, n50519 );
nand U81372 ( n49878, n50264, n50265 );
nand U81373 ( n50264, n50269, n50268 );
nand U81374 ( n50265, n50266, n50267 );
or U81375 ( n50266, n50268, n50269 );
nand U81376 ( n50299, n50305, n50306 );
nand U81377 ( n50306, n50307, n50308 );
nand U81378 ( n50305, n50314, n50315 );
nor U81379 ( n50308, n50309, n50310 );
nor U81380 ( n50314, n49925, n50307 );
or U81381 ( n49903, n50299, n50298 );
buf U81382 ( n76648, n8232 );
nor U81383 ( n15673, n15368, n5179 );
nand U81384 ( n49905, n50298, n50299 );
nor U81385 ( n16413, n15368, n16347 );
nor U81386 ( n16310, n15368, n16242 );
nor U81387 ( n16099, n15368, n16039 );
nor U81388 ( n15992, n15368, n15932 );
nor U81389 ( n15893, n15368, n15827 );
nor U81390 ( n15578, n15368, n15518 );
nor U81391 ( n15472, n15368, n15412 );
nor U81392 ( n15784, n15368, n15717 );
nor U81393 ( n16200, n15368, n16135 );
and U81394 ( n16719, n16728, n16729 );
nand U81395 ( n16728, n16734, n16735 );
nand U81396 ( n16729, n2363, n16730 );
nand U81397 ( n16735, n16733, n16736 );
not U81398 ( n2363, n16734 );
nor U81399 ( n16687, n15368, n5168 );
nand U81400 ( n8111, n16660, n16662 );
nor U81401 ( n16662, n16663, n16664 );
nor U81402 ( n16660, n16687, n16688 );
nand U81403 ( n16664, n16665, n16667 );
nand U81404 ( n16730, n16731, n16732 );
nand U81405 ( n16732, n2393, n16733 );
xnor U81406 ( n17563, n17348, n17571 );
xor U81407 ( n17571, n17346, n17347 );
nand U81408 ( n17327, n17333, n17334 );
nand U81409 ( n17334, n17335, n17336 );
nand U81410 ( n16736, n16731, n16737 );
not U81411 ( n2873, n17845 );
nand U81412 ( n17336, n17565, n17566 );
nand U81413 ( n17565, n17569, n17570 );
nand U81414 ( n17566, n17567, n17568 );
or U81415 ( n17568, n17569, n17570 );
xor U81416 ( n20626, n20637, n20701 );
xor U81417 ( n20701, n20635, n20636 );
nand U81418 ( n20448, n20687, n20688 );
nand U81419 ( n20688, n20629, n2688 );
nor U81420 ( n20687, n20689, n20690 );
nor U81421 ( n20689, n2688, n20694 );
nand U81422 ( n17384, n17626, n17627 );
nand U81423 ( n17626, n17633, n17637 );
nand U81424 ( n17627, n17628, n17629 );
nand U81425 ( n17629, n17630, n2364 );
nand U81426 ( n17915, n18186, n18187 );
nand U81427 ( n18187, n17963, n18188 );
nor U81428 ( n18186, n18190, n18191 );
nor U81429 ( n18190, n2480, n18194 );
xor U81430 ( n16694, n2355, n2353 );
not U81431 ( n2554, n19845 );
nor U81432 ( n20427, n20452, n8215 );
not U81433 ( n2555, n20101 );
nor U81434 ( n20094, n76159, n2555 );
nand U81435 ( n20720, n20772, n20773 );
nand U81436 ( n20773, n20753, n20774 );
nor U81437 ( n20772, n20775, n20776 );
nor U81438 ( n20775, n20774, n20780 );
not U81439 ( n2395, n17690 );
not U81440 ( n2702, n20704 );
nor U81441 ( n17406, n17404, n17407 );
xor U81442 ( n17407, n17384, n17385 );
nand U81443 ( n18914, n19248, n19249 );
nand U81444 ( n19249, n18926, n2524 );
nor U81445 ( n19251, n19250, n19253 );
xor U81446 ( n18207, n18203, n18208 );
not U81447 ( n2738, n20774 );
nor U81448 ( n20776, n20777, n20751 );
nor U81449 ( n20777, n20778, n20752 );
nor U81450 ( n20778, n2722, n2738 );
nor U81451 ( n20690, n20691, n20627 );
nor U81452 ( n20691, n20692, n20628 );
nor U81453 ( n20692, n2665, n20626 );
and U81454 ( n17687, n17625, n75760 );
nor U81455 ( n75760, n17623, n2395 );
nor U81456 ( n20110, n20111, n20112 );
nor U81457 ( n20111, n20113, n20114 );
nor U81458 ( n20113, n2597, n2613 );
not U81459 ( n2524, n18925 );
nand U81460 ( n20635, n20702, n20703 );
nand U81461 ( n19396, n19967, n19968 );
nor U81462 ( n19967, n19843, n19837 );
nand U81463 ( n19964, n20099, n20100 );
nand U81464 ( n20100, n20097, n20101 );
nor U81465 ( n20099, n20091, n20094 );
not U81466 ( n2353, n16724 );
nor U81467 ( n19252, n18924, n2522 );
nor U81468 ( n18188, n18159, n18195 );
and U81469 ( n18195, n2444, n18196 );
nand U81470 ( n18196, n2447, n18166 );
nand U81471 ( n18163, n18197, n18198 );
nand U81472 ( n18198, n18181, n18185 );
nor U81473 ( n18197, n18178, n2473 );
not U81474 ( n2473, n18182 );
and U81475 ( n18564, n18904, n18905 );
and U81476 ( n17635, n17685, n17686 );
nand U81477 ( n17686, n17621, n17623 );
nor U81478 ( n17685, n17687, n17688 );
nor U81479 ( n17688, n17689, n17690 );
and U81480 ( n20087, n20105, n20106 );
nor U81481 ( n20105, n20109, n20110 );
nand U81482 ( n17165, n17042, n17040 );
xor U81483 ( n50501, n50507, n50269 );
xnor U81484 ( n50507, n50268, n50267 );
nand U81485 ( n50257, n50501, n50500 );
nand U81486 ( n17683, n17908, n17909 );
nand U81487 ( n17909, n17910, n17911 );
nor U81488 ( n17912, n17911, n17916 );
nand U81489 ( n16585, n17651, n17652 );
nand U81490 ( n17651, n16547, n16548 );
nand U81491 ( n17652, n16549, n17653 );
or U81492 ( n17653, n16548, n16547 );
nand U81493 ( n16655, n17393, n17638 );
nand U81494 ( n17638, n16623, n17639 );
xor U81495 ( n17914, n17915, n17911 );
nand U81496 ( n16622, n17640, n17641 );
nand U81497 ( n17640, n16583, n16585 );
nand U81498 ( n17641, n17642, n16587 );
or U81499 ( n17642, n16585, n16583 );
nor U81500 ( n17678, n17679, n17680 );
and U81501 ( n16547, n17674, n17675 );
nand U81502 ( n17675, n17676, n2397 );
nor U81503 ( n17674, n17677, n17678 );
nor U81504 ( n17677, n17681, n17682 );
nor U81505 ( n18159, n18166, n2447 );
xnor U81506 ( n20522, n20700, n20756 );
xnor U81507 ( n20756, n20698, n20699 );
nor U81508 ( n20889, n20890, n20797 );
nor U81509 ( n20890, n20891, n20798 );
nor U81510 ( n20891, n2707, n2723 );
nor U81511 ( n20760, n20761, n20704 );
nor U81512 ( n20761, n20762, n20706 );
and U81513 ( n20449, n20754, n20755 );
nor U81514 ( n20754, n20524, n20518 );
nand U81515 ( n20770, n20885, n20886 );
nor U81516 ( n20885, n20888, n20889 );
xor U81517 ( n53497, n53546, n53547 );
xor U81518 ( n53547, n53548, n53549 );
xor U81519 ( n52674, n53041, n53042 );
xor U81520 ( n53042, n53043, n53044 );
nand U81521 ( n50871, n51142, n51143 );
nor U81522 ( n51142, n51146, n51147 );
nor U81523 ( n51146, n1364, n51150 );
nand U81524 ( n53271, n53313, n53314 );
nand U81525 ( n53313, n53188, n53191 );
nand U81526 ( n53314, n53315, n53190 );
or U81527 ( n53315, n53191, n53188 );
nor U81528 ( n53281, n53310, n8237 );
nand U81529 ( n53370, n53488, n53489 );
nand U81530 ( n53489, n53490, n1567 );
nor U81531 ( n53488, n53491, n53492 );
nor U81532 ( n53491, n1567, n53498 );
nand U81533 ( n51870, n52363, n52364 );
nand U81534 ( n52364, n51882, n1404 );
nor U81535 ( n52363, n52366, n52367 );
nor U81536 ( n52366, n52365, n52368 );
nor U81537 ( n51144, n51116, n51151 );
and U81538 ( n51151, n1327, n51152 );
xor U81539 ( n50604, n1248, n50605 );
and U81540 ( n51520, n51860, n51861 );
nand U81541 ( n53385, n53448, n53449 );
or U81542 ( n53448, n53370, n53373 );
nand U81543 ( n53449, n53450, n53372 );
nand U81544 ( n53450, n53373, n53370 );
nor U81545 ( n53615, n53616, n53617 );
nor U81546 ( n53618, n1589, n1602 );
nor U81547 ( n53492, n53493, n53494 );
nor U81548 ( n53493, n53495, n53496 );
nor U81549 ( n53495, n1549, n53497 );
nor U81550 ( n53066, n53067, n53068 );
nor U81551 ( n53067, n53069, n53070 );
not U81552 ( n1404, n51881 );
nand U81553 ( n52511, n52923, n52924 );
nand U81554 ( n50600, n50860, n50861 );
nand U81555 ( n50861, n50635, n50862 );
nor U81556 ( n50860, n50632, n1273 );
not U81557 ( n1273, n50636 );
nand U81558 ( n50351, n50595, n50596 );
nand U81559 ( n50595, n49558, n49561 );
nand U81560 ( n50596, n50597, n49560 );
or U81561 ( n50597, n49561, n49558 );
nand U81562 ( n50862, n50864, n50865 );
nand U81563 ( n53546, n53610, n53611 );
nor U81564 ( n53610, n53614, n53615 );
and U81565 ( n53191, n53374, n53375 );
nand U81566 ( n53375, n53376, n1518 );
nor U81567 ( n53374, n53377, n53378 );
nor U81568 ( n53377, n1544, n53384 );
nand U81569 ( n51120, n51153, n51154 );
nand U81570 ( n51154, n51137, n51141 );
nor U81571 ( n51153, n51134, n1354 );
not U81572 ( n1354, n51138 );
nand U81573 ( n50344, n50347, n50348 );
nor U81574 ( n50347, n1214, n50349 );
nor U81575 ( n50349, n50350, n1215 );
not U81576 ( n1215, n49605 );
and U81577 ( n53043, n53061, n53062 );
nor U81578 ( n53061, n53065, n53066 );
and U81579 ( n53267, n53274, n53271 );
and U81580 ( n52793, n52800, n52797 );
nand U81581 ( n50909, n51114, n51115 );
nand U81582 ( n51115, n51116, n1327 );
nor U81583 ( n51114, n51117, n51118 );
nand U81584 ( n50867, n51111, n51112 );
nand U81585 ( n51112, n50905, n50909 );
nor U81586 ( n51111, n50902, n1314 );
not U81587 ( n1314, n50906 );
xor U81588 ( n50513, n50784, n50525 );
xor U81589 ( n50784, n50523, n50526 );
nand U81590 ( n50267, n50509, n50510 );
nand U81591 ( n50509, n50514, n50513 );
nand U81592 ( n50510, n50511, n50512 );
or U81593 ( n50511, n50513, n50514 );
nand U81594 ( n17631, n17905, n17906 );
nand U81595 ( n17906, n17679, n17683 );
nor U81596 ( n17905, n17676, n2388 );
not U81597 ( n2388, n17680 );
nand U81598 ( n17637, n2387, n17903 );
not U81599 ( n2387, n17632 );
nand U81600 ( n17904, n17650, n17648 );
nand U81601 ( n17916, n2400, n17915 );
nor U81602 ( n53048, n53051, n53052 );
xor U81603 ( n53052, n1434, n1464 );
nand U81604 ( n53057, n53058, n53059 );
nand U81605 ( n53058, n53044, n53041 );
nand U81606 ( n53059, n53043, n53060 );
or U81607 ( n53060, n53041, n53044 );
nand U81608 ( n51843, n52050, n52051 );
nand U81609 ( n52050, n51833, n51836 );
nand U81610 ( n52051, n51835, n52052 );
or U81611 ( n52052, n51836, n51833 );
not U81612 ( n1405, n52650 );
nand U81613 ( n51836, n52053, n52054 );
nand U81614 ( n52054, n51827, n51831 );
nor U81615 ( n52053, n51823, n51829 );
nand U81616 ( n49469, n50616, n50617 );
nand U81617 ( n50616, n50621, n50620 );
nand U81618 ( n50617, n50618, n50619 );
or U81619 ( n50618, n50620, n50621 );
nand U81620 ( n49561, n50607, n50608 );
or U81621 ( n50607, n49528, n49531 );
nand U81622 ( n50608, n49530, n50609 );
nand U81623 ( n50609, n49531, n49528 );
not U81624 ( n1332, n52181 );
not U81625 ( n1288, n51827 );
nor U81626 ( n52644, n52645, n52646 );
nor U81627 ( n52645, n52647, n52648 );
nor U81628 ( n52647, n52649, n52650 );
nor U81629 ( n51852, n1253, n51853 );
xor U81630 ( n51853, n50882, n50883 );
nand U81631 ( n50882, n52048, n52049 );
nand U81632 ( n52049, n51846, n51843 );
nor U81633 ( n52048, n51845, n51839 );
and U81634 ( n52190, n52202, n52203 );
nand U81635 ( n52203, n52181, n52185 );
nor U81636 ( n52202, n52177, n52183 );
and U81637 ( n49531, n50610, n50611 );
nand U81638 ( n50610, n49499, n49501 );
nand U81639 ( n50611, n49502, n50612 );
or U81640 ( n50612, n49501, n49499 );
and U81641 ( n51839, n1262, n51843 );
not U81642 ( n2687, n20802 );
nand U81643 ( n20527, n20806, n20807 );
or U81644 ( n20806, n20512, n20515 );
nand U81645 ( n20807, n20808, n20514 );
nand U81646 ( n20808, n20515, n20512 );
nor U81647 ( n20850, n20851, n20803 );
nor U81648 ( n20851, n20852, n20804 );
nor U81649 ( n20852, n20848, n20802 );
nand U81650 ( n20426, n8215, n20452 );
nand U81651 ( n17389, n17392, n17393 );
nor U81652 ( n17392, n2355, n17394 );
nor U81653 ( n17394, n17395, n2357 );
not U81654 ( n2357, n16623 );
nor U81655 ( n17391, n2355, n16659 );
nor U81656 ( n20092, n20095, n20096 );
xor U81657 ( n20096, n2555, n2587 );
nand U81658 ( n20219, n20327, n20328 );
nor U81659 ( n20327, n20114, n20107 );
not U81660 ( n2587, n20097 );
and U81661 ( n19837, n19844, n19841 );
xor U81662 ( n53556, n53587, n53588 );
xor U81663 ( n53588, n53589, n53590 );
xor U81664 ( n53439, n53562, n53563 );
xor U81665 ( n53563, n53564, n53565 );
nor U81666 ( n53683, n53684, n53685 );
nor U81667 ( n53684, n53686, n53687 );
nor U81668 ( n53686, n1603, n1615 );
nor U81669 ( n53434, n53435, n53436 );
nor U81670 ( n53435, n53437, n53438 );
nand U81671 ( n53564, n53585, n53586 );
nor U81672 ( n53585, n53558, n53552 );
nand U81673 ( n53307, n53430, n53431 );
nand U81674 ( n53431, n53432, n1564 );
nor U81675 ( n53430, n53433, n53434 );
nor U81676 ( n53433, n1564, n53440 );
nand U81677 ( n53590, n53678, n53679 );
nor U81678 ( n53678, n53682, n53683 );
nand U81679 ( n20417, n20455, n20456 );
or U81680 ( n20455, n20334, n20337 );
nand U81681 ( n20456, n20457, n20336 );
nand U81682 ( n20457, n20337, n20334 );
nand U81683 ( n20337, n20516, n20517 );
nand U81684 ( n20517, n20518, n2640 );
nor U81685 ( n20516, n20519, n20520 );
nor U81686 ( n20519, n2667, n20526 );
and U81687 ( n20413, n20420, n20417 );
nand U81688 ( n49631, n50348, n50593 );
nand U81689 ( n50593, n49605, n50594 );
not U81690 ( n1210, n49680 );
nand U81691 ( n49707, n1358, n49715 );
nand U81692 ( n49715, n49716, n49717 );
not U81693 ( n1358, n49709 );
nand U81694 ( n49716, n49719, n49713 );
nand U81695 ( n17952, n18157, n18158 );
nor U81696 ( n18157, n18160, n18161 );
nand U81697 ( n18158, n18159, n2444 );
nand U81698 ( n17911, n18154, n18155 );
nand U81699 ( n18155, n17948, n17952 );
nor U81700 ( n18154, n17945, n2432 );
not U81701 ( n2432, n17949 );
or U81702 ( n50255, n50500, n50501 );
xor U81703 ( n51164, n51356, n51521 );
xnor U81704 ( n51521, n51357, n51355 );
xor U81705 ( n53504, n52842, n53575 );
xnor U81706 ( n53575, n52843, n52841 );
xor U81707 ( n53702, n53750, n53751 );
xor U81708 ( n53751, n53752, n53753 );
xnor U81709 ( n52500, n52495, n52824 );
xnor U81710 ( n52824, n52493, n52494 );
nand U81711 ( n51512, n51528, n51529 );
nand U81712 ( n51528, n51533, n51532 );
nand U81713 ( n51529, n51530, n51531 );
or U81714 ( n51530, n51532, n51533 );
nand U81715 ( n53641, n53655, n53656 );
or U81716 ( n53655, n53634, n53637 );
nand U81717 ( n53656, n53657, n53636 );
nand U81718 ( n53657, n53637, n53634 );
not U81719 ( n1487, n51899 );
nand U81720 ( n53634, n53694, n53695 );
nand U81721 ( n53695, n53696, n1600 );
nor U81722 ( n53694, n53697, n53698 );
and U81723 ( n53698, n1614, n53699 );
nand U81724 ( n52034, n52496, n52497 );
nand U81725 ( n52496, n52500, n52501 );
nand U81726 ( n52497, n52498, n52499 );
or U81727 ( n52498, n52500, n52501 );
nand U81728 ( n52393, n52909, n52910 );
nand U81729 ( n52910, n52911, n52912 );
nor U81730 ( n53697, n53700, n53701 );
xor U81731 ( n53701, n1600, n1614 );
nor U81732 ( n52374, n52375, n51900 );
nor U81733 ( n52375, n52376, n51901 );
nor U81734 ( n52376, n52372, n51899 );
nand U81735 ( n52841, n53576, n53577 );
or U81736 ( n53576, n53571, n53574 );
nand U81737 ( n53577, n53573, n53578 );
nand U81738 ( n53578, n53574, n53571 );
nand U81739 ( n51355, n51522, n51523 );
nand U81740 ( n51523, n1428, n51512 );
nor U81741 ( n51522, n51524, n51525 );
not U81742 ( n1428, n51509 );
nor U81743 ( n51525, n1432, n51526 );
xor U81744 ( n51526, n51512, n51513 );
and U81745 ( n52494, n52825, n52826 );
nand U81746 ( n52826, n52394, n1538 );
nor U81747 ( n52825, n52828, n52829 );
nor U81748 ( n52828, n52830, n52831 );
and U81749 ( n52829, n1557, n52395 );
nand U81750 ( n17900, n17960, n17961 );
nand U81751 ( n17961, n17962, n2442 );
nor U81752 ( n17960, n17963, n17964 );
nand U81753 ( n18562, n18903, n18905 );
nor U81754 ( n53050, n76094, n1434 );
not U81755 ( n1654, n53858 );
nand U81756 ( n50339, n50583, n50584 );
nand U81757 ( n50583, n50588, n50592 );
nand U81758 ( n50584, n50585, n50586 );
nand U81759 ( n50586, n50587, n1248 );
not U81760 ( n1280, n50645 );
nor U81761 ( n50361, n50359, n50362 );
xor U81762 ( n50362, n50339, n50340 );
and U81763 ( n50642, n50582, n75761 );
nor U81764 ( n75761, n50580, n1280 );
nand U81765 ( n53548, n53594, n53595 );
nand U81766 ( n53595, n1588, n53541 );
nor U81767 ( n53594, n53543, n53536 );
and U81768 ( n50590, n50640, n50641 );
nand U81769 ( n50641, n50578, n50580 );
nor U81770 ( n50640, n50642, n50643 );
nor U81771 ( n50643, n50644, n50645 );
nor U81772 ( n17621, n17625, n2395 );
nand U81773 ( n52916, n53392, n53406 );
nand U81774 ( n53406, n1539, n53393 );
nand U81775 ( n52822, n53397, n53398 );
or U81776 ( n53398, n52913, n52916 );
nor U81777 ( n53397, n53401, n53402 );
nor U81778 ( n53401, n53400, n53405 );
nor U81779 ( n53420, n53388, n53305 );
nor U81780 ( n53402, n53403, n53404 );
xor U81781 ( n53404, n52916, n53400 );
nand U81782 ( n52499, n52818, n52819 );
or U81783 ( n52818, n52823, n52822 );
nand U81784 ( n52819, n52820, n52821 );
nand U81785 ( n52820, n52822, n52823 );
nand U81786 ( n53309, n53418, n53419 );
nor U81787 ( n53418, n53420, n53421 );
nor U81788 ( n53421, n53303, n53302 );
xnor U81789 ( n17385, n17409, n17098 );
xor U81790 ( n17409, n17097, n17096 );
nor U81791 ( n17097, n17621, n17622 );
and U81792 ( n17622, n17623, n17624 );
nand U81793 ( n17624, n2395, n17625 );
buf U81794 ( n76651, n8230 );
not U81795 ( n2557, n19718 );
nand U81796 ( n19833, n19972, n19973 );
nand U81797 ( n19973, n19718, n19714 );
nor U81798 ( n19972, n19716, n19710 );
not U81799 ( n2717, n20641 );
nor U81800 ( n20712, n20713, n20642 );
nor U81801 ( n20713, n20714, n20643 );
nor U81802 ( n20714, n20710, n20641 );
nand U81803 ( n20684, n20749, n20750 );
nand U81804 ( n20750, n2738, n20751 );
nor U81805 ( n20749, n20752, n20753 );
xnor U81806 ( n50340, n50364, n50052 );
xor U81807 ( n50364, n50051, n50050 );
nor U81808 ( n50051, n50578, n50579 );
and U81809 ( n50579, n50580, n50581 );
nand U81810 ( n50581, n1280, n50582 );
nor U81811 ( n50346, n1214, n49634 );
xor U81812 ( n19253, n18925, n18924 );
xor U81813 ( n52368, n51881, n51880 );
xor U81814 ( n20207, n20334, n20335 );
xor U81815 ( n20335, n20336, n20337 );
not U81816 ( n2588, n20082 );
and U81817 ( n20085, n20117, n20118 );
nand U81818 ( n20118, n20082, n20079 );
nor U81819 ( n20117, n20081, n20075 );
xor U81820 ( n53380, n53444, n53445 );
xor U81821 ( n53445, n53446, n53447 );
nand U81822 ( n53447, n53550, n53551 );
nand U81823 ( n53551, n53552, n1565 );
nor U81824 ( n53553, n1587, n53560 );
nand U81825 ( n53561, n53591, n53592 );
or U81826 ( n53591, n53546, n53549 );
nand U81827 ( n53592, n53593, n53548 );
nand U81828 ( n53593, n53549, n53546 );
nand U81829 ( n53387, n53442, n53443 );
nor U81830 ( n53442, n53382, n53376 );
nand U81831 ( n53645, n8234, n53641 );
nor U81832 ( n19839, n19840, n19841 );
nor U81833 ( n19840, n19842, n19843 );
nand U81834 ( n18913, n19242, n19243 );
nand U81835 ( n19242, n19246, n19247 );
nand U81836 ( n19243, n19244, n19245 );
or U81837 ( n19244, n19246, n19247 );
xnor U81838 ( n53163, n53188, n53189 );
xnor U81839 ( n53189, n53190, n53191 );
not U81840 ( n1465, n53038 );
nand U81841 ( n53041, n53073, n53074 );
nand U81842 ( n53074, n53038, n53035 );
nor U81843 ( n53073, n53037, n53031 );
nand U81844 ( n18903, n18916, n18917 );
nand U81845 ( n18916, n18921, n18700 );
nand U81846 ( n18917, n2523, n18918 );
nand U81847 ( n18921, n18697, n18699 );
nand U81848 ( n18700, n18922, n18923 );
nand U81849 ( n18923, n18924, n18925 );
and U81850 ( n18563, n18904, n18903 );
nand U81851 ( n53494, n53516, n53517 );
nand U81852 ( n53516, n53484, n53487 );
nand U81853 ( n53517, n53518, n53486 );
or U81854 ( n53518, n53487, n53484 );
not U81855 ( n1588, n53537 );
nor U81856 ( n53539, n53540, n53541 );
nor U81857 ( n53540, n53542, n53543 );
nor U81858 ( n53542, n1569, n1588 );
and U81859 ( n53484, n53534, n53535 );
nand U81860 ( n53535, n53536, n53537 );
nor U81861 ( n53534, n53538, n53539 );
nor U81862 ( n53538, n53537, n53544 );
nand U81863 ( n20686, n20723, n20724 );
nand U81864 ( n20724, n20680, n2754 );
nor U81865 ( n20723, n20728, n20729 );
not U81866 ( n2754, n20725 );
nor U81867 ( n20729, n20730, n20727 );
nor U81868 ( n20730, n20731, n20679 );
nor U81869 ( n20731, n20726, n20725 );
and U81870 ( n20679, n20726, n20725 );
nand U81871 ( n20768, n20907, n20908 );
nand U81872 ( n20908, n2708, n20879 );
nor U81873 ( n20907, n20881, n20874 );
nor U81874 ( n20077, n20078, n20079 );
nor U81875 ( n20078, n20080, n20081 );
nor U81876 ( n20080, n2567, n20082 );
and U81877 ( n19830, n20073, n20074 );
nand U81878 ( n20074, n20075, n2588 );
nor U81879 ( n20073, n20076, n20077 );
nor U81880 ( n20076, n2588, n20083 );
and U81881 ( n19710, n19717, n19714 );
xor U81882 ( n17682, n17683, n17679 );
xor U81883 ( n53413, n53571, n53572 );
xor U81884 ( n53572, n53573, n53574 );
xor U81885 ( n53053, n53173, n53174 );
xor U81886 ( n53174, n53175, n53176 );
nor U81887 ( n53411, n53415, n53416 );
xor U81888 ( n53416, n53417, n53413 );
nand U81889 ( n53175, n53181, n53182 );
nor U81890 ( n53181, n53070, n53063 );
nand U81891 ( n51869, n52357, n52358 );
nand U81892 ( n52357, n52361, n52362 );
nand U81893 ( n52358, n52359, n52360 );
or U81894 ( n52359, n52361, n52362 );
nand U81895 ( n52654, n52660, n52661 );
nand U81896 ( n52661, n52650, n52646 );
nor U81897 ( n52660, n52648, n52642 );
nand U81898 ( n17322, n17559, n17560 );
nand U81899 ( n17559, n17564, n17336 );
nand U81900 ( n17560, n2865, n17561 );
nand U81901 ( n17564, n17333, n17335 );
nand U81902 ( n16923, n17318, n17319 );
nand U81903 ( n17318, n17323, n17322 );
nand U81904 ( n17319, n17320, n17321 );
or U81905 ( n17320, n17322, n17323 );
not U81906 ( n1370, n52344 );
nand U81907 ( n52351, n52515, n52516 );
nand U81908 ( n52516, n52344, n52340 );
nor U81909 ( n52515, n52342, n52336 );
nand U81910 ( n51169, n52036, n52037 );
or U81911 ( n52036, n52041, n52040 );
nand U81912 ( n52037, n52038, n52039 );
nand U81913 ( n52039, n52040, n52041 );
and U81914 ( n52040, n52353, n52514 );
nand U81915 ( n52514, n52354, n52351 );
and U81916 ( n51134, n8235, n51137 );
nand U81917 ( n51137, n51166, n51167 );
nand U81918 ( n51166, n51171, n51170 );
nand U81919 ( n51167, n51168, n51169 );
or U81920 ( n51168, n51170, n51171 );
nand U81921 ( n53280, n8237, n53310 );
xor U81922 ( n51876, n51532, n51884 );
xnor U81923 ( n51884, n51533, n51531 );
nand U81924 ( n51859, n51872, n51873 );
nand U81925 ( n51873, n1403, n51874 );
nand U81926 ( n51872, n51877, n51656 );
not U81927 ( n1403, n51656 );
and U81928 ( n51519, n51860, n51859 );
nand U81929 ( n51877, n51653, n51655 );
nand U81930 ( n20715, n2709, n20642 );
nand U81931 ( n49528, n50630, n50631 );
nand U81932 ( n50631, n50632, n1282 );
nor U81933 ( n50630, n50633, n50634 );
nor U81934 ( n50633, n50637, n50638 );
nor U81935 ( n50634, n50635, n50636 );
nor U81936 ( n50578, n50582, n1280 );
nand U81937 ( n52670, n52930, n52931 );
nand U81938 ( n52930, n52786, n52783 );
nand U81939 ( n52931, n52785, n52932 );
or U81940 ( n52932, n52783, n52786 );
nor U81941 ( n53033, n53034, n53035 );
nor U81942 ( n53034, n53036, n53037 );
nor U81943 ( n53036, n1448, n53038 );
and U81944 ( n52786, n53029, n53030 );
nand U81945 ( n53030, n53031, n1465 );
nor U81946 ( n53029, n53032, n53033 );
nor U81947 ( n53032, n1465, n53039 );
and U81948 ( n52666, n52673, n52670 );
not U81949 ( n1249, n50635 );
xor U81950 ( n49603, n50592, n50639 );
xor U81951 ( n50639, n50588, n50590 );
nand U81952 ( n20079, n20119, n20120 );
nand U81953 ( n20119, n20072, n20069 );
nand U81954 ( n20120, n20071, n20121 );
or U81955 ( n20121, n20069, n20072 );
nand U81956 ( n20211, n20338, n20339 );
nand U81957 ( n20338, n20200, n20197 );
nand U81958 ( n20339, n20199, n20340 );
or U81959 ( n20340, n20197, n20200 );
not U81960 ( n2670, n20825 );
nand U81961 ( n20410, n20460, n20461 );
nand U81962 ( n20460, n20395, n20398 );
nand U81963 ( n20461, n20397, n20462 );
or U81964 ( n20462, n20398, n20395 );
nor U81965 ( n20504, n20505, n20506 );
nor U81966 ( n20505, n20507, n20508 );
nor U81967 ( n20507, n20509, n20510 );
nor U81968 ( n20205, n20206, n20207 );
nor U81969 ( n20206, n20208, n20209 );
nor U81970 ( n20208, n20210, n20211 );
and U81971 ( n20498, n20814, n20815 );
nand U81972 ( n20815, n20816, n2670 );
nor U81973 ( n20814, n20817, n20818 );
nor U81974 ( n20817, n20823, n20824 );
and U81975 ( n20200, n20399, n20400 );
nand U81976 ( n20400, n20401, n2617 );
nor U81977 ( n20399, n20402, n20403 );
nor U81978 ( n20402, n2642, n20409 );
and U81979 ( n20075, n2567, n20079 );
nand U81980 ( n50872, n1284, n50871 );
nand U81981 ( n50592, n50601, n50858 );
nand U81982 ( n50859, n50910, n1272 );
xor U81983 ( n49662, n1214, n1210 );
and U81984 ( n53410, n53415, n53413 );
nand U81985 ( n52646, n52635, n52662 );
nand U81986 ( n52662, n1407, n52636 );
nor U81987 ( n52668, n52669, n52670 );
nor U81988 ( n52669, n52671, n52672 );
nor U81989 ( n52671, n52673, n52674 );
and U81990 ( n52642, n52649, n52646 );
nand U81991 ( n52325, n52632, n52633 );
nand U81992 ( n52632, n52637, n52638 );
nand U81993 ( n52633, n1407, n52634 );
xor U81994 ( n52637, n52639, n1383 );
nand U81995 ( n52174, n52318, n52319 );
nand U81996 ( n52319, n52320, n1333 );
nor U81997 ( n52318, n52322, n52323 );
not U81998 ( n1333, n52321 );
nor U81999 ( n52322, n52328, n52329 );
nand U82000 ( n52329, n52321, n52325 );
not U82001 ( n1289, n52185 );
not U82002 ( n1254, n51831 );
nor U82003 ( n52179, n52180, n52181 );
nor U82004 ( n52180, n52182, n52183 );
nor U82005 ( n52182, n52184, n52185 );
nand U82006 ( n17408, n17385, n17404 );
nor U82007 ( n20415, n20416, n20417 );
nor U82008 ( n20416, n20418, n20419 );
xor U82009 ( n17689, n17625, n17623 );
nor U82010 ( n52338, n52339, n52340 );
nor U82011 ( n52339, n52341, n52342 );
nor U82012 ( n52341, n52343, n52344 );
xnor U82013 ( n16620, n17637, n17684 );
xor U82014 ( n17684, n17633, n17635 );
and U82015 ( n52336, n52343, n52340 );
nand U82016 ( n50855, n50918, n50919 );
nand U82017 ( n50919, n50920, n1324 );
nor U82018 ( n50918, n50921, n50922 );
nand U82019 ( n51656, n51878, n51879 );
nand U82020 ( n51879, n51880, n51881 );
nand U82021 ( n53400, n53500, n53501 );
nand U82022 ( n53501, n1535, n53502 );
nand U82023 ( n53500, n53505, n52912 );
not U82024 ( n1535, n52912 );
nand U82025 ( n53505, n52909, n52911 );
and U82026 ( n20107, n2597, n20112 );
nand U82027 ( n20843, n20872, n20873 );
nand U82028 ( n20873, n20874, n20875 );
nor U82029 ( n20872, n20876, n20877 );
nor U82030 ( n20876, n20875, n20882 );
not U82031 ( n2708, n20875 );
nor U82032 ( n20877, n20878, n20879 );
nor U82033 ( n20878, n20880, n20881 );
nor U82034 ( n20880, n2692, n2708 );
nand U82035 ( n20853, n2669, n20803 );
and U82036 ( n20091, n20095, n20097 );
nand U82037 ( n53446, n53514, n53515 );
nand U82038 ( n53515, n53497, n53494 );
nor U82039 ( n53514, n53496, n53490 );
and U82040 ( n53490, n1549, n53494 );
not U82041 ( n1277, n50910 );
nand U82042 ( n50601, n50605, n1277 );
nor U82043 ( n50587, n1270, n50588 );
nand U82044 ( n50512, n50804, n50805 );
nand U82045 ( n50804, n50809, n50808 );
nand U82046 ( n50805, n50806, n50807 );
or U82047 ( n50806, n50808, n50809 );
xnor U82048 ( n51513, n51370, n51534 );
xor U82049 ( n51534, n51368, n51369 );
nand U82050 ( n51652, n51897, n51898 );
nand U82051 ( n51898, n51899, n51900 );
nor U82052 ( n51897, n51901, n51902 );
nand U82053 ( n51368, n51649, n51650 );
nand U82054 ( n51650, n51651, n51652 );
nand U82055 ( n51532, n51891, n51892 );
nand U82056 ( n51891, n51896, n51652 );
nand U82057 ( n51892, n1462, n51893 );
nand U82058 ( n51896, n51649, n51651 );
xor U82059 ( n52530, n52783, n52784 );
xor U82060 ( n52784, n52785, n52786 );
nand U82061 ( n52634, n52635, n52636 );
xor U82062 ( n49722, n50012, n50013 );
nand U82063 ( n50013, n50014, n50015 );
nand U82064 ( n50012, n50020, n50021 );
or U82065 ( n50014, n50018, n50019 );
nand U82066 ( n50021, n50022, n50023 );
or U82067 ( n50023, n50024, n50025 );
buf U82068 ( n76324, n75778 );
not U82069 ( n2668, n20506 );
nand U82070 ( n20627, n20695, n20696 );
nand U82071 ( n20695, n20700, n20699 );
nand U82072 ( n20696, n20697, n20698 );
or U82073 ( n20697, n20699, n20700 );
xor U82074 ( n50499, n50500, n50501 );
nand U82075 ( n49956, n50242, n50243 );
nand U82076 ( n50242, n50247, n50246 );
nand U82077 ( n50243, n50244, n50245 );
or U82078 ( n50244, n50246, n50247 );
nand U82079 ( n53285, n53389, n53390 );
nand U82080 ( n53389, n53394, n53395 );
nand U82081 ( n53390, n1539, n53391 );
xor U82082 ( n53394, n53396, n1525 );
nor U82083 ( n53287, n53288, n53289 );
nor U82084 ( n53288, n53290, n53291 );
nor U82085 ( n53290, n53292, n53285 );
nand U82086 ( n53391, n53392, n53393 );
nand U82087 ( n51888, n52502, n52503 );
nand U82088 ( n52502, n52507, n52506 );
nand U82089 ( n52503, n52504, n52505 );
or U82090 ( n52504, n52506, n52507 );
not U82091 ( n2525, n19694 );
nand U82092 ( n19698, n19704, n19705 );
nand U82093 ( n19705, n19694, n19690 );
nor U82094 ( n19704, n19692, n19686 );
nor U82095 ( n53269, n53270, n53271 );
xnor U82096 ( n51045, n50809, n51046 );
xor U82097 ( n51046, n50807, n50808 );
nand U82098 ( n50810, n51037, n1735 );
or U82099 ( n50506, n50781, n50780 );
nand U82100 ( n20398, n20463, n20464 );
nand U82101 ( n20464, n20352, n20356 );
nor U82102 ( n20463, n20348, n20354 );
not U82103 ( n2644, n20352 );
and U82104 ( n53063, n1477, n53068 );
and U82105 ( n20508, n20509, n20510 );
nand U82106 ( n18932, n19255, n19256 );
nand U82107 ( n19255, n19260, n19259 );
nand U82108 ( n19256, n19257, n19258 );
or U82109 ( n19257, n19259, n19260 );
xor U82110 ( n52032, n52383, n51914 );
xor U82111 ( n52383, n51913, n51915 );
nand U82112 ( n51913, n52490, n52491 );
nand U82113 ( n52490, n52495, n52494 );
nand U82114 ( n52491, n52492, n52493 );
or U82115 ( n52492, n52494, n52495 );
nand U82116 ( n53405, n53403, n52916 );
nand U82117 ( n18181, n18210, n18211 );
nand U82118 ( n18210, n18215, n18214 );
nand U82119 ( n18211, n18212, n18213 );
or U82120 ( n18212, n18214, n18215 );
nor U82121 ( n18906, n18904, n18562 );
and U82122 ( n18178, n8218, n18181 );
nand U82123 ( n50812, n51045, n1732 );
not U82124 ( n1732, n51037 );
and U82125 ( n53291, n53292, n53285 );
xor U82126 ( n53631, n53690, n53691 );
xor U82127 ( n53691, n53692, n53693 );
nand U82128 ( n53562, n53622, n53623 );
nand U82129 ( n53623, n53624, n1601 );
nor U82130 ( n53622, n53625, n53626 );
nor U82131 ( n53625, n1601, n53632 );
nor U82132 ( n53626, n53627, n53628 );
nor U82133 ( n53627, n53629, n53630 );
nor U82134 ( n53629, n1590, n53631 );
nand U82135 ( n53692, n53722, n53723 );
nor U82136 ( n53722, n53687, n53680 );
nand U82137 ( n53392, n1525, n53396 );
nor U82138 ( n53789, n53790, n53791 );
nand U82139 ( n53690, n53738, n53739 );
nand U82140 ( n53739, n53740, n1634 );
nor U82141 ( n53738, n53742, n53743 );
not U82142 ( n1634, n53741 );
nor U82143 ( n53743, n53744, n53745 );
nor U82144 ( n53744, n53746, n53747 );
nor U82145 ( n53746, n53748, n53741 );
and U82146 ( n53747, n53748, n53741 );
nor U82147 ( n51851, n50882, n51854 );
nand U82148 ( n51854, n50883, n1253 );
nor U82149 ( n52795, n52796, n52797 );
not U82150 ( n2643, n20510 );
or U82151 ( n20511, n20509, n2643 );
xnor U82152 ( n52836, n52844, n52484 );
xor U82153 ( n52844, n52483, n52485 );
nand U82154 ( n52392, n52832, n52833 );
nand U82155 ( n52833, n1562, n52834 );
nand U82156 ( n52832, n52837, n52489 );
not U82157 ( n1562, n52489 );
nand U82158 ( n52483, n52905, n52906 );
nand U82159 ( n52906, n52907, n52908 );
nand U82160 ( n52837, n52486, n52488 );
nand U82161 ( n20698, n20800, n20801 );
nand U82162 ( n20801, n20802, n20803 );
nor U82163 ( n20800, n20804, n20805 );
and U82164 ( n20805, n20848, n20803 );
nand U82165 ( n20430, n20530, n20531 );
nand U82166 ( n20530, n20536, n20535 );
nand U82167 ( n20531, n2662, n20532 );
xor U82168 ( n20536, n20534, n2635 );
nor U82169 ( n20617, n20529, n20446 );
nor U82170 ( n20434, n20435, n20432 );
nor U82171 ( n20435, n20436, n20322 );
nor U82172 ( n20436, n20431, n20430 );
nand U82173 ( n20451, n20615, n20616 );
nand U82174 ( n20616, n20449, n20448 );
nor U82175 ( n20615, n20617, n20618 );
nor U82176 ( n20618, n20444, n20443 );
and U82177 ( n20322, n20431, n20430 );
nand U82178 ( n20532, n20232, n20234 );
nand U82179 ( n50626, n50900, n50901 );
nand U82180 ( n50901, n50902, n1325 );
nor U82181 ( n50900, n50903, n50904 );
nor U82182 ( n50903, n50907, n50908 );
nor U82183 ( n50904, n50905, n50906 );
and U82184 ( n20753, n2722, n20751 );
nand U82185 ( n50363, n50340, n50359 );
nor U82186 ( n17632, n17648, n17650 );
nor U82187 ( n17630, n17632, n17633 );
nand U82188 ( n52635, n1383, n52639 );
xor U82189 ( n53567, n53634, n53635 );
xor U82190 ( n53635, n53636, n53637 );
nor U82191 ( n53414, n76311, n1542 );
nand U82192 ( n53426, n53509, n53510 );
nor U82193 ( n53509, n53438, n53432 );
not U82194 ( n2392, n17650 );
xnor U82195 ( n53364, n53484, n53485 );
xnor U82196 ( n53485, n53486, n53487 );
nand U82197 ( n53035, n53075, n53076 );
nand U82198 ( n53075, n53028, n53025 );
nand U82199 ( n53076, n53027, n53077 );
or U82200 ( n53077, n53025, n53028 );
nand U82201 ( n53167, n53192, n53193 );
nand U82202 ( n53192, n53156, n53153 );
nand U82203 ( n53193, n53155, n53194 );
or U82204 ( n53194, n53153, n53156 );
nand U82205 ( n53264, n53318, n53319 );
or U82206 ( n53318, n53250, n53251 );
nand U82207 ( n53319, n53252, n53320 );
nand U82208 ( n53320, n53251, n53250 );
nor U82209 ( n53161, n53162, n53163 );
nor U82210 ( n53162, n53164, n53165 );
nor U82211 ( n53164, n53166, n53167 );
and U82212 ( n53361, n53364, n75762 );
nor U82213 ( n75762, n53367, n1520 );
and U82214 ( n53156, n53253, n53254 );
nand U82215 ( n53254, n53255, n1493 );
nor U82216 ( n53253, n53256, n53257 );
nor U82217 ( n53256, n1519, n53263 );
and U82218 ( n53031, n1448, n53035 );
and U82219 ( n53047, n53051, n53053 );
nor U82220 ( n20728, n20726, n20678 );
nand U82221 ( n20678, n20725, n20727 );
nand U82222 ( n50937, n51352, n51353 );
nand U82223 ( n51352, n51357, n51356 );
nand U82224 ( n51353, n51354, n51355 );
or U82225 ( n51354, n51356, n51357 );
nand U82226 ( n51356, n51653, n51654 );
nand U82227 ( n51654, n51655, n51656 );
nor U82228 ( n51349, n51347, n51350 );
xor U82229 ( n51350, n50937, n51341 );
not U82230 ( n1368, n51123 );
nor U82231 ( n20433, n20431, n20321 );
nand U82232 ( n20321, n20430, n20432 );
xnor U82233 ( n52512, n52506, n52804 );
xnor U82234 ( n52804, n52505, n52507 );
xnor U82235 ( n51846, n52046, n52195 );
xnor U82236 ( n52195, n52045, n52047 );
nand U82237 ( n52045, n52196, n52197 );
nand U82238 ( n52196, n52193, n52191 );
nand U82239 ( n52197, n52198, n52194 );
or U82240 ( n52198, n52191, n52193 );
nand U82241 ( n19690, n19679, n19706 );
nand U82242 ( n19706, n2527, n19680 );
nor U82243 ( n19712, n19713, n19714 );
nor U82244 ( n19713, n19715, n19716 );
nor U82245 ( n19715, n19717, n19718 );
and U82246 ( n19686, n19693, n19690 );
xor U82247 ( n50644, n50582, n50580 );
and U82248 ( n20644, n20710, n20642 );
and U82249 ( n20496, n20826, n20827 );
nand U82250 ( n20827, n2672, n20479 );
nor U82251 ( n20826, n20470, n20475 );
xor U82252 ( n53206, n53354, n53355 );
xor U82253 ( n53355, n53356, n53357 );
nor U82254 ( n53460, n53461, n1568 );
nor U82255 ( n53461, n53462, n53463 );
nor U82256 ( n53462, n53464, n53465 );
and U82257 ( n53251, n53321, n53322 );
nand U82258 ( n53322, n53206, n53211 );
nor U82259 ( n53321, n53202, n53208 );
and U82260 ( n53536, n1569, n53541 );
and U82261 ( n53356, n53456, n53457 );
nand U82262 ( n53457, n53458, n1547 );
nor U82263 ( n53456, n53459, n53460 );
nor U82264 ( n53459, n53466, n53467 );
and U82265 ( n53463, n53464, n53465 );
xor U82266 ( n52777, n53025, n53026 );
xor U82267 ( n53026, n53027, n53028 );
nand U82268 ( n52534, n52678, n52679 );
nand U82269 ( n52678, n52629, n52630 );
nand U82270 ( n52679, n52631, n52680 );
or U82271 ( n52680, n52630, n52629 );
nor U82272 ( n52528, n52529, n52530 );
nor U82273 ( n52529, n52531, n52532 );
nor U82274 ( n52531, n52533, n52534 );
nor U82275 ( n52323, n52324, n52325 );
nor U82276 ( n52324, n52326, n52327 );
nor U82277 ( n52326, n52328, n52321 );
and U82278 ( n52327, n52328, n52321 );
and U82279 ( n52629, n52771, n52772 );
nor U82280 ( n52771, n52774, n52775 );
nand U82281 ( n52772, n52773, n1409 );
nor U82282 ( n52774, n1437, n52781 );
nor U82283 ( n18907, n18908, n18905 );
nor U82284 ( n18908, n18909, n18563 );
nor U82285 ( n18909, n18904, n18903 );
not U82286 ( n2690, n20823 );
nand U82287 ( n19402, n19559, n19560 );
nand U82288 ( n19560, n19551, n19547 );
nor U82289 ( n19559, n19549, n19543 );
nor U82290 ( n19688, n19689, n19690 );
nor U82291 ( n19689, n19691, n19692 );
nor U82292 ( n19691, n19693, n19694 );
nand U82293 ( n18213, n19080, n19081 );
or U82294 ( n19080, n19085, n19084 );
nand U82295 ( n19081, n19082, n19083 );
nand U82296 ( n19083, n19084, n19085 );
and U82297 ( n19084, n19399, n19400 );
nand U82298 ( n19400, n19401, n19402 );
and U82299 ( n19543, n19550, n19547 );
nand U82300 ( n20232, n2635, n20534 );
xor U82301 ( n52961, n53149, n53150 );
xor U82302 ( n53150, n53151, n53152 );
nand U82303 ( n52948, n53080, n53081 );
nand U82304 ( n53080, n53023, n53022 );
nand U82305 ( n53081, n53024, n53082 );
or U82306 ( n53082, n53022, n53023 );
nand U82307 ( n53022, n53095, n53096 );
nand U82308 ( n53096, n52961, n52966 );
nor U82309 ( n53095, n52957, n52963 );
not U82310 ( n1523, n53337 );
nand U82311 ( n53211, n53323, n53324 );
nand U82312 ( n53323, n53248, n53245 );
nand U82313 ( n53324, n53247, n53325 );
or U82314 ( n53325, n53245, n53248 );
nand U82315 ( n52782, n52935, n52936 );
nand U82316 ( n52935, n52769, n52768 );
nand U82317 ( n52936, n52770, n52937 );
or U82318 ( n52937, n52768, n52769 );
nor U82319 ( n52942, n52943, n52944 );
nor U82320 ( n52943, n52945, n52946 );
nor U82321 ( n52945, n52947, n52948 );
and U82322 ( n53247, n53326, n53327 );
nand U82323 ( n53327, n53328, n1523 );
nor U82324 ( n53326, n53329, n53330 );
nor U82325 ( n53329, n53335, n53336 );
and U82326 ( n53151, n53200, n53201 );
nand U82327 ( n53201, n53202, n1495 );
nor U82328 ( n53200, n53203, n53204 );
nor U82329 ( n53203, n1522, n53210 );
xnor U82330 ( n51833, n52191, n52192 );
xnor U82331 ( n52192, n52193, n52194 );
nand U82332 ( n51900, n52378, n52379 );
nand U82333 ( n52379, n52380, n52381 );
nand U82334 ( n52815, n53178, n53179 );
or U82335 ( n53178, n53173, n53176 );
nand U82336 ( n53179, n53180, n53175 );
nand U82337 ( n53180, n53176, n53173 );
nand U82338 ( n52381, n52811, n52812 );
nand U82339 ( n52811, n52816, n52815 );
nand U82340 ( n52812, n52813, n52814 );
or U82341 ( n52814, n52815, n52816 );
and U82342 ( n51902, n52372, n51900 );
xor U82343 ( n52809, n52500, n52817 );
xnor U82344 ( n52817, n52501, n52499 );
not U82345 ( n1547, n53465 );
or U82346 ( n53467, n53464, n1547 );
and U82347 ( n20502, n20509, n20506 );
and U82348 ( n53277, n53298, n53299 );
nand U82349 ( n53299, n53300, n53301 );
nand U82350 ( n53298, n1514, n53308 );
xnor U82351 ( n53301, n53302, n53303 );
nand U82352 ( n50899, n51132, n51133 );
nand U82353 ( n51133, n51134, n1369 );
nor U82354 ( n51132, n51135, n51136 );
nor U82355 ( n51136, n51137, n51138 );
and U82356 ( n50902, n8239, n50905 );
nor U82357 ( n51864, n51865, n51519 );
nor U82358 ( n51865, n51860, n51859 );
xor U82359 ( n18208, n18400, n18565 );
xnor U82360 ( n18565, n18401, n18399 );
nand U82361 ( n18400, n18697, n18698 );
nand U82362 ( n18698, n18699, n18700 );
and U82363 ( n53284, n53292, n53289 );
not U82364 ( n79, n15357 );
and U82365 ( n49734, n50010, n50009 );
nor U82366 ( n49728, n49732, n49733 );
nor U82367 ( n49732, n1452, n49734 );
not U82368 ( n2645, n20479 );
not U82369 ( n2619, n20356 );
and U82370 ( n20393, n20468, n20469 );
nand U82371 ( n20469, n20470, n2645 );
nor U82372 ( n20468, n20471, n20472 );
nor U82373 ( n20471, n20477, n20478 );
nand U82374 ( n52802, n1422, n52797 );
nand U82375 ( n53368, n53453, n53454 );
nand U82376 ( n53453, n53357, n53354 );
nand U82377 ( n53454, n53356, n53455 );
or U82378 ( n53455, n53354, n53357 );
nor U82379 ( n53363, n53365, n53366 );
nor U82380 ( n53365, n53367, n53368 );
nand U82381 ( n53354, n53468, n53469 );
nand U82382 ( n53469, n1548, n53337 );
nor U82383 ( n53468, n53328, n53333 );
xor U82384 ( n53424, n53425, n1563 );
nand U82385 ( n53570, n53582, n53583 );
or U82386 ( n53582, n53562, n53565 );
nand U82387 ( n53583, n53584, n53564 );
nand U82388 ( n53584, n53565, n53562 );
not U82389 ( n1563, n53566 );
and U82390 ( n49653, n51837, n51838 );
nand U82391 ( n51838, n51839, n1287 );
nor U82392 ( n51837, n51840, n51841 );
nor U82393 ( n51841, n51842, n51843 );
nand U82394 ( n50020, n50025, n50024 );
nand U82395 ( n52842, n53648, n53649 );
nand U82396 ( n53648, n53652, n52908 );
nand U82397 ( n53649, n1580, n53650 );
nand U82398 ( n53652, n52905, n52907 );
not U82399 ( n1580, n52908 );
and U82400 ( n53366, n53367, n53368 );
xnor U82401 ( n19397, n19259, n19848 );
xnor U82402 ( n19848, n19258, n19260 );
xnor U82403 ( n17557, n17323, n17558 );
xor U82404 ( n17558, n17321, n17322 );
nand U82405 ( n17309, n17551, n2854 );
nand U82406 ( n50504, n50780, n50781 );
xor U82407 ( n50505, n50783, n50513 );
xor U82408 ( n50783, n50514, n50512 );
nand U82409 ( n17311, n17557, n2850 );
not U82410 ( n2850, n17551 );
and U82411 ( n20423, n20439, n20440 );
nand U82412 ( n20440, n20441, n20442 );
nand U82413 ( n20439, n2638, n20450 );
xnor U82414 ( n20442, n20443, n20444 );
nand U82415 ( n20719, n20795, n20796 );
nand U82416 ( n20796, n2723, n20797 );
nor U82417 ( n20795, n20798, n20799 );
and U82418 ( n53680, n1603, n53685 );
and U82419 ( n20874, n2692, n20879 );
and U82420 ( n52320, n52328, n52325 );
xor U82421 ( n50908, n50909, n50905 );
not U82422 ( n2484, n18166 );
nand U82423 ( n53428, n53425, n1563 );
not U82424 ( n1568, n53466 );
nand U82425 ( n52489, n52838, n52839 );
nand U82426 ( n52838, n52843, n52842 );
nand U82427 ( n52839, n52840, n52841 );
or U82428 ( n52840, n52842, n52843 );
nand U82429 ( n19683, n19720, n19721 );
nand U82430 ( n19721, n19574, n19578 );
nor U82431 ( n19720, n19570, n19576 );
not U82432 ( n2528, n19574 );
not U82433 ( n1334, n52069 );
and U82434 ( n52171, n52207, n52208 );
nand U82435 ( n52208, n52069, n52073 );
nor U82436 ( n52207, n52065, n52071 );
nand U82437 ( n53709, n53716, n53717 );
nand U82438 ( n53717, n53702, n53718 );
nor U82439 ( n53716, n53696, n53699 );
and U82440 ( n53696, n53700, n53702 );
nor U82441 ( n51862, n51860, n51518 );
nand U82442 ( n52505, n52805, n52806 );
nand U82443 ( n52805, n52810, n52381 );
nand U82444 ( n52806, n1463, n52807 );
nand U82445 ( n52810, n52378, n52380 );
nand U82446 ( n17979, n18396, n18397 );
nand U82447 ( n18396, n18401, n18400 );
nand U82448 ( n18397, n18398, n18399 );
or U82449 ( n18398, n18400, n18401 );
nor U82450 ( n18393, n18391, n18394 );
xor U82451 ( n18394, n17979, n18385 );
xor U82452 ( n20405, n20512, n20513 );
xor U82453 ( n20513, n20514, n20515 );
nand U82454 ( n20336, n20458, n20459 );
nand U82455 ( n20459, n20405, n20410 );
nor U82456 ( n20458, n20401, n20407 );
nand U82457 ( n17670, n17943, n17944 );
nand U82458 ( n17944, n17945, n2443 );
nor U82459 ( n17943, n17946, n17947 );
nor U82460 ( n17946, n17950, n17951 );
nor U82461 ( n17947, n17948, n17949 );
and U82462 ( n20629, n2665, n20627 );
xor U82463 ( n52921, n52813, n53177 );
xnor U82464 ( n53177, n52816, n52815 );
nand U82465 ( n51509, n1432, n1459 );
and U82466 ( n53360, n53367, n53364 );
nand U82467 ( n19954, n20232, n20233 );
nand U82468 ( n20233, n2662, n20234 );
nand U82469 ( n18556, n18572, n18573 );
nand U82470 ( n18572, n18577, n18576 );
nand U82471 ( n18573, n18574, n18575 );
or U82472 ( n18574, n18576, n18577 );
not U82473 ( n2610, n18943 );
nand U82474 ( n19959, n20223, n20224 );
or U82475 ( n20224, n19951, n19954 );
nor U82476 ( n20223, n20227, n20228 );
nor U82477 ( n20227, n20226, n20231 );
nor U82478 ( n20228, n20229, n20230 );
xor U82479 ( n20230, n19954, n20226 );
nor U82480 ( n19265, n19266, n18944 );
nor U82481 ( n19266, n19267, n18945 );
nor U82482 ( n19267, n19263, n18943 );
nand U82483 ( n18399, n18566, n18567 );
nand U82484 ( n18567, n2549, n18556 );
nor U82485 ( n18566, n18568, n18569 );
not U82486 ( n2549, n18553 );
nor U82487 ( n18569, n2553, n18570 );
xor U82488 ( n18570, n18556, n18557 );
and U82489 ( n19078, n19274, n19275 );
or U82490 ( n19274, n19278, n19279 );
nand U82491 ( n19275, n19276, n19277 );
nand U82492 ( n19276, n19278, n19279 );
xor U82493 ( n20239, n19880, n20247 );
xnor U82494 ( n20247, n19881, n19879 );
nand U82495 ( n20263, n20605, n20606 );
or U82496 ( n20605, n20610, n20609 );
nand U82497 ( n20606, n20607, n20608 );
nand U82498 ( n20607, n20609, n20610 );
nand U82499 ( n20610, n20645, n20646 );
nand U82500 ( n20646, n20566, n2720 );
nor U82501 ( n20645, n20648, n20649 );
nor U82502 ( n20649, n20564, n2718 );
nand U82503 ( n19289, n19947, n19948 );
nand U82504 ( n19948, n19949, n19950 );
nand U82505 ( n19391, n19863, n19864 );
nand U82506 ( n19864, n19290, n2659 );
nor U82507 ( n19863, n19866, n19867 );
nor U82508 ( n19866, n19868, n19869 );
nor U82509 ( n20648, n20647, n20650 );
xor U82510 ( n20650, n20565, n20564 );
nand U82511 ( n19879, n20248, n20249 );
or U82512 ( n20248, n20253, n20252 );
nand U82513 ( n20249, n20250, n20251 );
nand U82514 ( n20251, n20252, n20253 );
not U82515 ( n2775, n20664 );
and U82516 ( n19867, n2678, n19291 );
not U82517 ( n1290, n51811 );
and U82518 ( n51818, n52058, n52059 );
nand U82519 ( n52059, n51811, n51815 );
nor U82520 ( n52058, n51807, n51813 );
xor U82521 ( n19821, n20069, n20070 );
xor U82522 ( n20070, n20071, n20072 );
nand U82523 ( n19827, n19977, n19978 );
nand U82524 ( n19978, n19821, n19826 );
nor U82525 ( n19977, n19817, n19823 );
nand U82526 ( n53628, n53660, n53661 );
or U82527 ( n53660, n53587, n53590 );
nand U82528 ( n53661, n53662, n53589 );
nand U82529 ( n53662, n53590, n53587 );
xor U82530 ( n20243, n20253, n20543 );
xor U82531 ( n20543, n20250, n20252 );
nor U82532 ( n20540, n20539, n20542 );
xor U82533 ( n20542, n2664, n2683 );
xnor U82534 ( n53708, n53754, n53755 );
xor U82535 ( n53754, n53756, n53757 );
nand U82536 ( n53756, n53762, n53763 );
or U82537 ( n53762, n53750, n53753 );
nand U82538 ( n53763, n53764, n53752 );
nand U82539 ( n53764, n53753, n53750 );
or U82540 ( n53711, n53707, n53708 );
not U82541 ( n2487, n19551 );
nor U82542 ( n53742, n53748, n53749 );
nand U82543 ( n53749, n53741, n53745 );
nand U82544 ( n52783, n52933, n52934 );
nand U82545 ( n52934, n52777, n52782 );
nor U82546 ( n52933, n52773, n52779 );
xnor U82547 ( n51895, n51546, n51903 );
xor U82548 ( n51903, n51544, n51545 );
not U82549 ( n342, n48492 );
xor U82550 ( n53706, n53707, n53708 );
xor U82551 ( n18920, n18576, n18928 );
xnor U82552 ( n18928, n18577, n18575 );
nand U82553 ( n17926, n19092, n19093 );
nand U82554 ( n19093, n18890, n18887 );
nor U82555 ( n19092, n18889, n18883 );
nand U82556 ( n18887, n19094, n19095 );
nand U82557 ( n19094, n18877, n18880 );
nand U82558 ( n19095, n18879, n19096 );
or U82559 ( n19096, n18880, n18877 );
nand U82560 ( n18880, n19097, n19098 );
nand U82561 ( n19098, n18871, n18875 );
nor U82562 ( n19097, n18867, n18873 );
nand U82563 ( n16472, n17660, n17661 );
nand U82564 ( n17660, n17665, n17664 );
nand U82565 ( n17661, n17662, n17663 );
or U82566 ( n17662, n17664, n17665 );
nand U82567 ( n16548, n17654, n17655 );
nand U82568 ( n17654, n16509, n16512 );
nand U82569 ( n17655, n16513, n17656 );
or U82570 ( n17656, n16512, n16509 );
not U82571 ( n2449, n19225 );
not U82572 ( n2404, n18871 );
nor U82573 ( n18896, n2368, n18897 );
xor U82574 ( n18897, n17926, n17927 );
and U82575 ( n19234, n19409, n19410 );
nand U82576 ( n19410, n19225, n19229 );
nor U82577 ( n19409, n19221, n19227 );
and U82578 ( n18883, n2377, n18887 );
not U82579 ( n2672, n20477 );
nand U82580 ( n53718, n53719, n53720 );
or U82581 ( n53719, n53690, n53693 );
nand U82582 ( n53720, n53721, n53692 );
nand U82583 ( n53721, n53693, n53690 );
xnor U82584 ( n17591, n17569, n17835 );
xnor U82585 ( n17835, n17567, n17570 );
nand U82586 ( n53712, n53708, n53707 );
and U82587 ( n50625, n50890, n50891 );
nand U82588 ( n50891, n50892, n50893 );
nor U82589 ( n50890, n50894, n50895 );
nor U82590 ( n50895, n1329, n50896 );
nand U82591 ( n52345, n1350, n52340 );
xor U82592 ( n19988, n20197, n20198 );
xor U82593 ( n20198, n20199, n20200 );
nor U82594 ( n53286, n53292, n53293 );
nand U82595 ( n53293, n53285, n53289 );
nand U82596 ( n19846, n2542, n19841 );
nand U82597 ( n20614, n20624, n20625 );
nand U82598 ( n20625, n20626, n20627 );
nor U82599 ( n20624, n20628, n20629 );
not U82600 ( n1548, n53335 );
nor U82601 ( n18180, n18181, n18182 );
nand U82602 ( n18175, n18176, n18177 );
nand U82603 ( n18177, n18178, n2485 );
nor U82604 ( n18176, n18179, n18180 );
nor U82605 ( n18179, n18183, n18184 );
and U82606 ( n17945, n8213, n17948 );
nand U82607 ( n53245, n53338, n53339 );
nand U82608 ( n53339, n1524, n53228 );
nor U82609 ( n53338, n53219, n53224 );
nand U82610 ( n53429, n53566, n1552 );
not U82611 ( n1552, n53425 );
xor U82612 ( n53259, n53370, n53371 );
xor U82613 ( n53371, n53372, n53373 );
nand U82614 ( n20265, n8219, n20263 );
and U82615 ( n53458, n53464, n1568 );
nand U82616 ( n19532, n19676, n19677 );
nand U82617 ( n19676, n19681, n19682 );
nand U82618 ( n19677, n2527, n19678 );
xor U82619 ( n19681, n19683, n2502 );
nand U82620 ( n19218, n19525, n19526 );
nand U82621 ( n19526, n19527, n2450 );
nor U82622 ( n19525, n19529, n19530 );
not U82623 ( n2450, n19528 );
nor U82624 ( n19529, n19535, n19536 );
nand U82625 ( n19536, n19528, n19532 );
nor U82626 ( n19223, n19224, n19225 );
nor U82627 ( n19224, n19226, n19227 );
nor U82628 ( n19226, n19228, n19229 );
not U82629 ( n2405, n19229 );
not U82630 ( n2369, n18875 );
nand U82631 ( n19678, n19679, n19680 );
and U82632 ( n51882, n52365, n51880 );
and U82633 ( n18926, n19250, n18924 );
nand U82634 ( n20514, n20809, n20810 );
nand U82635 ( n20810, n20506, n20510 );
nor U82636 ( n20809, n20502, n20508 );
nand U82637 ( n53791, n8233, n53787 );
nand U82638 ( n17353, n17359, n17360 );
nand U82639 ( n17360, n17361, n17362 );
nand U82640 ( n17359, n17368, n16984 );
nor U82641 ( n17362, n17363, n17364 );
nor U82642 ( n17368, n16987, n17361 );
or U82643 ( n16948, n17353, n17352 );
buf U82644 ( n76590, n75779 );
xor U82645 ( n52350, n52361, n52656 );
xnor U82646 ( n52656, n52362, n52360 );
nand U82647 ( n16950, n17352, n17353 );
xor U82648 ( n53106, n53245, n53246 );
xor U82649 ( n53246, n53247, n53248 );
nand U82650 ( n53093, n53197, n53198 );
nand U82651 ( n53197, n53152, n53149 );
nand U82652 ( n53198, n53151, n53199 );
or U82653 ( n53199, n53149, n53152 );
nand U82654 ( n53149, n53212, n53213 );
nand U82655 ( n53213, n53106, n53111 );
nor U82656 ( n53212, n53102, n53108 );
nor U82657 ( n53087, n53088, n53089 );
nor U82658 ( n53088, n53090, n53091 );
nor U82659 ( n53090, n53092, n53093 );
xor U82660 ( n52978, n53145, n53146 );
xor U82661 ( n53146, n53147, n53148 );
nand U82662 ( n53017, n53112, n53113 );
nand U82663 ( n53113, n52978, n52983 );
nor U82664 ( n53112, n52974, n52980 );
nand U82665 ( n53228, n53244, n53340 );
nand U82666 ( n53340, n53242, n53243 );
nand U82667 ( n52966, n53097, n53098 );
nand U82668 ( n53097, n53020, n53017 );
nand U82669 ( n53098, n53019, n53099 );
or U82670 ( n53099, n53017, n53020 );
and U82671 ( n53147, n53217, n53218 );
nand U82672 ( n53218, n53219, n1498 );
nor U82673 ( n53217, n53220, n53221 );
nor U82674 ( n53220, n53226, n53227 );
nand U82675 ( n49625, n51682, n51683 );
or U82676 ( n51682, n49594, n49597 );
nand U82677 ( n51683, n49596, n51684 );
nand U82678 ( n51684, n49597, n49594 );
nor U82679 ( n51825, n51826, n51827 );
nor U82680 ( n51826, n51828, n51829 );
nor U82681 ( n51828, n51830, n51831 );
nand U82682 ( n49654, n51679, n51680 );
nand U82683 ( n51679, n49622, n49625 );
nand U82684 ( n51680, n49624, n51681 );
or U82685 ( n51681, n49625, n49622 );
nor U82686 ( n51842, n51844, n51845 );
nor U82687 ( n51844, n1262, n51846 );
nand U82688 ( n53589, n53663, n53664 );
nand U82689 ( n53664, n1602, n53617 );
and U82690 ( n20680, n20726, n20727 );
nand U82691 ( n52191, n52346, n52347 );
nand U82692 ( n52346, n52352, n52351 );
nand U82693 ( n52347, n1330, n52348 );
nand U82694 ( n52352, n52353, n52354 );
and U82695 ( n53091, n53092, n53093 );
xor U82696 ( n17951, n17952, n17948 );
xor U82697 ( n19557, n19246, n19700 );
xnor U82698 ( n19700, n19247, n19245 );
nor U82699 ( n19545, n19546, n19547 );
nor U82700 ( n19546, n19548, n19549 );
nor U82701 ( n19548, n19550, n19551 );
and U82702 ( n20323, n20431, n20432 );
nand U82703 ( n53190, n53316, n53317 );
nand U82704 ( n53317, n53259, n53264 );
nor U82705 ( n53316, n53255, n53261 );
nand U82706 ( n53436, n53511, n53512 );
or U82707 ( n53511, n53444, n53447 );
nand U82708 ( n53512, n53513, n53446 );
nand U82709 ( n53513, n53447, n53444 );
and U82710 ( n53432, n1550, n53436 );
and U82711 ( n20391, n20480, n20481 );
nand U82712 ( n20481, n2647, n20374 );
nor U82713 ( n20480, n20365, n20370 );
xnor U82714 ( n52547, n52767, n52768 );
xnor U82715 ( n52767, n52769, n52770 );
nand U82716 ( n52630, n52681, n52682 );
nand U82717 ( n52682, n52547, n52552 );
nor U82718 ( n52681, n52543, n52549 );
nor U82719 ( n49733, n50009, n50010 );
nand U82720 ( n20845, n20857, n20858 );
nand U82721 ( n20858, n2690, n20825 );
nor U82722 ( n20857, n20816, n20821 );
xor U82723 ( n17550, n17551, n2854 );
nand U82724 ( n17001, n17296, n17297 );
nand U82725 ( n17296, n17301, n17300 );
nand U82726 ( n17297, n17298, n17299 );
or U82727 ( n17298, n17300, n17301 );
nand U82728 ( n17649, n2392, n17648 );
xnor U82729 ( n19965, n20221, n19857 );
xor U82730 ( n20221, n19860, n19859 );
xor U82731 ( n52944, n53153, n53154 );
xor U82732 ( n53154, n53155, n53156 );
nand U82733 ( n19679, n2502, n19683 );
nand U82734 ( n53486, n53519, n53520 );
nand U82735 ( n53520, n1568, n53465 );
nor U82736 ( n53519, n53458, n53463 );
and U82737 ( n20799, n2707, n20797 );
xor U82738 ( n20621, n20622, n2682 );
nand U82739 ( n20547, n20632, n20633 );
or U82740 ( n20632, n20637, n20636 );
nand U82741 ( n20633, n20634, n20635 );
nand U82742 ( n20634, n20636, n20637 );
not U82743 ( n2682, n20630 );
nand U82744 ( n20226, n20235, n20236 );
nand U82745 ( n20236, n2663, n20237 );
nand U82746 ( n20235, n20240, n19950 );
not U82747 ( n2663, n19950 );
nand U82748 ( n20240, n19947, n19949 );
nand U82749 ( n20231, n20229, n19954 );
nand U82750 ( n16751, n2475, n16759 );
nand U82751 ( n16759, n16760, n16761 );
not U82752 ( n2475, n16753 );
nand U82753 ( n16760, n16763, n16757 );
or U82754 ( n53094, n53092, n1469 );
xnor U82755 ( n49622, n51833, n51834 );
xnor U82756 ( n51834, n51835, n51836 );
nand U82757 ( n20611, n20622, n2682 );
xnor U82758 ( n51908, n51644, n51916 );
xor U82759 ( n51916, n51642, n51643 );
nand U82760 ( n51545, n51904, n51905 );
nand U82761 ( n51904, n51909, n51648 );
nand U82762 ( n51905, n1510, n51906 );
nand U82763 ( n51909, n51645, n51647 );
nand U82764 ( n52029, n52390, n52391 );
nand U82765 ( n52391, n52392, n52393 );
nor U82766 ( n52390, n52394, n52395 );
xor U82767 ( n20549, n20610, n20638 );
xor U82768 ( n20638, n20608, n20609 );
and U82769 ( n17676, n8212, n17679 );
xor U82770 ( n51130, n51171, n51856 );
xnor U82771 ( n51856, n51169, n51170 );
nand U82772 ( n50769, n50777, n50778 );
nand U82773 ( n50777, n50782, n50505 );
nand U82774 ( n50778, n1737, n50779 );
xor U82775 ( n50782, n50781, n50780 );
nand U82776 ( n50494, n50768, n50769 );
xor U82777 ( n51036, n51037, n1735 );
nand U82778 ( n50495, n50771, n50772 );
nand U82779 ( n50771, n50775, n50776 );
nand U82780 ( n50772, n50773, n50774 );
or U82781 ( n50774, n50775, n50776 );
nand U82782 ( n52186, n1309, n52185 );
nor U82783 ( n20246, n76569, n2664 );
and U82784 ( n53624, n1590, n53628 );
xor U82785 ( n52218, n52628, n52629 );
xor U82786 ( n52628, n52630, n52631 );
not U82787 ( n1524, n53226 );
xnor U82788 ( n51539, n51547, n51380 );
xor U82789 ( n51547, n51382, n51383 );
nand U82790 ( n51369, n51535, n51536 );
nand U82791 ( n51536, n1488, n51537 );
nand U82792 ( n51535, n51540, n51508 );
not U82793 ( n1488, n51508 );
nand U82794 ( n51382, n51645, n51646 );
nand U82795 ( n51646, n51647, n51648 );
nand U82796 ( n51540, n51505, n51507 );
xnor U82797 ( n51341, n51338, n51358 );
xor U82798 ( n51358, n51336, n51337 );
xnor U82799 ( n18557, n18414, n18578 );
xor U82800 ( n18578, n18412, n18413 );
nand U82801 ( n18696, n18941, n18942 );
nand U82802 ( n18942, n18943, n18944 );
nor U82803 ( n18941, n18945, n18946 );
nand U82804 ( n18412, n18693, n18694 );
nand U82805 ( n18694, n18695, n18696 );
nand U82806 ( n18576, n18935, n18936 );
nand U82807 ( n18935, n18940, n18696 );
nand U82808 ( n18936, n2584, n18937 );
nand U82809 ( n18940, n18693, n18695 );
and U82810 ( n53740, n53748, n53745 );
nor U82811 ( n19530, n19531, n19532 );
nor U82812 ( n19531, n19533, n19534 );
nor U82813 ( n19533, n19535, n19528 );
and U82814 ( n53612, n1589, n53617 );
xor U82815 ( n50483, n50246, n50491 );
xnor U82816 ( n50491, n50247, n50245 );
nand U82817 ( n50234, n50483, n50482 );
nand U82818 ( n17590, n17829, n17830 );
nand U82819 ( n17829, n17834, n17833 );
nand U82820 ( n17830, n17831, n17832 );
or U82821 ( n17831, n17833, n17834 );
nor U82822 ( n15663, n15357, n5179 );
xnor U82823 ( n18084, n17834, n18092 );
xor U82824 ( n18092, n17832, n17833 );
nand U82825 ( n17826, n17855, n17856 );
nand U82826 ( n17856, n17857, n17858 );
nand U82827 ( n17312, n17553, n17554 );
nand U82828 ( n17553, n17555, n17556 );
or U82829 ( n17556, n17826, n17825 );
nand U82830 ( n53636, n53658, n53659 );
nand U82831 ( n53659, n53631, n53628 );
nor U82832 ( n53658, n53630, n53624 );
nand U82833 ( n53111, n53214, n53215 );
nand U82834 ( n53214, n53148, n53145 );
nand U82835 ( n53215, n53147, n53216 );
or U82836 ( n53216, n53145, n53148 );
and U82837 ( n53019, n53100, n53101 );
nand U82838 ( n53101, n53102, n1472 );
nor U82839 ( n53100, n53103, n53104 );
nor U82840 ( n53103, n1497, n53110 );
xor U82841 ( n19853, n19861, n19278 );
xnor U82842 ( n19861, n19277, n19279 );
nand U82843 ( n19258, n19849, n19850 );
nand U82844 ( n19850, n2585, n19851 );
nand U82845 ( n19849, n19854, n19272 );
not U82846 ( n2585, n19272 );
nand U82847 ( n19854, n19269, n19271 );
xor U82848 ( n18890, n19239, n19090 );
xor U82849 ( n19239, n19089, n19091 );
nand U82850 ( n19089, n19403, n19404 );
nand U82851 ( n19403, n19238, n19236 );
nand U82852 ( n19404, n19405, n19237 );
or U82853 ( n19405, n19236, n19238 );
nor U82854 ( n16402, n15357, n16347 );
nor U82855 ( n16299, n15357, n16242 );
nor U82856 ( n16190, n15357, n16135 );
nor U82857 ( n16088, n15357, n16039 );
nor U82858 ( n15980, n15357, n15932 );
nor U82859 ( n15882, n15357, n15827 );
nor U82860 ( n15774, n15357, n15717 );
nor U82861 ( n15567, n15357, n15518 );
nor U82862 ( n15460, n15357, n15412 );
nor U82863 ( n16649, n15357, n5168 );
nand U82864 ( n8116, n16624, n16625 );
nor U82865 ( n16625, n16627, n16628 );
nor U82866 ( n16624, n16649, n16650 );
nand U82867 ( n16628, n16629, n16630 );
and U82868 ( n20245, n20539, n20243 );
nand U82869 ( n51129, n52042, n52043 );
nand U82870 ( n52042, n52047, n52046 );
nand U82871 ( n52043, n52044, n52045 );
or U82872 ( n52044, n52046, n52047 );
xnor U82873 ( n19874, n19301, n19882 );
xor U82874 ( n19882, n19302, n19300 );
nand U82875 ( n19288, n19870, n19871 );
nand U82876 ( n19871, n2684, n19872 );
nand U82877 ( n19870, n19875, n19386 );
not U82878 ( n2684, n19386 );
nand U82879 ( n19300, n19883, n19884 );
nand U82880 ( n19884, n19885, n19886 );
nand U82881 ( n19875, n19383, n19385 );
nor U82882 ( n20656, n20584, n20587 );
and U82883 ( n19523, n19568, n19569 );
nor U82884 ( n19568, n19571, n19572 );
nand U82885 ( n19569, n19570, n2489 );
nor U82886 ( n19572, n19573, n19574 );
nand U82887 ( n19272, n19855, n19856 );
nand U82888 ( n19855, n19860, n19859 );
nand U82889 ( n19856, n19857, n19858 );
or U82890 ( n19858, n19859, n19860 );
and U82891 ( n19534, n19535, n19528 );
xor U82892 ( n20568, n20314, n20569 );
xnor U82893 ( n20569, n20315, n20313 );
xor U82894 ( n20559, n20560, n2733 );
nand U82895 ( n50879, n1253, n1285 );
not U82896 ( n1285, n50883 );
nor U82897 ( n19571, n2528, n19579 );
nand U82898 ( n19579, n2507, n19578 );
not U82899 ( n2452, n19113 );
and U82900 ( n19215, n19414, n19415 );
nand U82901 ( n19415, n19113, n19117 );
nor U82902 ( n19414, n19109, n19115 );
nand U82903 ( n18944, n19269, n19270 );
nand U82904 ( n19270, n19271, n19272 );
and U82905 ( n18946, n19263, n18944 );
or U82906 ( n50492, n50769, n50768 );
xnor U82907 ( n52692, n53021, n53022 );
xnor U82908 ( n53021, n53023, n53024 );
not U82909 ( n2647, n20372 );
and U82910 ( n52688, n52695, n52692 );
nand U82911 ( n19672, n19815, n19816 );
nor U82912 ( n19815, n19818, n19819 );
nand U82913 ( n19816, n19817, n2529 );
nor U82914 ( n19819, n19820, n19821 );
not U82915 ( n2489, n19578 );
nor U82916 ( n19573, n19575, n19576 );
nor U82917 ( n19575, n19577, n19578 );
xnor U82918 ( n20133, n20395, n20396 );
xnor U82919 ( n20396, n20397, n20398 );
and U82920 ( n20129, n20136, n20133 );
xor U82921 ( n18877, n19235, n19236 );
xor U82922 ( n19235, n19237, n19238 );
nand U82923 ( n20319, n20562, n20563 );
nand U82924 ( n20563, n20564, n20565 );
nor U82925 ( n20562, n20566, n20567 );
and U82926 ( n20566, n20647, n20564 );
nand U82927 ( n53308, n53303, n53302 );
xor U82928 ( n52709, n53017, n53018 );
xor U82929 ( n53018, n53019, n53020 );
nand U82930 ( n52696, n52952, n52953 );
nand U82931 ( n52952, n52765, n52764 );
nand U82932 ( n52953, n52766, n52954 );
or U82933 ( n52954, n52764, n52765 );
nand U82934 ( n52764, n52967, n52968 );
nand U82935 ( n52968, n52709, n52714 );
nor U82936 ( n52967, n52705, n52711 );
and U82937 ( n52694, n52695, n52696 );
nand U82938 ( n19719, n2543, n19714 );
not U82939 ( n2624, n20374 );
xnor U82940 ( n51928, n51556, n51929 );
xor U82941 ( n51929, n51554, n51555 );
xor U82942 ( n51919, n51920, n1579 );
nand U82943 ( n52403, n52411, n52412 );
nand U82944 ( n52412, n51956, n1648 );
nor U82945 ( n52411, n52415, n52416 );
nor U82946 ( n52415, n1628, n52418 );
nand U82947 ( n51934, n51942, n51943 );
or U82948 ( n51943, n51632, n51631 );
nor U82949 ( n51942, n51944, n51945 );
nor U82950 ( n51944, n51634, n51947 );
nand U82951 ( n51555, n51930, n51931 );
nand U82952 ( n51930, n51935, n51561 );
nand U82953 ( n51931, n1598, n51932 );
nand U82954 ( n51935, n51558, n51560 );
nand U82955 ( n52856, n53801, n53841 );
nand U82956 ( n53841, n53802, n53799 );
nand U82957 ( n52471, n52853, n52854 );
nand U82958 ( n52854, n52855, n52856 );
nor U82959 ( n52853, n52857, n52858 );
and U82960 ( n51945, n51634, n75763 );
xor U82961 ( n75763, n51631, n51633 );
nand U82962 ( n52020, n52402, n52403 );
nand U82963 ( n50813, n51039, n51040 );
nand U82964 ( n51039, n51044, n51043 );
nand U82965 ( n51040, n51041, n51042 );
or U82966 ( n51041, n51043, n51044 );
and U82967 ( n17669, n17934, n17935 );
nand U82968 ( n17935, n2398, n17936 );
nor U82969 ( n17934, n17938, n17939 );
not U82970 ( n2398, n17937 );
or U82971 ( n50232, n50482, n50483 );
nor U82972 ( n20567, n76586, n2720 );
not U82973 ( n2720, n20565 );
nor U82974 ( n48757, n48492, n48719 );
nand U82975 ( n51648, n51910, n51911 );
nand U82976 ( n51910, n51915, n51914 );
nand U82977 ( n51911, n51912, n51913 );
or U82978 ( n51912, n51914, n51915 );
xnor U82979 ( n52813, n53294, n52823 );
xnor U82980 ( n53294, n52822, n52821 );
nand U82981 ( n20608, n20639, n20640 );
nand U82982 ( n20640, n20641, n20642 );
nor U82983 ( n20639, n20643, n20644 );
xor U82984 ( n52868, n52876, n52443 );
xnor U82985 ( n52876, n52442, n52441 );
xor U82986 ( n52851, n52859, n52430 );
xnor U82987 ( n52859, n52429, n52428 );
xor U82988 ( n52866, n52867, n52868 );
nand U82989 ( n52470, n52851, n52850 );
nor U82990 ( n49319, n48492, n49280 );
nor U82991 ( n49128, n48492, n7834 );
nor U82992 ( n49050, n48492, n48995 );
nor U82993 ( n48955, n48492, n48896 );
nor U82994 ( n48668, n48492, n48629 );
nor U82995 ( n48590, n48492, n48535 );
nor U82996 ( n49412, n48492, n49358 );
nor U82997 ( n49223, n48492, n49184 );
nor U82998 ( n48854, n48492, n48815 );
nand U82999 ( n20316, n20560, n2733 );
nand U83000 ( n49703, n50047, n50048 );
or U83001 ( n50047, n50052, n50051 );
nand U83002 ( n50048, n50049, n50050 );
nand U83003 ( n50049, n50051, n50052 );
nor U83004 ( n49626, n48492, n49462 );
nand U83005 ( n14851, n49606, n49607 );
nor U83006 ( n49607, n49608, n49609 );
nor U83007 ( n49606, n49626, n49627 );
nand U83008 ( n49609, n49610, n49611 );
and U83009 ( n52766, n52955, n52956 );
nand U83010 ( n52956, n52957, n1440 );
nor U83011 ( n52955, n52958, n52959 );
nor U83012 ( n52958, n1470, n52965 );
xnor U83013 ( n53814, n53822, n52874 );
xor U83014 ( n53822, n52875, n52873 );
xor U83015 ( n53812, n53813, n53814 );
nand U83016 ( n52466, n52868, n52867 );
nand U83017 ( n20613, n20630, n2673 );
not U83018 ( n2673, n20622 );
and U83019 ( n19527, n19535, n19532 );
nand U83020 ( n20137, n20343, n20344 );
nand U83021 ( n20343, n20195, n20194 );
nand U83022 ( n20344, n20196, n20345 );
or U83023 ( n20345, n20194, n20195 );
nor U83024 ( n20350, n20351, n20352 );
nor U83025 ( n20351, n20353, n20354 );
nor U83026 ( n20353, n20355, n20356 );
and U83027 ( n20135, n20136, n20137 );
xnor U83028 ( n53089, n53249, n53250 );
xnor U83029 ( n53249, n53251, n53252 );
and U83030 ( n53085, n53092, n53089 );
xor U83031 ( n19076, n19280, n18958 );
xor U83032 ( n19280, n18957, n18959 );
not U83033 ( n1684, n53828 );
nand U83034 ( n17096, n17410, n17411 );
nand U83035 ( n17410, n17415, n17111 );
nand U83036 ( n17411, n2437, n17412 );
nand U83037 ( n17415, n17108, n17110 );
not U83038 ( n2437, n17111 );
nand U83039 ( n51635, n51920, n1579 );
nand U83040 ( n52862, n53814, n53813 );
nor U83041 ( n18895, n17926, n18898 );
nand U83042 ( n18898, n17927, n2368 );
nand U83043 ( n18105, n76655, n8222 );
buf U83044 ( n76655, n8224 );
xnor U83045 ( n52046, n52355, n52041 );
xnor U83046 ( n52355, n52040, n52038 );
nand U83047 ( n51508, n51541, n51542 );
nand U83048 ( n51541, n51546, n51545 );
nand U83049 ( n51542, n51543, n51544 );
or U83050 ( n51543, n51545, n51546 );
xnor U83051 ( n52564, n52763, n52764 );
xnor U83052 ( n52763, n52765, n52766 );
nand U83053 ( n52222, n52538, n52539 );
nand U83054 ( n52538, n52312, n52311 );
nand U83055 ( n52539, n52313, n52540 );
or U83056 ( n52540, n52311, n52312 );
nand U83057 ( n52552, n52683, n52684 );
nand U83058 ( n52683, n52626, n52625 );
nand U83059 ( n52684, n52627, n52685 );
or U83060 ( n52685, n52625, n52626 );
and U83061 ( n52313, n52541, n52542 );
nand U83062 ( n52542, n52543, n1375 );
nor U83063 ( n52541, n52544, n52545 );
nor U83064 ( n52544, n1410, n52551 );
or U83065 ( n52860, n53813, n53814 );
xor U83066 ( n50767, n50768, n50769 );
nand U83067 ( n50235, n50485, n50486 );
nand U83068 ( n50485, n50489, n50490 );
nand U83069 ( n50486, n50487, n50488 );
or U83070 ( n50488, n50489, n50490 );
not U83071 ( n339, n48483 );
not U83072 ( n1474, n53128 );
nand U83073 ( n52983, n53114, n53115 );
nand U83074 ( n53114, n53016, n53013 );
nand U83075 ( n53115, n53015, n53116 );
or U83076 ( n53116, n53013, n53016 );
and U83077 ( n53015, n53117, n53118 );
nand U83078 ( n53118, n53119, n1474 );
nor U83079 ( n53117, n53120, n53121 );
nor U83080 ( n53120, n53126, n53127 );
or U83081 ( n52464, n52867, n52868 );
nand U83082 ( n20194, n20358, n20359 );
nand U83083 ( n20359, n20150, n20154 );
nor U83084 ( n20358, n20146, n20152 );
not U83085 ( n2620, n20150 );
xor U83086 ( n53650, n53651, n1597 );
not U83087 ( n1597, n53713 );
nand U83088 ( n53755, n53794, n53795 );
nand U83089 ( n53794, n53800, n53799 );
nand U83090 ( n53795, n1630, n53796 );
nand U83091 ( n53800, n53801, n53802 );
not U83092 ( n1630, n53799 );
not U83093 ( n1364, n50920 );
nand U83094 ( n52905, n53651, n1597 );
or U83095 ( n52018, n52403, n52402 );
nand U83096 ( n16684, n18723, n18724 );
nand U83097 ( n18723, n16644, n16647 );
nand U83098 ( n18724, n16648, n18725 );
or U83099 ( n18725, n16647, n16644 );
nor U83100 ( n18869, n18870, n18871 );
nor U83101 ( n18870, n18872, n18873 );
nor U83102 ( n18872, n18874, n18875 );
nand U83103 ( n16647, n18726, n18727 );
nand U83104 ( n18726, n16609, n16610 );
nand U83105 ( n18727, n16612, n18728 );
or U83106 ( n18728, n16610, n16609 );
nand U83107 ( n17663, n18720, n18721 );
nand U83108 ( n18720, n16683, n16684 );
nand U83109 ( n18721, n16685, n18722 );
or U83110 ( n18722, n16684, n16683 );
nand U83111 ( n17554, n17825, n17826 );
nand U83112 ( n52907, n53713, n1592 );
not U83113 ( n1592, n53651 );
not U83114 ( n1292, n52073 );
nor U83115 ( n52216, n52217, n52218 );
nor U83116 ( n52217, n52219, n52220 );
nor U83117 ( n52219, n52221, n52222 );
nand U83118 ( n50940, n51347, n1429 );
nand U83119 ( n53145, n53229, n53230 );
nand U83120 ( n53230, n1499, n53128 );
nor U83121 ( n53229, n53119, n53124 );
xor U83122 ( n53126, n53241, n53242 );
nand U83123 ( n53241, n53243, n53244 );
not U83124 ( n1293, n51703 );
not U83125 ( n1255, n51815 );
and U83126 ( n51802, n52075, n52076 );
nand U83127 ( n52076, n51703, n51707 );
nor U83128 ( n52075, n51699, n51705 );
xor U83129 ( n52581, n52759, n52760 );
xor U83130 ( n52760, n52761, n52762 );
xor U83131 ( n52091, n52306, n52307 );
xor U83132 ( n52307, n52308, n52309 );
nand U83133 ( n52568, n52700, n52701 );
nand U83134 ( n52700, n52622, n52621 );
nand U83135 ( n52701, n52623, n52702 );
or U83136 ( n52702, n52621, n52622 );
nand U83137 ( n52165, n52226, n52227 );
nand U83138 ( n52226, n52153, n52152 );
nand U83139 ( n52227, n52154, n52228 );
or U83140 ( n52228, n52152, n52153 );
nand U83141 ( n52621, n52715, n52716 );
nand U83142 ( n52716, n52581, n52586 );
nor U83143 ( n52715, n52577, n52583 );
nand U83144 ( n52152, n52241, n52242 );
nand U83145 ( n52242, n52091, n52096 );
nor U83146 ( n52241, n52087, n52093 );
nor U83147 ( n52562, n52563, n52564 );
nor U83148 ( n52563, n52565, n52566 );
nor U83149 ( n52565, n52567, n52568 );
nor U83150 ( n52159, n52160, n52161 );
nor U83151 ( n52160, n52162, n52163 );
nor U83152 ( n52162, n52164, n52165 );
not U83153 ( n1257, n51707 );
and U83154 ( n52761, n52972, n52973 );
nand U83155 ( n52973, n52974, n1443 );
nor U83156 ( n52972, n52975, n52976 );
nor U83157 ( n52975, n1473, n52982 );
nand U83158 ( n19880, n20254, n20255 );
nand U83159 ( n20254, n20259, n19886 );
nand U83160 ( n20255, n2700, n20256 );
nand U83161 ( n20259, n19883, n19885 );
not U83162 ( n2700, n19886 );
nand U83163 ( n18862, n19102, n19103 );
nand U83164 ( n19103, n18855, n18859 );
nor U83165 ( n19102, n18851, n18857 );
not U83166 ( n2407, n18855 );
or U83167 ( n52468, n52850, n52851 );
xor U83168 ( n53798, n53863, n53821 );
xnor U83169 ( n53863, n53820, n53819 );
nand U83170 ( n53802, n53798, n53797 );
xor U83171 ( n17962, n18220, n18150 );
xor U83172 ( n18220, n18151, n18148 );
xnor U83173 ( n18939, n18590, n18947 );
xor U83174 ( n18947, n18588, n18589 );
xor U83175 ( n16766, n17058, n17059 );
nand U83176 ( n17059, n17060, n17061 );
nand U83177 ( n17058, n17066, n17067 );
or U83178 ( n17060, n17064, n17065 );
nand U83179 ( n17067, n17068, n17069 );
nand U83180 ( n17069, n17070, n17071 );
nand U83181 ( n50050, n50365, n50366 );
nand U83182 ( n50365, n50369, n50065 );
nand U83183 ( n50366, n1319, n50367 );
nand U83184 ( n50369, n50062, n50064 );
not U83185 ( n1319, n50065 );
nand U83186 ( n19386, n19876, n19877 );
nand U83187 ( n19876, n19881, n19880 );
nand U83188 ( n19877, n19878, n19879 );
or U83189 ( n19878, n19880, n19881 );
xnor U83190 ( n20005, n20193, n20194 );
xnor U83191 ( n20193, n20195, n20196 );
nand U83192 ( n19992, n20124, n20125 );
nand U83193 ( n20124, n20067, n20066 );
nand U83194 ( n20125, n20068, n20126 );
or U83195 ( n20126, n20066, n20067 );
nand U83196 ( n20066, n20139, n20140 );
nand U83197 ( n20140, n20005, n20010 );
nor U83198 ( n20139, n20001, n20007 );
xor U83199 ( n52726, n53013, n53014 );
xor U83200 ( n53014, n53015, n53016 );
nand U83201 ( n52759, n52984, n52985 );
nand U83202 ( n52985, n52726, n52731 );
nor U83203 ( n52984, n52722, n52728 );
nand U83204 ( n52714, n52969, n52970 );
nand U83205 ( n52969, n52762, n52759 );
nand U83206 ( n52970, n52761, n52971 );
or U83207 ( n52971, n52759, n52762 );
and U83208 ( n52623, n52703, n52704 );
nand U83209 ( n52704, n52705, n1414 );
nor U83210 ( n52703, n52706, n52707 );
nor U83211 ( n52706, n1442, n52713 );
nand U83212 ( n20318, n20568, n2724 );
not U83213 ( n2724, n20560 );
nand U83214 ( n18553, n2553, n2582 );
xnor U83215 ( n52436, n51987, n52444 );
xor U83216 ( n52444, n51985, n51986 );
xnor U83217 ( n52423, n51974, n52431 );
xor U83218 ( n52431, n51972, n51973 );
or U83219 ( n52010, n52435, n52436 );
or U83220 ( n52014, n52422, n52423 );
xnor U83221 ( n52161, n52310, n52311 );
xnor U83222 ( n52310, n52312, n52313 );
xor U83223 ( n52387, n52396, n51924 );
xor U83224 ( n52396, n51926, n51927 );
nand U83225 ( n51926, n52486, n52487 );
nand U83226 ( n52487, n52488, n52489 );
or U83227 ( n52028, n52387, n52388 );
nand U83228 ( n20450, n20444, n20443 );
or U83229 ( n53801, n53797, n53798 );
nand U83230 ( n16747, n17093, n17094 );
or U83231 ( n17093, n17098, n17097 );
nand U83232 ( n17094, n17095, n17096 );
nand U83233 ( n17095, n17097, n17098 );
xor U83234 ( n53796, n53797, n53798 );
xor U83235 ( n52421, n52422, n52423 );
nand U83236 ( n19826, n19979, n19980 );
nand U83237 ( n19979, n19813, n19812 );
nand U83238 ( n19980, n19814, n19981 );
or U83239 ( n19981, n19812, n19813 );
nor U83240 ( n19986, n19987, n19988 );
nor U83241 ( n19987, n19989, n19990 );
nor U83242 ( n19989, n19991, n19992 );
nand U83243 ( n19236, n19553, n19554 );
nand U83244 ( n19553, n19558, n19402 );
nand U83245 ( n19554, n2445, n19555 );
nand U83246 ( n19558, n19399, n19401 );
nor U83247 ( n18885, n18886, n18887 );
nor U83248 ( n18886, n18888, n18889 );
nor U83249 ( n18888, n2377, n18890 );
and U83250 ( n16683, n18881, n18882 );
nand U83251 ( n18882, n18883, n2403 );
nor U83252 ( n18881, n18884, n18885 );
nor U83253 ( n18884, n2403, n18891 );
not U83254 ( n76, n15339 );
nand U83255 ( n51637, n51928, n1572 );
not U83256 ( n1572, n51920 );
nor U83257 ( n52690, n52691, n52692 );
nor U83258 ( n52691, n52693, n52694 );
nor U83259 ( n52693, n52695, n52696 );
xor U83260 ( n52434, n52435, n52436 );
nand U83261 ( n52016, n52423, n52422 );
nand U83262 ( n19552, n2468, n19547 );
nand U83263 ( n52012, n52436, n52435 );
nand U83264 ( n20062, n20156, n20157 );
nand U83265 ( n20157, n20022, n20026 );
nor U83266 ( n20156, n20018, n20024 );
not U83267 ( n2595, n20022 );
nand U83268 ( n20010, n20141, n20142 );
nand U83269 ( n20141, n20063, n20062 );
nand U83270 ( n20142, n20064, n20143 );
or U83271 ( n20143, n20062, n20063 );
and U83272 ( n20191, n20363, n20364 );
nand U83273 ( n20364, n20365, n2624 );
nor U83274 ( n20363, n20366, n20367 );
nor U83275 ( n20366, n20372, n20373 );
or U83276 ( n49748, n49755, n49756 );
xor U83277 ( n51021, n50775, n51029 );
xnor U83278 ( n51029, n50773, n50776 );
nand U83279 ( n50816, n51021, n51020 );
or U83280 ( n52697, n52695, n1412 );
nand U83281 ( n52478, n52480, n52481 );
nand U83282 ( n52480, n52484, n52485 );
nand U83283 ( n52481, n52482, n52483 );
or U83284 ( n52482, n52484, n52485 );
buf U83285 ( n76649, n8232 );
xnor U83286 ( n51273, n51044, n51281 );
xor U83287 ( n51281, n51042, n51043 );
nand U83288 ( n51032, n51273, n51272 );
or U83289 ( n17066, n17071, n17070 );
xor U83290 ( n51950, n51951, n51952 );
nand U83291 ( n51952, n51958, n51959 );
nand U83292 ( n51958, n51963, n51573 );
nand U83293 ( n51959, n1660, n51960 );
xor U83294 ( n51963, n51962, n51961 );
or U83295 ( n51572, n51962, n51961 );
xor U83296 ( n52401, n52402, n52403 );
nand U83297 ( n51561, n51936, n51937 );
nand U83298 ( n51936, n51940, n51941 );
nand U83299 ( n51937, n51938, n51939 );
or U83300 ( n51939, n51940, n51941 );
nand U83301 ( n49750, n49756, n49755 );
nor U83302 ( n52067, n52068, n52069 );
nor U83303 ( n52068, n52070, n52071 );
nor U83304 ( n52070, n52072, n52073 );
xor U83305 ( n52484, n52845, n52476 );
xor U83306 ( n52845, n52477, n52474 );
xor U83307 ( n52476, n52846, n52409 );
xor U83308 ( n52846, n52408, n52410 );
nand U83309 ( n52408, n52893, n52894 );
nand U83310 ( n52893, n52898, n52897 );
nand U83311 ( n52894, n52895, n52896 );
or U83312 ( n52896, n52897, n52898 );
and U83313 ( n52898, n53803, n53804 );
nand U83314 ( n53804, n52857, n1629 );
nor U83315 ( n53803, n53806, n53807 );
nor U83316 ( n53806, n53808, n53809 );
and U83317 ( n53807, n1645, n52858 );
nand U83318 ( n16768, n16770, n16771 );
nand U83319 ( n16770, n16780, n16781 );
nand U83320 ( n16771, n16772, n16773 );
nor U83321 ( n16780, n17055, n16778 );
nand U83322 ( n51627, n51951, n51952 );
xor U83323 ( n52269, n52616, n52617 );
xor U83324 ( n52617, n52618, n52619 );
nand U83325 ( n52256, n52572, n52573 );
nand U83326 ( n52572, n52304, n52303 );
nand U83327 ( n52573, n52305, n52574 );
or U83328 ( n52574, n52303, n52304 );
nand U83329 ( n52303, n52587, n52588 );
nand U83330 ( n52588, n52269, n52274 );
nor U83331 ( n52587, n52265, n52271 );
not U83332 ( n1445, n53012 );
nand U83333 ( n52731, n52986, n52987 );
or U83334 ( n52986, n52756, n52758 );
nand U83335 ( n52987, n52757, n52988 );
nand U83336 ( n52988, n52758, n52756 );
nand U83337 ( n52096, n52243, n52244 );
nand U83338 ( n52243, n52150, n52147 );
nand U83339 ( n52244, n52149, n52245 );
or U83340 ( n52245, n52147, n52150 );
nor U83341 ( n52250, n52251, n52252 );
nor U83342 ( n52251, n52253, n52254 );
nor U83343 ( n52253, n52255, n52256 );
nand U83344 ( n52756, n53001, n53002 );
nand U83345 ( n53002, n53003, n1445 );
nor U83346 ( n53001, n53004, n53005 );
nor U83347 ( n53004, n1475, n53011 );
and U83348 ( n52618, n52720, n52721 );
nand U83349 ( n52721, n52722, n1417 );
nor U83350 ( n52720, n52723, n52724 );
nor U83351 ( n52723, n1444, n52730 );
nand U83352 ( n51571, n51961, n51962 );
or U83353 ( n51625, n51952, n51951 );
nand U83354 ( n51832, n1265, n51831 );
nand U83355 ( n52863, n53816, n53817 );
nand U83356 ( n53816, n53821, n53820 );
nand U83357 ( n53817, n53818, n53819 );
or U83358 ( n53818, n53820, n53821 );
nand U83359 ( n49966, n50220, n50221 );
nand U83360 ( n50220, n50224, n50225 );
nand U83361 ( n50221, n50222, n50223 );
or U83362 ( n50223, n50224, n50225 );
or U83363 ( n50814, n51020, n51021 );
nand U83364 ( n19230, n2427, n19229 );
nand U83365 ( n20587, n8225, n20585 );
nor U83366 ( n20131, n20132, n20133 );
nor U83367 ( n20132, n20134, n20135 );
nor U83368 ( n20134, n20136, n20137 );
nand U83369 ( n52467, n52870, n52871 );
nand U83370 ( n52870, n52875, n52874 );
nand U83371 ( n52871, n52872, n52873 );
or U83372 ( n52872, n52874, n52875 );
xor U83373 ( n50481, n50482, n50483 );
xor U83374 ( n20258, n20266, n2734 );
xor U83375 ( n20266, n19891, n2715 );
nand U83376 ( n19885, n20258, n20257 );
nand U83377 ( n51503, n51639, n51640 );
nand U83378 ( n51639, n51644, n51643 );
nand U83379 ( n51640, n51641, n51642 );
or U83380 ( n51641, n51643, n51644 );
xnor U83381 ( n18952, n18688, n18960 );
xor U83382 ( n18960, n18686, n18687 );
nand U83383 ( n18589, n18948, n18949 );
nand U83384 ( n18948, n18953, n18692 );
nand U83385 ( n18949, n2633, n18950 );
nand U83386 ( n18953, n18689, n18691 );
nand U83387 ( n19073, n19286, n19287 );
nand U83388 ( n19287, n19288, n19289 );
nor U83389 ( n19286, n19290, n19291 );
nand U83390 ( n18686, n19070, n19071 );
nand U83391 ( n19071, n19072, n19073 );
or U83392 ( n20138, n20136, n2592 );
xor U83393 ( n52386, n52387, n52388 );
and U83394 ( n49597, n51685, n51686 );
nand U83395 ( n51685, n49549, n49551 );
nand U83396 ( n51686, n49552, n51687 );
or U83397 ( n51687, n49551, n49549 );
nand U83398 ( n52586, n52717, n52718 );
nand U83399 ( n52717, n52619, n52616 );
nand U83400 ( n52718, n52618, n52719 );
or U83401 ( n52719, n52616, n52619 );
xor U83402 ( n50856, n50923, n50665 );
xnor U83403 ( n50923, n50664, n50663 );
xor U83404 ( n52903, n52898, n53758 );
xnor U83405 ( n53758, n52895, n52897 );
nand U83406 ( n52026, n52388, n52387 );
nand U83407 ( n51337, n51359, n51360 );
nand U83408 ( n51359, n51364, n51332 );
nand U83409 ( n51360, n1460, n51361 );
nand U83410 ( n51364, n51329, n51331 );
nand U83411 ( n51332, n51365, n51366 );
nand U83412 ( n51365, n51370, n51369 );
nand U83413 ( n51366, n51367, n51368 );
or U83414 ( n51367, n51369, n51370 );
xnor U83415 ( n18583, n18591, n18424 );
xor U83416 ( n18591, n18426, n18427 );
nand U83417 ( n18413, n18579, n18580 );
nand U83418 ( n18580, n2612, n18581 );
nand U83419 ( n18579, n18584, n18552 );
not U83420 ( n2612, n18552 );
nand U83421 ( n18426, n18689, n18690 );
nand U83422 ( n18690, n18691, n18692 );
nand U83423 ( n18584, n18549, n18551 );
or U83424 ( n51030, n51272, n51273 );
nor U83425 ( n48749, n48483, n48719 );
not U83426 ( n2490, n19425 );
and U83427 ( n19521, n19580, n19581 );
nand U83428 ( n19581, n19425, n19429 );
nor U83429 ( n19580, n19421, n19427 );
nor U83430 ( n49311, n48483, n49280 );
nor U83431 ( n49120, n48483, n7834 );
nor U83432 ( n49042, n48483, n48995 );
nor U83433 ( n48947, n48483, n48896 );
nor U83434 ( n48660, n48483, n48629 );
nor U83435 ( n48582, n48483, n48535 );
nor U83436 ( n49404, n48483, n49358 );
nor U83437 ( n49215, n48483, n49184 );
nor U83438 ( n48846, n48483, n48815 );
nor U83439 ( n49598, n48483, n49462 );
nand U83440 ( n14856, n49578, n49579 );
nor U83441 ( n49579, n49580, n49581 );
nor U83442 ( n49578, n49598, n49599 );
nand U83443 ( n49581, n49582, n49583 );
nand U83444 ( n17814, n17822, n17823 );
nand U83445 ( n17822, n17827, n17555 );
nand U83446 ( n17823, n2853, n17824 );
xor U83447 ( n17827, n17826, n17825 );
nand U83448 ( n17546, n17813, n17814 );
nand U83449 ( n17923, n2368, n2402 );
not U83450 ( n2402, n17927 );
nand U83451 ( n18172, n19086, n19087 );
nand U83452 ( n19086, n19091, n19090 );
nand U83453 ( n19087, n19088, n19089 );
or U83454 ( n19088, n19090, n19091 );
not U83455 ( n335, n48474 );
nand U83456 ( n51628, n51954, n51955 );
nand U83457 ( n51954, n1625, n51957 );
or U83458 ( n51955, n51956, n1648 );
nor U83459 ( n51956, n51957, n1625 );
xnor U83460 ( n17901, n17710, n17965 );
xor U83461 ( n17965, n17709, n17708 );
nand U83462 ( n17709, n18146, n18147 );
nand U83463 ( n18146, n18150, n18151 );
nand U83464 ( n18147, n18148, n18149 );
or U83465 ( n18149, n18150, n18151 );
nand U83466 ( n52239, n52555, n52556 );
nand U83467 ( n52555, n52309, n52306 );
nand U83468 ( n52556, n52308, n52557 );
or U83469 ( n52557, n52306, n52309 );
nor U83470 ( n52233, n52234, n52235 );
nor U83471 ( n52234, n52236, n52237 );
nor U83472 ( n52236, n52238, n52239 );
and U83473 ( n52237, n52238, n52239 );
xnor U83474 ( n52024, n51940, n52398 );
xnor U83475 ( n52398, n51941, n51938 );
xor U83476 ( n18173, n18215, n18900 );
xnor U83477 ( n18900, n18213, n18214 );
not U83478 ( n2594, n20154 );
xor U83479 ( n17542, n17300, n17543 );
xnor U83480 ( n17543, n17301, n17299 );
nand U83481 ( n17286, n17534, n2833 );
nand U83482 ( n51947, n51631, n51633 );
nor U83483 ( n20148, n20149, n20150 );
nor U83484 ( n20149, n20151, n20152 );
nor U83485 ( n20151, n20153, n20154 );
xnor U83486 ( n52235, n52624, n52625 );
xnor U83487 ( n52624, n52626, n52627 );
and U83488 ( n52231, n52238, n52235 );
nand U83489 ( n52013, n52438, n52439 );
nand U83490 ( n52438, n52443, n52442 );
nand U83491 ( n52439, n52440, n52441 );
or U83492 ( n52440, n52442, n52443 );
nand U83493 ( n52017, n52425, n52426 );
nand U83494 ( n52425, n52430, n52429 );
nand U83495 ( n52426, n52427, n52428 );
or U83496 ( n52427, n52429, n52430 );
nand U83497 ( n53013, n53129, n53130 );
nand U83498 ( n53130, n53007, n53012 );
nor U83499 ( n53129, n53003, n53009 );
xnor U83500 ( n19591, n19811, n19812 );
xnor U83501 ( n19811, n19813, n19814 );
and U83502 ( n19675, n19725, n19726 );
nand U83503 ( n19726, n19591, n19596 );
nor U83504 ( n19725, n19587, n19593 );
nand U83505 ( n17288, n17542, n2828 );
not U83506 ( n2828, n17534 );
and U83507 ( n52305, n52575, n52576 );
nand U83508 ( n52576, n52577, n1380 );
nor U83509 ( n52575, n52578, n52579 );
nor U83510 ( n52578, n1415, n52585 );
xnor U83511 ( n50756, n50764, n50489 );
xor U83512 ( n50764, n50490, n50487 );
nand U83513 ( n49973, n50208, n50209 );
nand U83514 ( n50208, n50212, n50213 );
nand U83515 ( n50209, n50210, n50211 );
or U83516 ( n50211, n50212, n50213 );
nand U83517 ( n50213, n50544, n50545 );
nand U83518 ( n50544, n50549, n50548 );
nand U83519 ( n50545, n50546, n50547 );
or U83520 ( n50546, n50548, n50549 );
or U83521 ( n50475, n50755, n50756 );
or U83522 ( n19883, n20257, n20258 );
xor U83523 ( n50754, n50755, n50756 );
nand U83524 ( n20314, n20576, n20577 );
nand U83525 ( n20576, n20581, n20309 );
nand U83526 ( n20577, n2753, n20578 );
nand U83527 ( n20581, n20306, n20308 );
not U83528 ( n2753, n20309 );
xor U83529 ( n20279, n19924, n20287 );
xnor U83530 ( n20287, n19925, n19923 );
xnor U83531 ( n18965, n18600, n18973 );
xor U83532 ( n18973, n18598, n18599 );
nand U83533 ( n19001, n19379, n19380 );
nand U83534 ( n19380, n19381, n19382 );
nand U83535 ( n19314, n19322, n19323 );
nand U83536 ( n19323, n19000, n2768 );
nor U83537 ( n19322, n19326, n19327 );
nor U83538 ( n19326, n2750, n19329 );
nand U83539 ( n18978, n18986, n18987 );
or U83540 ( n18987, n18676, n18675 );
nor U83541 ( n18986, n18988, n18989 );
nor U83542 ( n18988, n18678, n18991 );
nand U83543 ( n18599, n18974, n18975 );
nand U83544 ( n18974, n18979, n18605 );
nand U83545 ( n18975, n2714, n18976 );
nand U83546 ( n18979, n18602, n18604 );
nand U83547 ( n18687, n18961, n18962 );
nand U83548 ( n18961, n18966, n18682 );
nand U83549 ( n18962, n2680, n18963 );
nand U83550 ( n18966, n18679, n18681 );
and U83551 ( n18989, n18678, n75764 );
xor U83552 ( n75764, n18675, n18677 );
nand U83553 ( n19064, n19313, n19314 );
nand U83554 ( n19909, n20275, n20276 );
nand U83555 ( n20275, n20280, n19946 );
nand U83556 ( n20276, n2773, n20277 );
nand U83557 ( n20280, n19943, n19945 );
xnor U83558 ( n20580, n20286, n20588 );
xor U83559 ( n20588, n20284, n20285 );
xnor U83560 ( n51975, n51590, n51976 );
xor U83561 ( n51976, n51588, n51589 );
xor U83562 ( n51966, n51967, n1678 );
xnor U83563 ( n19090, n19240, n19085 );
xnor U83564 ( n19240, n19084, n19082 );
nor U83565 ( n16785, n16786, n16787 );
nor U83566 ( n16786, n16788, n16789 );
nand U83567 ( n51638, n51922, n51923 );
nand U83568 ( n51922, n51927, n51926 );
nand U83569 ( n51923, n51924, n51925 );
or U83570 ( n51925, n51926, n51927 );
xor U83571 ( n20256, n20257, n20258 );
nand U83572 ( n51033, n51275, n51276 );
nand U83573 ( n51275, n51280, n51279 );
nand U83574 ( n51276, n51277, n51278 );
or U83575 ( n51277, n51279, n51280 );
nand U83576 ( n50817, n51023, n51024 );
nand U83577 ( n51023, n51028, n51027 );
nand U83578 ( n51024, n51025, n51026 );
or U83579 ( n51025, n51027, n51028 );
xnor U83580 ( n52141, n52302, n52303 );
xnor U83581 ( n52302, n52304, n52305 );
nand U83582 ( n50056, n50062, n50063 );
nand U83583 ( n50063, n50064, n50065 );
not U83584 ( n2802, n20297 );
nand U83585 ( n50477, n50756, n50755 );
xnor U83586 ( n52252, n52620, n52621 );
xnor U83587 ( n52620, n52622, n52623 );
nand U83588 ( n51940, n52472, n52473 );
nand U83589 ( n52472, n52476, n52477 );
nand U83590 ( n52473, n52474, n52475 );
or U83591 ( n52475, n52476, n52477 );
nand U83592 ( n51575, n51967, n1678 );
xnor U83593 ( n16644, n18877, n18878 );
xnor U83594 ( n18878, n18879, n18880 );
xnor U83595 ( n19608, n19807, n19808 );
xnor U83596 ( n19807, n19809, n19810 );
not U83597 ( n2454, n19205 );
nand U83598 ( n19596, n19727, n19728 );
nand U83599 ( n19727, n19670, n19669 );
nand U83600 ( n19728, n19671, n19729 );
or U83601 ( n19729, n19669, n19670 );
not U83602 ( n2408, n19117 );
and U83603 ( n19212, n19431, n19432 );
nand U83604 ( n19432, n19205, n19209 );
nor U83605 ( n19431, n19201, n19207 );
and U83606 ( n19810, n19999, n20000 );
nand U83607 ( n20000, n20001, n2562 );
nor U83608 ( n19999, n20002, n20003 );
nor U83609 ( n20002, n2593, n20009 );
and U83610 ( n19520, n19585, n19586 );
nand U83611 ( n19586, n19587, n2492 );
nor U83612 ( n19585, n19588, n19589 );
nor U83613 ( n19588, n2530, n19595 );
nand U83614 ( n52145, n52260, n52261 );
nand U83615 ( n52260, n52133, n52132 );
nand U83616 ( n52261, n52134, n52262 );
or U83617 ( n52262, n52132, n52133 );
not U83618 ( n1420, n52754 );
nand U83619 ( n52277, n52604, n52605 );
nand U83620 ( n52605, n52606, n1384 );
nor U83621 ( n52604, n52607, n52608 );
nor U83622 ( n52607, n1418, n52614 );
nand U83623 ( n52274, n52589, n52590 );
or U83624 ( n52589, n52277, n52280 );
nand U83625 ( n52590, n52279, n52591 );
nand U83626 ( n52591, n52280, n52277 );
nand U83627 ( n52615, n52734, n52735 );
or U83628 ( n52734, n52601, n52603 );
nand U83629 ( n52735, n52602, n52736 );
nand U83630 ( n52736, n52603, n52601 );
nand U83631 ( n52601, n52743, n52744 );
nand U83632 ( n52744, n52745, n1420 );
nor U83633 ( n52743, n52746, n52747 );
nor U83634 ( n52746, n1447, n52753 );
and U83635 ( n52134, n52263, n52264 );
nand U83636 ( n52264, n52265, n1343 );
nor U83637 ( n52263, n52266, n52267 );
nor U83638 ( n52266, n1382, n52273 );
nand U83639 ( n52022, n8237, n52478 );
or U83640 ( n17544, n17814, n17813 );
nor U83641 ( n19912, n76586, n2752 );
nand U83642 ( n19910, n20306, n20307 );
nand U83643 ( n20307, n20308, n20309 );
nand U83644 ( n17102, n17108, n17109 );
nand U83645 ( n17109, n17110, n17111 );
nand U83646 ( n52897, n53759, n53760 );
nand U83647 ( n53759, n53757, n53755 );
nand U83648 ( n53760, n53761, n53756 );
or U83649 ( n53761, n53755, n53757 );
xor U83650 ( n51271, n51272, n51273 );
nand U83651 ( n52616, n52732, n52733 );
nand U83652 ( n52733, n52610, n52615 );
nor U83653 ( n52732, n52606, n52612 );
not U83654 ( n2453, n19429 );
nor U83655 ( n19423, n19424, n19425 );
nor U83656 ( n19424, n19426, n19427 );
nor U83657 ( n19426, n19428, n19429 );
not U83658 ( n1475, n53007 );
nand U83659 ( n18958, n19281, n19282 );
nand U83660 ( n19281, n19285, n19073 );
nand U83661 ( n19282, n19283, n2658 );
nand U83662 ( n19285, n19070, n19072 );
xnor U83663 ( n18385, n18382, n18402 );
xor U83664 ( n18402, n18380, n18381 );
nand U83665 ( n52021, n52405, n52406 );
nand U83666 ( n52405, n52410, n52409 );
nand U83667 ( n52406, n52407, n52408 );
or U83668 ( n52407, n52409, n52410 );
xnor U83669 ( n19918, n19358, n19926 );
xor U83670 ( n19926, n19356, n19357 );
xnor U83671 ( n19905, n19341, n19913 );
xor U83672 ( n19913, n19339, n19340 );
nand U83673 ( n19381, n19905, n19904 );
nand U83674 ( n19919, n19343, n19345 );
nand U83675 ( n19340, n19914, n19915 );
nand U83676 ( n19915, n2787, n19916 );
nand U83677 ( n19914, n19919, n19346 );
not U83678 ( n2787, n19346 );
or U83679 ( n52240, n52238, n1338 );
not U83680 ( n2600, n20172 );
not U83681 ( n2564, n20026 );
and U83682 ( n20059, n20161, n20162 );
nand U83683 ( n20162, n20163, n2600 );
nor U83684 ( n20161, n20164, n20165 );
nor U83685 ( n20164, n20170, n20171 );
nor U83686 ( n15653, n15339, n5179 );
nand U83687 ( n18692, n18954, n18955 );
nand U83688 ( n18954, n18959, n18958 );
nand U83689 ( n18955, n18956, n18957 );
or U83690 ( n18956, n18958, n18959 );
nand U83691 ( n18552, n18585, n18586 );
nand U83692 ( n18585, n18590, n18589 );
nand U83693 ( n18586, n18587, n18588 );
or U83694 ( n18587, n18589, n18590 );
nand U83695 ( n20189, n20375, n20376 );
nand U83696 ( n20376, n2625, n20172 );
nor U83697 ( n20375, n20163, n20168 );
nand U83698 ( n49773, n49983, n49984 );
nand U83699 ( n49984, n49985, n49986 );
xor U83700 ( n51019, n51020, n51021 );
nand U83701 ( n50478, n50758, n50759 );
nand U83702 ( n50758, n50763, n50762 );
nand U83703 ( n50759, n50760, n50761 );
or U83704 ( n50760, n50762, n50763 );
nand U83705 ( n17858, n18086, n18087 );
nand U83706 ( n18086, n18091, n18090 );
nand U83707 ( n18087, n18088, n18089 );
or U83708 ( n18088, n18090, n18091 );
nor U83709 ( n16289, n15339, n16242 );
nor U83710 ( n16180, n15339, n16135 );
nor U83711 ( n16078, n15339, n16039 );
nor U83712 ( n15970, n15339, n15932 );
nor U83713 ( n15865, n15339, n15827 );
nor U83714 ( n15764, n15339, n15717 );
nor U83715 ( n15557, n15339, n15518 );
nor U83716 ( n15450, n15339, n15412 );
nor U83717 ( n16385, n15339, n16347 );
nor U83718 ( n16613, n15339, n5168 );
nand U83719 ( n8121, n16588, n16589 );
nor U83720 ( n16589, n16590, n16592 );
nor U83721 ( n16588, n16613, n16614 );
nand U83722 ( n16592, n16593, n16594 );
or U83723 ( n19379, n19904, n19905 );
nand U83724 ( n17820, n18080, n18081 );
nand U83725 ( n18080, n18085, n17858 );
nand U83726 ( n18081, n2848, n18082 );
nand U83727 ( n18085, n17855, n17857 );
nand U83728 ( n17547, n17816, n17817 );
nand U83729 ( n17816, n17820, n17821 );
nand U83730 ( n17817, n17818, n17819 );
or U83731 ( n17819, n17820, n17821 );
xnor U83732 ( n50212, n50224, n50474 );
xnor U83733 ( n50474, n50222, n50225 );
xor U83734 ( n51363, n51196, n51371 );
xnor U83735 ( n51371, n51194, n51197 );
xnor U83736 ( n51376, n51210, n51384 );
xor U83737 ( n51384, n51208, n51209 );
nand U83738 ( n51197, n51372, n51373 );
nand U83739 ( n51373, n1509, n51374 );
nand U83740 ( n51372, n51377, n51328 );
not U83741 ( n1509, n51328 );
nand U83742 ( n51377, n51325, n51327 );
nand U83743 ( n19740, n19996, n19997 );
nand U83744 ( n19996, n19809, n19808 );
nand U83745 ( n19997, n19810, n19998 );
or U83746 ( n19998, n19808, n19809 );
and U83747 ( n19738, n19739, n19740 );
or U83748 ( n19062, n19314, n19313 );
xor U83749 ( n17812, n17813, n17814 );
nand U83750 ( n17289, n17536, n17537 );
nand U83751 ( n17536, n17540, n17541 );
nand U83752 ( n17537, n17538, n17539 );
or U83753 ( n17539, n17540, n17541 );
xor U83754 ( n19284, n19293, n18969 );
xor U83755 ( n19293, n18971, n18972 );
nand U83756 ( n18971, n19383, n19384 );
nand U83757 ( n19384, n19385, n19386 );
nand U83758 ( n18876, n2382, n18875 );
not U83759 ( n2409, n18747 );
not U83760 ( n2370, n18859 );
and U83761 ( n18846, n19119, n19120 );
nand U83762 ( n19120, n18747, n18751 );
nor U83763 ( n19119, n18743, n18749 );
xnor U83764 ( n19736, n20065, n20066 );
xnor U83765 ( n20065, n20067, n20068 );
and U83766 ( n19732, n19739, n19736 );
nand U83767 ( n52409, n52847, n52848 );
nand U83768 ( n52848, n1627, n52849 );
nand U83769 ( n52847, n52852, n52471 );
xor U83770 ( n52849, n52850, n52851 );
nand U83771 ( n20357, n2623, n20356 );
nand U83772 ( n51577, n51975, n1667 );
not U83773 ( n1667, n51967 );
nor U83774 ( n19734, n19735, n19736 );
nor U83775 ( n19735, n19737, n19738 );
nor U83776 ( n19737, n19739, n19740 );
xor U83777 ( n51256, n51264, n51028 );
xnor U83778 ( n51264, n51027, n51026 );
nand U83779 ( n50822, n51067, n51068 );
nand U83780 ( n51067, n51072, n51071 );
nand U83781 ( n51068, n51069, n51070 );
or U83782 ( n51069, n51071, n51072 );
nand U83783 ( n50547, n50818, n50819 );
nand U83784 ( n50818, n50823, n50822 );
nand U83785 ( n50819, n50820, n50821 );
or U83786 ( n50821, n50822, n50823 );
or U83787 ( n51063, n51255, n51256 );
not U83788 ( n73, n15328 );
xor U83789 ( n17533, n17534, n2833 );
nand U83790 ( n17011, n17274, n17275 );
nand U83791 ( n17274, n17278, n17279 );
nand U83792 ( n17275, n17276, n17277 );
or U83793 ( n17277, n17278, n17279 );
and U83794 ( n49843, n49972, n49973 );
nor U83795 ( n49770, n49991, n49992 );
nor U83796 ( n49992, n49993, n49994 );
nor U83797 ( n49991, n49995, n49996 );
nand U83798 ( n51328, n51378, n51379 );
nand U83799 ( n51378, n51383, n51382 );
nand U83800 ( n51379, n51380, n51381 );
or U83801 ( n51381, n51382, n51383 );
nor U83802 ( n19111, n19112, n19113 );
nor U83803 ( n19112, n19114, n19115 );
nor U83804 ( n19114, n19116, n19117 );
or U83805 ( n19741, n19739, n2532 );
xnor U83806 ( n51389, n51319, n51397 );
xor U83807 ( n51397, n51318, n51320 );
nand U83808 ( n51402, n51551, n51552 );
nand U83809 ( n51551, n51556, n51555 );
nand U83810 ( n51552, n51553, n51554 );
or U83811 ( n51553, n51555, n51556 );
nand U83812 ( n51209, n51385, n51386 );
nand U83813 ( n51385, n51390, n51324 );
nand U83814 ( n51386, n1560, n51387 );
nand U83815 ( n51390, n51321, n51323 );
nand U83816 ( n51318, n51398, n51399 );
nand U83817 ( n51398, n51403, n51402 );
nand U83818 ( n51399, n51400, n51401 );
or U83819 ( n51401, n51402, n51403 );
xor U83820 ( n51457, n51465, n51280 );
xnor U83821 ( n51465, n51279, n51278 );
nand U83822 ( n51267, n51457, n51456 );
xnor U83823 ( n19753, n20061, n20062 );
xnor U83824 ( n20061, n20063, n20064 );
nand U83825 ( n19808, n20011, n20012 );
nand U83826 ( n20012, n19753, n19758 );
nor U83827 ( n20011, n19749, n19755 );
xor U83828 ( n19334, n19342, n19019 );
xnor U83829 ( n19342, n19018, n19017 );
xnor U83830 ( n19351, n19036, n19359 );
xor U83831 ( n19359, n19034, n19035 );
nand U83832 ( n19018, n19347, n19348 );
nand U83833 ( n19347, n19352, n19024 );
nand U83834 ( n19348, n2800, n19349 );
nand U83835 ( n19352, n19021, n19023 );
or U83836 ( n19058, n19333, n19334 );
xor U83837 ( n51787, n52147, n52148 );
xor U83838 ( n52148, n52149, n52150 );
nand U83839 ( n51725, n52082, n52083 );
nand U83840 ( n52082, n51795, n51794 );
nand U83841 ( n52083, n51796, n52084 );
or U83842 ( n52084, n51794, n51795 );
nand U83843 ( n51794, n52097, n52098 );
nand U83844 ( n52098, n51787, n51792 );
nor U83845 ( n52097, n51783, n51789 );
and U83846 ( n51723, n51724, n51725 );
xor U83847 ( n51254, n51255, n51256 );
xor U83848 ( n19332, n19333, n19334 );
nand U83849 ( n51578, n51969, n51970 );
nand U83850 ( n51969, n51974, n51973 );
nand U83851 ( n51970, n51971, n51972 );
or U83852 ( n51971, n51973, n51974 );
nand U83853 ( n19612, n19744, n19745 );
nand U83854 ( n19744, n19666, n19665 );
nand U83855 ( n19745, n19667, n19746 );
or U83856 ( n19746, n19665, n19666 );
nand U83857 ( n19758, n20013, n20014 );
nand U83858 ( n20013, n19805, n19804 );
nand U83859 ( n20014, n19806, n20015 );
or U83860 ( n20015, n19804, n19805 );
nor U83861 ( n20020, n20021, n20022 );
nor U83862 ( n20021, n20023, n20024 );
nor U83863 ( n20023, n20025, n20026 );
and U83864 ( n19667, n19747, n19748 );
nand U83865 ( n19748, n19749, n2534 );
nor U83866 ( n19747, n19750, n19751 );
nor U83867 ( n19750, n2563, n19757 );
nand U83868 ( n19060, n19334, n19333 );
xor U83869 ( n18994, n18995, n18996 );
nand U83870 ( n18996, n19002, n19003 );
nand U83871 ( n19002, n19007, n18621 );
nand U83872 ( n19003, n2782, n19004 );
xor U83873 ( n19007, n19006, n19005 );
or U83874 ( n18620, n19006, n19005 );
xor U83875 ( n50820, n50763, n51016 );
xor U83876 ( n51016, n50761, n50762 );
nand U83877 ( n19017, n19343, n19344 );
nand U83878 ( n19344, n19345, n19346 );
nand U83879 ( n17982, n18391, n2550 );
and U83880 ( n51796, n52085, n52086 );
nand U83881 ( n52086, n52087, n1297 );
nor U83882 ( n52085, n52088, n52089 );
nor U83883 ( n52088, n1339, n52095 );
xor U83884 ( n51107, n51177, n50934 );
xor U83885 ( n51177, n50932, n1398 );
xnor U83886 ( n19893, n20267, n19900 );
xnor U83887 ( n20267, n19899, n19897 );
not U83888 ( n2853, n17555 );
nor U83889 ( n48741, n48474, n48719 );
and U83890 ( n52758, n52989, n52990 );
nand U83891 ( n52990, n52749, n52754 );
nor U83892 ( n52989, n52745, n52751 );
nand U83893 ( n18610, n18995, n18996 );
nand U83894 ( n18619, n19005, n19006 );
or U83895 ( n18608, n18996, n18995 );
nand U83896 ( n51065, n51256, n51255 );
nor U83897 ( n49396, n48474, n49358 );
nor U83898 ( n49303, n48474, n49280 );
nor U83899 ( n49112, n48474, n7834 );
nor U83900 ( n49018, n48474, n48995 );
nor U83901 ( n48935, n48474, n48896 );
nor U83902 ( n48838, n48474, n48815 );
nor U83903 ( n48652, n48474, n48629 );
nor U83904 ( n48558, n48474, n48535 );
nor U83905 ( n49553, n48474, n49462 );
nor U83906 ( n49207, n48474, n49184 );
nand U83907 ( n14861, n49532, n49533 );
nor U83908 ( n49533, n49534, n49535 );
nor U83909 ( n49532, n49553, n49554 );
nand U83910 ( n49535, n49536, n49537 );
nand U83911 ( n19804, n20028, n20029 );
nand U83912 ( n20029, n19770, n19774 );
nor U83913 ( n20028, n19766, n19772 );
not U83914 ( n2565, n19770 );
not U83915 ( n2625, n20170 );
xor U83916 ( n19312, n19313, n19314 );
nand U83917 ( n18605, n18980, n18981 );
nand U83918 ( n18980, n18984, n18985 );
nand U83919 ( n18981, n18982, n18983 );
or U83920 ( n18983, n18984, n18985 );
nand U83921 ( n51792, n52099, n52100 );
nand U83922 ( n52099, n51778, n51779 );
nand U83923 ( n52100, n51780, n52101 );
or U83924 ( n52101, n51779, n51778 );
nor U83925 ( n52139, n52140, n52141 );
nor U83926 ( n52140, n52142, n52143 );
nor U83927 ( n52142, n52144, n52145 );
nand U83928 ( n18547, n18683, n18684 );
nand U83929 ( n18683, n18688, n18687 );
nand U83930 ( n18684, n18685, n18686 );
or U83931 ( n18685, n18687, n18688 );
nand U83932 ( n52074, n1310, n52073 );
nand U83933 ( n51624, n51982, n51983 );
nand U83934 ( n51982, n51987, n51986 );
nand U83935 ( n51983, n51984, n51985 );
or U83936 ( n51984, n51986, n51987 );
nand U83937 ( n19346, n19920, n19921 );
nand U83938 ( n19920, n19925, n19924 );
nand U83939 ( n19921, n19922, n19923 );
or U83940 ( n19922, n19924, n19925 );
xor U83941 ( n51501, n51549, n51393 );
xor U83942 ( n51549, n51395, n51396 );
xor U83943 ( n19301, n19308, n19887 );
xnor U83944 ( n19887, n19306, n19309 );
xnor U83945 ( n19625, n19803, n19804 );
xnor U83946 ( n19803, n19805, n19806 );
nand U83947 ( n19665, n19759, n19760 );
nand U83948 ( n19760, n19625, n19630 );
nor U83949 ( n19759, n19621, n19627 );
xnor U83950 ( n52610, n52755, n52756 );
xnor U83951 ( n52755, n52757, n52758 );
xor U83952 ( n52116, n52277, n52278 );
xor U83953 ( n52278, n52279, n52280 );
nand U83954 ( n52132, n52275, n52276 );
nand U83955 ( n52276, n52116, n52113 );
nor U83956 ( n52275, n52109, n52115 );
or U83957 ( n51265, n51456, n51457 );
xnor U83958 ( n18317, n18091, n18325 );
xor U83959 ( n18325, n18089, n18090 );
nand U83960 ( n17821, n18076, n18077 );
nand U83961 ( n18077, n18078, n18079 );
xnor U83962 ( n19135, n19513, n19514 );
xnor U83963 ( n19513, n19515, n19516 );
nand U83964 ( n19196, n19448, n19449 );
nand U83965 ( n19449, n19135, n19140 );
nor U83966 ( n19448, n19131, n19137 );
nor U83967 ( n19606, n19607, n19608 );
nor U83968 ( n19607, n19609, n19610 );
nor U83969 ( n19609, n19611, n19612 );
not U83970 ( n2410, n19209 );
not U83971 ( n2372, n18751 );
nor U83972 ( n19203, n19204, n19205 );
nor U83973 ( n19204, n19206, n19207 );
nor U83974 ( n19206, n19208, n19209 );
nand U83975 ( n19946, n20281, n20282 );
nand U83976 ( n20281, n20286, n20285 );
nand U83977 ( n20282, n20283, n20284 );
or U83978 ( n20283, n20285, n20286 );
nor U83979 ( n51809, n51810, n51811 );
nor U83980 ( n51810, n51812, n51813 );
nor U83981 ( n51812, n51814, n51815 );
xor U83982 ( n19068, n19303, n18984 );
xor U83983 ( n19303, n18985, n18982 );
nand U83984 ( n19339, n19943, n19944 );
nand U83985 ( n19944, n19945, n19946 );
nand U83986 ( n19070, n2655, n19284 );
nand U83987 ( n51196, n51505, n51506 );
nand U83988 ( n51506, n51507, n51508 );
xnor U83989 ( n50928, n50678, n50942 );
xor U83990 ( n50942, n50676, n50677 );
nand U83991 ( n50952, n51329, n51330 );
nand U83992 ( n51330, n51331, n51332 );
nor U83993 ( n51183, n50951, n1457 );
not U83994 ( n1457, n50954 );
nand U83995 ( n50663, n50924, n50925 );
nand U83996 ( n50925, n1397, n50926 );
nand U83997 ( n50924, n50929, n50851 );
not U83998 ( n1397, n50851 );
nand U83999 ( n50929, n50848, n50850 );
nand U84000 ( n50676, n51097, n51098 );
nand U84001 ( n51097, n51102, n51101 );
nand U84002 ( n51098, n51099, n51100 );
or U84003 ( n51099, n51101, n51102 );
xor U84004 ( n18067, n17820, n18075 );
xnor U84005 ( n18075, n17818, n17821 );
nand U84006 ( n17808, n18067, n18066 );
buf U84007 ( n76650, n8232 );
xnor U84008 ( n51721, n52151, n52152 );
xnor U84009 ( n52151, n52153, n52154 );
and U84010 ( n51717, n51724, n51721 );
xor U84011 ( n18150, n18221, n17976 );
xor U84012 ( n18221, n17974, n2518 );
not U84013 ( n2570, n20056 );
not U84014 ( n2537, n19774 );
nand U84015 ( n19800, n20045, n20046 );
nand U84016 ( n20046, n20047, n2570 );
nor U84017 ( n20045, n20048, n20049 );
nor U84018 ( n20048, n2602, n20055 );
not U84019 ( n1447, n52749 );
nand U84020 ( n18611, n18998, n18999 );
nand U84021 ( n18998, n2748, n19001 );
or U84022 ( n18999, n19000, n2768 );
nor U84023 ( n19000, n19001, n2748 );
xor U84024 ( n19283, n19284, n2655 );
nand U84025 ( n18682, n18967, n18968 );
nand U84026 ( n18967, n18972, n18971 );
nand U84027 ( n18968, n18969, n18970 );
or U84028 ( n18970, n18971, n18972 );
nand U84029 ( n17019, n17262, n17263 );
nand U84030 ( n17262, n17266, n17267 );
nand U84031 ( n17263, n17264, n17265 );
or U84032 ( n17265, n17266, n17267 );
xor U84033 ( n17804, n17540, n17805 );
xnor U84034 ( n17805, n17538, n17541 );
xor U84035 ( n17795, n17796, n2822 );
nand U84036 ( n17267, n17519, n17520 );
nand U84037 ( n17519, n17524, n17523 );
nand U84038 ( n17520, n17521, n17522 );
or U84039 ( n17521, n17523, n17524 );
xnor U84040 ( n19476, n19660, n19661 );
xnor U84041 ( n19660, n19662, n19663 );
nand U84042 ( n19463, n19616, n19617 );
nand U84043 ( n19616, n19511, n19510 );
nand U84044 ( n19617, n19512, n19618 );
or U84045 ( n19618, n19510, n19511 );
nand U84046 ( n19510, n19631, n19632 );
nand U84047 ( n19632, n19476, n19481 );
nor U84048 ( n19631, n19472, n19478 );
nand U84049 ( n19140, n19450, n19451 );
nand U84050 ( n19450, n19193, n19192 );
nand U84051 ( n19451, n19194, n19452 );
or U84052 ( n19452, n19192, n19193 );
nor U84053 ( n19768, n19769, n19770 );
nor U84054 ( n19769, n19771, n19772 );
nor U84055 ( n19771, n19773, n19774 );
nor U84056 ( n19457, n19458, n19459 );
nor U84057 ( n19458, n19460, n19461 );
nor U84058 ( n19460, n19462, n19463 );
nand U84059 ( n19630, n19761, n19762 );
nand U84060 ( n19761, n19662, n19661 );
nand U84061 ( n19762, n19663, n19763 );
or U84062 ( n19763, n19661, n19662 );
and U84063 ( n19295, n19297, n19298 );
or U84064 ( n19297, n19301, n19302 );
nand U84065 ( n19298, n19299, n19300 );
nand U84066 ( n19299, n19301, n19302 );
nand U84067 ( n17620, n17705, n17706 );
nand U84068 ( n17705, n17710, n17709 );
nand U84069 ( n17706, n17707, n17708 );
or U84070 ( n17707, n17709, n17710 );
nand U84071 ( n17419, n17699, n17700 );
nand U84072 ( n17699, n17704, n17620 );
nand U84073 ( n17700, n2483, n17701 );
nand U84074 ( n17704, n17617, n17619 );
and U84075 ( n19512, n19619, n19620 );
nand U84076 ( n19620, n19621, n2497 );
nor U84077 ( n19619, n19622, n19623 );
nor U84078 ( n19622, n2535, n19629 );
nand U84079 ( n19189, n19467, n19468 );
nand U84080 ( n19467, n19178, n19175 );
nand U84081 ( n19468, n19177, n19469 );
or U84082 ( n19469, n19175, n19178 );
nand U84083 ( n19645, n19787, n19788 );
nand U84084 ( n19788, n19789, n2540 );
nor U84085 ( n19787, n19790, n19791 );
nor U84086 ( n19790, n2572, n19797 );
not U84087 ( n2540, n19798 );
nand U84088 ( n19481, n19633, n19634 );
nand U84089 ( n19633, n19485, n19486 );
nand U84090 ( n19634, n19487, n19635 );
or U84091 ( n19635, n19486, n19485 );
nor U84092 ( n19652, n19653, n19654 );
nor U84093 ( n19653, n19655, n19656 );
nor U84094 ( n19655, n19657, n19658 );
not U84095 ( n2499, n19658 );
and U84096 ( n19177, n19470, n19471 );
nand U84097 ( n19471, n19472, n2462 );
nor U84098 ( n19470, n19473, n19474 );
nor U84099 ( n19473, n2498, n19480 );
and U84100 ( n19899, n20310, n20311 );
nand U84101 ( n20310, n20315, n20314 );
nand U84102 ( n20311, n20312, n20313 );
or U84103 ( n20312, n20314, n20315 );
nand U84104 ( n20155, n2599, n20154 );
nand U84105 ( n18991, n18675, n18677 );
nand U84106 ( n19061, n19336, n19337 );
nand U84107 ( n19336, n19341, n19340 );
nand U84108 ( n19337, n19338, n19339 );
or U84109 ( n19338, n19340, n19341 );
or U84110 ( n16793, n16800, n16801 );
nand U84111 ( n16610, n18729, n18730 );
nand U84112 ( n18729, n16572, n16574 );
nand U84113 ( n18730, n16575, n18731 );
or U84114 ( n18731, n16574, n16572 );
nand U84115 ( n50373, n50654, n50655 );
nand U84116 ( n50654, n50659, n50577 );
nand U84117 ( n50655, n1367, n50656 );
nand U84118 ( n50659, n50574, n50576 );
nand U84119 ( n50577, n50660, n50661 );
nand U84120 ( n50660, n50665, n50664 );
nand U84121 ( n50661, n50662, n50663 );
or U84122 ( n50662, n50664, n50665 );
xnor U84123 ( n19308, n19320, n19894 );
xnor U84124 ( n19894, n19321, n19319 );
nand U84125 ( n19319, n19895, n19896 );
or U84126 ( n19895, n19900, n19899 );
nand U84127 ( n19896, n19897, n19898 );
nand U84128 ( n19898, n19899, n19900 );
xnor U84129 ( n51440, n51448, n51262 );
xor U84130 ( n51448, n51261, n51263 );
xor U84131 ( n51455, n51456, n51457 );
nand U84132 ( n51250, n51440, n51439 );
xnor U84133 ( n19442, n19668, n19669 );
xnor U84134 ( n19668, n19670, n19671 );
and U84135 ( n19438, n19445, n19442 );
nand U84136 ( n17527, n17796, n2822 );
nand U84137 ( n16795, n16801, n16800 );
nand U84138 ( n50851, n50930, n50931 );
nand U84139 ( n50931, n1398, n50932 );
nand U84140 ( n50930, n50933, n50934 );
nor U84141 ( n50933, n50935, n50936 );
xnor U84142 ( n19185, n19509, n19510 );
xnor U84143 ( n19509, n19511, n19512 );
not U84144 ( n1388, n52740 );
nand U84145 ( n52295, n52594, n52595 );
or U84146 ( n52594, n52599, n52598 );
nand U84147 ( n52595, n52596, n52597 );
nand U84148 ( n52597, n52598, n52599 );
nand U84149 ( n52599, n53960, n53961 );
nand U84150 ( n53961, n52741, n1388 );
nor U84151 ( n53960, n53963, n53964 );
nor U84152 ( n53963, n1419, n53967 );
and U84153 ( n52280, n52592, n52593 );
nand U84154 ( n52593, n52290, n52295 );
nor U84155 ( n52592, n52286, n52292 );
or U84156 ( n17806, n18066, n18067 );
nand U84157 ( n51324, n51391, n51392 );
nand U84158 ( n51391, n51396, n51395 );
nand U84159 ( n51392, n51393, n51394 );
or U84160 ( n51394, n51395, n51396 );
and U84161 ( n52603, n52737, n52738 );
nand U84162 ( n52738, n52739, n52740 );
nor U84163 ( n52737, n52741, n52742 );
nor U84164 ( n15643, n15328, n5179 );
nand U84165 ( n19024, n19353, n19354 );
nand U84166 ( n19353, n19358, n19357 );
nand U84167 ( n19354, n19355, n19356 );
or U84168 ( n19355, n19357, n19358 );
nand U84169 ( n18381, n18403, n18404 );
nand U84170 ( n18403, n18408, n18376 );
nand U84171 ( n18404, n2583, n18405 );
nand U84172 ( n18408, n18373, n18375 );
nand U84173 ( n18376, n18409, n18410 );
nand U84174 ( n18409, n18414, n18413 );
nand U84175 ( n18410, n18411, n18412 );
or U84176 ( n18411, n18413, n18414 );
nand U84177 ( n51496, n51558, n51559 );
nand U84178 ( n51559, n51560, n51561 );
and U84179 ( n20057, n20173, n20174 );
nand U84180 ( n20174, n20051, n20056 );
nor U84181 ( n20173, n20047, n20053 );
nor U84182 ( n16375, n15328, n16347 );
nor U84183 ( n16279, n15328, n16242 );
nor U84184 ( n16068, n15328, n16039 );
nor U84185 ( n15960, n15328, n15932 );
nor U84186 ( n15855, n15328, n15827 );
nor U84187 ( n15547, n15328, n15518 );
nor U84188 ( n15440, n15328, n15412 );
nor U84189 ( n16170, n15328, n16135 );
nor U84190 ( n15754, n15328, n15717 );
nand U84191 ( n19446, n19599, n19600 );
nand U84192 ( n19599, n19515, n19514 );
nand U84193 ( n19600, n19516, n19601 );
or U84194 ( n19601, n19514, n19515 );
nor U84195 ( n19440, n19441, n19442 );
nor U84196 ( n19441, n19443, n19444 );
nor U84197 ( n19443, n19445, n19446 );
nor U84198 ( n16577, n15328, n5168 );
nand U84199 ( n8126, n16550, n16552 );
nor U84200 ( n16552, n16553, n16554 );
nor U84201 ( n16550, n16577, n16578 );
nand U84202 ( n16554, n16555, n16557 );
and U84203 ( n19444, n19445, n19446 );
xnor U84204 ( n17266, n17278, n17526 );
xnor U84205 ( n17526, n17276, n17279 );
xor U84206 ( n19012, n19020, n18634 );
xnor U84207 ( n19020, n18633, n18632 );
nand U84208 ( n18632, n19021, n19022 );
nand U84209 ( n19022, n19023, n19024 );
or U84210 ( n18669, n19011, n19012 );
nand U84211 ( n19661, n19776, n19777 );
nand U84212 ( n19777, n19654, n19658 );
nor U84213 ( n19776, n19650, n19656 );
nand U84214 ( n51268, n51459, n51460 );
nand U84215 ( n51459, n51464, n51463 );
nand U84216 ( n51460, n51461, n51462 );
or U84217 ( n51461, n51463, n51464 );
xor U84218 ( n19010, n19011, n19012 );
nand U84219 ( n18079, n18319, n18320 );
nand U84220 ( n18319, n18324, n18323 );
nand U84221 ( n18320, n18321, n18322 );
or U84222 ( n18321, n18323, n18324 );
nand U84223 ( n17809, n18069, n18070 );
nand U84224 ( n18069, n18074, n18073 );
nand U84225 ( n18070, n18071, n18072 );
or U84226 ( n18071, n18073, n18074 );
nand U84227 ( n18318, n18076, n18078 );
nand U84228 ( n18073, n18313, n18314 );
nand U84229 ( n18314, n2838, n18315 );
nand U84230 ( n18313, n18318, n18079 );
not U84231 ( n2838, n18079 );
nand U84232 ( n18671, n19012, n19011 );
xnor U84233 ( n50200, n50473, n50212 );
xor U84234 ( n50473, n50213, n50210 );
not U84235 ( n1675, n49977 );
xnor U84236 ( n51745, n52131, n52132 );
xnor U84237 ( n52131, n52133, n52134 );
xnor U84238 ( n19459, n19664, n19665 );
xnor U84239 ( n19664, n19666, n19667 );
or U84240 ( n51248, n51439, n51440 );
xnor U84241 ( n52290, n52600, n52601 );
xnor U84242 ( n52600, n52602, n52603 );
or U84243 ( n19447, n19445, n2455 );
nand U84244 ( n19430, n2469, n19429 );
xnor U84245 ( n50376, n50077, n50377 );
xor U84246 ( n50377, n50075, n50076 );
xor U84247 ( n50367, n50368, n1360 );
nand U84248 ( n50075, n50574, n50575 );
nand U84249 ( n50575, n50576, n50577 );
xor U84250 ( n20738, n20739, n2758 );
nand U84251 ( n51066, n51258, n51259 );
nand U84252 ( n51258, n51263, n51262 );
nand U84253 ( n51259, n51260, n51261 );
or U84254 ( n51260, n51262, n51263 );
not U84255 ( n1419, n52739 );
and U84256 ( n16888, n17018, n17019 );
not U84257 ( n2602, n20051 );
nand U84258 ( n17529, n17804, n2818 );
not U84259 ( n2818, n17796 );
xor U84260 ( n18407, n18240, n18415 );
xnor U84261 ( n18415, n18238, n18241 );
xnor U84262 ( n18420, n18258, n18428 );
xor U84263 ( n18428, n18256, n18257 );
xnor U84264 ( n18433, n18367, n18441 );
xor U84265 ( n18441, n18366, n18368 );
nand U84266 ( n18241, n18416, n18417 );
nand U84267 ( n18417, n2632, n18418 );
nand U84268 ( n18416, n18421, n18246 );
not U84269 ( n2632, n18246 );
nand U84270 ( n18446, n18595, n18596 );
nand U84271 ( n18595, n18600, n18599 );
nand U84272 ( n18596, n18597, n18598 );
or U84273 ( n18597, n18599, n18600 );
nand U84274 ( n18257, n18429, n18430 );
nand U84275 ( n18429, n18434, n18372 );
nand U84276 ( n18430, n2677, n18431 );
nand U84277 ( n18434, n18369, n18371 );
nand U84278 ( n18421, n18243, n18245 );
xor U84279 ( n19903, n19904, n19905 );
nand U84280 ( n19320, n19901, n19902 );
nand U84281 ( n19901, n19906, n19382 );
nand U84282 ( n19902, n2749, n19903 );
nand U84283 ( n19906, n19379, n19381 );
nand U84284 ( n19065, n19316, n19317 );
nand U84285 ( n19316, n19321, n19320 );
nand U84286 ( n19317, n19318, n19319 );
or U84287 ( n19318, n19320, n19321 );
nand U84288 ( n20673, n2758, n20739 );
xor U84289 ( n51596, n51604, n51464 );
xnor U84290 ( n51604, n51463, n51462 );
nand U84291 ( n51451, n51596, n51595 );
xor U84292 ( n18545, n18593, n18437 );
xor U84293 ( n18593, n18439, n18440 );
nand U84294 ( n18439, n18679, n18680 );
nand U84295 ( n18680, n18681, n18682 );
not U84296 ( n2749, n19382 );
nand U84297 ( n50062, n50368, n1360 );
buf U84298 ( n76656, n8224 );
xnor U84299 ( n51393, n51400, n51550 );
xnor U84300 ( n51550, n51403, n51402 );
nand U84301 ( n17930, n17931, n17927 );
nor U84302 ( n17931, n8214, n8213 );
xor U84303 ( n51185, n50952, n50951 );
xnor U84304 ( n50743, n50549, n50751 );
xor U84305 ( n50751, n50547, n50548 );
nand U84306 ( n50199, n50469, n50470 );
nand U84307 ( n50470, n50471, n50472 );
nand U84308 ( n51251, n51442, n51443 );
nand U84309 ( n51442, n51447, n51446 );
nand U84310 ( n51443, n51444, n51445 );
or U84311 ( n51444, n51446, n51447 );
or U84312 ( n51449, n51595, n51596 );
xnor U84313 ( n50934, n51102, n51178 );
xnor U84314 ( n51178, n51100, n51101 );
nand U84315 ( n52113, n52281, n52282 );
nand U84316 ( n52281, n52129, n52128 );
nand U84317 ( n52282, n52130, n52283 );
or U84318 ( n52283, n52128, n52129 );
and U84319 ( n52109, n1302, n52113 );
and U84320 ( n52130, n52284, n52285 );
nand U84321 ( n52285, n52286, n1347 );
nor U84322 ( n52284, n52287, n52288 );
nor U84323 ( n52287, n1385, n52294 );
nand U84324 ( n18672, n19014, n19015 );
nand U84325 ( n19014, n19019, n19018 );
nand U84326 ( n19015, n19016, n19017 );
or U84327 ( n19016, n19018, n19019 );
buf U84328 ( n76652, n8230 );
not U84329 ( n330, n48465 );
xor U84330 ( n49529, n49530, n49531 );
nand U84331 ( n18246, n18422, n18423 );
nand U84332 ( n18422, n18427, n18426 );
nand U84333 ( n18423, n18424, n18425 );
or U84334 ( n18425, n18426, n18427 );
xor U84335 ( n18300, n18308, n18074 );
xnor U84336 ( n18308, n18073, n18072 );
nand U84337 ( n17863, n18114, n18115 );
nand U84338 ( n18114, n18119, n18118 );
nand U84339 ( n18115, n18116, n18117 );
or U84340 ( n18116, n18118, n18119 );
nand U84341 ( n17522, n17859, n17860 );
nand U84342 ( n17859, n17864, n17863 );
nand U84343 ( n17860, n17861, n17862 );
or U84344 ( n17862, n17863, n17864 );
or U84345 ( n18110, n18299, n18300 );
nand U84346 ( n18984, n19304, n19305 );
nand U84347 ( n19304, n19308, n19309 );
nand U84348 ( n19305, n19306, n19307 );
or U84349 ( n19307, n19308, n19309 );
nand U84350 ( n17530, n17798, n17799 );
nand U84351 ( n17798, n17803, n17802 );
nand U84352 ( n17799, n17800, n17801 );
or U84353 ( n17800, n17802, n17803 );
xnor U84354 ( n50658, n50389, n50666 );
xor U84355 ( n50666, n50387, n50388 );
nand U84356 ( n50387, n50848, n50849 );
nand U84357 ( n50849, n50850, n50851 );
xor U84358 ( n18065, n18066, n18067 );
nand U84359 ( n19118, n2428, n19117 );
xnor U84360 ( n51497, n51562, n51491 );
xor U84361 ( n51562, n51492, n51489 );
xnor U84362 ( n51319, n51404, n51216 );
xor U84363 ( n51404, n51218, n51219 );
nand U84364 ( n51492, n51629, n51630 );
nand U84365 ( n51629, n51633, n51634 );
nand U84366 ( n51630, n51631, n51632 );
and U84367 ( n19802, n20033, n20034 );
nand U84368 ( n20034, n19793, n19798 );
nor U84369 ( n20033, n19789, n19795 );
nand U84370 ( n16818, n17029, n17030 );
nand U84371 ( n17030, n17031, n17032 );
nand U84372 ( n50807, n51059, n51060 );
nand U84373 ( n51060, n51061, n1740 );
not U84374 ( n1740, n51062 );
xnor U84375 ( n18497, n18324, n18505 );
xor U84376 ( n18505, n18322, n18323 );
nand U84377 ( n18072, n18309, n18310 );
nand U84378 ( n18310, n18311, n18312 );
xor U84379 ( n18298, n18299, n18300 );
xnor U84380 ( n17414, n17122, n17422 );
xor U84381 ( n17422, n17120, n17121 );
xor U84382 ( n17412, n17413, n17414 );
nand U84383 ( n17120, n17617, n17618 );
nand U84384 ( n17618, n17619, n17620 );
nor U84385 ( n51290, n51061, n51062 );
nand U84386 ( n51043, n51282, n51283 );
nand U84387 ( n51283, n51061, n51284 );
nand U84388 ( n51282, n51290, n51059 );
nand U84389 ( n51284, n51285, n51286 );
nand U84390 ( n17896, n17972, n17973 );
nand U84391 ( n17973, n2518, n17974 );
nand U84392 ( n17972, n17975, n17976 );
nor U84393 ( n17975, n17977, n17978 );
nand U84394 ( n17708, n17966, n17967 );
nand U84395 ( n17966, n17971, n17896 );
nand U84396 ( n17967, n2517, n17968 );
nand U84397 ( n17971, n17893, n17895 );
or U84398 ( n17108, n17413, n17414 );
nand U84399 ( n50677, n50943, n50944 );
nand U84400 ( n50943, n50948, n50847 );
nand U84401 ( n50944, n1454, n50945 );
nand U84402 ( n50948, n50844, n50846 );
not U84403 ( n1454, n50847 );
nand U84404 ( n50064, n50376, n1355 );
not U84405 ( n1355, n50368 );
nand U84406 ( n18843, n19124, n19125 );
nand U84407 ( n19125, n18765, n18769 );
nor U84408 ( n19124, n18761, n18767 );
nand U84409 ( n18836, n19143, n19144 );
or U84410 ( n19143, n18821, n18824 );
nand U84411 ( n19144, n18823, n19145 );
nand U84412 ( n19145, n18824, n18821 );
nor U84413 ( n19183, n19184, n19185 );
nor U84414 ( n19184, n19186, n19187 );
nor U84415 ( n19186, n19188, n19189 );
and U84416 ( n18767, n18768, n18769 );
and U84417 ( n18838, n19141, n19142 );
nand U84418 ( n19142, n18831, n18836 );
nor U84419 ( n19141, n18827, n18833 );
nor U84420 ( n18853, n18854, n18855 );
nor U84421 ( n18854, n18856, n18857 );
nor U84422 ( n18856, n18858, n18859 );
xor U84423 ( n51594, n51595, n51596 );
xnor U84424 ( n51988, n51603, n51989 );
xor U84425 ( n51989, n51601, n51602 );
xor U84426 ( n51979, n51980, n1694 );
nor U84427 ( n51999, n51608, n51992 );
nand U84428 ( n51602, n51990, n51991 );
nand U84429 ( n51991, n51992, n51993 );
nand U84430 ( n51990, n51999, n51605 );
nor U84431 ( n51993, n51994, n51995 );
nand U84432 ( n20027, n2569, n20026 );
not U84433 ( n2504, n19784 );
and U84434 ( n19647, n19781, n19782 );
nand U84435 ( n19782, n19783, n19784 );
nor U84436 ( n19781, n19785, n19786 );
not U84437 ( n2538, n19654 );
nand U84438 ( n19210, n2429, n19209 );
xor U84439 ( n19160, n19484, n19485 );
xor U84440 ( n19484, n19486, n19487 );
nand U84441 ( n19175, n19482, n19483 );
nand U84442 ( n19483, n19160, n19157 );
nor U84443 ( n19482, n19153, n19159 );
nor U84444 ( n52454, n52009, n52447 );
nand U84445 ( n51986, n52445, n52446 );
nand U84446 ( n52446, n52447, n52448 );
nand U84447 ( n52445, n52454, n52006 );
nor U84448 ( n52448, n52449, n52450 );
nand U84449 ( n51816, n1267, n51815 );
nand U84450 ( n18112, n18300, n18299 );
nand U84451 ( n17110, n17414, n17413 );
nand U84452 ( n51749, n52104, n52105 );
or U84453 ( n52104, n51775, n51774 );
nand U84454 ( n52105, n51776, n52106 );
nand U84455 ( n52106, n51774, n51775 );
nor U84456 ( n52111, n52112, n52113 );
nor U84457 ( n52112, n52114, n52115 );
nor U84458 ( n52114, n1302, n52116 );
and U84459 ( n51776, n52107, n52108 );
nand U84460 ( n52108, n52109, n1344 );
nor U84461 ( n52107, n52110, n52111 );
nor U84462 ( n52110, n1344, n52117 );
nand U84463 ( n50186, n50459, n1673 );
not U84464 ( n1673, n50467 );
not U84465 ( n1348, n53985 );
and U84466 ( n52598, n53982, n53983 );
nand U84467 ( n53983, n53984, n53985 );
nor U84468 ( n53982, n53986, n53987 );
nor U84469 ( n16815, n17037, n17038 );
nor U84470 ( n17038, n17039, n17040 );
nor U84471 ( n17037, n17041, n17042 );
nand U84472 ( n51621, n51980, n1694 );
nand U84473 ( n18372, n18435, n18436 );
nand U84474 ( n18435, n18440, n18439 );
nand U84475 ( n18436, n18437, n18438 );
or U84476 ( n18438, n18439, n18440 );
and U84477 ( n18840, n19129, n19130 );
nand U84478 ( n19130, n19131, n2413 );
nor U84479 ( n19129, n19132, n19133 );
nor U84480 ( n19132, n2457, n19139 );
nand U84481 ( n52128, n52296, n52297 );
nand U84482 ( n52297, n52298, n52299 );
nor U84483 ( n52296, n52300, n52301 );
nand U84484 ( n53958, n54037, n54038 );
nand U84485 ( n54038, n53986, n1348 );
nor U84486 ( n54037, n54040, n54041 );
nor U84487 ( n54040, n1387, n54044 );
nand U84488 ( n52299, n53953, n53954 );
or U84489 ( n53953, n53958, n53957 );
nand U84490 ( n53954, n53955, n53956 );
nand U84491 ( n53956, n53957, n53958 );
nand U84492 ( n50188, n50467, n1669 );
not U84493 ( n1669, n50459 );
nand U84494 ( n19486, n19636, n19637 );
nand U84495 ( n19637, n19497, n19501 );
nor U84496 ( n19636, n19493, n19499 );
not U84497 ( n2464, n19501 );
nand U84498 ( n19643, n21065, n21066 );
nand U84499 ( n21066, n19785, n2504 );
nor U84500 ( n21065, n21068, n21069 );
nor U84501 ( n21068, n2539, n21072 );
nand U84502 ( n18240, n18549, n18550 );
nand U84503 ( n18550, n18551, n18552 );
nand U84504 ( n49774, n49775, n49776 );
nand U84505 ( n49776, n1608, n49777 );
nand U84506 ( n49775, n49782, n49783 );
nand U84507 ( n49777, n49778, n49779 );
nand U84508 ( n49783, n49784, n49785 );
nand U84509 ( n49784, n49787, n49780 );
or U84510 ( n49785, n49786, n1594 );
xor U84511 ( n18789, n19175, n19176 );
xor U84512 ( n19176, n19177, n19178 );
xnor U84513 ( n18831, n19191, n19192 );
xnor U84514 ( n19191, n19193, n19194 );
xor U84515 ( n51239, n51247, n51072 );
xnor U84516 ( n51247, n51071, n51070 );
nand U84517 ( n50472, n50745, n50746 );
nand U84518 ( n50745, n50750, n50749 );
nand U84519 ( n50746, n50747, n50748 );
or U84520 ( n50748, n50749, n50750 );
nand U84521 ( n51075, n51239, n51238 );
nand U84522 ( n50465, n50739, n50740 );
nand U84523 ( n50739, n50744, n50472 );
nand U84524 ( n50740, n1683, n50741 );
nand U84525 ( n50744, n50469, n50471 );
nand U84526 ( n50189, n50461, n50462 );
nand U84527 ( n50461, n50466, n50465 );
nand U84528 ( n50462, n50463, n50464 );
or U84529 ( n50463, n50465, n50466 );
nand U84530 ( n51100, n51333, n51334 );
nand U84531 ( n51333, n51338, n51337 );
nand U84532 ( n51334, n51335, n51336 );
or U84533 ( n51335, n51337, n51338 );
nand U84534 ( n18633, n19025, n19026 );
nand U84535 ( n19025, n19030, n18668 );
nand U84536 ( n19026, n2808, n19027 );
nand U84537 ( n19030, n18665, n18667 );
nand U84538 ( n18668, n19031, n19032 );
nand U84539 ( n19031, n19036, n19035 );
nand U84540 ( n19032, n19033, n19034 );
or U84541 ( n19033, n19035, n19036 );
xor U84542 ( n17861, n17803, n18062 );
xor U84543 ( n18062, n17801, n17802 );
nand U84544 ( n19775, n2544, n19774 );
nand U84545 ( n18540, n18602, n18603 );
nand U84546 ( n18603, n18604, n18605 );
not U84547 ( n2572, n19793 );
xor U84548 ( n17254, n17266, n17518 );
xnor U84549 ( n17518, n17264, n17267 );
not U84550 ( n2794, n17023 );
not U84551 ( n1387, n53984 );
xor U84552 ( n18484, n18306, n18492 );
xnor U84553 ( n18492, n18307, n18305 );
nand U84554 ( n18347, n18484, n18483 );
nand U84555 ( n18305, n18493, n18494 );
nand U84556 ( n18493, n18498, n18312 );
nand U84557 ( n18494, n2825, n18495 );
nand U84558 ( n18498, n18309, n18311 );
nor U84559 ( n51701, n51702, n51703 );
nor U84560 ( n51702, n51704, n51705 );
nor U84561 ( n51704, n51706, n51707 );
nand U84562 ( n49521, n51691, n51692 );
or U84563 ( n51691, n49490, n49493 );
nand U84564 ( n51692, n49492, n51693 );
nand U84565 ( n51693, n49493, n49490 );
xnor U84566 ( n17703, n17434, n17711 );
xor U84567 ( n17711, n17432, n17433 );
nand U84568 ( n17432, n17893, n17894 );
nand U84569 ( n17894, n17895, n17896 );
and U84570 ( n18761, n18768, n18765 );
nand U84571 ( n19659, n2509, n19658 );
not U84572 ( n2539, n19783 );
nand U84573 ( n50037, n50072, n50073 );
nand U84574 ( n50072, n50077, n50076 );
nand U84575 ( n50073, n50074, n50075 );
or U84576 ( n50074, n50076, n50077 );
nand U84577 ( n51623, n51988, n1690 );
not U84578 ( n1690, n51980 );
or U84579 ( n51073, n51238, n51239 );
xnor U84580 ( n51203, n51211, n50976 );
xor U84581 ( n51211, n50978, n50979 );
xor U84582 ( n51190, n50966, n51198 );
xnor U84583 ( n51198, n50965, n50967 );
nand U84584 ( n50978, n51321, n51322 );
nand U84585 ( n51322, n51323, n51324 );
nand U84586 ( n50965, n51199, n51200 );
nand U84587 ( n51200, n1533, n51201 );
nand U84588 ( n51199, n51204, n50972 );
not U84589 ( n1533, n50972 );
nand U84590 ( n51191, n51093, n51095 );
nand U84591 ( n51204, n50969, n50971 );
xnor U84592 ( n17970, n17723, n17984 );
xor U84593 ( n17984, n17721, n17722 );
nand U84594 ( n17994, n18373, n18374 );
nand U84595 ( n18374, n18375, n18376 );
nor U84596 ( n18227, n17993, n2579 );
not U84597 ( n2579, n17996 );
nand U84598 ( n17721, n18140, n18141 );
nand U84599 ( n18140, n18145, n18144 );
nand U84600 ( n18141, n18142, n18143 );
or U84601 ( n18142, n18144, n18145 );
nor U84602 ( n48733, n48465, n48719 );
xor U84603 ( n50747, n51015, n50820 );
xor U84604 ( n51015, n50822, n50823 );
nand U84605 ( n51096, n51192, n51193 );
nand U84606 ( n51192, n51196, n51197 );
nand U84607 ( n51193, n51194, n51195 );
or U84608 ( n51195, n51196, n51197 );
nor U84609 ( n49388, n48465, n49358 );
nor U84610 ( n49295, n48465, n49280 );
nor U84611 ( n49104, n48465, n7834 );
nor U84612 ( n49010, n48465, n48995 );
nor U84613 ( n48927, n48465, n48896 );
nor U84614 ( n48644, n48465, n48629 );
nor U84615 ( n48550, n48465, n48535 );
nor U84616 ( n49199, n48465, n49184 );
nor U84617 ( n48830, n48465, n48815 );
nor U84618 ( n49523, n48465, n49462 );
nand U84619 ( n14866, n49503, n49504 );
nor U84620 ( n49504, n49505, n49506 );
nor U84621 ( n49503, n49523, n49524 );
nand U84622 ( n49506, n49507, n49508 );
nand U84623 ( n49790, n49978, n49979 );
nand U84624 ( n49979, n49980, n49981 );
not U84625 ( n1608, n49782 );
xor U84626 ( n51410, n51418, n51233 );
xnor U84627 ( n51418, n51231, n51232 );
xnor U84628 ( n51216, n51313, n51405 );
xnor U84629 ( n51405, n51312, n51314 );
xor U84630 ( n51434, n51245, n51435 );
xnor U84631 ( n51435, n51246, n51243 );
xor U84632 ( n51425, n51426, n1680 );
nand U84633 ( n51312, n51406, n51407 );
nand U84634 ( n51407, n1624, n51408 );
nand U84635 ( n51406, n51411, n51308 );
not U84636 ( n1624, n51308 );
nand U84637 ( n51411, n51305, n51307 );
xor U84638 ( n51438, n51439, n51440 );
or U84639 ( n18345, n18483, n18484 );
nand U84640 ( n18312, n18499, n18500 );
nand U84641 ( n18499, n18504, n18503 );
nand U84642 ( n18500, n18501, n18502 );
or U84643 ( n18501, n18503, n18504 );
not U84644 ( n2500, n19497 );
xnor U84645 ( n51769, n52127, n52128 );
xnor U84646 ( n52127, n52129, n52130 );
xor U84647 ( n50458, n50459, n1673 );
nand U84648 ( n49813, n50172, n50173 );
nand U84649 ( n50172, n50177, n50176 );
nand U84650 ( n50173, n50174, n50175 );
or U84651 ( n50174, n50176, n50177 );
nand U84652 ( n51076, n51241, n51242 );
nand U84653 ( n51241, n51245, n51246 );
nand U84654 ( n51242, n51243, n51244 );
or U84655 ( n51244, n51245, n51246 );
not U84656 ( n70, n15317 );
nand U84657 ( n50388, n50667, n50668 );
nand U84658 ( n50667, n50672, n50394 );
nand U84659 ( n50668, n1430, n50669 );
nand U84660 ( n50672, n50391, n50393 );
nand U84661 ( n50394, n50673, n50674 );
nand U84662 ( n50673, n50678, n50677 );
nand U84663 ( n50674, n50675, n50676 );
or U84664 ( n50675, n50677, n50678 );
and U84665 ( n17363, n17365, n17367 );
nand U84666 ( n51301, n51426, n1680 );
xnor U84667 ( n17784, n17524, n17792 );
xor U84668 ( n17792, n17522, n17523 );
nand U84669 ( n17253, n17514, n17515 );
nand U84670 ( n17515, n17516, n17517 );
xnor U84671 ( n50671, n50679, n50406 );
xor U84672 ( n50679, n50407, n50404 );
nand U84673 ( n50407, n50844, n50845 );
nand U84674 ( n50845, n50846, n50847 );
xnor U84675 ( n52298, n53959, n52599 );
xnor U84676 ( n53959, n52596, n52598 );
nand U84677 ( n18113, n18302, n18303 );
nand U84678 ( n18302, n18307, n18306 );
nand U84679 ( n18303, n18304, n18305 );
or U84680 ( n18304, n18306, n18307 );
nand U84681 ( n50966, n51325, n51326 );
nand U84682 ( n51326, n51327, n51328 );
xor U84683 ( n18640, n18648, n18504 );
xnor U84684 ( n18648, n18502, n18503 );
nand U84685 ( n18306, n18523, n18524 );
nand U84686 ( n18524, n18525, n18526 );
xnor U84687 ( n18541, n18606, n18535 );
xor U84688 ( n18606, n18536, n18533 );
nand U84689 ( n19157, n19488, n19489 );
nand U84690 ( n19488, n19174, n19172 );
nand U84691 ( n19489, n19173, n19490 );
or U84692 ( n19490, n19172, n19174 );
nand U84693 ( n18536, n18673, n18674 );
nand U84694 ( n18673, n18677, n18678 );
nand U84695 ( n18674, n18675, n18676 );
nor U84696 ( n19495, n19496, n19497 );
nor U84697 ( n19496, n19498, n19499 );
nor U84698 ( n19498, n19500, n19501 );
and U84699 ( n19153, n2418, n19157 );
xor U84700 ( n51568, n51574, n51433 );
xnor U84701 ( n51574, n51432, n51431 );
xnor U84702 ( n51583, n51447, n51591 );
xor U84703 ( n51591, n51445, n51446 );
nand U84704 ( n51421, n51568, n51567 );
or U84705 ( n51483, n51582, n51583 );
not U84706 ( n327, n48440 );
xor U84707 ( n49500, n49501, n49502 );
xor U84708 ( n51581, n51582, n51583 );
nand U84709 ( n51485, n51583, n51582 );
xnor U84710 ( n51006, n51014, n50747 );
xor U84711 ( n51014, n50749, n50750 );
nand U84712 ( n50464, n50824, n50825 );
nand U84713 ( n50825, n50826, n50827 );
nand U84714 ( n17234, n17240, n17241 );
nand U84715 ( n17241, n17242, n17243 );
xor U84716 ( n50382, n50329, n50390 );
xnor U84717 ( n50390, n50327, n50330 );
nand U84718 ( n50330, n50391, n50392 );
nand U84719 ( n50392, n50393, n50394 );
nand U84720 ( n50076, n50378, n50379 );
nand U84721 ( n50379, n1395, n50380 );
nand U84722 ( n50378, n50383, n50335 );
not U84723 ( n1395, n50335 );
nand U84724 ( n50383, n50332, n50334 );
nand U84725 ( n50972, n51205, n51206 );
nand U84726 ( n51205, n51210, n51209 );
nand U84727 ( n51206, n51207, n51208 );
or U84728 ( n51207, n51209, n51210 );
nand U84729 ( n18641, n18523, n18525 );
nand U84730 ( n18348, n18486, n18487 );
nand U84731 ( n18486, n18491, n18490 );
nand U84732 ( n18487, n18488, n18489 );
or U84733 ( n18488, n18490, n18491 );
nand U84734 ( n18490, n18636, n18637 );
nand U84735 ( n18637, n2817, n18638 );
nand U84736 ( n18636, n18641, n18526 );
not U84737 ( n2817, n18526 );
nand U84738 ( n51303, n51434, n1668 );
not U84739 ( n1668, n51426 );
nand U84740 ( n17083, n17117, n17118 );
nand U84741 ( n17117, n17122, n17121 );
nand U84742 ( n17118, n17119, n17120 );
or U84743 ( n17119, n17121, n17122 );
nand U84744 ( n51313, n51487, n51488 );
nand U84745 ( n51487, n51491, n51492 );
nand U84746 ( n51488, n51489, n51490 );
or U84747 ( n51490, n51491, n51492 );
nand U84748 ( n50024, n50332, n50333 );
nand U84749 ( n50333, n50334, n50335 );
nand U84750 ( n18860, n2383, n18859 );
nand U84751 ( n50335, n50384, n50385 );
nand U84752 ( n50384, n50389, n50388 );
nand U84753 ( n50385, n50386, n50387 );
or U84754 ( n50386, n50388, n50389 );
or U84755 ( n51419, n51567, n51568 );
nand U84756 ( n18793, n19148, n19149 );
or U84757 ( n19148, n18819, n18818 );
nand U84758 ( n19149, n18820, n19150 );
nand U84759 ( n19150, n18818, n18819 );
nor U84760 ( n19155, n19156, n19157 );
nor U84761 ( n19156, n19158, n19159 );
nor U84762 ( n19158, n2418, n19160 );
and U84763 ( n18820, n19151, n19152 );
nand U84764 ( n19152, n19153, n2463 );
nor U84765 ( n19151, n19154, n19155 );
nor U84766 ( n19154, n2463, n19161 );
xnor U84767 ( n50447, n50177, n50455 );
xor U84768 ( n50455, n50175, n50176 );
nand U84769 ( n50156, n50162, n50163 );
nand U84770 ( n50163, n50164, n50165 );
xnor U84771 ( n50947, n50690, n50955 );
xor U84772 ( n50955, n50688, n50689 );
xor U84773 ( n50945, n50946, n50947 );
nand U84774 ( n50688, n51093, n51094 );
nand U84775 ( n51094, n51095, n51096 );
nand U84776 ( n19172, n19503, n19504 );
nand U84777 ( n19504, n19505, n19506 );
nor U84778 ( n19503, n19507, n19508 );
not U84779 ( n2465, n21063 );
not U84780 ( n2420, n19506 );
nand U84781 ( n21023, n21052, n21053 );
nand U84782 ( n21053, n21054, n2465 );
nor U84783 ( n21052, n21055, n21056 );
nor U84784 ( n21055, n2503, n21062 );
nand U84785 ( n17511, n17780, n17781 );
nand U84786 ( n17780, n17785, n17517 );
nand U84787 ( n17781, n2799, n17782 );
nand U84788 ( n17785, n17514, n17516 );
nand U84789 ( n17243, n17507, n17508 );
nand U84790 ( n17507, n17512, n17511 );
nand U84791 ( n17508, n17509, n17510 );
or U84792 ( n17509, n17511, n17512 );
nand U84793 ( n50827, n51008, n51009 );
nand U84794 ( n51008, n51013, n51012 );
nand U84795 ( n51009, n51010, n51011 );
or U84796 ( n51010, n51012, n51013 );
or U84797 ( n50844, n50946, n50947 );
xnor U84798 ( n50730, n50466, n50738 );
xor U84799 ( n50738, n50464, n50465 );
nand U84800 ( n50552, n50730, n50729 );
and U84801 ( n19642, n21087, n21088 );
nand U84802 ( n21088, n21058, n21063 );
nor U84803 ( n21087, n21054, n21060 );
xor U84804 ( n51237, n51238, n51239 );
xnor U84805 ( n17976, n18145, n18222 );
xnor U84806 ( n18222, n18143, n18144 );
or U84807 ( n50550, n50729, n50730 );
xor U84808 ( n51491, n51563, n51416 );
xor U84809 ( n51563, n51415, n51417 );
xor U84810 ( n51566, n51567, n51568 );
nand U84811 ( n50846, n50947, n50946 );
nand U84812 ( n51766, n52121, n52122 );
nand U84813 ( n52121, n52126, n52125 );
nand U84814 ( n52122, n52123, n52124 );
or U84815 ( n52124, n52125, n52126 );
and U84816 ( n52126, n53945, n53946 );
nand U84817 ( n53946, n52300, n1305 );
nor U84818 ( n53945, n53948, n53949 );
nor U84819 ( n53948, n1345, n53952 );
nand U84820 ( n51308, n51412, n51413 );
nand U84821 ( n51412, n51417, n51416 );
nand U84822 ( n51413, n51414, n51415 );
or U84823 ( n51414, n51416, n51417 );
nand U84824 ( n16537, n18735, n18736 );
or U84825 ( n18735, n16498, n16502 );
nand U84826 ( n18736, n16500, n18737 );
nand U84827 ( n18737, n16502, n16498 );
xnor U84828 ( n50960, n50842, n50968 );
xor U84829 ( n50968, n50841, n50843 );
nand U84830 ( n50689, n50956, n50957 );
nand U84831 ( n50956, n50961, n50696 );
nand U84832 ( n50957, n1508, n50958 );
nand U84833 ( n50961, n50693, n50695 );
nand U84834 ( n50841, n50969, n50970 );
nand U84835 ( n50970, n50971, n50972 );
nand U84836 ( n50696, n50962, n50963 );
nand U84837 ( n50962, n50967, n50966 );
nand U84838 ( n50963, n50964, n50965 );
or U84839 ( n50964, n50966, n50967 );
nand U84840 ( n51304, n51428, n51429 );
nand U84841 ( n51428, n51433, n51432 );
nand U84842 ( n51429, n51430, n51431 );
or U84843 ( n51430, n51432, n51433 );
nor U84844 ( n15633, n15317, n5179 );
nand U84845 ( n51708, n1268, n51707 );
xor U84846 ( n18454, n18462, n18281 );
xnor U84847 ( n18462, n18279, n18280 );
xnor U84848 ( n18264, n18361, n18449 );
xnor U84849 ( n18449, n18360, n18362 );
xor U84850 ( n18478, n18292, n18479 );
xnor U84851 ( n18479, n18293, n18290 );
xor U84852 ( n18482, n18483, n18484 );
xor U84853 ( n18469, n18470, n2797 );
nand U84854 ( n18360, n18450, n18451 );
nand U84855 ( n18451, n2747, n18452 );
nand U84856 ( n18450, n18455, n18356 );
not U84857 ( n2747, n18356 );
nand U84858 ( n18455, n18353, n18355 );
not U84859 ( n1307, n54004 );
and U84860 ( n53957, n54022, n54023 );
nand U84861 ( n54023, n53999, n54004 );
nor U84862 ( n54022, n53995, n54001 );
nor U84863 ( n16539, n15317, n5168 );
nor U84864 ( n16365, n15317, n16347 );
nor U84865 ( n16260, n15317, n16242 );
nor U84866 ( n16160, n15317, n16135 );
nor U84867 ( n16058, n15317, n16039 );
nor U84868 ( n15950, n15317, n15932 );
nor U84869 ( n15845, n15317, n15827 );
nor U84870 ( n15735, n15317, n15717 );
nor U84871 ( n15537, n15317, n15518 );
nor U84872 ( n15430, n15317, n15412 );
nand U84873 ( n8131, n16514, n16515 );
nor U84874 ( n16515, n16517, n16518 );
nor U84875 ( n16514, n16539, n16540 );
nand U84876 ( n16518, n16519, n16520 );
xnor U84877 ( n18294, n18119, n18295 );
xor U84878 ( n18295, n18117, n18118 );
nand U84879 ( n17517, n17786, n17787 );
nand U84880 ( n17786, n17791, n17790 );
nand U84881 ( n17787, n17788, n17789 );
or U84882 ( n17789, n17790, n17791 );
nand U84883 ( n18057, n18286, n2807 );
xor U84884 ( n16545, n16548, n16549 );
nand U84885 ( n17722, n17985, n17986 );
nand U84886 ( n17985, n17990, n17892 );
nand U84887 ( n17986, n2577, n17987 );
nand U84888 ( n17990, n17889, n17891 );
not U84889 ( n2577, n17892 );
nand U84890 ( n18059, n18294, n2803 );
not U84891 ( n2803, n18286 );
nand U84892 ( n51091, n51315, n51316 );
or U84893 ( n51315, n51319, n51320 );
nand U84894 ( n51316, n51317, n51318 );
nand U84895 ( n51317, n51319, n51320 );
nand U84896 ( n18349, n18470, n2797 );
nand U84897 ( n50019, n50325, n50326 );
nand U84898 ( n50325, n50329, n50330 );
nand U84899 ( n50326, n50327, n50328 );
or U84900 ( n50328, n50329, n50330 );
not U84901 ( n2503, n21058 );
not U84902 ( n1349, n53999 );
nor U84903 ( n48725, n48440, n48719 );
xor U84904 ( n50728, n50729, n50730 );
nand U84905 ( n50165, n50449, n50450 );
nand U84906 ( n50449, n50454, n50453 );
nand U84907 ( n50450, n50451, n50452 );
or U84908 ( n50451, n50453, n50454 );
xnor U84909 ( n18234, n18242, n18008 );
xor U84910 ( n18242, n18007, n18009 );
xnor U84911 ( n18251, n18259, n18132 );
xor U84912 ( n18259, n18134, n18135 );
nand U84913 ( n17993, n18230, n18231 );
nand U84914 ( n18231, n2609, n18232 );
nand U84915 ( n18230, n18235, n18139 );
not U84916 ( n2609, n18139 );
nand U84917 ( n18134, n18369, n18370 );
nand U84918 ( n18370, n18371, n18372 );
nand U84919 ( n18007, n18247, n18248 );
nand U84920 ( n18248, n2654, n18249 );
nand U84921 ( n18247, n18252, n18014 );
not U84922 ( n2654, n18014 );
nand U84923 ( n18235, n18136, n18138 );
nand U84924 ( n18252, n18011, n18013 );
nor U84925 ( n49287, n48440, n49280 );
nor U84926 ( n49191, n48440, n49184 );
nor U84927 ( n49096, n48440, n7834 );
nor U84928 ( n49002, n48440, n48995 );
nor U84929 ( n48903, n48440, n48896 );
nor U84930 ( n48822, n48440, n48815 );
nor U84931 ( n48636, n48440, n48629 );
nor U84932 ( n48542, n48440, n48535 );
nor U84933 ( n49365, n48440, n49358 );
nor U84934 ( n49494, n48440, n49462 );
nand U84935 ( n14871, n49470, n49471 );
nor U84936 ( n49471, n49472, n49473 );
nor U84937 ( n49470, n49494, n49495 );
nand U84938 ( n49473, n49474, n49475 );
nand U84939 ( n16819, n16820, n16821 );
nand U84940 ( n16821, n2729, n16822 );
nand U84941 ( n16820, n16827, n16828 );
nand U84942 ( n16822, n16823, n16824 );
nand U84943 ( n16828, n16829, n16830 );
nand U84944 ( n16829, n16832, n16825 );
or U84945 ( n16830, n16831, n2712 );
xnor U84946 ( n51226, n51013, n51234 );
xor U84947 ( n51234, n51011, n51012 );
nand U84948 ( n50736, n51077, n51078 );
nand U84949 ( n51078, n51079, n51080 );
nand U84950 ( n50553, n50732, n50733 );
nand U84951 ( n50732, n50737, n50736 );
nand U84952 ( n50733, n50734, n50735 );
or U84953 ( n50734, n50736, n50737 );
nand U84954 ( n17230, n17501, n17502 );
nand U84955 ( n17502, n2780, n17503 );
nand U84956 ( n17501, n17506, n17243 );
not U84957 ( n2780, n17243 );
nand U84958 ( n16858, n17226, n17227 );
nand U84959 ( n17226, n17231, n17230 );
nand U84960 ( n17227, n17228, n17229 );
or U84961 ( n17228, n17230, n17231 );
nand U84962 ( n17506, n17240, n17242 );
nand U84963 ( n17128, n17429, n17430 );
nand U84964 ( n17429, n17434, n17433 );
nand U84965 ( n17430, n17431, n17432 );
or U84966 ( n17431, n17433, n17434 );
and U84967 ( n17070, n17125, n17126 );
nand U84968 ( n17126, n17127, n17128 );
xor U84969 ( n17788, n18061, n17861 );
xor U84970 ( n18061, n17863, n17864 );
xnor U84971 ( n18616, n18477, n18622 );
xor U84972 ( n18622, n18475, n18476 );
xnor U84973 ( n18627, n18491, n18635 );
xor U84974 ( n18635, n18489, n18490 );
nand U84975 ( n18465, n18616, n18615 );
or U84976 ( n18527, n18626, n18627 );
nand U84977 ( n18143, n18377, n18378 );
nand U84978 ( n18377, n18382, n18381 );
nand U84979 ( n18378, n18379, n18380 );
or U84980 ( n18379, n18381, n18382 );
nand U84981 ( n18060, n18288, n18289 );
nand U84982 ( n18288, n18292, n18293 );
nand U84983 ( n18289, n18290, n18291 );
or U84984 ( n18291, n18292, n18293 );
xor U84985 ( n18625, n18626, n18627 );
not U84986 ( n2460, n19505 );
nand U84987 ( n18351, n18478, n2789 );
not U84988 ( n2789, n18470 );
nand U84989 ( n50703, n50974, n50975 );
nand U84990 ( n50974, n50979, n50978 );
nand U84991 ( n50975, n50976, n50977 );
or U84992 ( n50977, n50978, n50979 );
nand U84993 ( n18529, n18627, n18626 );
nand U84994 ( n18139, n18236, n18237 );
nand U84995 ( n18236, n18240, n18241 );
nand U84996 ( n18237, n18238, n18239 );
or U84997 ( n18239, n18240, n18241 );
xnor U84998 ( n18813, n19171, n19172 );
xnor U84999 ( n19171, n19173, n19174 );
nand U85000 ( n16296, n43976, n43977 );
nor U85001 ( n43977, n43978, n43979 );
nor U85002 ( n43976, n44017, n44018 );
nor U85003 ( n43978, n43457, n76362 );
or U85004 ( n18463, n18615, n18616 );
nand U85005 ( n17433, n17712, n17713 );
nand U85006 ( n17712, n17717, n17439 );
nand U85007 ( n17713, n2552, n17714 );
nand U85008 ( n17717, n17436, n17438 );
nand U85009 ( n17439, n17718, n17719 );
nand U85010 ( n17718, n17723, n17722 );
nand U85011 ( n17719, n17720, n17721 );
or U85012 ( n17720, n17722, n17723 );
nor U85013 ( n18745, n18746, n18747 );
nor U85014 ( n18746, n18748, n18749 );
nor U85015 ( n18748, n18750, n18751 );
nand U85016 ( n18361, n18531, n18532 );
nand U85017 ( n18531, n18535, n18536 );
nand U85018 ( n18532, n18533, n18534 );
or U85019 ( n18534, n18535, n18536 );
nand U85020 ( n50152, n50443, n50444 );
nand U85021 ( n50444, n1622, n50445 );
nand U85022 ( n50443, n50448, n50165 );
not U85023 ( n1622, n50165 );
nand U85024 ( n49981, n50148, n50149 );
nand U85025 ( n50148, n50153, n50152 );
nand U85026 ( n50149, n50150, n50151 );
or U85027 ( n50150, n50152, n50153 );
nand U85028 ( n50448, n50162, n50164 );
xnor U85029 ( n17716, n17724, n17451 );
xor U85030 ( n17724, n17452, n17449 );
nand U85031 ( n17452, n17889, n17890 );
nand U85032 ( n17890, n17891, n17892 );
nand U85033 ( n19502, n2472, n19501 );
and U85034 ( n49456, n51709, n51710 );
nand U85035 ( n51709, n45513, n45515 );
nand U85036 ( n51710, n45516, n51711 );
or U85037 ( n51711, n45515, n45513 );
nand U85038 ( n50735, n51002, n51003 );
nand U85039 ( n51003, n1664, n51004 );
nand U85040 ( n51002, n51007, n50827 );
not U85041 ( n1664, n50827 );
nand U85042 ( n51007, n50824, n50826 );
nand U85043 ( n16835, n17024, n17025 );
nand U85044 ( n17025, n17026, n17027 );
not U85045 ( n2729, n16827 );
nand U85046 ( n18014, n18253, n18254 );
nand U85047 ( n18253, n18258, n18257 );
nand U85048 ( n18254, n18255, n18256 );
or U85049 ( n18255, n18257, n18258 );
xor U85050 ( n18285, n18286, n2807 );
nand U85051 ( n17868, n18050, n18051 );
nand U85052 ( n18050, n18055, n18054 );
nand U85053 ( n18051, n18052, n18053 );
or U85054 ( n18052, n18054, n18055 );
nand U85055 ( n17510, n17865, n17866 );
nand U85056 ( n17866, n17867, n17868 );
xnor U85057 ( n17771, n17512, n17779 );
xor U85058 ( n17779, n17510, n17511 );
nand U85059 ( n17229, n17593, n17594 );
nand U85060 ( n17594, n17595, n17596 );
and U85061 ( n45474, n51781, n51782 );
nand U85062 ( n51782, n51783, n1259 );
nor U85063 ( n51781, n51784, n51785 );
nor U85064 ( n51784, n1298, n51791 );
xor U85065 ( n18048, n17788, n18056 );
xnor U85066 ( n18056, n17790, n17791 );
nor U85067 ( n19369, n19057, n19362 );
nand U85068 ( n19035, n19360, n19361 );
nand U85069 ( n19361, n19362, n19363 );
nand U85070 ( n19360, n19369, n19054 );
nor U85071 ( n19363, n19364, n19365 );
nand U85072 ( n18008, n18243, n18244 );
nand U85073 ( n18244, n18245, n18246 );
nand U85074 ( n17121, n17423, n17424 );
nand U85075 ( n17423, n17428, n17128 );
nand U85076 ( n17424, n2515, n17425 );
nand U85077 ( n17428, n17125, n17127 );
nand U85078 ( n50329, n50396, n50397 );
nand U85079 ( n50396, n50401, n50324 );
nand U85080 ( n50397, n1455, n50398 );
nand U85081 ( n50401, n50321, n50323 );
nand U85082 ( n50324, n50402, n50403 );
nand U85083 ( n50402, n50406, n50407 );
nand U85084 ( n50403, n50404, n50405 );
or U85085 ( n50405, n50406, n50407 );
xor U85086 ( n18614, n18615, n18616 );
nand U85087 ( n18356, n18456, n18457 );
nand U85088 ( n18456, n18461, n18460 );
nand U85089 ( n18457, n18458, n18459 );
or U85090 ( n18458, n18460, n18461 );
nand U85091 ( n49792, n49799, n49800 );
nand U85092 ( n49800, n49801, n49802 );
nand U85093 ( n49801, n49804, n49797 );
or U85094 ( n49802, n49803, n1619 );
nor U85095 ( n51719, n51720, n51721 );
nor U85096 ( n51720, n51722, n51723 );
nor U85097 ( n51722, n51724, n51725 );
nand U85098 ( n18352, n18472, n18473 );
nand U85099 ( n18472, n18477, n18476 );
nand U85100 ( n18473, n18474, n18475 );
or U85101 ( n18474, n18476, n18477 );
xnor U85102 ( n17492, n17231, n17500 );
xor U85103 ( n17500, n17229, n17230 );
nand U85104 ( n17210, n17216, n17217 );
nand U85105 ( n17217, n17218, n17219 );
nand U85106 ( n51080, n51228, n51229 );
nand U85107 ( n51228, n51233, n51232 );
nand U85108 ( n51229, n51230, n51231 );
or U85109 ( n51230, n51232, n51233 );
not U85110 ( n324, n48428 );
xnor U85111 ( n18535, n18460, n18607 );
xnor U85112 ( n18607, n18461, n18459 );
xor U85113 ( n51000, n50736, n51001 );
xnor U85114 ( n51001, n50737, n50735 );
nand U85115 ( n50828, n50992, n1640 );
xnor U85116 ( n51089, n51085, n51213 );
xnor U85117 ( n51213, n51084, n51086 );
nand U85118 ( n51084, n51214, n51215 );
nand U85119 ( n51214, n51219, n51218 );
nand U85120 ( n51215, n51216, n51217 );
or U85121 ( n51217, n51218, n51219 );
not U85122 ( n2424, n21005 );
and U85123 ( n21025, n21037, n21038 );
nand U85124 ( n21038, n21000, n21005 );
nor U85125 ( n21037, n20996, n21002 );
xor U85126 ( n17427, n17379, n17435 );
xnor U85127 ( n17435, n17377, n17380 );
nand U85128 ( n17380, n17436, n17437 );
nand U85129 ( n17437, n17438, n17439 );
nand U85130 ( n50830, n51000, n1635 );
not U85131 ( n1635, n50992 );
xnor U85132 ( n19029, n18647, n19037 );
xor U85133 ( n19037, n18645, n18646 );
nand U85134 ( n18646, n19038, n19039 );
nand U85135 ( n19039, n19040, n19041 );
nand U85136 ( n19038, n19047, n18661 );
nor U85137 ( n19041, n19042, n19043 );
nor U85138 ( n19047, n18664, n19040 );
xnor U85139 ( n17989, n17736, n17997 );
xor U85140 ( n17997, n17734, n17735 );
xnor U85141 ( n18002, n17883, n18010 );
xor U85142 ( n18010, n17882, n17884 );
xor U85143 ( n17987, n17988, n17989 );
nand U85144 ( n17735, n17998, n17999 );
nand U85145 ( n17998, n18003, n17888 );
nand U85146 ( n17999, n2630, n18000 );
nand U85147 ( n18003, n17885, n17887 );
nand U85148 ( n17882, n18011, n18012 );
nand U85149 ( n18012, n18013, n18014 );
or U85150 ( n17889, n17988, n17989 );
or U85151 ( n51726, n51724, n1258 );
nand U85152 ( n17734, n18136, n18137 );
nand U85153 ( n18137, n18138, n18139 );
nand U85154 ( n49807, n49810, n49811 );
nand U85155 ( n49811, n49812, n49813 );
nand U85156 ( n49793, n1618, n49794 );
nand U85157 ( n49794, n49795, n49796 );
not U85158 ( n1618, n49799 );
nand U85159 ( n49795, n1619, n1637 );
nand U85160 ( n50010, n50321, n50322 );
nand U85161 ( n50322, n50323, n50324 );
nand U85162 ( n17891, n17989, n17988 );
nand U85163 ( n52125, n53988, n53989 );
nand U85164 ( n53989, n53938, n53943 );
nor U85165 ( n53988, n53934, n53940 );
nand U85166 ( n53943, n53990, n53991 );
nand U85167 ( n53990, n53930, n53929 );
nand U85168 ( n53991, n53931, n53992 );
or U85169 ( n53992, n53929, n53930 );
and U85170 ( n53931, n53993, n53994 );
nand U85171 ( n53994, n53995, n1307 );
nor U85172 ( n53993, n53996, n53997 );
nor U85173 ( n53996, n1349, n54003 );
xnor U85174 ( n50420, n50105, n50421 );
xor U85175 ( n50421, n50102, n50104 );
xnor U85176 ( n50400, n50087, n50408 );
xor U85177 ( n50408, n50085, n50086 );
xor U85178 ( n50411, n50412, n1530 );
nand U85179 ( n50426, n50838, n50839 );
or U85180 ( n50838, n50842, n50843 );
nand U85181 ( n50839, n50840, n50841 );
nand U85182 ( n50840, n50842, n50843 );
nand U85183 ( n50999, n51305, n51306 );
nand U85184 ( n51306, n51307, n51308 );
nand U85185 ( n50831, n50994, n50995 );
nand U85186 ( n50994, n50998, n50999 );
nand U85187 ( n50995, n50996, n50997 );
or U85188 ( n50997, n50998, n50999 );
nand U85189 ( n50998, n51222, n51223 );
nand U85190 ( n51222, n51227, n51080 );
nand U85191 ( n51223, n1652, n51224 );
nand U85192 ( n51227, n51077, n51079 );
xnor U85193 ( n50434, n50153, n50442 );
xor U85194 ( n50442, n50151, n50152 );
nand U85195 ( n50132, n50138, n50139 );
nand U85196 ( n50139, n50140, n50141 );
nand U85197 ( n17498, n17767, n17768 );
nand U85198 ( n17767, n17772, n17596 );
nand U85199 ( n17768, n2765, n17769 );
nand U85200 ( n17772, n17593, n17595 );
nand U85201 ( n17219, n17494, n17495 );
nand U85202 ( n17494, n17499, n17498 );
nand U85203 ( n17495, n17496, n17497 );
or U85204 ( n17496, n17498, n17499 );
xnor U85205 ( n50691, n50418, n50692 );
xor U85206 ( n50692, n50417, n50419 );
xor U85207 ( n50682, n50683, n1504 );
nand U85208 ( n50417, n50693, n50694 );
nand U85209 ( n50694, n50695, n50696 );
xnor U85210 ( n50717, n50454, n50725 );
xor U85211 ( n50725, n50452, n50453 );
nand U85212 ( n50151, n50554, n50555 );
nand U85213 ( n50555, n50556, n50557 );
xnor U85214 ( n18274, n18055, n18282 );
xor U85215 ( n18282, n18053, n18054 );
nand U85216 ( n17777, n18120, n18121 );
nand U85217 ( n18121, n18122, n18123 );
nand U85218 ( n17596, n17773, n17774 );
nand U85219 ( n17773, n17778, n17777 );
nand U85220 ( n17774, n17775, n17776 );
or U85221 ( n17775, n17777, n17778 );
nand U85222 ( n18810, n19165, n19166 );
or U85223 ( n19165, n19170, n19169 );
nand U85224 ( n19166, n19167, n19168 );
nand U85225 ( n19168, n19169, n19170 );
nor U85226 ( n21029, n21030, n19505 );
nor U85227 ( n21030, n21031, n19508 );
nor U85228 ( n21031, n21032, n19506 );
not U85229 ( n67, n15305 );
xor U85230 ( n16510, n16512, n16513 );
xor U85231 ( n53938, n53958, n54021 );
xor U85232 ( n54021, n53955, n53957 );
nand U85233 ( n50090, n50412, n1530 );
nand U85234 ( n51486, n51585, n51586 );
nand U85235 ( n51585, n51590, n51589 );
nand U85236 ( n51586, n51587, n51588 );
or U85237 ( n51587, n51589, n51590 );
nand U85238 ( n17888, n18004, n18005 );
nand U85239 ( n18004, n18009, n18008 );
nand U85240 ( n18005, n18006, n18007 );
or U85241 ( n18006, n18008, n18009 );
nand U85242 ( n18128, n18363, n18364 );
or U85243 ( n18363, n18367, n18368 );
nand U85244 ( n18364, n18365, n18366 );
nand U85245 ( n18365, n18367, n18368 );
xnor U85246 ( n45481, n51793, n51794 );
xnor U85247 ( n51793, n51795, n51796 );
nand U85248 ( n50570, n50683, n1504 );
xnor U85249 ( n51085, n51220, n50987 );
xnor U85250 ( n51220, n50988, n50985 );
and U85251 ( n50988, n51309, n51310 );
nand U85252 ( n51309, n51314, n51313 );
nand U85253 ( n51310, n51311, n51312 );
or U85254 ( n51311, n51313, n51314 );
not U85255 ( n2467, n21000 );
nand U85256 ( n9561, n10060, n10062 );
nor U85257 ( n10062, n10063, n10064 );
nor U85258 ( n10060, n10112, n10113 );
nor U85259 ( n10063, n9497, n76632 );
xor U85260 ( n50701, n50980, n50708 );
xor U85261 ( n50980, n50710, n50711 );
nand U85262 ( n50723, n50983, n50984 );
or U85263 ( n50983, n50987, n50988 );
nand U85264 ( n50984, n50985, n50986 );
nand U85265 ( n50986, n50987, n50988 );
nand U85266 ( n50557, n50719, n50720 );
nand U85267 ( n50719, n50724, n50723 );
nand U85268 ( n50720, n50721, n50722 );
or U85269 ( n50721, n50723, n50724 );
nand U85270 ( n53929, n54005, n54006 );
nand U85271 ( n54006, n1308, n53927 );
nor U85272 ( n54005, n53918, n53923 );
nand U85273 ( n18752, n2384, n18751 );
nand U85274 ( n17744, n18130, n18131 );
nand U85275 ( n18130, n18135, n18134 );
nand U85276 ( n18131, n18132, n18133 );
or U85277 ( n18133, n18134, n18135 );
nand U85278 ( n50572, n50691, n1502 );
not U85279 ( n1502, n50683 );
nand U85280 ( n50440, n50713, n50714 );
nand U85281 ( n50713, n50718, n50557 );
nand U85282 ( n50714, n1613, n50715 );
nand U85283 ( n50718, n50554, n50556 );
nand U85284 ( n50141, n50436, n50437 );
nand U85285 ( n50436, n50441, n50440 );
nand U85286 ( n50437, n50438, n50439 );
or U85287 ( n50438, n50440, n50441 );
nand U85288 ( n50092, n50420, n1528 );
not U85289 ( n1528, n50412 );
nand U85290 ( n17206, n17488, n17489 );
nand U85291 ( n17489, n2743, n17490 );
nand U85292 ( n17488, n17493, n17219 );
not U85293 ( n2743, n17219 );
nand U85294 ( n17027, n17202, n17203 );
nand U85295 ( n17202, n17207, n17206 );
nand U85296 ( n17203, n17204, n17205 );
or U85297 ( n17204, n17206, n17207 );
nand U85298 ( n17493, n17216, n17218 );
nand U85299 ( n51452, n51598, n51599 );
nand U85300 ( n51598, n51603, n51602 );
nand U85301 ( n51599, n51600, n51601 );
or U85302 ( n51600, n51602, n51603 );
nor U85303 ( n48714, n48428, n48719 );
xnor U85304 ( n50424, n50568, n50698 );
xnor U85305 ( n50698, n50567, n50569 );
nor U85306 ( n49355, n48428, n49358 );
nor U85307 ( n49277, n48428, n49280 );
nor U85308 ( n49181, n48428, n49184 );
nor U85309 ( n49087, n48428, n7834 );
nor U85310 ( n48992, n48428, n48995 );
nor U85311 ( n48893, n48428, n48896 );
nor U85312 ( n48812, n48428, n48815 );
nor U85313 ( n48626, n48428, n48629 );
nor U85314 ( n48532, n48428, n48535 );
nor U85315 ( n49459, n48428, n49462 );
nand U85316 ( n14876, n49439, n49440 );
nor U85317 ( n49440, n49441, n49442 );
nor U85318 ( n49439, n49459, n49460 );
nand U85319 ( n49442, n49443, n49444 );
nand U85320 ( n11724, n18771, n18772 );
nand U85321 ( n18771, n11710, n11713 );
nand U85322 ( n18772, n11714, n18773 );
or U85323 ( n18773, n11713, n11710 );
and U85324 ( n11702, n18825, n18826 );
nand U85325 ( n18826, n18827, n2374 );
nor U85326 ( n18825, n18828, n18829 );
nor U85327 ( n18828, n2414, n18835 );
and U85328 ( n16457, n18753, n18754 );
or U85329 ( n18753, n11738, n11742 );
nand U85330 ( n18754, n11740, n18755 );
nand U85331 ( n18755, n11742, n11738 );
nand U85332 ( n17065, n17375, n17376 );
nand U85333 ( n17375, n17379, n17380 );
nand U85334 ( n17376, n17377, n17378 );
or U85335 ( n17378, n17379, n17380 );
nor U85336 ( n48118, n48134, n48135 );
nor U85337 ( n48134, n48032, n48139 );
nor U85338 ( n48135, n48030, n48136 );
not U85339 ( n1308, n53925 );
nand U85340 ( n17776, n18044, n18045 );
nand U85341 ( n18045, n2785, n18046 );
nand U85342 ( n18044, n18049, n17868 );
not U85343 ( n2785, n17868 );
nand U85344 ( n18049, n17865, n17867 );
nand U85345 ( n50573, n50685, n50686 );
nand U85346 ( n50685, n50690, n50689 );
nand U85347 ( n50686, n50687, n50688 );
or U85348 ( n50687, n50689, n50690 );
xor U85349 ( n50562, n50441, n50712 );
xor U85350 ( n50712, n50439, n50440 );
nand U85351 ( n49986, n50124, n50125 );
nand U85352 ( n50124, n50129, n50128 );
nand U85353 ( n50125, n50126, n50127 );
or U85354 ( n50126, n50128, n50129 );
not U85355 ( n1264, n53927 );
nor U85356 ( n48775, n48786, n48787 );
nor U85357 ( n48786, n47941, n48122 );
nor U85358 ( n48787, n48136, n48722 );
nor U85359 ( n48710, n48136, n48628 );
nor U85360 ( n48616, n48136, n48534 );
nor U85361 ( n49076, n48136, n48994 );
nor U85362 ( n49250, n48136, n49183 );
nor U85363 ( n48881, n48136, n48814 );
nor U85364 ( n48981, n48136, n48895 );
nor U85365 ( n49345, n48136, n49279 );
nor U85366 ( n49438, n48136, n49357 );
nor U85367 ( n51670, n48136, n49450 );
nand U85368 ( n49665, n51658, n51659 );
nor U85369 ( n51659, n51660, n51661 );
nor U85370 ( n51658, n51669, n51670 );
nor U85371 ( n51660, n48122, n51665 );
nor U85372 ( n49159, n49170, n49171 );
nor U85373 ( n49170, n48122, n49086 );
nor U85374 ( n49171, n48136, n49089 );
nor U85375 ( n48507, n48520, n48521 );
nor U85376 ( n48520, n48139, n48433 );
nor U85377 ( n48521, n48136, n48432 );
nor U85378 ( n48222, n48235, n48236 );
nor U85379 ( n48235, n48122, n48155 );
nor U85380 ( n48236, n48136, n48154 );
nor U85381 ( n48402, n48415, n48416 );
nor U85382 ( n48415, n48122, n48350 );
nor U85383 ( n48416, n48136, n48349 );
xnor U85384 ( n50987, n51221, n50998 );
xor U85385 ( n51221, n50999, n50996 );
nand U85386 ( n18489, n18665, n18666 );
nand U85387 ( n18666, n18667, n18668 );
xor U85388 ( n50991, n50992, n1640 );
nor U85389 ( n15623, n15305, n5179 );
xnor U85390 ( n51675, n50619, n50621 );
nor U85391 ( n16150, n15305, n16135 );
nor U85392 ( n15725, n15305, n15717 );
nor U85393 ( n16355, n15305, n16347 );
nor U85394 ( n16250, n15305, n16242 );
nor U85395 ( n16048, n15305, n16039 );
nor U85396 ( n15940, n15305, n15932 );
nor U85397 ( n15835, n15305, n15827 );
nor U85398 ( n15527, n15305, n15518 );
nor U85399 ( n15420, n15305, n15412 );
nor U85400 ( n16503, n15305, n5168 );
nand U85401 ( n8136, n16473, n16474 );
nor U85402 ( n16474, n16475, n16477 );
nor U85403 ( n16473, n16503, n16504 );
nand U85404 ( n16477, n16478, n16479 );
nand U85405 ( n18041, n18270, n18271 );
nand U85406 ( n18270, n18275, n18123 );
nand U85407 ( n18271, n2772, n18272 );
nand U85408 ( n18275, n18120, n18122 );
nand U85409 ( n17872, n18037, n18038 );
nand U85410 ( n18037, n18041, n18042 );
nand U85411 ( n18038, n18039, n18040 );
or U85412 ( n18040, n18041, n18042 );
nand U85413 ( n17497, n17869, n17870 );
nand U85414 ( n17870, n17871, n17872 );
nand U85415 ( n18123, n18276, n18277 );
nand U85416 ( n18276, n18281, n18280 );
nand U85417 ( n18277, n18278, n18279 );
or U85418 ( n18278, n18280, n18281 );
and U85419 ( n50837, n51081, n51082 );
nand U85420 ( n51081, n51085, n51086 );
nand U85421 ( n51082, n51083, n51084 );
or U85422 ( n51083, n51085, n51086 );
xnor U85423 ( n17758, n17499, n17766 );
xor U85424 ( n17766, n17497, n17498 );
nand U85425 ( n17205, n17597, n17598 );
nand U85426 ( n17598, n17599, n17600 );
xor U85427 ( n18035, n17777, n18043 );
xnor U85428 ( n18043, n17778, n17776 );
xnor U85429 ( n18126, n18022, n18261 );
xnor U85430 ( n18261, n18021, n18023 );
nand U85431 ( n50563, n50706, n50707 );
nand U85432 ( n50706, n50711, n50710 );
nand U85433 ( n50707, n50708, n50709 );
or U85434 ( n50709, n50710, n50711 );
nand U85435 ( n17379, n17441, n17442 );
nand U85436 ( n17441, n17446, n17135 );
nand U85437 ( n17442, n2578, n17443 );
nand U85438 ( n17446, n17132, n17134 );
nand U85439 ( n17135, n17447, n17448 );
nand U85440 ( n17447, n17451, n17452 );
nand U85441 ( n17448, n17449, n17450 );
or U85442 ( n17450, n17451, n17452 );
xnor U85443 ( n50836, n50982, n50723 );
xor U85444 ( n50982, n50722, n50724 );
xnor U85445 ( n17465, n17159, n17466 );
xor U85446 ( n17466, n17156, n17158 );
xnor U85447 ( n17445, n17142, n17453 );
xor U85448 ( n17453, n17140, n17141 );
xor U85449 ( n17456, n17457, n2652 );
nand U85450 ( n17471, n17879, n17880 );
or U85451 ( n17879, n17883, n17884 );
nand U85452 ( n17880, n17881, n17882 );
nand U85453 ( n17881, n17883, n17884 );
nand U85454 ( n49744, n50082, n50083 );
nand U85455 ( n50082, n50087, n50086 );
nand U85456 ( n50083, n50084, n50085 );
or U85457 ( n50084, n50086, n50087 );
nand U85458 ( n18042, n18353, n18354 );
nand U85459 ( n18354, n18355, n18356 );
nor U85460 ( n18763, n18764, n18765 );
nor U85461 ( n18764, n18766, n18767 );
nor U85462 ( n18766, n18768, n18769 );
nand U85463 ( n50093, n50414, n50415 );
or U85464 ( n50414, n50418, n50419 );
nand U85465 ( n50415, n50416, n50417 );
nand U85466 ( n50416, n50418, n50419 );
xnor U85467 ( n17479, n17207, n17487 );
xor U85468 ( n17487, n17205, n17206 );
nand U85469 ( n17186, n17192, n17193 );
nand U85470 ( n17193, n17194, n17195 );
nand U85471 ( n50127, n50430, n50431 );
nand U85472 ( n50431, n1595, n50432 );
nand U85473 ( n50430, n50435, n50141 );
not U85474 ( n1595, n50141 );
nand U85475 ( n50435, n50138, n50140 );
nand U85476 ( n50116, n50564, n50565 );
nand U85477 ( n50564, n50568, n50569 );
nand U85478 ( n50565, n50566, n50567 );
or U85479 ( n50566, n50568, n50569 );
nand U85480 ( n17144, n17457, n2652 );
not U85481 ( n2373, n18769 );
or U85482 ( n18770, n18768, n2373 );
nand U85483 ( n16837, n16844, n16845 );
nand U85484 ( n16845, n16846, n16847 );
nand U85485 ( n16846, n16849, n16842 );
or U85486 ( n16847, n16848, n2742 );
nand U85487 ( n18530, n18629, n18630 );
nand U85488 ( n18629, n18634, n18633 );
nand U85489 ( n18630, n18631, n18632 );
or U85490 ( n18631, n18633, n18634 );
xnor U85491 ( n17729, n17737, n17463 );
xor U85492 ( n17737, n17462, n17464 );
nand U85493 ( n17462, n17885, n17886 );
nand U85494 ( n17886, n17887, n17888 );
or U85495 ( n17613, n17728, n17729 );
nand U85496 ( n21033, n2423, n19506 );
xor U85497 ( n17727, n17728, n17729 );
not U85498 ( n2378, n20986 );
and U85499 ( n20975, n20994, n20995 );
nand U85500 ( n20995, n20996, n2424 );
nor U85501 ( n20994, n20997, n20998 );
nor U85502 ( n20997, n2467, n21004 );
and U85503 ( n19169, n20989, n20990 );
nand U85504 ( n20990, n20982, n20986 );
nor U85505 ( n20989, n20978, n20984 );
and U85506 ( n18030, n18357, n18358 );
nand U85507 ( n18357, n18362, n18361 );
nand U85508 ( n18358, n18359, n18360 );
or U85509 ( n18359, n18361, n18362 );
nand U85510 ( n17615, n17729, n17728 );
nand U85511 ( n16852, n16855, n16856 );
nand U85512 ( n16856, n16857, n16858 );
nand U85513 ( n16838, n2740, n16839 );
nand U85514 ( n16839, n16840, n16841 );
not U85515 ( n2740, n16844 );
nand U85516 ( n16840, n2742, n2760 );
nand U85517 ( n17485, n17754, n17755 );
nand U85518 ( n17754, n17759, n17600 );
nand U85519 ( n17755, n2732, n17756 );
nand U85520 ( n17759, n17597, n17599 );
nand U85521 ( n17195, n17481, n17482 );
nand U85522 ( n17481, n17486, n17485 );
nand U85523 ( n17482, n17483, n17484 );
or U85524 ( n17483, n17485, n17486 );
not U85525 ( n2422, n20982 );
xor U85526 ( n17742, n18016, n17749 );
xor U85527 ( n18016, n17751, n17752 );
nand U85528 ( n17600, n17760, n17761 );
nand U85529 ( n17760, n17765, n17764 );
nand U85530 ( n17761, n17762, n17763 );
or U85531 ( n17762, n17764, n17765 );
xnor U85532 ( n50114, n50128, n50429 );
xnor U85533 ( n50429, n50127, n50129 );
nand U85534 ( n17616, n17731, n17732 );
nand U85535 ( n17731, n17736, n17735 );
nand U85536 ( n17732, n17733, n17734 );
or U85537 ( n17733, n17735, n17736 );
nand U85538 ( n17146, n17465, n2649 );
not U85539 ( n2649, n17457 );
not U85540 ( n64, n15290 );
xnor U85541 ( n17469, n17611, n17739 );
xnor U85542 ( n17739, n17610, n17612 );
nand U85543 ( n17056, n17132, n17133 );
nand U85544 ( n17133, n17134, n17135 );
xor U85545 ( n17605, n17486, n17753 );
xor U85546 ( n17753, n17484, n17485 );
nand U85547 ( n17032, n17178, n17179 );
nand U85548 ( n17178, n17183, n17182 );
nand U85549 ( n17179, n17180, n17181 );
or U85550 ( n17180, n17182, n17183 );
xor U85551 ( n45461, n51777, n51778 );
xor U85552 ( n51777, n51779, n51780 );
nand U85553 ( n45472, n51733, n51734 );
nand U85554 ( n51733, n45461, n45463 );
nand U85555 ( n51734, n45464, n51735 );
or U85556 ( n51735, n45463, n45461 );
nand U85557 ( n49814, n49817, n49818 );
nand U85558 ( n49818, n1655, n49819 );
nand U85559 ( n49817, n49824, n49825 );
nand U85560 ( n49819, n49820, n49821 );
nand U85561 ( n49825, n49826, n49827 );
nand U85562 ( n49826, n49829, n49822 );
or U85563 ( n49827, n49828, n1658 );
and U85564 ( n20973, n21006, n21007 );
nand U85565 ( n21007, n2425, n20971 );
nor U85566 ( n21006, n20962, n20967 );
not U85567 ( n1555, n49994 );
nand U85568 ( n17147, n17459, n17460 );
nand U85569 ( n17459, n17463, n17464 );
nand U85570 ( n17460, n17461, n17462 );
or U85571 ( n17461, n17463, n17464 );
xnor U85572 ( n18029, n18269, n18041 );
xor U85573 ( n18269, n18042, n18039 );
nand U85574 ( n45463, n51736, n51737 );
nand U85575 ( n51736, n45454, n45452 );
nand U85576 ( n51737, n45453, n51738 );
or U85577 ( n51738, n45452, n45454 );
nor U85578 ( n51743, n51744, n51745 );
nor U85579 ( n51744, n51746, n51747 );
nor U85580 ( n51746, n51748, n51749 );
nand U85581 ( n17878, n18018, n18019 );
nand U85582 ( n18018, n18022, n18023 );
nand U85583 ( n18019, n18020, n18021 );
or U85584 ( n18020, n18022, n18023 );
xor U85585 ( n11685, n18821, n18822 );
xor U85586 ( n18822, n18823, n18824 );
nand U85587 ( n11699, n18777, n18778 );
nand U85588 ( n18777, n11685, n11688 );
nand U85589 ( n18778, n11689, n18779 );
or U85590 ( n18779, n11688, n11685 );
not U85591 ( n2379, n20971 );
not U85592 ( n2425, n20969 );
nand U85593 ( n16789, n17137, n17138 );
nand U85594 ( n17137, n17142, n17141 );
nand U85595 ( n17138, n17139, n17140 );
or U85596 ( n17139, n17141, n17142 );
nand U85597 ( n17170, n17607, n17608 );
nand U85598 ( n17607, n17611, n17612 );
nand U85599 ( n17608, n17609, n17610 );
or U85600 ( n17609, n17611, n17612 );
nand U85601 ( n17606, n17747, n17748 );
nand U85602 ( n17747, n17752, n17751 );
nand U85603 ( n17748, n17749, n17750 );
or U85604 ( n17750, n17751, n17752 );
nand U85605 ( n17763, n18031, n18032 );
nand U85606 ( n18031, n18036, n17872 );
nand U85607 ( n18032, n2744, n18033 );
nand U85608 ( n18036, n17869, n17871 );
not U85609 ( n2412, n18765 );
xor U85610 ( n49850, n49851, n49852 );
nor U85611 ( n49852, n49853, n49854 );
nand U85612 ( n49851, n49963, n49964 );
nor U85613 ( n49853, n49860, n49856 );
xor U85614 ( n49838, n49839, n49840 );
nand U85615 ( n49964, n49965, n49966 );
not U85616 ( n1655, n49824 );
xor U85617 ( n17877, n18024, n17764 );
xor U85618 ( n18024, n17763, n17765 );
nand U85619 ( n17181, n17475, n17476 );
nand U85620 ( n17476, n2713, n17477 );
nand U85621 ( n17475, n17480, n17195 );
not U85622 ( n2713, n17195 );
nand U85623 ( n17480, n17192, n17194 );
nor U85624 ( n15604, n15290, n5179 );
xnor U85625 ( n49846, n49840, n49839 );
nor U85626 ( n16343, n15290, n16347 );
nor U85627 ( n16238, n15290, n16242 );
nor U85628 ( n16132, n15290, n16135 );
nor U85629 ( n16035, n15290, n16039 );
nor U85630 ( n15928, n15290, n15932 );
nor U85631 ( n15823, n15290, n15827 );
nor U85632 ( n15713, n15290, n15717 );
nor U85633 ( n15514, n15290, n15518 );
nor U85634 ( n15408, n15290, n15412 );
nor U85635 ( n16460, n15290, n5168 );
nand U85636 ( n8141, n16435, n16437 );
nor U85637 ( n16437, n16438, n16439 );
nor U85638 ( n16435, n16460, n16462 );
nand U85639 ( n16439, n16440, n16442 );
xnor U85640 ( n18719, n17663, n17665 );
nor U85641 ( n14929, n14948, n14949 );
nor U85642 ( n14948, n14830, n14954 );
nor U85643 ( n14949, n14828, n14950 );
nand U85644 ( n50000, n50100, n50101 );
or U85645 ( n50100, n50105, n50104 );
nand U85646 ( n50101, n50102, n50103 );
nand U85647 ( n50103, n50104, n50105 );
nor U85648 ( n16120, n14950, n16038 );
nor U85649 ( n16022, n14950, n15930 );
nor U85650 ( n15914, n14950, n15825 );
nor U85651 ( n15808, n14950, n15715 );
nor U85652 ( n16224, n14950, n16134 );
nor U85653 ( n15599, n14950, n15517 );
nor U85654 ( n15502, n14950, n15410 );
nor U85655 ( n16330, n14950, n16240 );
nor U85656 ( n16434, n14950, n16345 );
nor U85657 ( n15259, n15275, n15277 );
nor U85658 ( n15275, n14934, n15185 );
nor U85659 ( n15277, n14950, n15184 );
nor U85660 ( n15039, n15055, n15057 );
nor U85661 ( n15055, n14934, n14974 );
nor U85662 ( n15057, n14950, n14973 );
nor U85663 ( n15375, n15393, n15394 );
nor U85664 ( n15393, n14954, n15297 );
nor U85665 ( n15394, n14950, n15295 );
nor U85666 ( n18702, n18713, n18714 );
nor U85667 ( n18713, n14954, n16677 );
nor U85668 ( n18714, n14950, n16449 );
xnor U85669 ( n17168, n17182, n17474 );
xnor U85670 ( n17474, n17181, n17183 );
nand U85671 ( n18526, n18642, n18643 );
nand U85672 ( n18642, n18647, n18646 );
nand U85673 ( n18643, n18644, n18645 );
or U85674 ( n18644, n18646, n18647 );
xnor U85675 ( n45441, n51773, n51774 );
xor U85676 ( n51773, n51775, n51776 );
not U85677 ( n2868, n16936 );
nor U85678 ( n15687, n15700, n15702 );
nor U85679 ( n15700, n14735, n14934 );
nor U85680 ( n15702, n14950, n15613 );
not U85681 ( n2675, n17040 );
nand U85682 ( n11688, n18780, n18781 );
nand U85683 ( n18780, n11675, n11674 );
nand U85684 ( n18781, n11677, n18782 );
or U85685 ( n18782, n11674, n11675 );
nand U85686 ( n45431, n51763, n51764 );
nand U85687 ( n51764, n51765, n51766 );
nor U85688 ( n51763, n51767, n51768 );
nor U85689 ( n51767, n51766, n51772 );
nand U85690 ( n16859, n16862, n16863 );
nand U85691 ( n16863, n2778, n16864 );
nand U85692 ( n16862, n16869, n16870 );
nand U85693 ( n16864, n16865, n16866 );
nand U85694 ( n16870, n16871, n16872 );
nand U85695 ( n16871, n16874, n16867 );
or U85696 ( n16872, n16873, n2779 );
nor U85697 ( n18788, n18790, n18791 );
nor U85698 ( n18790, n18792, n18793 );
nor U85699 ( n48111, n48030, n48112 );
nor U85700 ( n48771, n48112, n48722 );
nor U85701 ( n48398, n48112, n48349 );
nor U85702 ( n48301, n48112, n48252 );
nor U85703 ( n48218, n48112, n48154 );
nor U85704 ( n49329, n48112, n49279 );
nor U85705 ( n49422, n48112, n49357 );
nor U85706 ( n49232, n48112, n49183 );
nor U85707 ( n49154, n48112, n49089 );
nor U85708 ( n49060, n48112, n48994 );
nor U85709 ( n48965, n48112, n48895 );
nor U85710 ( n48863, n48112, n48814 );
nor U85711 ( n48694, n48112, n48628 );
nor U85712 ( n48600, n48112, n48534 );
nor U85713 ( n48503, n48112, n48432 );
xor U85714 ( n11660, n18817, n18818 );
xor U85715 ( n18817, n18819, n18820 );
nor U85716 ( n49637, n48112, n49450 );
and U85717 ( n19364, n19366, n19368 );
nand U85718 ( n17046, n17154, n17155 );
or U85719 ( n17154, n17159, n17158 );
nand U85720 ( n17155, n17156, n17157 );
nand U85721 ( n17157, n17158, n17159 );
xor U85722 ( n16895, n16896, n16897 );
nor U85723 ( n16897, n16898, n16899 );
nand U85724 ( n16896, n17008, n17009 );
nor U85725 ( n16898, n16905, n16901 );
nand U85726 ( n16877, n16880, n16881 );
nand U85727 ( n16880, n16890, n16891 );
nand U85728 ( n16881, n16882, n16883 );
nor U85729 ( n16890, n16888, n17017 );
nand U85730 ( n17009, n17010, n17011 );
not U85731 ( n2778, n16869 );
nand U85732 ( n16281, n44114, n44115 );
nor U85733 ( n44115, n44116, n44117 );
nor U85734 ( n44114, n44208, n44209 );
nor U85735 ( n44116, n43486, n76361 );
and U85736 ( n19042, n19044, n19046 );
nor U85737 ( n49860, n49957, n49958 );
nor U85738 ( n49958, n49959, n49960 );
nor U85739 ( n49957, n49961, n49962 );
xor U85740 ( n51762, n52125, n53944 );
xor U85741 ( n53944, n52123, n52126 );
nand U85742 ( n45433, n51757, n51758 );
nand U85743 ( n51757, n51762, n51761 );
nand U85744 ( n51758, n51759, n51760 );
or U85745 ( n51760, n51761, n51762 );
nand U85746 ( n11648, n18807, n18808 );
nand U85747 ( n18808, n18809, n18810 );
nor U85748 ( n18807, n18811, n18812 );
nor U85749 ( n18811, n18810, n18816 );
nor U85750 ( n48100, n48030, n48101 );
xor U85751 ( n49623, n49624, n49625 );
xor U85752 ( n49856, n49861, n49862 );
nor U85753 ( n49862, n49863, n49864 );
nand U85754 ( n49861, n49953, n49954 );
nor U85755 ( n49863, n49870, n49866 );
nor U85756 ( n14912, n14828, n14913 );
xor U85757 ( n16682, n16684, n16685 );
nor U85758 ( n48390, n48101, n48349 );
nor U85759 ( n48293, n48101, n48252 );
nor U85760 ( n48195, n48101, n48154 );
nor U85761 ( n48762, n48101, n48722 );
nor U85762 ( n49224, n48101, n49183 );
nor U85763 ( n48855, n48101, n48814 );
nor U85764 ( n48494, n48101, n48432 );
nor U85765 ( n49320, n48101, n49279 );
nor U85766 ( n49129, n48101, n49089 );
nor U85767 ( n49051, n48101, n48994 );
nor U85768 ( n48956, n48101, n48895 );
nor U85769 ( n48669, n48101, n48628 );
nor U85770 ( n48591, n48101, n48534 );
nor U85771 ( n49413, n48101, n49357 );
nor U85772 ( n15682, n14913, n15613 );
nor U85773 ( n15254, n14913, n15184 );
nor U85774 ( n15144, n14913, n15077 );
nor U85775 ( n15034, n14913, n14973 );
nor U85776 ( n16414, n14913, n16345 );
nor U85777 ( n16312, n14913, n16240 );
nor U85778 ( n16100, n14913, n16038 );
nor U85779 ( n15993, n14913, n15930 );
nor U85780 ( n15894, n14913, n15825 );
nor U85781 ( n15785, n14913, n15715 );
nor U85782 ( n15579, n14913, n15517 );
nor U85783 ( n15473, n14913, n15410 );
nor U85784 ( n15370, n14913, n15295 );
nor U85785 ( n16202, n14913, n16134 );
nor U85786 ( n49608, n48101, n49450 );
nor U85787 ( n16663, n14913, n16449 );
and U85788 ( n49645, n53932, n53933 );
nand U85789 ( n53933, n53934, n1263 );
nor U85790 ( n53932, n53935, n53936 );
nor U85791 ( n53935, n1304, n53942 );
xor U85792 ( n18806, n20988, n19169 );
xor U85793 ( n20988, n19170, n19167 );
nand U85794 ( n11650, n18801, n18802 );
nand U85795 ( n18801, n18806, n18805 );
nand U85796 ( n18802, n18803, n18804 );
or U85797 ( n18804, n18805, n18806 );
not U85798 ( n2709, n20710 );
not U85799 ( n2693, n20763 );
not U85800 ( n2669, n20848 );
nand U85801 ( n9546, n10238, n10239 );
nor U85802 ( n10239, n10240, n10242 );
nor U85803 ( n10238, n10355, n10357 );
nor U85804 ( n10240, n9533, n76631 );
nor U85805 ( n16905, n17002, n17003 );
nor U85806 ( n17003, n17004, n17005 );
nor U85807 ( n17002, n17006, n17007 );
nor U85808 ( n14898, n14828, n14899 );
xor U85809 ( n16645, n16647, n16648 );
nor U85810 ( n15669, n14899, n15613 );
nor U85811 ( n15244, n14899, n15184 );
nor U85812 ( n15134, n14899, n15077 );
nor U85813 ( n15024, n14899, n14973 );
nor U85814 ( n16403, n14899, n16345 );
nor U85815 ( n16300, n14899, n16240 );
nor U85816 ( n16192, n14899, n16134 );
nor U85817 ( n16089, n14899, n16038 );
nor U85818 ( n15982, n14899, n15930 );
nor U85819 ( n15883, n14899, n15825 );
nor U85820 ( n15775, n14899, n15715 );
nor U85821 ( n15568, n14899, n15517 );
nor U85822 ( n15462, n14899, n15410 );
nor U85823 ( n15359, n14899, n15295 );
nor U85824 ( n49864, n49865, n1722 );
not U85825 ( n1722, n49866 );
nor U85826 ( n49865, n49867, n49868 );
nor U85827 ( n49867, n1729, n49869 );
nor U85828 ( n16627, n14899, n16449 );
xnor U85829 ( n49615, n53928, n53929 );
xnor U85830 ( n53928, n53930, n53931 );
nand U85831 ( n49646, n53893, n53894 );
nand U85832 ( n53893, n49615, n49617 );
nand U85833 ( n53894, n49618, n53895 );
or U85834 ( n53895, n49617, n49615 );
xor U85835 ( n16901, n16906, n16907 );
nor U85836 ( n16907, n16908, n16909 );
nand U85837 ( n16906, n16998, n16999 );
nor U85838 ( n16908, n16915, n16911 );
nor U85839 ( n20980, n20981, n20982 );
nor U85840 ( n20981, n20983, n20984 );
nor U85841 ( n20983, n20985, n20986 );
nand U85842 ( n49587, n53916, n53917 );
nand U85843 ( n53917, n53918, n1264 );
nor U85844 ( n53916, n53919, n53920 );
nor U85845 ( n53919, n53925, n53926 );
not U85846 ( n2623, n20355 );
nor U85847 ( n48089, n48030, n48090 );
nor U85848 ( n49870, n49948, n49949 );
nor U85849 ( n49949, n1725, n49950 );
nor U85850 ( n49948, n49951, n49952 );
nor U85851 ( n48754, n48090, n48722 );
nor U85852 ( n48382, n48090, n48349 );
nor U85853 ( n48285, n48090, n48252 );
nor U85854 ( n48187, n48090, n48154 );
nor U85855 ( n49312, n48090, n49279 );
nor U85856 ( n49216, n48090, n49183 );
nor U85857 ( n49121, n48090, n49089 );
nor U85858 ( n49043, n48090, n48994 );
nor U85859 ( n48948, n48090, n48895 );
nor U85860 ( n48847, n48090, n48814 );
nor U85861 ( n48661, n48090, n48628 );
nor U85862 ( n48583, n48090, n48534 );
nor U85863 ( n48485, n48090, n48432 );
nor U85864 ( n49405, n48090, n49357 );
nor U85865 ( n49580, n48090, n49450 );
and U85866 ( n16675, n20937, n20938 );
nand U85867 ( n20937, n16635, n16638 );
nand U85868 ( n20938, n16639, n20939 );
or U85869 ( n20939, n16638, n16635 );
xor U85870 ( n49595, n49596, n49597 );
nand U85871 ( n20987, n2380, n20986 );
nor U85872 ( n16909, n16910, n2842 );
not U85873 ( n2842, n16911 );
nor U85874 ( n16910, n16912, n16913 );
nor U85875 ( n16912, n2847, n16914 );
nand U85876 ( n16600, n20960, n20961 );
nand U85877 ( n20961, n20962, n2379 );
nor U85878 ( n20960, n20963, n20964 );
nor U85879 ( n20963, n20969, n20970 );
nand U85880 ( n49873, n49879, n49880 );
nand U85881 ( n49879, n1734, n49888 );
nand U85882 ( n49880, n49881, n49882 );
not U85883 ( n1734, n49881 );
and U85884 ( n16784, n16789, n16788 );
and U85885 ( n49590, n53899, n53900 );
nand U85886 ( n53899, n49542, n49544 );
nand U85887 ( n53900, n49543, n53901 );
or U85888 ( n53901, n49544, n49542 );
nor U85889 ( n14884, n14828, n14885 );
nor U85890 ( n15659, n14885, n15613 );
nor U85891 ( n15234, n14885, n15184 );
nor U85892 ( n15124, n14885, n15077 );
nor U85893 ( n15014, n14885, n14973 );
nor U85894 ( n16290, n14885, n16240 );
nor U85895 ( n16182, n14885, n16134 );
nor U85896 ( n16079, n14885, n16038 );
nor U85897 ( n15972, n14885, n15930 );
nor U85898 ( n15867, n14885, n15825 );
nor U85899 ( n15765, n14885, n15715 );
nor U85900 ( n15558, n14885, n15517 );
nor U85901 ( n15452, n14885, n15410 );
nor U85902 ( n15342, n14885, n15295 );
nor U85903 ( n16387, n14885, n16345 );
nor U85904 ( n16590, n14885, n16449 );
not U85905 ( n1712, n49959 );
nor U85906 ( n16915, n16993, n16994 );
nor U85907 ( n16994, n2844, n16995 );
nor U85908 ( n16993, n16996, n16997 );
nand U85909 ( n16266, n44298, n44299 );
nor U85910 ( n44298, n44308, n44309 );
nor U85911 ( n44299, n44300, n44301 );
nor U85912 ( n44308, n7587, n76361 );
not U85913 ( n2599, n20153 );
nand U85914 ( n49888, n49889, n49890 );
nand U85915 ( n49889, n1747, n49885 );
or U85916 ( n49890, n49891, n1749 );
nor U85917 ( n49842, n49972, n49973 );
not U85918 ( n2569, n20025 );
not U85919 ( n1527, n53388 );
and U85920 ( n16603, n20943, n20944 );
nand U85921 ( n20943, n16563, n16564 );
nand U85922 ( n20944, n16565, n20945 );
or U85923 ( n20945, n16564, n16563 );
xor U85924 ( n16608, n16610, n16612 );
nor U85925 ( n48064, n48030, n48065 );
nor U85926 ( n48746, n48065, n48722 );
nor U85927 ( n48374, n48065, n48349 );
nor U85928 ( n48277, n48065, n48252 );
nor U85929 ( n48179, n48065, n48154 );
nor U85930 ( n49397, n48065, n49357 );
nor U85931 ( n49304, n48065, n49279 );
nor U85932 ( n49113, n48065, n49089 );
nor U85933 ( n49019, n48065, n48994 );
nor U85934 ( n48936, n48065, n48895 );
nor U85935 ( n48839, n48065, n48814 );
nor U85936 ( n48653, n48065, n48628 );
nor U85937 ( n48559, n48065, n48534 );
nor U85938 ( n48476, n48065, n48432 );
nor U85939 ( n49208, n48065, n49183 );
nor U85940 ( n49534, n48065, n49450 );
xor U85941 ( n49550, n49551, n49552 );
nand U85942 ( n9531, n10468, n10469 );
nor U85943 ( n10468, n10480, n10482 );
nor U85944 ( n10469, n10470, n10472 );
nor U85945 ( n10480, n4933, n76631 );
not U85946 ( n2544, n19773 );
nor U85947 ( n16887, n17018, n17019 );
not U85948 ( n2509, n19657 );
nand U85949 ( n16932, n16933, n16934 );
nand U85950 ( n16933, n16936, n16930 );
or U85951 ( n16934, n16935, n2864 );
xor U85952 ( n16926, n16937, n16938 );
xor U85953 ( n16937, n16962, n16963 );
xor U85954 ( n16938, n16939, n16940 );
xor U85955 ( n16963, n16964, n16965 );
nand U85956 ( n16939, n16958, n16959 );
nand U85957 ( n16959, n16960, n16961 );
not U85958 ( n1500, n53274 );
not U85959 ( n2472, n19500 );
nor U85960 ( n14870, n14828, n14872 );
xor U85961 ( n16573, n16574, n16575 );
nor U85962 ( n16553, n14872, n16449 );
nor U85963 ( n15649, n14872, n15613 );
nor U85964 ( n15224, n14872, n15184 );
nor U85965 ( n15114, n14872, n15077 );
nor U85966 ( n15004, n14872, n14973 );
nor U85967 ( n16377, n14872, n16345 );
nor U85968 ( n16280, n14872, n16240 );
nor U85969 ( n16172, n14872, n16134 );
nor U85970 ( n16069, n14872, n16038 );
nor U85971 ( n15962, n14872, n15930 );
nor U85972 ( n15857, n14872, n15825 );
nor U85973 ( n15755, n14872, n15715 );
nor U85974 ( n15548, n14872, n15517 );
nor U85975 ( n15442, n14872, n15410 );
nor U85976 ( n15330, n14872, n15295 );
not U85977 ( n1449, n52947 );
not U85978 ( n1478, n53166 );
nor U85979 ( n48053, n48030, n48054 );
nor U85980 ( n48738, n48054, n48722 );
nor U85981 ( n48366, n48054, n48349 );
nor U85982 ( n48269, n48054, n48252 );
nor U85983 ( n48171, n48054, n48154 );
nor U85984 ( n49389, n48054, n49357 );
nor U85985 ( n49296, n48054, n49279 );
nor U85986 ( n49200, n48054, n49183 );
nor U85987 ( n49105, n48054, n49089 );
nor U85988 ( n49011, n48054, n48994 );
nor U85989 ( n48928, n48054, n48895 );
nor U85990 ( n48831, n48054, n48814 );
nor U85991 ( n48645, n48054, n48628 );
nor U85992 ( n48551, n48054, n48534 );
nor U85993 ( n48467, n48054, n48432 );
nor U85994 ( n49505, n48054, n49450 );
not U85995 ( n2648, n20529 );
not U85996 ( n2423, n21032 );
not U85997 ( n2829, n17004 );
not U85998 ( n1392, n52567 );
nor U85999 ( n14857, n14828, n14858 );
nor U86000 ( n48042, n48030, n48043 );
xor U86001 ( n49491, n49492, n49493 );
nor U86002 ( n15639, n14858, n15613 );
nor U86003 ( n15205, n14858, n15184 );
nor U86004 ( n15104, n14858, n15077 );
nor U86005 ( n14994, n14858, n14973 );
nor U86006 ( n16367, n14858, n16345 );
nor U86007 ( n16262, n14858, n16240 );
nor U86008 ( n16162, n14858, n16134 );
nor U86009 ( n16059, n14858, n16038 );
nor U86010 ( n15952, n14858, n15930 );
nor U86011 ( n15847, n14858, n15825 );
nor U86012 ( n15737, n14858, n15715 );
nor U86013 ( n15538, n14858, n15517 );
nor U86014 ( n15432, n14858, n15410 );
nor U86015 ( n15319, n14858, n15295 );
nor U86016 ( n48730, n48043, n48722 );
nor U86017 ( n48358, n48043, n48349 );
nor U86018 ( n48261, n48043, n48252 );
nor U86019 ( n48163, n48043, n48154 );
nor U86020 ( n49288, n48043, n49279 );
nor U86021 ( n49192, n48043, n49183 );
nor U86022 ( n49097, n48043, n49089 );
nor U86023 ( n49003, n48043, n48994 );
nor U86024 ( n48904, n48043, n48895 );
nor U86025 ( n48823, n48043, n48814 );
nor U86026 ( n48637, n48043, n48628 );
nor U86027 ( n48543, n48043, n48534 );
nor U86028 ( n48442, n48043, n48432 );
nor U86029 ( n49366, n48043, n49357 );
nor U86030 ( n16517, n14858, n16449 );
nor U86031 ( n49472, n48043, n49450 );
not U86032 ( n1353, n52255 );
not U86033 ( n2622, n20420 );
not U86034 ( n1313, n52144 );
nor U86035 ( n48029, n48030, n48031 );
nor U86036 ( n48721, n48031, n48722 );
nor U86037 ( n48348, n48031, n48349 );
nor U86038 ( n48251, n48031, n48252 );
nor U86039 ( n48153, n48031, n48154 );
nor U86040 ( n49356, n48031, n49357 );
nor U86041 ( n49278, n48031, n49279 );
nor U86042 ( n49182, n48031, n49183 );
nor U86043 ( n49088, n48031, n49089 );
nor U86044 ( n48993, n48031, n48994 );
nor U86045 ( n48894, n48031, n48895 );
nor U86046 ( n48813, n48031, n48814 );
nor U86047 ( n48627, n48031, n48628 );
nor U86048 ( n48533, n48031, n48534 );
nor U86049 ( n48431, n48031, n48432 );
not U86050 ( n2380, n20985 );
nor U86051 ( n49441, n48031, n49450 );
nand U86052 ( n40799, n41250, n41251 );
nand U86053 ( n41250, n41174, n41176 );
nand U86054 ( n41251, n41252, n41177 );
or U86055 ( n41252, n41176, n41174 );
nor U86056 ( n42285, n552, n40825 );
nand U86057 ( n41053, n41343, n41344 );
nand U86058 ( n41343, n40860, n40862 );
nand U86059 ( n41344, n41345, n40863 );
or U86060 ( n41345, n40862, n40860 );
nand U86061 ( n41034, n41360, n41361 );
nand U86062 ( n41361, n590, n40783 );
nor U86063 ( n41360, n41362, n41363 );
nor U86064 ( n41363, n607, n41364 );
nand U86065 ( n41176, n41255, n41256 );
nand U86066 ( n41256, n592, n41005 );
nor U86067 ( n41255, n41257, n41258 );
nor U86068 ( n41258, n609, n41259 );
nand U86069 ( n40982, n41355, n41356 );
nand U86070 ( n41355, n41032, n41034 );
nand U86071 ( n41356, n41357, n41035 );
or U86072 ( n41357, n41034, n41032 );
nand U86073 ( n40758, n41338, n41339 );
nand U86074 ( n41338, n41050, n41053 );
nand U86075 ( n41339, n41340, n41052 );
or U86076 ( n41340, n41053, n41050 );
nand U86077 ( n41194, n41350, n41351 );
nand U86078 ( n41350, n40980, n40982 );
nand U86079 ( n41351, n41352, n40983 );
or U86080 ( n41352, n40982, n40980 );
nand U86081 ( n41161, n41372, n41373 );
nand U86082 ( n41372, n40877, n40880 );
nand U86083 ( n41373, n41374, n40879 );
or U86084 ( n41374, n40880, n40877 );
nand U86085 ( n40964, n41267, n41268 );
nand U86086 ( n41267, n41272, n41271 );
nand U86087 ( n41268, n41269, n41270 );
or U86088 ( n41269, n41271, n41272 );
nor U86089 ( n41362, n41365, n40781 );
nor U86090 ( n41365, n40783, n40782 );
nor U86091 ( n41257, n41260, n41003 );
nor U86092 ( n41260, n41005, n41004 );
nor U86093 ( n41244, n41246, n41248 );
nand U86094 ( n41248, n41249, n40799 );
or U86095 ( n41249, n40800, n40797 );
nand U86096 ( n41270, n41324, n41325 );
nand U86097 ( n41324, n40723, n40725 );
nand U86098 ( n41325, n41326, n40726 );
or U86099 ( n41326, n40725, n40723 );
and U86100 ( n75765, n814, n812 );
and U86101 ( n41111, n41333, n41334 );
nand U86102 ( n41333, n40756, n40758 );
nand U86103 ( n41334, n41335, n40759 );
or U86104 ( n41335, n40758, n40756 );
not U86105 ( n2598, n20210 );
nand U86106 ( n41207, n41208, n41209 );
nand U86107 ( n41208, n584, n41024 );
nand U86108 ( n41209, n41210, n76850 );
nor U86109 ( n41210, n41211, n41212 );
and U86110 ( n75766, n2197, n2153 );
nor U86111 ( n37770, n1893, n36423 );
nand U86112 ( n36588, n36990, n36991 );
nand U86113 ( n36990, n36647, n36648 );
nand U86114 ( n36991, n36645, n36992 );
or U86115 ( n36992, n36648, n36647 );
nand U86116 ( n36727, n36965, n36966 );
nand U86117 ( n36965, n36351, n36353 );
nand U86118 ( n36966, n36967, n36354 );
or U86119 ( n36967, n36353, n36351 );
nand U86120 ( n36666, n36978, n36979 );
nand U86121 ( n36978, n36458, n36460 );
nand U86122 ( n36979, n36980, n36461 );
or U86123 ( n36980, n36460, n36458 );
nand U86124 ( n36795, n36869, n36870 );
nand U86125 ( n36870, n1984, n36612 );
nor U86126 ( n36869, n36871, n36872 );
nor U86127 ( n36872, n1989, n36873 );
nand U86128 ( n36647, n36998, n36999 );
nand U86129 ( n36999, n1912, n36380 );
nor U86130 ( n36998, n37000, n37001 );
nor U86131 ( n37001, n1917, n37002 );
nand U86132 ( n36813, n36985, n36986 );
nand U86133 ( n36985, n36585, n36588 );
nand U86134 ( n36986, n36987, n36587 );
or U86135 ( n36987, n36588, n36585 );
nand U86136 ( n36778, n37010, n37011 );
nand U86137 ( n37011, n36487, n36486 );
nor U86138 ( n37010, n37012, n37013 );
nor U86139 ( n37013, n37014, n37015 );
nand U86140 ( n36569, n36880, n36881 );
nand U86141 ( n36880, n36885, n36884 );
nand U86142 ( n36881, n36882, n36883 );
or U86143 ( n36882, n36884, n36885 );
nor U86144 ( n37012, n36485, n37017 );
nand U86145 ( n37017, n37018, n2008 );
not U86146 ( n2008, n37014 );
nand U86147 ( n37018, n1849, n2040 );
nor U86148 ( n37000, n37003, n36378 );
nor U86149 ( n37003, n36380, n36379 );
nor U86150 ( n36871, n36874, n36610 );
nor U86151 ( n36874, n36612, n36611 );
and U86152 ( n36397, n36864, n36865 );
nand U86153 ( n36864, n36793, n36795 );
nand U86154 ( n36865, n36866, n36796 );
or U86155 ( n36866, n36795, n36793 );
nand U86156 ( n36883, n36956, n36957 );
nand U86157 ( n36956, n36318, n36320 );
nand U86158 ( n36957, n36958, n36321 );
or U86159 ( n36958, n36320, n36318 );
nand U86160 ( n36407, n36408, n36409 );
nand U86161 ( n36408, n76821, n36442 );
nand U86162 ( n36409, n76831, n36410 );
nand U86163 ( n36410, n36411, n36412 );
nand U86164 ( n36353, n36970, n36971 );
nand U86165 ( n36970, n36666, n36665 );
nand U86166 ( n36971, n36663, n36972 );
or U86167 ( n36972, n36665, n36666 );
not U86168 ( n2154, n40489 );
nand U86169 ( n36297, n36298, n36299 );
nand U86170 ( n36298, n76821, n36305 );
nand U86171 ( n36299, n76830, n36300 );
xor U86172 ( n36300, n36301, n36302 );
nor U86173 ( n14843, n14828, n14844 );
xor U86174 ( n16499, n16500, n16502 );
nand U86175 ( n16251, n44441, n44442 );
nor U86176 ( n44442, n44443, n44444 );
nor U86177 ( n44441, n44480, n44481 );
nor U86178 ( n44443, n7627, n76361 );
nand U86179 ( n36826, n36827, n36828 );
nand U86180 ( n36827, n76823, n36925 );
nand U86181 ( n36828, n36829, n36830 );
nor U86182 ( n36829, n36842, n36843 );
nor U86183 ( n15195, n14844, n15184 );
nor U86184 ( n15094, n14844, n15077 );
nor U86185 ( n14984, n14844, n14973 );
nor U86186 ( n15629, n14844, n15613 );
nor U86187 ( n16152, n14844, n16134 );
nor U86188 ( n15727, n14844, n15715 );
nor U86189 ( n15308, n14844, n15295 );
nor U86190 ( n16357, n14844, n16345 );
nor U86191 ( n16252, n14844, n16240 );
nor U86192 ( n16049, n14844, n16038 );
nor U86193 ( n15942, n14844, n15930 );
nor U86194 ( n15837, n14844, n15825 );
nor U86195 ( n15528, n14844, n15517 );
nor U86196 ( n15422, n14844, n15410 );
nor U86197 ( n16475, n14844, n16449 );
not U86198 ( n2568, n19991 );
not U86199 ( n1269, n51748 );
nor U86200 ( n37014, n36486, n36487 );
nor U86201 ( n36424, n76807, n37765 );
nand U86202 ( n37766, n37772, n36265 );
nand U86203 ( n37772, n37773, n37104 );
nor U86204 ( n37773, n76801, n2064 );
not U86205 ( n2065, n37297 );
nor U86206 ( n49589, n76321, n76835 );
nor U86207 ( n14827, n14828, n14829 );
nor U86208 ( n16438, n14829, n16449 );
nor U86209 ( n16344, n14829, n16345 );
nor U86210 ( n16239, n14829, n16240 );
nor U86211 ( n16133, n14829, n16134 );
nor U86212 ( n16037, n14829, n16038 );
nor U86213 ( n15929, n14829, n15930 );
nor U86214 ( n15824, n14829, n15825 );
nor U86215 ( n15714, n14829, n15715 );
nor U86216 ( n15612, n14829, n15613 );
nor U86217 ( n15515, n14829, n15517 );
nor U86218 ( n15409, n14829, n15410 );
nor U86219 ( n15294, n14829, n15295 );
nor U86220 ( n15183, n14829, n15184 );
nor U86221 ( n15075, n14829, n15077 );
nor U86222 ( n14972, n14829, n14973 );
nor U86223 ( n37287, n37288, n1893 );
nor U86224 ( n37243, n37247, n37248 );
nor U86225 ( n37247, n37246, n37245 );
nand U86226 ( n37248, n37249, n37250 );
or U86227 ( n37249, n37254, n37253 );
nor U86228 ( n37231, n37235, n37236 );
nor U86229 ( n37235, n37234, n37233 );
nand U86230 ( n37236, n37237, n37238 );
or U86231 ( n37237, n37242, n37241 );
nor U86232 ( n37270, n37272, n37273 );
nor U86233 ( n37272, n37274, n37275 );
nand U86234 ( n37275, n37276, n37277 );
nand U86235 ( n37277, n37278, n37279 );
nor U86236 ( n37255, n37258, n37259 );
nor U86237 ( n37258, n37257, n36667 );
nand U86238 ( n37259, n37260, n37261 );
nand U86239 ( n37261, n37262, n37263 );
nor U86240 ( n37262, n37264, n37265 );
nor U86241 ( n37264, n37266, n37267 );
nand U86242 ( n37267, n37268, n37269 );
nand U86243 ( n37269, n37270, n37271 );
nand U86244 ( n37250, n37251, n37252 );
nand U86245 ( n37252, n37253, n37254 );
nor U86246 ( n37251, n37255, n37256 );
and U86247 ( n37256, n36667, n37257 );
nor U86248 ( n37219, n37223, n37224 );
nor U86249 ( n37223, n37222, n37221 );
nand U86250 ( n37224, n37225, n37226 );
or U86251 ( n37225, n37230, n37229 );
nor U86252 ( n37207, n37211, n37212 );
nor U86253 ( n37211, n37210, n37209 );
nand U86254 ( n37212, n37213, n37214 );
or U86255 ( n37213, n37218, n37217 );
nor U86256 ( n37195, n37199, n37200 );
nor U86257 ( n37199, n37198, n37197 );
nand U86258 ( n37200, n37201, n37202 );
or U86259 ( n37201, n37206, n37205 );
nor U86260 ( n37183, n37187, n37188 );
nor U86261 ( n37187, n37186, n37185 );
nand U86262 ( n37188, n37189, n37190 );
or U86263 ( n37189, n37194, n37193 );
nor U86264 ( n37172, n37175, n37176 );
nor U86265 ( n37175, n37174, n36339 );
nand U86266 ( n37176, n37177, n37178 );
or U86267 ( n37177, n37182, n37181 );
nand U86268 ( n37214, n37215, n37216 );
nand U86269 ( n37216, n37217, n37218 );
nor U86270 ( n37215, n37219, n37220 );
and U86271 ( n37220, n37221, n37222 );
nand U86272 ( n37202, n37203, n37204 );
nand U86273 ( n37204, n37205, n37206 );
nor U86274 ( n37203, n37207, n37208 );
and U86275 ( n37208, n37209, n37210 );
nand U86276 ( n37238, n37239, n37240 );
nand U86277 ( n37240, n37241, n37242 );
nor U86278 ( n37239, n37243, n37244 );
and U86279 ( n37244, n37245, n37246 );
nand U86280 ( n37190, n37191, n37192 );
nand U86281 ( n37192, n37193, n37194 );
nor U86282 ( n37191, n37195, n37196 );
and U86283 ( n37196, n37197, n37198 );
nand U86284 ( n37226, n37227, n37228 );
nand U86285 ( n37228, n37229, n37230 );
nor U86286 ( n37227, n37231, n37232 );
and U86287 ( n37232, n37233, n37234 );
nand U86288 ( n37168, n37169, n37170 );
nand U86289 ( n37170, n37171, n36633 );
nor U86290 ( n37169, n37172, n37173 );
and U86291 ( n37173, n36339, n37174 );
nor U86292 ( n37128, n37139, n37140 );
nand U86293 ( n37140, n37141, n37142 );
nand U86294 ( n37139, n37144, n37145 );
nand U86295 ( n37142, n2190, n37143 );
nor U86296 ( n37161, n37165, n37166 );
nor U86297 ( n37165, n37164, n37163 );
nand U86298 ( n37166, n37167, n37168 );
or U86299 ( n37167, n36633, n37171 );
nor U86300 ( n37150, n37154, n37155 );
nor U86301 ( n37154, n37153, n37152 );
nand U86302 ( n37155, n37156, n37157 );
or U86303 ( n37156, n36925, n37160 );
nand U86304 ( n37157, n37158, n37159 );
nand U86305 ( n37159, n37160, n36925 );
nor U86306 ( n37158, n37161, n37162 );
and U86307 ( n37162, n37163, n37164 );
nand U86308 ( n37118, n37119, n37120 );
nor U86309 ( n37119, n37309, n37310 );
nor U86310 ( n37120, n37121, n37122 );
nand U86311 ( n37310, n37311, n37312 );
nand U86312 ( n36541, n36542, n36543 );
nand U86313 ( n36542, n76821, n36551 );
nand U86314 ( n36543, n76831, n36544 );
nand U86315 ( n36544, n36545, n36546 );
not U86316 ( n2508, n19611 );
nand U86317 ( n39127, n37456, n39315 );
nand U86318 ( n39315, n39316, n37557 );
nand U86319 ( n39104, n39124, n37594 );
nand U86320 ( n39124, n39125, n39126 );
and U86321 ( n39125, n39128, n37512 );
nand U86322 ( n39126, n37503, n39127 );
nand U86323 ( n39378, n37593, n39429 );
nand U86324 ( n39429, n39430, n37553 );
nand U86325 ( n39554, n37573, n39730 );
nand U86326 ( n39730, n39731, n37567 );
nand U86327 ( n39020, n37595, n39068 );
nand U86328 ( n39068, n1903, n37596 );
nor U86329 ( n39009, n1900, n38865 );
nand U86330 ( n39848, n37579, n39981 );
nand U86331 ( n39981, n39982, n37583 );
nand U86332 ( n37591, n40196, n40197 );
nor U86333 ( n40196, n37412, n40199 );
nand U86334 ( n40197, n40198, n37276 );
nor U86335 ( n40199, n37411, n1914 );
nor U86336 ( n40198, n1905, n1910 );
not U86337 ( n1910, n37472 );
nand U86338 ( n38172, n38914, n38915 );
nor U86339 ( n38914, n38950, n38951 );
nor U86340 ( n38915, n38916, n38917 );
nor U86341 ( n38950, n2188, n38822 );
nand U86342 ( n40273, n37398, n40279 );
nand U86343 ( n40279, n37384, n37401 );
nand U86344 ( n39982, n37263, n40013 );
nand U86345 ( n40013, n40014, n37260 );
nand U86346 ( n39482, n39551, n37453 );
nand U86347 ( n39551, n39552, n39553 );
and U86348 ( n39552, n39555, n39556 );
nand U86349 ( n39553, n37563, n39554 );
nand U86350 ( n37398, n2098, n37023 );
nor U86351 ( n38929, n2132, n38931 );
nor U86352 ( n38931, n38932, n38933 );
nor U86353 ( n38932, n2034, n37532 );
nand U86354 ( n39316, n37554, n39377 );
nand U86355 ( n39377, n39378, n37555 );
nand U86356 ( n38933, n39006, n39007 );
nor U86357 ( n39006, n39010, n39011 );
nor U86358 ( n39007, n39008, n39009 );
nor U86359 ( n39010, n1900, n37513 );
nand U86360 ( n39731, n37574, n39797 );
nand U86361 ( n39797, n39798, n37569 );
nand U86362 ( n38633, n38890, n38891 );
nor U86363 ( n38891, n38892, n38893 );
nor U86364 ( n38890, n38913, n38172 );
nor U86365 ( n38892, n2190, n38604 );
nand U86366 ( n38886, n37535, n39019 );
nand U86367 ( n39019, n39020, n37460 );
nand U86368 ( n38926, n38927, n38928 );
nor U86369 ( n38927, n38934, n38935 );
nor U86370 ( n38928, n38929, n38930 );
nor U86371 ( n38934, n38875, n38877 );
and U86372 ( n39798, n39843, n37420 );
nand U86373 ( n39843, n39844, n37577 );
nor U86374 ( n39844, n39846, n39847 );
nor U86375 ( n39846, n1948, n37442 );
nor U86376 ( n39008, n1900, n38866 );
nand U86377 ( n38169, n38170, n38171 );
nand U86378 ( n38171, n76815, n2138 );
nand U86379 ( n38170, n76811, n38172 );
nand U86380 ( n2801, n38157, n38158 );
nor U86381 ( n38158, n38159, n38160 );
nor U86382 ( n38157, n38168, n38169 );
nand U86383 ( n38160, n38161, n38162 );
nor U86384 ( n16529, n76575, n76789 );
nand U86385 ( n40778, n41163, n41162 );
nor U86386 ( n41364, n590, n40783 );
nand U86387 ( n38818, n38883, n38884 );
and U86388 ( n38883, n37507, n38887 );
nand U86389 ( n38884, n38885, n38886 );
nand U86390 ( n38887, n2134, n37389 );
nand U86391 ( n38627, n38760, n38761 );
nor U86392 ( n38761, n38762, n38763 );
nor U86393 ( n38760, n38774, n38136 );
nor U86394 ( n38762, n38601, n38135 );
nand U86395 ( n38778, n38779, n38780 );
nand U86396 ( n38779, n37361, n38789 );
nand U86397 ( n38780, n38781, n37361 );
nand U86398 ( n38789, n38790, n38791 );
nand U86399 ( n9516, n10629, n10630 );
nor U86400 ( n10630, n10632, n10633 );
nor U86401 ( n10629, n10678, n10679 );
nor U86402 ( n10632, n4973, n76631 );
nor U86403 ( n38806, n38808, n38809 );
nor U86404 ( n38809, n38773, n38810 );
nor U86405 ( n38808, n2144, n38811 );
nor U86406 ( n38811, n38812, n38813 );
nand U86407 ( n38132, n38133, n38134 );
or U86408 ( n38134, n38135, n38109 );
nand U86409 ( n38133, n76811, n38136 );
nand U86410 ( n36375, n36780, n36779 );
nor U86411 ( n37002, n1912, n36380 );
nand U86412 ( n37411, n1909, n36381 );
nand U86413 ( n36622, n36623, n36624 );
nand U86414 ( n36623, n76822, n36633 );
nand U86415 ( n36624, n76831, n36625 );
nand U86416 ( n36625, n36626, n36627 );
or U86417 ( n36627, n75767, n36629 );
xnor U86418 ( n75767, n36630, n2021 );
or U86419 ( n40777, n41162, n41163 );
nor U86420 ( n38880, n38881, n38882 );
nor U86421 ( n38881, n1902, n38866 );
nor U86422 ( n38882, n1902, n38865 );
nand U86423 ( n38630, n38826, n38827 );
nor U86424 ( n38827, n38828, n38829 );
nor U86425 ( n38826, n38847, n38156 );
nor U86426 ( n38828, n2192, n38604 );
nand U86427 ( n38156, n38848, n38849 );
nand U86428 ( n38849, n2074, n36442 );
nor U86429 ( n38848, n38850, n38851 );
nor U86430 ( n38851, n38834, n38852 );
nand U86431 ( n39488, n39609, n39610 );
nand U86432 ( n39610, n39611, n39612 );
nand U86433 ( n39419, n39485, n39486 );
nand U86434 ( n39486, n39487, n39488 );
nor U86435 ( n40028, n40103, n40104 );
nor U86436 ( n40104, n40105, n40106 );
nor U86437 ( n40105, n40107, n40108 );
and U86438 ( n40108, n40109, n40110 );
nand U86439 ( n39369, n39417, n39418 );
nand U86440 ( n39418, n39419, n39420 );
nor U86441 ( n40282, n2155, n1893 );
nand U86442 ( n38857, n38835, n38876 );
nand U86443 ( n38876, n38877, n38838 );
nand U86444 ( n39742, n39888, n39889 );
nand U86445 ( n39889, n39890, n39891 );
and U86446 ( n39888, n39892, n39893 );
nand U86447 ( n39611, n39666, n39677 );
nand U86448 ( n39677, n39678, n39669 );
nor U86449 ( n38874, n38875, n38857 );
nand U86450 ( n40112, n40226, n40227 );
nand U86451 ( n40227, n40228, n40229 );
nand U86452 ( n40228, n40230, n40231 );
nand U86453 ( n39892, n39900, n39898 );
and U86454 ( n39900, n39901, n39902 );
nand U86455 ( n39072, n39132, n39133 );
nand U86456 ( n39133, n39134, n39135 );
nor U86457 ( n39254, n2104, n1887 );
not U86458 ( n2104, n39255 );
nand U86459 ( n39134, n39181, n39182 );
nand U86460 ( n39182, n39183, n39184 );
nand U86461 ( n40110, n1888, n40111 );
not U86462 ( n1888, n40112 );
nand U86463 ( n39183, n39252, n39253 );
and U86464 ( n39252, n39256, n39257 );
nand U86465 ( n39253, n39254, n2052 );
nand U86466 ( n39257, n2058, n39255 );
nor U86467 ( n40023, n40025, n40027 );
or U86468 ( n40027, n40028, n40029 );
nand U86469 ( n2806, n38140, n38141 );
nor U86470 ( n38141, n38142, n38143 );
nor U86471 ( n38140, n38152, n38153 );
nand U86472 ( n38143, n38144, n38145 );
nand U86473 ( n38153, n38154, n38155 );
nand U86474 ( n38155, n76815, n2145 );
nand U86475 ( n38154, n76811, n38156 );
or U86476 ( n36374, n36779, n36780 );
not U86477 ( n2470, n19462 );
nor U86478 ( n38862, n38863, n38864 );
nor U86479 ( n38863, n38818, n38866 );
nor U86480 ( n38864, n38818, n38865 );
not U86481 ( n1914, n37276 );
nand U86482 ( n62866, n41590, n62978 );
nand U86483 ( n62978, n62979, n41594 );
nand U86484 ( n62395, n62460, n62461 );
and U86485 ( n62460, n62467, n62468 );
nand U86486 ( n62461, n740, n62462 );
nand U86487 ( n62468, n41134, n76388 );
nand U86488 ( n62979, n42098, n63299 );
nand U86489 ( n63299, n63300, n41593 );
nand U86490 ( n64809, n41560, n65947 );
nand U86491 ( n65947, n65948, n42081 );
nand U86492 ( n65948, n41569, n65949 );
nand U86493 ( n66441, n42000, n66747 );
nand U86494 ( n66747, n41990, n42011 );
nand U86495 ( n64525, n64806, n64807 );
nand U86496 ( n64806, n64810, n42058 );
nand U86497 ( n64807, n64808, n670 );
nand U86498 ( n64810, n64811, n64812 );
nand U86499 ( n66219, n42087, n66299 );
nand U86500 ( n66299, n565, n42084 );
nand U86501 ( n64376, n41544, n64524 );
nand U86502 ( n64524, n64525, n42045 );
nor U86503 ( n66035, n66107, n41567 );
and U86504 ( n66107, n66108, n66109 );
nor U86505 ( n66108, n643, n41577 );
nand U86506 ( n66371, n42001, n66440 );
nand U86507 ( n66440, n66441, n41989 );
nor U86508 ( n45487, n45493, n45363 );
nand U86509 ( n42000, n785, n41377 );
nand U86510 ( n65949, n66035, n41578 );
nand U86511 ( n62776, n41586, n62865 );
nand U86512 ( n62865, n62866, n41595 );
nand U86513 ( n63300, n63703, n63704 );
nand U86514 ( n63703, n63708, n41596 );
nand U86515 ( n63704, n63705, n63706 );
nand U86516 ( n63708, n41532, n63709 );
not U86517 ( n565, n66367 );
nand U86518 ( n66109, n66219, n41562 );
nand U86519 ( n63706, n41546, n64375 );
nand U86520 ( n64375, n64376, n41542 );
and U86521 ( n64808, n42079, n64809 );
not U86522 ( n2430, n19188 );
nand U86523 ( n40283, n2157, n2098 );
nand U86524 ( n36331, n36332, n36333 );
nand U86525 ( n36332, n76821, n36339 );
nand U86526 ( n36333, n76832, n36334 );
xnor U86527 ( n36334, n36335, n36336 );
nand U86528 ( n55790, n61392, n45493 );
nor U86529 ( n61392, n61442, n61296 );
nor U86530 ( n61442, n45492, n61443 );
nand U86531 ( n45759, n61600, n61601 );
nand U86532 ( n61601, n813, n40834 );
nor U86533 ( n61600, n61602, n61603 );
nor U86534 ( n61603, n61586, n61604 );
nor U86535 ( n61629, n61630, n61631 );
nor U86536 ( n61630, n564, n61618 );
nor U86537 ( n61631, n564, n61617 );
nand U86538 ( n1581, n45742, n45743 );
nor U86539 ( n45743, n45744, n45745 );
nor U86540 ( n45742, n45755, n45756 );
nand U86541 ( n45745, n45746, n45747 );
nand U86542 ( n39291, n39417, n39425 );
nand U86543 ( n39425, n39426, n39420 );
nand U86544 ( n39490, n39609, n39613 );
nand U86545 ( n39613, n39614, n39612 );
nand U86546 ( n38905, n39132, n39136 );
nand U86547 ( n39136, n39137, n39135 );
nand U86548 ( n39614, n39666, n39667 );
nand U86549 ( n39667, n39668, n39669 );
nand U86550 ( n39426, n39485, n39489 );
nand U86551 ( n39489, n39487, n39490 );
nand U86552 ( n39137, n39181, n39185 );
nand U86553 ( n39185, n39186, n39184 );
nand U86554 ( n39186, n39256, n39258 );
nand U86555 ( n39258, n39259, n39255 );
nand U86556 ( n38860, n38835, n38878 );
nand U86557 ( n38878, n38879, n38838 );
nor U86558 ( n61614, n61615, n61616 );
nor U86559 ( n61615, n61438, n61618 );
nor U86560 ( n61616, n61438, n61617 );
nor U86561 ( n38920, n38922, n38866 );
nand U86562 ( n38917, n38918, n38919 );
nand U86563 ( n38918, n38923, n38921 );
nand U86564 ( n38919, n38920, n38921 );
nor U86565 ( n38923, n38922, n38865 );
nor U86566 ( n49647, n76316, n76835 );
nor U86567 ( n38954, n38922, n37513 );
nand U86568 ( n38790, n38793, n38771 );
nand U86569 ( n40904, n41083, n41084 );
nand U86570 ( n41083, n40797, n40799 );
nand U86571 ( n41084, n41085, n40800 );
or U86572 ( n41085, n40799, n40797 );
nor U86573 ( n37274, n1919, n36589 );
not U86574 ( n607, n40782 );
nand U86575 ( n42001, n786, n40784 );
nor U86576 ( n37592, n37265, n40070 );
and U86577 ( n40070, n40071, n37273 );
nor U86578 ( n40071, n1927, n37266 );
nand U86579 ( n38636, n38959, n38960 );
nor U86580 ( n38960, n38961, n38962 );
nor U86581 ( n38959, n38976, n38188 );
nand U86582 ( n38962, n38963, n38964 );
nand U86583 ( n40229, n2158, n1909 );
not U86584 ( n1927, n37268 );
nand U86585 ( n38184, n38185, n38186 );
nand U86586 ( n38186, n38187, n76818 );
nand U86587 ( n38185, n76811, n38188 );
nand U86588 ( n2796, n38173, n38174 );
nor U86589 ( n38174, n38175, n38176 );
nor U86590 ( n38173, n38183, n38184 );
nand U86591 ( n38175, n38180, n38181 );
not U86592 ( n1917, n36379 );
not U86593 ( n2043, n37513 );
nor U86594 ( n40327, n2072, n2069 );
nand U86595 ( n40825, n42286, n40665 );
nand U86596 ( n42286, n42287, n41472 );
nand U86597 ( n42279, n76844, n42184 );
nand U86598 ( n37279, n1913, n36649 );
nor U86599 ( n39014, n39015, n39016 );
nor U86600 ( n39015, n38866, n38886 );
nor U86601 ( n39016, n38865, n38886 );
nand U86602 ( n36496, n36497, n36498 );
nand U86603 ( n36497, n76821, n36512 );
nand U86604 ( n36498, n36499, n76830 );
nor U86605 ( n36499, n36500, n36501 );
nand U86606 ( n62677, n63303, n63304 );
and U86607 ( n63303, n63309, n63310 );
nand U86608 ( n63304, n63305, n63306 );
nand U86609 ( n63310, n63311, n41178 );
nand U86610 ( n64024, n64230, n64231 );
nand U86611 ( n64231, n64232, n64233 );
nand U86612 ( n64804, n65338, n65339 );
nand U86613 ( n65338, n65342, n673 );
nand U86614 ( n65339, n65340, n65341 );
not U86615 ( n673, n65343 );
nor U86616 ( n66752, n624, n552 );
nand U86617 ( n66205, n66750, n66751 );
nand U86618 ( n66751, n66752, n66753 );
nor U86619 ( n66195, n66197, n66199 );
nand U86620 ( n66199, n66200, n66201 );
nand U86621 ( n66200, n66202, n66203 );
nor U86622 ( n66202, n66208, n66209 );
not U86623 ( n543, n66116 );
nand U86624 ( n63306, n64022, n64023 );
nand U86625 ( n64023, n64024, n64025 );
and U86626 ( n65340, n65945, n65946 );
nand U86627 ( n64232, n64377, n64378 );
nand U86628 ( n64377, n64381, n690 );
nand U86629 ( n64378, n64379, n64380 );
not U86630 ( n690, n64382 );
nor U86631 ( n39013, n39017, n39018 );
nor U86632 ( n39017, n37513, n38886 );
nor U86633 ( n39018, n38956, n38886 );
xor U86634 ( n45514, n45515, n45516 );
nor U86635 ( n36500, n36506, n36507 );
xor U86636 ( n36506, n36511, n2020 );
nand U86637 ( n36507, n36508, n2018 );
nand U86638 ( n36508, n36509, n36510 );
nand U86639 ( n37271, n1925, n36817 );
nand U86640 ( n36739, n36740, n36741 );
nand U86641 ( n36740, n76822, n36747 );
nand U86642 ( n36741, n76830, n36742 );
xnor U86643 ( n36742, n36743, n36744 );
not U86644 ( n1670, n49829 );
nor U86645 ( n62269, n61617, n61633 );
nand U86646 ( n46003, n62255, n62256 );
nand U86647 ( n62256, n813, n40950 );
nor U86648 ( n62255, n62257, n62258 );
nor U86649 ( n62257, n62276, n41926 );
nand U86650 ( n62260, n62266, n62267 );
nor U86651 ( n62266, n62270, n62271 );
nor U86652 ( n62267, n62268, n62269 );
nor U86653 ( n62270, n41487, n61633 );
not U86654 ( n624, n42184 );
buf U86655 ( n76248, n76247 );
nand U86656 ( n66206, n635, n787 );
nor U86657 ( n66209, n786, n66210 );
nand U86658 ( n66210, n40784, n66206 );
nand U86659 ( n40113, n2160, n1919 );
nand U86660 ( n40114, n2159, n1913 );
nor U86661 ( n39047, n39049, n39050 );
nor U86662 ( n39049, n1885, n38872 );
nor U86663 ( n39050, n37513, n39020 );
nand U86664 ( n38204, n39040, n39041 );
nand U86665 ( n39041, n2074, n36551 );
nor U86666 ( n39040, n39042, n39043 );
nor U86667 ( n39042, n39057, n37342 );
nand U86668 ( n38639, n39024, n39025 );
nor U86669 ( n39025, n39026, n39027 );
nor U86670 ( n39024, n39039, n38204 );
nor U86671 ( n39026, n2188, n38604 );
nor U86672 ( n39052, n39053, n39054 );
nor U86673 ( n39053, n38866, n39020 );
nor U86674 ( n39054, n38865, n39020 );
buf U86675 ( n76793, n76790 );
nand U86676 ( n38201, n38202, n38203 );
nand U86677 ( n38203, n76815, n2128 );
nand U86678 ( n38202, n76812, n38204 );
nand U86679 ( n2791, n38189, n38190 );
nor U86680 ( n38190, n38191, n38192 );
nor U86681 ( n38189, n38200, n38201 );
nand U86682 ( n38192, n38193, n38194 );
buf U86683 ( n76241, n76240 );
not U86684 ( n2385, n18792 );
nor U86685 ( n40107, n2160, n1919 );
nand U86686 ( n38990, n38949, n39071 );
nand U86687 ( n39071, n39072, n38904 );
nand U86688 ( n66753, n623, n785 );
nor U86689 ( n39051, n39055, n39056 );
nor U86690 ( n39055, n1875, n2039 );
nor U86691 ( n39056, n1885, n38875 );
nand U86692 ( n39235, n37457, n39243 );
nor U86693 ( n39232, n39194, n38865 );
nand U86694 ( n38236, n39154, n39155 );
nor U86695 ( n39154, n39187, n39188 );
nor U86696 ( n39155, n39156, n39157 );
nor U86697 ( n39187, n2183, n38822 );
nand U86698 ( n38645, n39140, n39141 );
nor U86699 ( n39141, n39142, n39143 );
nor U86700 ( n39140, n39153, n38236 );
nor U86701 ( n39142, n2185, n38604 );
nand U86702 ( n39166, n39167, n39168 );
nor U86703 ( n39167, n39174, n39175 );
nor U86704 ( n39168, n39169, n39170 );
nor U86705 ( n39174, n38875, n39134 );
nand U86706 ( n36688, n36689, n36690 );
nand U86707 ( n36689, n76822, n36702 );
nand U86708 ( n36690, n76831, n36691 );
nand U86709 ( n36691, n36692, n36693 );
nand U86710 ( n41472, n54989, n842 );
nor U86711 ( n54989, n838, n845 );
nand U86712 ( n36693, n36694, n1843 );
xor U86713 ( n36694, n36695, n36696 );
nor U86714 ( n39231, n39194, n38866 );
nor U86715 ( n39233, n39194, n37513 );
nand U86716 ( n38232, n38233, n38234 );
nand U86717 ( n38234, n38235, n76818 );
nand U86718 ( n38233, n76811, n38236 );
nand U86719 ( n2781, n38221, n38222 );
nor U86720 ( n38222, n38223, n38224 );
nor U86721 ( n38221, n38231, n38232 );
nand U86722 ( n38224, n38225, n38226 );
xor U86723 ( n72502, n72519, n72698 );
xor U86724 ( n72698, n72517, n72518 );
nor U86725 ( n72537, n1205, n1228 );
nand U86726 ( n71345, n71656, n71657 );
nand U86727 ( n71656, n71661, n71660 );
nand U86728 ( n71657, n71658, n71659 );
or U86729 ( n71659, n71660, n71661 );
nand U86730 ( n71076, n71052, n71077 );
nand U86731 ( n71077, n71053, n71055 );
nand U86732 ( n71056, n71335, n71336 );
or U86733 ( n71335, n71340, n71339 );
nand U86734 ( n71336, n71337, n71338 );
nand U86735 ( n71338, n71339, n71340 );
nor U86736 ( n66208, n635, n787 );
xnor U86737 ( n71057, n71341, n71091 );
xor U86738 ( n71341, n71086, n71090 );
nor U86739 ( n71648, n72189, n1059 );
nand U86740 ( n71351, n71492, n71493 );
or U86741 ( n71492, n71497, n71496 );
nand U86742 ( n71493, n71494, n71495 );
nand U86743 ( n71494, n71496, n71497 );
nor U86744 ( n71363, n1044, n71311 );
xor U86745 ( n71344, n71497, n71527 );
xor U86746 ( n71527, n71495, n71496 );
or U86747 ( n41264, n76847, n42281 );
nand U86748 ( n40830, n42288, n40665 );
nand U86749 ( n42288, n829, n842 );
buf U86750 ( n76254, n76251 );
not U86751 ( n1227, n71429 );
nand U86752 ( n72540, n72764, n71265 );
nor U86753 ( n72764, n1228, n1227 );
nor U86754 ( n71114, n1033, n71325 );
nand U86755 ( n71078, n71080, n71081 );
nand U86756 ( n71080, n71087, n71088 );
nand U86757 ( n71081, n1019, n71082 );
nand U86758 ( n71088, n71085, n71089 );
not U86759 ( n1019, n71087 );
not U86760 ( n1228, n71303 );
nand U86761 ( n66207, n628, n786 );
nor U86762 ( n71347, n1030, n71325 );
nand U86763 ( n67226, n845, n842 );
nand U86764 ( n71276, n1209, n71278 );
nand U86765 ( n72775, n71276, n72782 );
nand U86766 ( n72782, n1225, n76043 );
and U86767 ( n72539, n72771, n72772 );
nand U86768 ( n72772, n72773, n71244 );
nand U86769 ( n72771, n72775, n71429 );
nand U86770 ( n72773, n71272, n72774 );
nand U86771 ( n42092, n789, n41198 );
not U86772 ( n2155, n37288 );
buf U86773 ( n76414, n76413 );
nand U86774 ( MUL_1411_U438, n71049, n71050 );
nand U86775 ( n71049, n71054, n71055 );
nand U86776 ( n71050, n1022, n71051 );
xor U86777 ( n71054, n71056, n71057 );
xnor U86778 ( n71807, n71931, n71932 );
xnor U86779 ( n71932, n71933, n71934 );
xor U86780 ( n36395, n36396, n36397 );
nand U86781 ( n36390, n36391, n36392 );
nand U86782 ( n36391, n76821, n36398 );
nand U86783 ( n36392, n76831, n36393 );
xnor U86784 ( n36393, n36394, n36395 );
nor U86785 ( n72720, n1205, n1229 );
not U86786 ( n1229, n71413 );
nand U86787 ( n38975, n38949, n39073 );
nand U86788 ( n39073, n38905, n38904 );
nand U86789 ( n72719, n72744, n71265 );
nor U86790 ( n72744, n1229, n1228 );
not U86791 ( n1225, n71244 );
or U86792 ( n71272, n76044, n1209 );
nor U86793 ( n39064, n39069, n39070 );
nor U86794 ( n39069, n2039, n38975 );
nor U86795 ( n39070, n38875, n38990 );
xor U86796 ( n71577, n71625, n72520 );
xor U86797 ( n72520, n71623, n71624 );
nor U86798 ( n71616, n1205, n1227 );
nand U86799 ( n72190, n72189, n71647 );
buf U86800 ( n76403, n76402 );
nand U86801 ( n38980, n38981, n38982 );
nand U86802 ( n38981, n38986, n38984 );
nand U86803 ( n38982, n38983, n38984 );
nor U86804 ( n38986, n38875, n38985 );
and U86805 ( n39194, n37457, n39243 );
xnor U86806 ( n40798, n40799, n40800 );
nand U86807 ( n40793, n40794, n40795 );
nand U86808 ( n40794, n584, n40801 );
nand U86809 ( n40795, n76851, n40796 );
xnor U86810 ( n40796, n40797, n40798 );
nor U86811 ( n62347, n61617, n62275 );
nand U86812 ( n62343, n62344, n62345 );
nor U86813 ( n62344, n62348, n62349 );
nor U86814 ( n62345, n62346, n62347 );
nor U86815 ( n62348, n41487, n62275 );
nor U86816 ( n38763, n38130, n38764 );
nand U86817 ( n38770, n38835, n38836 );
nand U86818 ( n38836, n38837, n38838 );
nand U86819 ( n38837, n38900, n38901 );
nand U86820 ( n38901, n38902, n38903 );
and U86821 ( n38902, n38904, n38905 );
nand U86822 ( n38769, n38770, n38771 );
nand U86823 ( n71531, n71943, n71944 );
nand U86824 ( n71943, n71931, n71933 );
nand U86825 ( n71944, n71934, n71945 );
or U86826 ( n71945, n71933, n71931 );
nand U86827 ( n72742, n71276, n72743 );
nand U86828 ( n72743, n1227, n76044 );
and U86829 ( n72717, n72738, n72739 );
nand U86830 ( n72739, n72740, n71429 );
nand U86831 ( n72738, n72742, n71303 );
nand U86832 ( n72740, n71272, n72741 );
xnor U86833 ( n71045, n71813, n71660 );
xnor U86834 ( n71813, n71661, n71658 );
xnor U86835 ( n71360, n71490, n71540 );
xnor U86836 ( n71540, n71488, n71491 );
nand U86837 ( n71619, n72542, n71265 );
nor U86838 ( n72542, n1227, n1225 );
not U86839 ( n2095, n40524 );
nor U86840 ( n39102, n39105, n39106 );
nor U86841 ( n39106, n1903, n37513 );
nor U86842 ( n39105, n1884, n38872 );
nand U86843 ( n38220, n39095, n39096 );
nand U86844 ( n39096, n2074, n36633 );
nor U86845 ( n39095, n39097, n39098 );
nor U86846 ( n39097, n39113, n37341 );
nand U86847 ( n38642, n39076, n39077 );
nor U86848 ( n39077, n39078, n39079 );
nor U86849 ( n39076, n39094, n38220 );
nand U86850 ( n39079, n39080, n39081 );
nor U86851 ( n39107, n39111, n39112 );
nor U86852 ( n39111, n1874, n2039 );
nor U86853 ( n39112, n1884, n38875 );
nand U86854 ( n72547, n71276, n72548 );
nand U86855 ( n72548, n1233, n76043 );
and U86856 ( n71618, n72543, n72544 );
nand U86857 ( n72544, n72545, n71246 );
nand U86858 ( n72543, n72547, n71244 );
nand U86859 ( n72545, n71272, n72546 );
nor U86860 ( n45434, n76314, n76835 );
buf U86861 ( n76246, n61295 );
nand U86862 ( n36423, n37771, n36265 );
nand U86863 ( n37771, n37106, n37103 );
nand U86864 ( n42087, n788, n40984 );
nand U86865 ( n38217, n38218, n38219 );
nand U86866 ( n38219, n76815, n2122 );
nand U86867 ( n38218, n76812, n38220 );
nand U86868 ( n2786, n38205, n38206 );
nor U86869 ( n38206, n38207, n38208 );
nor U86870 ( n38205, n38216, n38217 );
nand U86871 ( n38207, n38213, n38214 );
xor U86872 ( n11739, n11740, n11742 );
or U86873 ( n71085, n71091, n71090 );
nor U86874 ( n39108, n39109, n39110 );
nor U86875 ( n39109, n1903, n38866 );
nor U86876 ( n39110, n1903, n38865 );
nor U86877 ( n62654, n62586, n61617 );
nand U86878 ( n47420, n62548, n62549 );
nor U86879 ( n62548, n62579, n62580 );
nor U86880 ( n62549, n62550, n62551 );
nor U86881 ( n62579, n745, n61441 );
and U86882 ( n72670, n72710, n72711 );
nand U86883 ( n72710, n72714, n71413 );
nand U86884 ( n72711, n72712, n71303 );
nand U86885 ( n72714, n71276, n72715 );
nor U86886 ( n40103, n1925, n2162 );
nand U86887 ( n71083, n71090, n71091 );
nor U86888 ( n62655, n62586, n41487 );
nand U86889 ( n72715, n1228, n71278 );
nor U86890 ( n71322, n1048, n71311 );
nand U86891 ( n71320, n71486, n71487 );
or U86892 ( n71486, n71491, n71490 );
nand U86893 ( n71487, n71488, n71489 );
nand U86894 ( n71489, n71490, n71491 );
not U86895 ( n1233, n71246 );
nand U86896 ( n37762, n76827, n37288 );
nor U86897 ( n16639, n76586, n76789 );
buf U86898 ( n76420, n76417 );
not U86899 ( n2157, n37023 );
nand U86900 ( n72503, n72655, n72656 );
or U86901 ( n72655, n72612, n72615 );
nand U86902 ( n72656, n72657, n72614 );
nand U86903 ( n72657, n72615, n72612 );
or U86904 ( n40685, n41195, n41196 );
not U86905 ( n1230, n71574 );
nand U86906 ( n72672, n72716, n71265 );
nor U86907 ( n72716, n1230, n1229 );
buf U86908 ( n76840, n76836 );
nor U86909 ( n62373, n62375, n62376 );
nor U86910 ( n62375, n542, n61624 );
nor U86911 ( n62376, n41487, n62351 );
nand U86912 ( n46555, n62366, n62367 );
nand U86913 ( n62367, n813, n40747 );
nor U86914 ( n62366, n62368, n62369 );
nor U86915 ( n62368, n62383, n41936 );
nand U86916 ( n71047, n71671, n71672 );
or U86917 ( n71671, n71026, n71027 );
nand U86918 ( n71672, n71028, n71673 );
nand U86919 ( n71673, n71027, n71026 );
not U86920 ( n1234, n71312 );
nand U86921 ( n72163, n72230, n72231 );
or U86922 ( n72230, n72149, n72152 );
nand U86923 ( n72231, n72151, n72232 );
nand U86924 ( n72232, n72152, n72149 );
nor U86925 ( n71923, n71924, n1089 );
nor U86926 ( n71688, n71689, n1067 );
nor U86927 ( n71919, n71920, n71921 );
nor U86928 ( n71920, n71922, n71923 );
and U86929 ( n71922, n71924, n1089 );
nand U86930 ( n72245, n72337, n72338 );
nand U86931 ( n72337, n72341, n71312 );
nand U86932 ( n72338, n72339, n71308 );
nand U86933 ( n72341, n71276, n72342 );
nand U86934 ( n71811, n71816, n71817 );
or U86935 ( n71816, n71798, n71799 );
nand U86936 ( n71817, n71800, n71818 );
nand U86937 ( n71818, n71799, n71798 );
nor U86938 ( n41567, n40690, n790 );
nor U86939 ( n39116, n39118, n39119 );
nor U86940 ( n39119, n37513, n39104 );
nor U86941 ( n39118, n38872, n39072 );
nor U86942 ( n62378, n62379, n62380 );
nor U86943 ( n62379, n61618, n62351 );
nor U86944 ( n62380, n61617, n62351 );
nand U86945 ( n66201, n639, n788 );
nor U86946 ( n39120, n39130, n39131 );
nor U86947 ( n39130, n2039, n38905 );
nor U86948 ( n39131, n38875, n39072 );
nand U86949 ( n1566, n46543, n46544 );
nor U86950 ( n46544, n46545, n46546 );
nor U86951 ( n46543, n46552, n46553 );
nand U86952 ( n46546, n46547, n46548 );
not U86953 ( n2064, n37304 );
buf U86954 ( n76841, n76836 );
not U86955 ( n1223, n71308 );
nand U86956 ( n72342, n1223, n71278 );
nor U86957 ( n39160, n39162, n38866 );
nand U86958 ( n39157, n39158, n39159 );
nand U86959 ( n39158, n39163, n39161 );
nand U86960 ( n39159, n39160, n39161 );
nor U86961 ( n39163, n39162, n38865 );
nor U86962 ( n39191, n39162, n37513 );
xor U86963 ( n72469, n72593, n72594 );
xor U86964 ( n72594, n72595, n72596 );
nand U86965 ( n37263, n1933, n36462 );
nand U86966 ( n38829, n38830, n38831 );
nand U86967 ( n38831, n38150, n76797 );
nand U86968 ( n38830, n2033, n38151 );
nor U86969 ( n72673, n1205, n1230 );
nand U86970 ( n71578, n72514, n72515 );
or U86971 ( n72514, n72519, n72518 );
nand U86972 ( n72515, n72516, n72517 );
nand U86973 ( n72516, n72518, n72519 );
nand U86974 ( n38252, n39219, n39220 );
nor U86975 ( n39219, n39236, n39237 );
nor U86976 ( n39220, n39221, n39222 );
nor U86977 ( n39237, n2182, n38822 );
nand U86978 ( n38648, n39201, n39202 );
nor U86979 ( n39202, n39203, n39204 );
nor U86980 ( n39201, n39218, n38252 );
nor U86981 ( n39203, n2184, n38604 );
nand U86982 ( n38973, n38997, n38998 );
nor U86983 ( n38997, n2130, n2127 );
nand U86984 ( n38998, n38975, n38994 );
nand U86985 ( n40325, n2042, n2069 );
buf U86986 ( n76412, n38757 );
nand U86987 ( n40683, n41196, n41195 );
nor U86988 ( n39241, n39244, n39245 );
and U86989 ( n39244, n39183, n2005 );
nor U86990 ( n39245, n37513, n39235 );
nand U86991 ( n38249, n38250, n38251 );
nand U86992 ( n38251, n76815, n2113 );
nand U86993 ( n38250, n76812, n38252 );
nand U86994 ( n2776, n38237, n38238 );
nor U86995 ( n38238, n38239, n38240 );
nor U86996 ( n38237, n38248, n38249 );
nand U86997 ( n38240, n38241, n38242 );
nor U86998 ( n72090, n72093, n1084 );
xnor U86999 ( n36794, n36795, n36796 );
nand U87000 ( n36789, n36790, n36791 );
nand U87001 ( n36790, n76822, n36797 );
nand U87002 ( n36791, n76830, n36792 );
xnor U87003 ( n36792, n36793, n36794 );
nand U87004 ( n3106, n36786, n36787 );
nor U87005 ( n36786, n36798, n36799 );
nor U87006 ( n36787, n36788, n36789 );
nand U87007 ( n36799, n36800, n36801 );
or U87008 ( n36281, n36814, n36815 );
nand U87009 ( n72607, n72616, n72617 );
or U87010 ( n72616, n72593, n72596 );
nand U87011 ( n72617, n72618, n72595 );
nand U87012 ( n72618, n72596, n72593 );
nor U87013 ( n39247, n39248, n39249 );
nor U87014 ( n39248, n38866, n39235 );
nor U87015 ( n39249, n38865, n39235 );
or U87016 ( n40684, n40688, n40689 );
nand U87017 ( n37103, n38603, n2069 );
nor U87018 ( n38603, n2072, n2042 );
nor U87019 ( n72248, n1235, n1205 );
not U87020 ( n2159, n36649 );
nor U87021 ( n39123, n39104, n38865 );
nor U87022 ( n39122, n39104, n38866 );
not U87023 ( n1235, n71371 );
not U87024 ( n1224, n72453 );
xor U87025 ( n71974, n72165, n72166 );
xor U87026 ( n72166, n72167, n72168 );
nand U87027 ( n72226, n72328, n72329 );
or U87028 ( n72328, n72261, n72264 );
nand U87029 ( n72329, n72263, n72330 );
nand U87030 ( n72330, n72264, n72261 );
nand U87031 ( n72343, n72448, n72449 );
nand U87032 ( n72448, n72452, n72453 );
nand U87033 ( n72449, n72450, n71308 );
nand U87034 ( n72452, n71272, n72454 );
nand U87035 ( n72450, n71276, n72451 );
nand U87036 ( n72451, n1224, n76044 );
nor U87037 ( n45443, n76310, n76835 );
nand U87038 ( n72633, n72669, n71265 );
nor U87039 ( n72669, n1232, n1230 );
not U87040 ( n1232, n72499 );
nand U87041 ( n41170, n41171, n41172 );
nand U87042 ( n41171, n584, n41178 );
nand U87043 ( n41172, n76850, n41173 );
xnor U87044 ( n41173, n41174, n41175 );
xnor U87045 ( n41175, n41176, n41177 );
nand U87046 ( n1881, n41167, n41168 );
nor U87047 ( n41167, n41179, n41180 );
nor U87048 ( n41168, n41169, n41170 );
nand U87049 ( n41180, n41181, n41182 );
nor U87050 ( n72634, n1232, n1205 );
not U87051 ( n623, n41377 );
not U87052 ( n1479, n52372 );
and U87053 ( n72631, n72663, n72664 );
nand U87054 ( n72663, n72667, n71574 );
nand U87055 ( n72664, n72665, n71413 );
nand U87056 ( n72667, n71276, n72668 );
nor U87057 ( n71789, n71790, n1092 );
nor U87058 ( n71907, n1119, n71910 );
nor U87059 ( n71783, n71790, n1090 );
nor U87060 ( n72107, n72108, n1115 );
nand U87061 ( n72110, n72213, n72214 );
or U87062 ( n72213, n72165, n72167 );
nand U87063 ( n72214, n72168, n72215 );
nand U87064 ( n72215, n72167, n72165 );
nor U87065 ( n72103, n72104, n72105 );
nor U87066 ( n72104, n72106, n72107 );
and U87067 ( n72106, n72108, n1115 );
xor U87068 ( n72603, n72612, n72613 );
xor U87069 ( n72613, n72614, n72615 );
and U87070 ( n72247, n72336, n71265 );
nor U87071 ( n72336, n1235, n1234 );
not U87072 ( n2158, n36381 );
nand U87073 ( n72668, n1229, n76043 );
nand U87074 ( n71109, n71115, n71116 );
nand U87075 ( n71115, n71122, n71123 );
nand U87076 ( n71116, n1024, n71117 );
nand U87077 ( n71123, n71120, n71124 );
not U87078 ( n1390, n52533 );
not U87079 ( n1423, n52673 );
nand U87080 ( n36279, n36815, n36814 );
nor U87081 ( n71917, n71924, n1088 );
buf U87082 ( n76795, n76790 );
nor U87083 ( n71682, n71689, n1065 );
nor U87084 ( n72145, n72146, n1195 );
nand U87085 ( n72133, n72239, n72240 );
nand U87086 ( n72239, n72243, n71371 );
nand U87087 ( n72240, n72241, n71312 );
nand U87088 ( n72243, n71276, n72244 );
nor U87089 ( n72141, n72142, n72143 );
nor U87090 ( n72142, n72144, n72145 );
and U87091 ( n72144, n72146, n1195 );
nand U87092 ( n72036, n72118, n72119 );
or U87093 ( n72118, n71991, n71994 );
nand U87094 ( n72119, n71993, n72120 );
nand U87095 ( n72120, n71994, n71991 );
xnor U87096 ( MUL_1411_U10, n71520, n71340 );
xnor U87097 ( n71520, n71337, n71339 );
nor U87098 ( n72346, n1234, n1205 );
nand U87099 ( n72244, n1234, n76043 );
nand U87100 ( n72628, n71276, n72629 );
nand U87101 ( n72629, n1230, n76044 );
and U87102 ( n72577, n72624, n72625 );
nand U87103 ( n72625, n72626, n71574 );
nand U87104 ( n72624, n72628, n72499 );
nand U87105 ( n72626, n71272, n72627 );
nand U87106 ( n71153, n71155, n71307 );
nor U87107 ( n72139, n72146, n1194 );
nand U87108 ( n40681, n40689, n40688 );
nand U87109 ( n38893, n38894, n38895 );
nand U87110 ( n38895, n38166, n76797 );
nand U87111 ( n38894, n2033, n38167 );
nand U87112 ( n37579, n1937, n36667 );
nor U87113 ( n16674, n76579, n76789 );
nand U87114 ( n38142, n38148, n38149 );
nand U87115 ( n38149, n38150, n76818 );
nand U87116 ( n38148, n38151, n76442 );
nand U87117 ( n71905, n71986, n71987 );
or U87118 ( n71986, n71895, n71898 );
nand U87119 ( n71987, n71897, n71988 );
nand U87120 ( n71988, n71898, n71895 );
nor U87121 ( n62442, n41487, n62395 );
nand U87122 ( n37585, n37445, n37422 );
nand U87123 ( n46942, n62432, n62433 );
nand U87124 ( n62433, n813, n41134 );
nor U87125 ( n62432, n62434, n62435 );
nor U87126 ( n62434, n62449, n41920 );
nand U87127 ( n71043, n71677, n71678 );
or U87128 ( n71677, n71031, n71030 );
nand U87129 ( n71678, n71032, n71679 );
nand U87130 ( n71679, n71030, n71031 );
nor U87131 ( n71684, n71685, n71686 );
nor U87132 ( n71685, n71687, n71688 );
and U87133 ( n71687, n71689, n1067 );
or U87134 ( n36280, n36284, n36285 );
not U87135 ( n1024, n71122 );
nor U87136 ( n38961, n38179, n38764 );
and U87137 ( n71389, n71388, n71396 );
nand U87138 ( n71925, n71924, n71926 );
nor U87139 ( n62444, n62445, n62446 );
nor U87140 ( n62445, n61618, n62395 );
nor U87141 ( n62446, n61617, n62395 );
nand U87142 ( n41569, n792, n40864 );
nand U87143 ( n62551, n62552, n62553 );
nand U87144 ( n62552, n62557, n62555 );
nand U87145 ( n62553, n62554, n62555 );
nor U87146 ( n62557, n62556, n61617 );
nor U87147 ( n72101, n72108, n1114 );
nor U87148 ( n62583, n62556, n41487 );
xor U87149 ( n72032, n72149, n72150 );
xor U87150 ( n72150, n72151, n72152 );
nand U87151 ( n39027, n39028, n39029 );
nand U87152 ( n39029, n38198, n76797 );
nand U87153 ( n39028, n2033, n38199 );
and U87154 ( n72345, n72447, n71265 );
nor U87155 ( n72447, n1234, n1223 );
nand U87156 ( n37442, n1940, n36355 );
nand U87157 ( n72579, n72630, n71265 );
nor U87158 ( n72630, n1224, n1232 );
nand U87159 ( n47964, n62641, n62642 );
nor U87160 ( n62641, n62658, n62659 );
nor U87161 ( n62642, n62643, n62644 );
nor U87162 ( n62659, n743, n61441 );
nand U87163 ( n72465, n72562, n72563 );
or U87164 ( n72562, n72423, n72426 );
nand U87165 ( n72563, n72564, n72425 );
nand U87166 ( n72564, n72426, n72423 );
nor U87167 ( n66020, n650, n790 );
xor U87168 ( n72320, n72423, n72424 );
xor U87169 ( n72424, n72425, n72426 );
nand U87170 ( n72733, n71245, n71413 );
nand U87171 ( n1551, n47952, n47953 );
nor U87172 ( n47953, n47954, n47955 );
nor U87173 ( n47952, n47961, n47962 );
nand U87174 ( n47955, n47956, n47957 );
not U87175 ( n1352, n52221 );
xor U87176 ( n72159, n72261, n72262 );
xor U87177 ( n72262, n72263, n72264 );
nand U87178 ( n42077, n795, n41145 );
nor U87179 ( n39309, n39311, n39312 );
nor U87180 ( n39311, n38865, n39127 );
nor U87181 ( n39312, n37513, n39127 );
nand U87182 ( n38651, n39263, n39264 );
nor U87183 ( n39264, n39265, n39266 );
nor U87184 ( n39263, n39276, n38268 );
nor U87185 ( n39265, n2183, n38604 );
nor U87186 ( n62663, n62666, n62667 );
and U87187 ( n62666, n62577, n822 );
nor U87188 ( n62667, n41487, n62657 );
nand U87189 ( n38176, n38177, n38178 );
nand U87190 ( n38177, n76815, n2133 );
nand U87191 ( n38178, n1877, n76442 );
not U87192 ( n1877, n38179 );
nor U87193 ( n39246, n39250, n39251 );
nor U87194 ( n39250, n1872, n2039 );
nor U87195 ( n39251, n1883, n38875 );
nand U87196 ( n42082, n794, n40760 );
nand U87197 ( n72092, n72093, n72088 );
not U87198 ( n1948, n37422 );
nand U87199 ( n38264, n38265, n38266 );
nand U87200 ( n38266, n38267, n76818 );
nand U87201 ( n38265, n76812, n38268 );
nand U87202 ( n2771, n38253, n38254 );
nor U87203 ( n38254, n38255, n38256 );
nor U87204 ( n38253, n38263, n38264 );
nand U87205 ( n38256, n38257, n38258 );
nor U87206 ( n62669, n62670, n62671 );
nor U87207 ( n62670, n61618, n62657 );
nor U87208 ( n62671, n61617, n62657 );
xnor U87209 ( n71041, n71797, n71798 );
xnor U87210 ( n71797, n71799, n71800 );
nand U87211 ( n72324, n72427, n72428 );
or U87212 ( n72427, n72360, n72362 );
nand U87213 ( n72428, n72361, n72429 );
nand U87214 ( n72429, n72362, n72360 );
nand U87215 ( n72455, n72571, n72572 );
nand U87216 ( n72571, n72575, n72453 );
nand U87217 ( n72572, n72573, n72499 );
nand U87218 ( n72575, n71276, n72576 );
nor U87219 ( n72136, n1237, n1205 );
nand U87220 ( n36600, n36601, n36602 );
nand U87221 ( n36601, n76822, n36613 );
nand U87222 ( n36602, n36603, n76830 );
nor U87223 ( n36603, n36604, n36605 );
nand U87224 ( n3156, n36597, n36598 );
nor U87225 ( n36597, n36614, n36615 );
nor U87226 ( n36598, n36599, n36600 );
nand U87227 ( n36615, n36616, n36617 );
nand U87228 ( n72576, n1232, n71278 );
not U87229 ( n1637, n49804 );
nand U87230 ( n71909, n71910, n71905 );
not U87231 ( n628, n40784 );
nand U87232 ( n62684, n62779, n62780 );
nand U87233 ( n62780, n62781, n62782 );
nand U87234 ( n62782, n76386, n41297 );
nand U87235 ( n62683, n62684, n62685 );
or U87236 ( n62685, n62686, n62687 );
not U87237 ( n76386, n76387 );
and U87238 ( n72457, n72570, n71265 );
nor U87239 ( n72570, n1223, n1224 );
xnor U87240 ( n72222, n72359, n72360 );
xnor U87241 ( n72359, n72361, n72362 );
xor U87242 ( n11712, n11713, n11714 );
nand U87243 ( n72685, n71574, n71245 );
nand U87244 ( n71404, n71402, n71410 );
nand U87245 ( n36277, n36285, n36284 );
nand U87246 ( n41550, n64814, n42058 );
nand U87247 ( n40993, n40994, n40995 );
nand U87248 ( n40994, n584, n41006 );
nand U87249 ( n40995, n40996, n76850 );
nor U87250 ( n40996, n40997, n40998 );
nand U87251 ( n1931, n40990, n40991 );
nor U87252 ( n40990, n41007, n41008 );
nor U87253 ( n40991, n40992, n40993 );
nand U87254 ( n41008, n41009, n41010 );
not U87255 ( n2162, n36817 );
nor U87256 ( n71419, n1148, n71247 );
nand U87257 ( n71417, n71620, n71621 );
or U87258 ( n71620, n71625, n71624 );
nand U87259 ( n71621, n71622, n71623 );
nand U87260 ( n71622, n71624, n71625 );
and U87261 ( n72135, n72238, n71265 );
nor U87262 ( n72238, n1235, n1237 );
nand U87263 ( n62760, n62687, n62975 );
nand U87264 ( n62975, n62677, n62680 );
nand U87265 ( n48079, n62742, n62743 );
nor U87266 ( n62742, n62764, n62765 );
nor U87267 ( n62743, n62744, n62745 );
nor U87268 ( n62765, n737, n61441 );
nor U87269 ( n72580, n1224, n1205 );
not U87270 ( n1312, n52164 );
nand U87271 ( n37466, n1947, n36762 );
and U87272 ( n37577, n37466, n39845 );
nand U87273 ( n39845, n1953, n36532 );
nor U87274 ( n72458, n1205, n1223 );
nand U87275 ( n71176, n71178, n71396 );
nand U87276 ( n38159, n38164, n38165 );
nand U87277 ( n38165, n38166, n76818 );
nand U87278 ( n38164, n38167, n76442 );
nand U87279 ( n72533, n71245, n71303 );
nand U87280 ( n41560, n793, n41054 );
nand U87281 ( n72109, n72108, n72110 );
nand U87282 ( n72009, n72123, n72124 );
nand U87283 ( n72123, n72025, n72022 );
nand U87284 ( n72124, n72024, n72125 );
or U87285 ( n72125, n72022, n72025 );
xor U87286 ( n71136, n71145, n71146 );
xor U87287 ( n71145, n71309, n71310 );
xor U87288 ( n71146, n71147, n71148 );
nand U87289 ( n71309, n71312, n71313 );
xor U87290 ( n71134, n71135, n71136 );
nand U87291 ( n72132, n1235, n76044 );
nand U87292 ( n39891, n2168, n1947 );
nand U87293 ( n39890, n39896, n39897 );
nand U87294 ( n39897, n39898, n1938 );
not U87295 ( n1938, n39899 );
xor U87296 ( n71771, n71895, n71896 );
xor U87297 ( n71896, n71897, n71898 );
nor U87298 ( n71767, n71774, n1120 );
nor U87299 ( n71785, n71786, n71787 );
nor U87300 ( n71786, n71788, n71789 );
and U87301 ( n71788, n71790, n1092 );
xnor U87302 ( n71142, n71136, n71135 );
not U87303 ( n604, n40665 );
nand U87304 ( n72147, n72146, n72148 );
nand U87305 ( n38191, n38196, n38197 );
nand U87306 ( n38197, n38198, n76818 );
nand U87307 ( n38196, n38199, n76442 );
buf U87308 ( n76405, n76402 );
nand U87309 ( n41665, n41672, n41673 );
nor U87310 ( n41672, n41786, n41787 );
nor U87311 ( n41673, n41674, n41675 );
nor U87312 ( n41787, n41788, n41789 );
nand U87313 ( n41628, n41636, n41637 );
nand U87314 ( n41636, n41830, n41831 );
nand U87315 ( n41637, n41638, n41639 );
nor U87316 ( n41638, n41828, n41829 );
nor U87317 ( n41666, n41665, n41664 );
nor U87318 ( n41686, n41692, n41693 );
nor U87319 ( n41693, n41694, n41695 );
nor U87320 ( n41692, n41698, n41699 );
nand U87321 ( n41695, n41696, n41697 );
nor U87322 ( n41720, n41722, n41723 );
nor U87323 ( n41722, n41736, n41737 );
nand U87324 ( n41723, n41724, n41725 );
nand U87325 ( n41724, n41734, n41735 );
nand U87326 ( n41698, n41714, n41715 );
nand U87327 ( n41714, n41772, n41773 );
nand U87328 ( n41715, n41716, n41717 );
nor U87329 ( n41716, n41770, n41771 );
nand U87330 ( n41606, n41607, n41608 );
nand U87331 ( n41607, n41862, n41863 );
nand U87332 ( n41608, n41609, n41610 );
nor U87333 ( n41609, n41854, n41855 );
nor U87334 ( n41639, n41640, n41641 );
nor U87335 ( n41640, n41811, n41816 );
nand U87336 ( n41641, n41642, n41643 );
nand U87337 ( n41816, n715, n41810 );
nor U87338 ( n41656, n41662, n41663 );
and U87339 ( n41663, n41664, n41665 );
nor U87340 ( n41662, n41666, n41667 );
nand U87341 ( n41667, n41668, n41669 );
and U87342 ( n41648, n41652, n41653 );
nand U87343 ( n41653, n41654, n41655 );
nand U87344 ( n41652, n41656, n41657 );
or U87345 ( n41657, n41655, n41654 );
nand U87346 ( n41725, n41726, n41727 );
nand U87347 ( n41727, n41728, n41729 );
nand U87348 ( n41728, n41732, n41733 );
nand U87349 ( n41729, n41730, n41731 );
nand U87350 ( n41643, n41644, n41645 );
nor U87351 ( n41644, n41808, n41809 );
nor U87352 ( n41645, n41646, n41647 );
nor U87353 ( n41808, n710, n41810 );
nor U87354 ( n41646, n41650, n41651 );
nor U87355 ( n41650, n41806, n41807 );
and U87356 ( n41651, n41649, n41648 );
nor U87357 ( n41806, n76010, n700 );
nor U87358 ( n41726, n75768, n75769 );
nor U87359 ( n75768, n41735, n41734 );
nor U87360 ( n75769, n41733, n41732 );
nand U87361 ( n39943, n2167, n1940 );
xor U87362 ( n71856, n71991, n71992 );
xor U87363 ( n71992, n71993, n71994 );
nor U87364 ( n71773, n71774, n1122 );
nand U87365 ( n71776, n71843, n71844 );
or U87366 ( n71843, n71763, n71762 );
nand U87367 ( n71844, n71764, n71845 );
nand U87368 ( n71845, n71762, n71763 );
or U87369 ( n39314, n39127, n38866 );
not U87370 ( n2790, n16874 );
nand U87371 ( n71690, n71689, n71691 );
not U87372 ( n2088, n36265 );
not U87373 ( n635, n41036 );
nand U87374 ( n41738, n41758, n41759 );
or U87375 ( n41759, n41731, n41730 );
nor U87376 ( n41758, n41764, n41765 );
nor U87377 ( n41764, n552, n41767 );
nor U87378 ( n41765, n41766, n76378 );
and U87379 ( n41766, n41767, n624 );
nor U87380 ( n62769, n62771, n62772 );
nor U87381 ( n62771, n61617, n62462 );
nor U87382 ( n62772, n41487, n62462 );
not U87383 ( n1238, n71357 );
nor U87384 ( n72025, n1238, n1205 );
nand U87385 ( n71199, n71201, n71410 );
nand U87386 ( n41721, n41740, n41741 );
nand U87387 ( n41740, n41736, n41737 );
nand U87388 ( n41741, n41742, n41743 );
nand U87389 ( n39901, n2165, n1937 );
nand U87390 ( n3166, n36556, n36557 );
nor U87391 ( n36556, n36573, n36574 );
nor U87392 ( n36557, n36558, n36559 );
nand U87393 ( n36574, n36575, n36576 );
nand U87394 ( n36559, n36560, n36561 );
nand U87395 ( n36560, n76822, n36572 );
nand U87396 ( n36561, n76831, n36562 );
nand U87397 ( n36562, n36563, n36564 );
nand U87398 ( n36564, n36565, n1844 );
xor U87399 ( n36565, n36566, n36567 );
nor U87400 ( n41647, n41648, n41649 );
not U87401 ( n2160, n36589 );
xor U87402 ( n36952, n36883, n36884 );
nand U87403 ( n36948, n36949, n36950 );
nand U87404 ( n36949, n76823, n36961 );
nand U87405 ( n36950, n76831, n36951 );
xor U87406 ( n36951, n36885, n36952 );
nand U87407 ( n3091, n36945, n36946 );
nor U87408 ( n36945, n37081, n37082 );
nor U87409 ( n36946, n36947, n36948 );
nand U87410 ( n37082, n37083, n37084 );
xnor U87411 ( n71716, n71891, n71892 );
xnor U87412 ( n71892, n71893, n71894 );
nand U87413 ( n40954, n40955, n40956 );
nand U87414 ( n40955, n584, n40967 );
nand U87415 ( n40956, n76851, n40957 );
nand U87416 ( n40957, n40958, n40959 );
nand U87417 ( n1941, n40951, n40952 );
nor U87418 ( n40951, n40968, n40969 );
nor U87419 ( n40952, n40953, n40954 );
nand U87420 ( n40969, n40970, n40971 );
nand U87421 ( n40959, n40960, n518 );
xor U87422 ( n40960, n40961, n40962 );
nand U87423 ( n37522, n37527, n37528 );
nor U87424 ( n37527, n2137, n37529 );
nor U87425 ( n37529, n37530, n37531 );
nand U87426 ( n37531, n37507, n37532 );
nand U87427 ( n37586, n37587, n37263 );
nand U87428 ( n37587, n37588, n37268 );
nand U87429 ( n37588, n1923, n37589 );
not U87430 ( n1923, n37403 );
nand U87431 ( n37559, n1993, n37560 );
nand U87432 ( n37560, n37561, n37453 );
nand U87433 ( n37561, n37562, n37492 );
nand U87434 ( n37562, n37563, n37564 );
nand U87435 ( n37524, n37525, n37526 );
nand U87436 ( n37525, n37597, n37598 );
or U87437 ( n37526, n37522, n2145 );
nor U87438 ( n37597, n2149, n37521 );
nand U87439 ( n37537, n37538, n37512 );
nor U87440 ( n37538, n2123, n37539 );
nor U87441 ( n37539, n2115, n37540 );
nand U87442 ( n37540, n37541, n37542 );
nand U87443 ( n37541, n37543, n37544 );
nor U87444 ( n37543, n37402, n2108 );
nand U87445 ( n37544, n37545, n37546 );
nand U87446 ( n37545, n37456, n37547 );
nand U87447 ( n37547, n37548, n37450 );
nor U87448 ( n37548, n37556, n2100 );
nor U87449 ( n37556, n37558, n37559 );
or U87450 ( n37558, n37496, n1985 );
and U87451 ( n72024, n72126, n71265 );
nor U87452 ( n72126, n1237, n1238 );
xor U87453 ( n71416, n71467, n71587 );
xor U87454 ( n71587, n71465, n71466 );
nand U87455 ( n64812, n797, n40930 );
nor U87456 ( n40140, n38508, n76405 );
xor U87457 ( n41320, n41270, n41271 );
nand U87458 ( n41316, n41317, n41318 );
nand U87459 ( n41317, n584, n41329 );
nand U87460 ( n41318, n76851, n41319 );
xor U87461 ( n41319, n41272, n41320 );
nand U87462 ( n1866, n41313, n41314 );
nor U87463 ( n41313, n41450, n41451 );
nor U87464 ( n41314, n41315, n41316 );
nand U87465 ( n41451, n41452, n41453 );
nand U87466 ( n45996, n45997, n45998 );
nand U87467 ( n45997, n76340, n40713 );
or U87468 ( n45998, n45999, n573 );
not U87469 ( n1422, n52800 );
nor U87470 ( n37309, n37308, n37513 );
nand U87471 ( n71720, n71860, n71861 );
nand U87472 ( n71860, n71760, n71758 );
nand U87473 ( n71861, n71759, n71862 );
or U87474 ( n71862, n71758, n71760 );
nor U87475 ( n71871, n71872, n1200 );
nand U87476 ( n71874, n72012, n72013 );
or U87477 ( n72012, n71889, n71887 );
nand U87478 ( n72013, n71890, n72014 );
nand U87479 ( n72014, n71887, n71889 );
nor U87480 ( n71867, n71868, n71869 );
nor U87481 ( n71868, n71870, n71871 );
and U87482 ( n71870, n71872, n1200 );
nand U87483 ( n38208, n38209, n38210 );
nand U87484 ( n38210, n76448, n2899 );
nand U87485 ( n38209, n38212, n76442 );
nor U87486 ( n65348, n667, n794 );
nand U87487 ( n71852, n71995, n71996 );
or U87488 ( n71995, n71894, n71891 );
nand U87489 ( n71996, n71893, n71997 );
nand U87490 ( n71997, n71891, n71894 );
nor U87491 ( n41245, n41246, n41247 );
nand U87492 ( n41247, n40797, n40800 );
xor U87493 ( n40905, n40826, n41294 );
nor U87494 ( n41294, n41295, n40824 );
nor U87495 ( n41295, n737, n40825 );
nand U87496 ( n72646, n72499, n71245 );
nand U87497 ( n39143, n39144, n39145 );
nand U87498 ( n39144, n38235, n76797 );
nand U87499 ( n39145, n2033, n38230 );
nand U87500 ( n72020, n1237, n71278 );
buf U87501 ( n76419, n76417 );
nor U87502 ( n71458, n1205, n1225 );
nand U87503 ( n48337, n62949, n62950 );
nand U87504 ( n62950, n813, n40801 );
nor U87505 ( n62949, n62951, n62952 );
nor U87506 ( n62952, n724, n62953 );
nor U87507 ( n65347, n795, n672 );
nor U87508 ( n65341, n65824, n65343 );
nand U87509 ( n1536, n48322, n48323 );
nor U87510 ( n48323, n48324, n48325 );
nor U87511 ( n48322, n48332, n48333 );
nand U87512 ( n48324, n48329, n48330 );
nand U87513 ( n39792, n2170, n1959 );
nand U87514 ( n39734, n39743, n39744 );
nand U87515 ( n39743, n39745, n39746 );
and U87516 ( n39745, n39748, n39749 );
nand U87517 ( n39746, n1954, n39737 );
nand U87518 ( n72258, n71371, n71245 );
nand U87519 ( n62681, n76386, n41090 );
nor U87520 ( n39402, n39405, n39406 );
nor U87521 ( n39405, n37513, n39378 );
nor U87522 ( n39406, n38956, n39378 );
nand U87523 ( n38300, n39395, n39396 );
nand U87524 ( n39396, n2074, n36398 );
nor U87525 ( n39395, n39397, n39398 );
nor U87526 ( n39397, n39411, n37338 );
nand U87527 ( n72592, n72453, n71245 );
nand U87528 ( n71791, n71790, n71792 );
buf U87529 ( n76839, n76836 );
xor U87530 ( n40907, n40826, n41291 );
nor U87531 ( n41291, n41292, n40824 );
nor U87532 ( n41292, n743, n40825 );
nor U87533 ( n39407, n39409, n39410 );
nor U87534 ( n39409, n38866, n39378 );
nor U87535 ( n39410, n38865, n39378 );
nand U87536 ( n38658, n39326, n39327 );
nor U87537 ( n39327, n39328, n39329 );
nor U87538 ( n39326, n39350, n38284 );
nand U87539 ( n39329, n39330, n39331 );
nand U87540 ( n2761, n38285, n38286 );
nor U87541 ( n38286, n38287, n38288 );
nor U87542 ( n38285, n38295, n38296 );
nand U87543 ( n38287, n38292, n38293 );
nand U87544 ( n47381, n47856, n7812 );
nand U87545 ( n44985, n47749, n47750 );
nor U87546 ( n47750, n47751, n47752 );
nor U87547 ( n47749, n47765, n47766 );
nand U87548 ( n47751, n47759, n47760 );
nand U87549 ( n48005, n7799, n7805 );
not U87550 ( n7797, n43287 );
nor U87551 ( n47856, n47849, n7797 );
nor U87552 ( n46296, n46299, n76330 );
nor U87553 ( n46299, n46301, n46302 );
nand U87554 ( n46301, n46322, n46323 );
nand U87555 ( n46302, n46303, n46304 );
not U87556 ( n7537, n46871 );
not U87557 ( n2163, n36286 );
nand U87558 ( n39744, n2172, n1967 );
nand U87559 ( n47391, n47863, n7812 );
buf U87560 ( n76243, n76240 );
nand U87561 ( n47386, n47856, n7807 );
nand U87562 ( n71435, n71433, n71245 );
nand U87563 ( n47396, n47863, n7807 );
nand U87564 ( n38281, n38282, n38283 );
nand U87565 ( n38283, n76815, n2102 );
nand U87566 ( n38282, n76812, n38284 );
nand U87567 ( n2766, n38269, n38270 );
nor U87568 ( n38270, n38271, n38272 );
nor U87569 ( n38269, n38280, n38281 );
nand U87570 ( n38271, n38277, n38278 );
nand U87571 ( n71606, n71276, n71607 );
nand U87572 ( n71607, n1240, n71278 );
and U87573 ( n71460, n71602, n71603 );
nand U87574 ( n71603, n71604, n71267 );
nand U87575 ( n71602, n71606, n71246 );
nand U87576 ( n71604, n71272, n71605 );
nand U87577 ( n71461, n71601, n71265 );
nor U87578 ( n71601, n1225, n1233 );
xor U87579 ( n71422, n71306, n71428 );
xor U87580 ( n71428, n71234, n71305 );
nand U87581 ( n71423, n71462, n71463 );
or U87582 ( n71462, n71467, n71466 );
nand U87583 ( n71463, n71464, n71465 );
nand U87584 ( n71464, n71466, n71467 );
nand U87585 ( n37574, n1959, n36730 );
nor U87586 ( n65346, n793, n660 );
xor U87587 ( n71164, n71169, n71170 );
nor U87588 ( n71170, n71171, n1224 );
xor U87589 ( n71169, n71172, n71173 );
nand U87590 ( n71172, n71180, n71181 );
nand U87591 ( n1541, n48196, n48197 );
nor U87592 ( n48197, n48198, n48199 );
nor U87593 ( n48196, n48205, n48206 );
nand U87594 ( n48199, n48200, n48201 );
nand U87595 ( n47359, n47839, n7812 );
not U87596 ( n7803, n47849 );
nor U87597 ( n47839, n7803, n43287 );
nand U87598 ( n71889, n72021, n71265 );
nor U87599 ( n72021, n1239, n1238 );
not U87600 ( n1173, n71245 );
nand U87601 ( n47364, n47839, n7807 );
not U87602 ( n1949, n39893 );
nand U87603 ( n37492, n1975, n36572 );
nor U87604 ( n39555, n37496, n1974 );
nand U87605 ( n39372, n39373, n39374 );
nand U87606 ( n39373, n2074, n36702 );
nand U87607 ( n39374, n2038, n39362 );
nand U87608 ( n68413, n68876, n6024 );
nand U87609 ( n65893, n68770, n68771 );
nor U87610 ( n68771, n68772, n68773 );
nor U87611 ( n68770, n68786, n68787 );
nand U87612 ( n68772, n68780, n68781 );
nand U87613 ( n69013, n6012, n6018 );
not U87614 ( n6009, n63972 );
nor U87615 ( n68876, n68869, n6009 );
nand U87616 ( n26412, n26877, n4247 );
nand U87617 ( n59551, n60017, n6879 );
nand U87618 ( n24311, n26771, n26772 );
nor U87619 ( n26772, n26773, n26774 );
nor U87620 ( n26771, n26787, n26788 );
nand U87621 ( n26773, n26781, n26782 );
nand U87622 ( n57434, n59911, n59912 );
nor U87623 ( n59912, n59913, n59914 );
nor U87624 ( n59911, n59927, n59928 );
nand U87625 ( n59913, n59921, n59922 );
nand U87626 ( n27016, n4234, n4240 );
nand U87627 ( n60157, n6867, n6873 );
not U87628 ( n4232, n22693 );
not U87629 ( n6864, n55809 );
nor U87630 ( n26877, n26870, n4232 );
nor U87631 ( n60017, n60010, n6864 );
not U87632 ( n5750, n67918 );
not U87633 ( n3993, n25915 );
not U87634 ( n6625, n59053 );
nand U87635 ( n68423, n68883, n6024 );
nand U87636 ( n26422, n26884, n4247 );
nand U87637 ( n59561, n60024, n6879 );
nor U87638 ( n71753, n71754, n1203 );
nor U87639 ( n11652, n76572, n76789 );
nand U87640 ( n71756, n71877, n71878 );
or U87641 ( n71877, n71743, n71741 );
nand U87642 ( n71878, n71744, n71879 );
nand U87643 ( n71879, n71741, n71743 );
not U87644 ( n1240, n71267 );
nand U87645 ( n71885, n1238, n76043 );
nand U87646 ( n68418, n68876, n6019 );
nand U87647 ( n26417, n26877, n4242 );
nand U87648 ( n59556, n60017, n6874 );
nand U87649 ( n26427, n26884, n4242 );
nand U87650 ( n59566, n60024, n6874 );
nand U87651 ( n68428, n68883, n6019 );
xor U87652 ( n71869, n72022, n72023 );
xor U87653 ( n72023, n72024, n72025 );
nor U87654 ( n71865, n71872, n1199 );
nand U87655 ( n72356, n71312, n71245 );
nor U87656 ( n37563, n1970, n37500 );
not U87657 ( n1970, n37501 );
nand U87658 ( n47683, n47696, n47697 );
nor U87659 ( n47697, n47698, n47699 );
nor U87660 ( n47696, n47712, n47713 );
nand U87661 ( n47698, n47706, n47707 );
not U87662 ( n1389, n52649 );
nand U87663 ( n47369, n47846, n7812 );
nor U87664 ( n47846, n43287, n47849 );
nand U87665 ( n68391, n68859, n6024 );
not U87666 ( n6015, n68869 );
nor U87667 ( n68859, n6015, n63972 );
nand U87668 ( n26390, n26860, n4247 );
nand U87669 ( n59529, n60000, n6879 );
not U87670 ( n4238, n26870 );
not U87671 ( n6870, n60010 );
nor U87672 ( n26860, n4238, n22693 );
nor U87673 ( n60000, n6870, n55809 );
xnor U87674 ( n71298, n71292, n71442 );
xor U87675 ( n71442, n71293, n71295 );
nand U87676 ( n71293, n71443, n71265 );
nor U87677 ( n71443, n1233, n1240 );
not U87678 ( n639, n40984 );
nand U87679 ( n47374, n47846, n7807 );
nand U87680 ( n26395, n26860, n4242 );
nand U87681 ( n59534, n60000, n6874 );
nand U87682 ( n68396, n68859, n6019 );
nand U87683 ( n36710, n36711, n36712 );
nand U87684 ( n36711, n76822, n36730 );
nand U87685 ( n36712, n36713, n76830 );
nor U87686 ( n36713, n36714, n36715 );
nand U87687 ( n3126, n36707, n36708 );
nor U87688 ( n36707, n36731, n36732 );
nor U87689 ( n36708, n36709, n36710 );
nand U87690 ( n36732, n36733, n36734 );
or U87691 ( n41418, n41112, n41113 );
nor U87692 ( n41770, n41742, n41743 );
nand U87693 ( n40929, n40925, n40926 );
nand U87694 ( n38354, n39583, n39584 );
nor U87695 ( n39583, n39615, n39616 );
nor U87696 ( n39584, n39585, n39586 );
nor U87697 ( n39615, n2174, n38822 );
nand U87698 ( n39604, n39652, n39653 );
nor U87699 ( n39653, n39654, n39655 );
nor U87700 ( n39652, n39656, n39657 );
nor U87701 ( n39655, n39594, n38865 );
nand U87702 ( n39674, n39554, n37501 );
nand U87703 ( n65946, n660, n793 );
nor U87704 ( n39654, n39594, n38866 );
nor U87705 ( n41771, n41772, n41773 );
nor U87706 ( n39656, n39594, n37513 );
nand U87707 ( n26703, n26716, n26717 );
nor U87708 ( n26717, n26718, n26719 );
nor U87709 ( n26716, n26732, n26733 );
nand U87710 ( n26718, n26726, n26727 );
nand U87711 ( n68704, n68717, n68718 );
nor U87712 ( n68718, n68719, n68720 );
nor U87713 ( n68717, n68733, n68734 );
nand U87714 ( n68719, n68727, n68728 );
nand U87715 ( n59845, n59858, n59859 );
nor U87716 ( n59859, n59860, n59861 );
nor U87717 ( n59858, n59874, n59875 );
nand U87718 ( n59860, n59868, n59869 );
nand U87719 ( n71743, n71886, n71265 );
nor U87720 ( n71886, n1239, n1222 );
nand U87721 ( n38223, n38228, n38229 );
nand U87722 ( n38228, n76439, n36551 );
nand U87723 ( n38229, n38230, n76443 );
xnor U87724 ( n71751, n71887, n71888 );
xnor U87725 ( n71888, n71889, n71890 );
nor U87726 ( n71747, n71754, n1202 );
nand U87727 ( n2746, n38339, n38340 );
nor U87728 ( n38340, n38341, n38342 );
nor U87729 ( n38339, n38350, n38351 );
nand U87730 ( n38341, n38347, n38348 );
nand U87731 ( n71301, n71299, n71245 );
nand U87732 ( n39204, n39205, n39206 );
nand U87733 ( n39206, n38246, n76797 );
nand U87734 ( n39205, n2033, n38247 );
nand U87735 ( n71448, n71276, n71449 );
nand U87736 ( n71449, n1242, n76044 );
and U87737 ( n71292, n71444, n71445 );
nand U87738 ( n71445, n71446, n71266 );
nand U87739 ( n71444, n71448, n71267 );
nand U87740 ( n71446, n71272, n71447 );
nand U87741 ( n40906, n40829, n41296 );
nand U87742 ( n41296, n76848, n41297 );
nand U87743 ( n68401, n68866, n6024 );
nand U87744 ( n26400, n26867, n4247 );
nand U87745 ( n59539, n60007, n6879 );
nor U87746 ( n68866, n63972, n68869 );
nor U87747 ( n26867, n22693, n26870 );
nor U87748 ( n60007, n55809, n60010 );
nor U87749 ( n36714, n36720, n36721 );
xor U87750 ( n36720, n36728, n36729 );
nand U87751 ( n36721, n36722, n1963 );
nand U87752 ( n36722, n36530, n36531 );
nor U87753 ( n71222, n1162, n71247 );
nand U87754 ( n41544, n798, n41114 );
nand U87755 ( n68406, n68866, n6019 );
nand U87756 ( n26405, n26867, n4242 );
nand U87757 ( n59544, n60007, n6874 );
nand U87758 ( n41094, n41095, n41096 );
nand U87759 ( n41095, n584, n41114 );
nand U87760 ( n41096, n41097, n76850 );
nor U87761 ( n41097, n41098, n41099 );
nand U87762 ( n1901, n41091, n41092 );
nor U87763 ( n41091, n41115, n41116 );
nor U87764 ( n41092, n41093, n41094 );
nand U87765 ( n41116, n41117, n41118 );
not U87766 ( n1954, n39747 );
nand U87767 ( n37573, n1967, n36322 );
nand U87768 ( n39738, n2169, n1953 );
nand U87769 ( n41691, n41696, n41705 );
nand U87770 ( n41705, n664, n41694 );
not U87771 ( n664, n41697 );
or U87772 ( n41699, n41691, n75770 );
and U87773 ( n75770, n41690, n41689 );
nand U87774 ( n41696, n41684, n41685 );
nand U87775 ( n71873, n71872, n71874 );
nand U87776 ( n36314, n36315, n36316 );
nand U87777 ( n36315, n76821, n36322 );
nand U87778 ( n36316, n76832, n36317 );
xnor U87779 ( n36317, n36318, n36319 );
xnor U87780 ( n36319, n36320, n36321 );
nand U87781 ( n3221, n36311, n36312 );
nor U87782 ( n36311, n36323, n36324 );
nor U87783 ( n36312, n36313, n36314 );
nand U87784 ( n36324, n36325, n36326 );
not U87785 ( n650, n40690 );
nor U87786 ( n71890, n1239, n1205 );
nor U87787 ( n41098, n41104, n41105 );
xor U87788 ( n41104, n41112, n41113 );
nand U87789 ( n41105, n41106, n588 );
nand U87790 ( n41106, n40928, n40929 );
nor U87791 ( n62956, n62959, n62960 );
nor U87792 ( n62959, n41487, n62866 );
nor U87793 ( n62960, n62272, n62866 );
nand U87794 ( n36531, n36527, n36528 );
not U87795 ( n2543, n19717 );
nand U87796 ( n40719, n40720, n40721 );
nand U87797 ( n40720, n584, n40727 );
nand U87798 ( n40721, n76852, n40722 );
xnor U87799 ( n40722, n40723, n40724 );
xnor U87800 ( n40724, n40725, n40726 );
nand U87801 ( n1996, n40716, n40717 );
nor U87802 ( n40716, n40728, n40729 );
nor U87803 ( n40717, n40718, n40719 );
nand U87804 ( n40729, n40730, n40731 );
nand U87805 ( n47533, n47619, n47620 );
nor U87806 ( n47620, n47621, n47622 );
nor U87807 ( n47619, n47635, n47636 );
nand U87808 ( n47621, n47629, n47630 );
not U87809 ( n7809, n47864 );
nor U87810 ( n64387, n684, n798 );
nor U87811 ( n62961, n62963, n62964 );
nor U87812 ( n62963, n61618, n62866 );
nor U87813 ( n62964, n61617, n62866 );
not U87814 ( n7808, n44517 );
or U87815 ( n37051, n36728, n36729 );
and U87816 ( n40908, n40829, n41293 );
nand U87817 ( n41293, n76848, n41090 );
nor U87818 ( n39460, n39462, n39463 );
and U87819 ( n39462, n39419, n2005 );
nor U87820 ( n39463, n37513, n39430 );
nand U87821 ( n38322, n39453, n39454 );
nand U87822 ( n39454, n2074, n36797 );
nor U87823 ( n39453, n39455, n39456 );
nor U87824 ( n39455, n39470, n37367 );
nand U87825 ( n37491, n1969, n36961 );
nand U87826 ( n41108, n41142, n41144 );
nor U87827 ( n39465, n39466, n39467 );
nor U87828 ( n39466, n38866, n39430 );
nor U87829 ( n39467, n38865, n39430 );
not U87830 ( n648, n41198 );
nand U87831 ( n39266, n39267, n39268 );
nand U87832 ( n39267, n38267, n76797 );
nand U87833 ( n39268, n38262, n2033 );
nand U87834 ( n2756, n38307, n38308 );
nor U87835 ( n38308, n38309, n38310 );
nor U87836 ( n38307, n38318, n38319 );
nand U87837 ( n38309, n38315, n38316 );
nor U87838 ( n72649, n71247, n1232 );
not U87839 ( n1242, n71266 );
buf U87840 ( n76253, n76251 );
nor U87841 ( n71769, n71770, n71771 );
nor U87842 ( n71770, n71772, n71773 );
and U87843 ( n71772, n71774, n1122 );
not U87844 ( n1310, n52072 );
nor U87845 ( n64380, n64382, n64514 );
nor U87846 ( n64386, n799, n689 );
nand U87847 ( n62575, n76386, n40913 );
nand U87848 ( n68554, n68640, n68641 );
nor U87849 ( n68641, n68642, n68643 );
nor U87850 ( n68640, n68656, n68657 );
nand U87851 ( n68642, n68650, n68651 );
nand U87852 ( n26553, n26639, n26640 );
nor U87853 ( n26640, n26641, n26642 );
nor U87854 ( n26639, n26655, n26656 );
nand U87855 ( n26641, n26649, n26650 );
nand U87856 ( n59695, n59781, n59782 );
nor U87857 ( n59782, n59783, n59784 );
nor U87858 ( n59781, n59797, n59798 );
nand U87859 ( n59783, n59791, n59792 );
not U87860 ( n6022, n68884 );
not U87861 ( n4244, n26885 );
not U87862 ( n6877, n60025 );
nor U87863 ( n66276, n54645, n76243 );
not U87864 ( n6020, n65392 );
nand U87865 ( n62860, n62861, n62862 );
nand U87866 ( n62861, n813, n41284 );
nand U87867 ( n62862, n837, n62848 );
not U87868 ( n4243, n23846 );
not U87869 ( n6875, n56970 );
not U87870 ( n2603, n19263 );
xnor U87871 ( MUL_1411_U9, n71025, n71026 );
xnor U87872 ( n71025, n71027, n71028 );
nor U87873 ( n71744, n1205, n1222 );
nor U87874 ( n39477, n39483, n39484 );
nor U87875 ( n39483, n2039, n39426 );
nor U87876 ( n39484, n38875, n39419 );
nor U87877 ( n41107, n40926, n40925 );
nand U87878 ( n41546, n799, n40727 );
nand U87879 ( n3176, n36517, n36518 );
nor U87880 ( n36517, n36533, n36534 );
nor U87881 ( n36518, n36519, n36520 );
nand U87882 ( n36534, n36535, n36536 );
nand U87883 ( n36520, n36521, n36522 );
nand U87884 ( n36521, n76821, n36532 );
nand U87885 ( n36522, n76831, n36523 );
nand U87886 ( n36523, n36524, n36525 );
nand U87887 ( n36525, n36526, n1845 );
xor U87888 ( n36526, n36527, n36528 );
nor U87889 ( n64385, n797, n679 );
nor U87890 ( n46441, n46453, n45623 );
nor U87891 ( n67505, n67369, n66548 );
nor U87892 ( n25500, n25364, n24713 );
nor U87893 ( n58637, n58501, n57847 );
nand U87894 ( n38239, n38244, n38245 );
nand U87895 ( n38245, n38246, n76818 );
nand U87896 ( n38244, n38247, n76442 );
not U87897 ( n2164, n36462 );
nand U87898 ( n41540, n800, n41329 );
nand U87899 ( n63709, n697, n42042 );
or U87900 ( n41687, n75771, n41689 );
or U87901 ( n75771, n41690, n41691 );
nor U87902 ( n11664, n76569, n76789 );
nor U87903 ( n64211, n64032, n61617 );
nand U87904 ( n64226, n63706, n41535 );
nand U87905 ( n48685, n63994, n63995 );
nor U87906 ( n63994, n64026, n64027 );
nor U87907 ( n63995, n63996, n63997 );
nor U87908 ( n64026, n700, n61441 );
nand U87909 ( n64014, n64208, n64209 );
nor U87910 ( n64208, n64213, n64214 );
nor U87911 ( n64209, n64210, n64211 );
nor U87912 ( n64213, n64032, n41487 );
nor U87913 ( n64010, n699, n64012 );
nor U87914 ( n64012, n64013, n64014 );
and U87915 ( n64013, n61410, n42049 );
nand U87916 ( n62833, n535, n62781 );
not U87917 ( n7810, n44509 );
nor U87918 ( n41532, n42049, n42099 );
nand U87919 ( n48458, n63271, n63272 );
nand U87920 ( n63272, n813, n41178 );
nor U87921 ( n63271, n63273, n63274 );
nor U87922 ( n63274, n718, n63275 );
xor U87923 ( n36760, n36727, n36761 );
nand U87924 ( n36755, n36756, n36757 );
nand U87925 ( n36756, n76822, n36762 );
nand U87926 ( n36757, n76830, n36758 );
xor U87927 ( n36758, n36759, n36760 );
nand U87928 ( n3116, n36752, n36753 );
nor U87929 ( n36752, n36763, n36764 );
nor U87930 ( n36753, n36754, n36755 );
nand U87931 ( n36764, n36765, n36766 );
nand U87932 ( n1521, n48670, n48671 );
nor U87933 ( n48671, n48672, n48673 );
nor U87934 ( n48670, n48680, n48681 );
nand U87935 ( n48672, n48677, n48678 );
nand U87936 ( n1531, n48443, n48444 );
nor U87937 ( n48444, n48445, n48446 );
nor U87938 ( n48443, n48454, n48455 );
nand U87939 ( n48446, n48447, n48448 );
nand U87940 ( n40918, n40919, n40920 );
nand U87941 ( n40919, n584, n40930 );
nand U87942 ( n40920, n76851, n40921 );
nand U87943 ( n40921, n40922, n40923 );
nand U87944 ( n1951, n40915, n40916 );
nor U87945 ( n40915, n40931, n40932 );
nor U87946 ( n40916, n40917, n40918 );
nand U87947 ( n40932, n40933, n40934 );
nand U87948 ( n40923, n40924, n519 );
xor U87949 ( n40924, n40925, n40926 );
nand U87950 ( n36724, n36759, n36761 );
nor U87951 ( n72508, n71247, n1230 );
nor U87952 ( n41110, n41144, n41142 );
not U87953 ( n6023, n65384 );
not U87954 ( n4245, n23838 );
not U87955 ( n6878, n56962 );
not U87956 ( n2507, n19577 );
nand U87957 ( n64805, n679, n797 );
xor U87958 ( n45462, n45463, n45464 );
nand U87959 ( n72007, n71357, n71245 );
nand U87960 ( n47479, n47541, n47542 );
nor U87961 ( n47542, n47543, n47544 );
nor U87962 ( n47541, n47557, n47558 );
nand U87963 ( n47543, n47551, n47552 );
nor U87964 ( n41681, n675, n41682 );
not U87965 ( n675, n41683 );
nand U87966 ( n38255, n38260, n38261 );
nand U87967 ( n38260, n76439, n36339 );
nand U87968 ( n38261, n38262, n76442 );
nor U87969 ( n63278, n63280, n63281 );
nor U87970 ( n63281, n41487, n62979 );
and U87971 ( n63280, n62677, n822 );
nand U87972 ( n47413, n47414, n47415 );
nand U87973 ( n47414, n76339, n40747 );
or U87974 ( n47415, n47416, n573 );
and U87975 ( n63705, n63707, n41535 );
and U87976 ( n63707, n41596, n42042 );
nor U87977 ( n36723, n36528, n36527 );
nand U87978 ( n48070, n48071, n48072 );
nand U87979 ( n48071, n76339, n40913 );
nand U87980 ( n48072, n48073, n45754 );
and U87981 ( n48073, n48074, n48075 );
nor U87982 ( n39328, n38276, n38764 );
not U87983 ( n654, n40864 );
nand U87984 ( n39669, n2173, n1969 );
xnor U87985 ( n41143, n41144, n41111 );
nand U87986 ( n41138, n41139, n41140 );
nand U87987 ( n41139, n584, n41145 );
nand U87988 ( n41140, n76850, n41141 );
xor U87989 ( n41141, n41142, n41143 );
nand U87990 ( n1891, n41135, n41136 );
nor U87991 ( n41135, n41146, n41147 );
nor U87992 ( n41136, n41137, n41138 );
nand U87993 ( n41147, n41148, n41149 );
nor U87994 ( n41680, n41684, n41685 );
nor U87995 ( n63285, n61617, n62979 );
not U87996 ( n2168, n36762 );
nand U87997 ( n68500, n68562, n68563 );
nor U87998 ( n68563, n68564, n68565 );
nor U87999 ( n68562, n68578, n68579 );
nand U88000 ( n68564, n68572, n68573 );
nand U88001 ( n26499, n26561, n26562 );
nor U88002 ( n26562, n26563, n26564 );
nor U88003 ( n26561, n26577, n26578 );
nand U88004 ( n26563, n26571, n26572 );
nand U88005 ( n59638, n59703, n59704 );
nor U88006 ( n59704, n59705, n59706 );
nor U88007 ( n59703, n59719, n59720 );
nand U88008 ( n59705, n59713, n59714 );
nand U88009 ( n2751, n38323, n38324 );
nor U88010 ( n38324, n38325, n38326 );
nor U88011 ( n38323, n38333, n38334 );
nand U88012 ( n38325, n38330, n38331 );
nand U88013 ( n41102, n41113, n41112 );
and U88014 ( n41679, n41784, n41793 );
nand U88015 ( n41793, n680, n41782 );
not U88016 ( n680, n41785 );
xnor U88017 ( n71066, n71761, n71762 );
xor U88018 ( n71761, n71763, n71764 );
nand U88019 ( n62779, n737, n76388 );
nor U88020 ( n37551, n36797, n1987 );
nor U88021 ( n39589, n39591, n38866 );
nand U88022 ( n39586, n39587, n39588 );
nand U88023 ( n39587, n39592, n39590 );
nand U88024 ( n39588, n39589, n39590 );
nor U88025 ( n39592, n39593, n38865 );
nand U88026 ( n41784, n41788, n41789 );
not U88027 ( n2167, n36355 );
nand U88028 ( n71775, n71774, n71776 );
nor U88029 ( n39619, n39591, n37513 );
not U88030 ( n2469, n19428 );
nand U88031 ( n62938, n62939, n62940 );
nand U88032 ( n62939, n784, n41297 );
nand U88033 ( n62940, n48328, n827 );
nor U88034 ( n41786, n41683, n41790 );
nand U88035 ( n41790, n41679, n41682 );
not U88036 ( n1268, n51706 );
nand U88037 ( n38370, n39644, n39645 );
nor U88038 ( n39644, n39659, n39660 );
nor U88039 ( n39645, n39646, n39647 );
nor U88040 ( n39660, n2173, n38822 );
xnor U88041 ( n41126, n40826, n41298 );
nor U88042 ( n41298, n41299, n40824 );
nor U88043 ( n41299, n745, n40825 );
nand U88044 ( n62471, n76386, n41134 );
nand U88045 ( n47333, n47449, n47450 );
nor U88046 ( n47450, n47451, n47452 );
nor U88047 ( n47449, n47465, n47466 );
nand U88048 ( n47451, n47459, n47460 );
nand U88049 ( n38272, n38273, n38274 );
nand U88050 ( n38274, n76447, n2894 );
nand U88051 ( n38273, n1870, n76442 );
not U88052 ( n1870, n38276 );
or U88053 ( n36726, n36761, n36759 );
nand U88054 ( n2741, n38355, n38356 );
nor U88055 ( n38356, n38357, n38358 );
nor U88056 ( n38355, n38365, n38366 );
nand U88057 ( n38358, n38359, n38360 );
not U88058 ( n2542, n19844 );
not U88059 ( n2165, n36667 );
nor U88060 ( n39968, n38440, n76404 );
buf U88061 ( n76404, n76402 );
nor U88062 ( n39664, n39670, n39671 );
nor U88063 ( n39670, n37513, n39658 );
nor U88064 ( n39671, n38956, n39658 );
nor U88065 ( n39672, n39675, n39676 );
and U88066 ( n39675, n37100, n39611 );
nor U88067 ( n39676, n38866, n39658 );
and U88068 ( n41627, n41634, n41635 );
nand U88069 ( n41634, n76011, n41297 );
not U88070 ( n679, n40930 );
not U88071 ( n2760, n16849 );
nand U88072 ( n68365, n68470, n68471 );
nor U88073 ( n68471, n68472, n68473 );
nor U88074 ( n68470, n68486, n68487 );
nand U88075 ( n68472, n68480, n68481 );
nand U88076 ( n26364, n26469, n26470 );
nor U88077 ( n26470, n26471, n26472 );
nor U88078 ( n26469, n26485, n26486 );
nand U88079 ( n26471, n26479, n26480 );
nand U88080 ( n59503, n59608, n59609 );
nor U88081 ( n59609, n59610, n59611 );
nor U88082 ( n59608, n59624, n59625 );
nand U88083 ( n59610, n59618, n59619 );
nand U88084 ( n39612, n2174, n1975 );
nand U88085 ( n1526, n48560, n48561 );
nor U88086 ( n48561, n48562, n48563 );
nor U88087 ( n48560, n48571, n48572 );
nand U88088 ( n48562, n48568, n48569 );
nor U88089 ( n72468, n71247, n1223 );
not U88090 ( n672, n41145 );
nand U88091 ( n36718, n36729, n36728 );
not U88092 ( n1604, n49787 );
nor U88093 ( n41674, n41782, n41783 );
nand U88094 ( n41783, n41784, n41785 );
nor U88095 ( n72606, n71247, n1224 );
nand U88096 ( n37498, n1987, n36797 );
not U88097 ( n2429, n19208 );
nor U88098 ( n72162, n1237, n71247 );
nor U88099 ( n40047, n38476, n76405 );
buf U88100 ( n76242, n76240 );
xnor U88101 ( n45451, n45453, n45454 );
nor U88102 ( n65928, n49373, n76242 );
and U88103 ( n71069, n71707, n71708 );
or U88104 ( n71707, n71510, n71509 );
nand U88105 ( n71708, n71511, n71709 );
nand U88106 ( n71709, n71509, n71510 );
nand U88107 ( n36347, n36348, n36349 );
nand U88108 ( n36348, n76821, n36355 );
nand U88109 ( n36349, n76831, n36350 );
xnor U88110 ( n36350, n36351, n36352 );
xnor U88111 ( n36352, n36353, n36354 );
nand U88112 ( n3211, n36344, n36345 );
nor U88113 ( n36344, n36356, n36357 );
nor U88114 ( n36345, n36346, n36347 );
nand U88115 ( n36357, n36358, n36359 );
nand U88116 ( n62679, n743, n76388 );
nor U88117 ( n72225, n1235, n71247 );
nand U88118 ( n48803, n64203, n64204 );
nor U88119 ( n64203, n64217, n64218 );
nor U88120 ( n64204, n64205, n64206 );
nor U88121 ( n64218, n695, n61441 );
and U88122 ( n64206, n64014, n75772 );
or U88123 ( n75772, n42049, n699 );
nand U88124 ( n39492, n2177, n1987 );
nand U88125 ( n39491, n2175, n1982 );
nand U88126 ( n47288, n47351, n47352 );
nor U88127 ( n47352, n47353, n47354 );
nor U88128 ( n47351, n47375, n47376 );
nand U88129 ( n47353, n47365, n47366 );
xor U88130 ( n71229, n71237, n71238 );
xor U88131 ( n71238, n71239, n71240 );
xor U88132 ( n71237, n71248, n71249 );
nor U88133 ( n71239, n1227, n71247 );
not U88134 ( n1934, n37260 );
nor U88135 ( n41556, n41557, n41558 );
nand U88136 ( n41557, n41568, n41569 );
nand U88137 ( n41558, n41559, n41560 );
nand U88138 ( n41559, n41561, n41562 );
nand U88139 ( n41566, n42084, n42085 );
nand U88140 ( n42085, n42086, n635 );
nor U88141 ( n42086, n787, n637 );
nor U88142 ( n41536, n41537, n41538 );
nand U88143 ( n41538, n41539, n41540 );
nand U88144 ( n41537, n41545, n41546 );
nand U88145 ( n41539, n41541, n41542 );
nor U88146 ( n41500, n41501, n41502 );
and U88147 ( n41502, n41503, n41504 );
nor U88148 ( n41501, n41505, n41506 );
nand U88149 ( n41506, n41507, n41503 );
nor U88150 ( n41526, n41530, n41531 );
nand U88151 ( n41531, n41532, n41533 );
nand U88152 ( n41533, n41534, n41535 );
nor U88153 ( n41534, n699, n41536 );
nand U88154 ( n64233, n695, n800 );
nand U88155 ( n1516, n48788, n48789 );
nor U88156 ( n48789, n48790, n48791 );
nor U88157 ( n48788, n48799, n48800 );
nand U88158 ( n48791, n48792, n48793 );
nor U88159 ( n64030, n64004, n41487 );
xor U88160 ( n39537, n39482, n37360 );
nor U88161 ( n64003, n64004, n61617 );
not U88162 ( n660, n41054 );
nand U88163 ( n39546, n39547, n39548 );
nand U88164 ( n39547, n2074, n36613 );
nand U88165 ( n39548, n39537, n2038 );
nor U88166 ( n72323, n71247, n1234 );
xor U88167 ( n11687, n11688, n11689 );
nand U88168 ( n42098, n804, n41178 );
not U88169 ( n1939, n37583 );
nor U88170 ( n39724, n39726, n39727 );
nor U88171 ( n39726, n38865, n39554 );
nor U88172 ( n39727, n37513, n39554 );
buf U88173 ( n76411, n38757 );
xnor U88174 ( n40739, n40826, n41300 );
nor U88175 ( n41300, n41301, n40824 );
nor U88176 ( n41301, n750, n40825 );
nand U88177 ( n68319, n68383, n68384 );
nor U88178 ( n68384, n68385, n68386 );
nor U88179 ( n68383, n68407, n68408 );
nand U88180 ( n68385, n68397, n68398 );
nand U88181 ( n26318, n26382, n26383 );
nor U88182 ( n26383, n26384, n26385 );
nor U88183 ( n26382, n26406, n26407 );
nand U88184 ( n26384, n26396, n26397 );
nand U88185 ( n59457, n59521, n59522 );
nor U88186 ( n59522, n59523, n59524 );
nor U88187 ( n59521, n59545, n59546 );
nand U88188 ( n59523, n59535, n59536 );
nand U88189 ( n33657, n34122, n3409 );
nand U88190 ( n31607, n34014, n34015 );
nor U88191 ( n34015, n34016, n34017 );
nor U88192 ( n34014, n34030, n34031 );
nand U88193 ( n34016, n34024, n34025 );
nand U88194 ( n34259, n3397, n3403 );
not U88195 ( n3394, n30016 );
nor U88196 ( n34122, n34115, n3394 );
nor U88197 ( n32776, n32817, n32818 );
and U88198 ( n32818, n32780, n76471 );
nand U88199 ( n33667, n34129, n3409 );
and U88200 ( n41623, n41849, n41632 );
nand U88201 ( n41849, n41090, n76379 );
nand U88202 ( n40752, n40753, n40754 );
nand U88203 ( n40753, n584, n40760 );
nand U88204 ( n40754, n76852, n40755 );
xnor U88205 ( n40755, n40756, n40757 );
xnor U88206 ( n40757, n40758, n40759 );
nand U88207 ( n1986, n40749, n40750 );
nor U88208 ( n40749, n40761, n40762 );
nor U88209 ( n40750, n40751, n40752 );
nand U88210 ( n40762, n40763, n40764 );
nand U88211 ( n33662, n34122, n3404 );
nand U88212 ( n2736, n38371, n38372 );
nor U88213 ( n38372, n38373, n38374 );
nor U88214 ( n38371, n38382, n38383 );
nand U88215 ( n38374, n38375, n38376 );
nand U88216 ( n33672, n34129, n3404 );
nor U88217 ( n41882, n41863, n41862 );
nor U88218 ( n72035, n1238, n71247 );
nand U88219 ( n41624, n41848, n41635 );
nand U88220 ( n41848, n76383, n41090 );
nand U88221 ( n41900, n41904, n41632 );
nand U88222 ( n41904, n40713, n76380 );
xor U88223 ( MUL_1411_U8, n71029, n71030 );
xor U88224 ( n71029, n71031, n71032 );
nand U88225 ( n33635, n34105, n3409 );
not U88226 ( n3400, n34115 );
nor U88227 ( n34105, n3400, n30016 );
nand U88228 ( n62291, n76386, n40950 );
and U88229 ( n41887, n41894, n41632 );
nand U88230 ( n41894, n40852, n76380 );
and U88231 ( n41885, n780, n41632 );
nand U88232 ( n62290, n76386, n40747 );
nand U88233 ( n33640, n34105, n3404 );
and U88234 ( n41899, n41903, n41635 );
nand U88235 ( n41903, n76383, n40713 );
and U88236 ( n71232, n71305, n71306 );
nand U88237 ( n41888, n41895, n41635 );
nand U88238 ( n41895, n76383, n40852 );
nand U88239 ( n37488, n37567, n37568 );
or U88240 ( n37568, n37569, n1965 );
nand U88241 ( n42016, n41297, n76388 );
nand U88242 ( n33948, n33961, n33962 );
nor U88243 ( n33962, n33963, n33964 );
nor U88244 ( n33961, n33977, n33978 );
nand U88245 ( n33963, n33971, n33972 );
nand U88246 ( n41563, n41579, n41578 );
nor U88247 ( n66094, n54614, n76243 );
nand U88248 ( n41886, n780, n41635 );
buf U88249 ( n76794, n76790 );
nand U88250 ( n41129, n40829, n41241 );
nand U88251 ( n41241, n76848, n40913 );
nor U88252 ( n37571, n37420, n37572 );
nand U88253 ( n37572, n37573, n37574 );
xnor U88254 ( n71062, n71757, n71758 );
xnor U88255 ( n71757, n71759, n71760 );
nand U88256 ( n33645, n34112, n3409 );
nor U88257 ( n34112, n30016, n34115 );
buf U88258 ( n76245, n61295 );
nand U88259 ( n41976, n41978, n41979 );
nor U88260 ( n41979, n41980, n41981 );
nor U88261 ( n41978, n42027, n42028 );
nand U88262 ( n41981, n41982, n41983 );
nor U88263 ( n41964, n41973, n41490 );
nor U88264 ( n41973, n41974, n41975 );
nor U88265 ( n41974, n41976, n41977 );
and U88266 ( n41975, n41976, n840 );
nand U88267 ( n33650, n34112, n3404 );
nand U88268 ( n62289, n76386, n41024 );
nand U88269 ( n46277, n47800, n47801 );
nor U88270 ( n47801, n47802, n47803 );
nor U88271 ( n47800, n47816, n47817 );
nand U88272 ( n47802, n47810, n47811 );
nand U88273 ( n41841, n41859, n41632 );
nand U88274 ( n41859, n40747, n76380 );
not U88275 ( n667, n40760 );
and U88276 ( n41840, n41858, n41635 );
nand U88277 ( n41858, n76383, n40747 );
nand U88278 ( n71064, n71725, n71726 );
or U88279 ( n71725, n71512, n71515 );
nand U88280 ( n71726, n71514, n71727 );
nand U88281 ( n71727, n71515, n71512 );
nor U88282 ( n71749, n71750, n71751 );
nor U88283 ( n71750, n71752, n71753 );
and U88284 ( n71752, n71754, n1203 );
nand U88285 ( n41843, n41850, n41635 );
nand U88286 ( n41850, n76383, n41134 );
and U88287 ( n41846, n41852, n41632 );
nand U88288 ( n41852, n40913, n76380 );
nand U88289 ( n64025, n700, n802 );
nand U88290 ( n41847, n41853, n41635 );
nand U88291 ( n41853, n76383, n40913 );
nand U88292 ( n48920, n64353, n64354 );
nand U88293 ( n64354, n813, n40727 );
nor U88294 ( n64353, n64355, n64356 );
nor U88295 ( n64355, n64366, n41963 );
nor U88296 ( n39508, n38329, n38764 );
nor U88297 ( n71233, n71305, n71306 );
xor U88298 ( n36664, n36665, n36666 );
nand U88299 ( n36659, n36660, n36661 );
nand U88300 ( n36660, n76822, n36667 );
nand U88301 ( n36661, n76830, n36662 );
xor U88302 ( n36662, n36663, n36664 );
nand U88303 ( n3141, n36656, n36657 );
nor U88304 ( n36656, n36668, n36669 );
nor U88305 ( n36657, n36658, n36659 );
nand U88306 ( n36669, n36670, n36671 );
and U88307 ( n41842, n41851, n41632 );
nand U88308 ( n41851, n41134, n76379 );
not U88309 ( n653, n41578 );
nor U88310 ( n45473, n76089, n76835 );
nand U88311 ( n1511, n48905, n48906 );
nor U88312 ( n48906, n48907, n48908 );
nor U88313 ( n48905, n48916, n48917 );
nand U88314 ( n48908, n48909, n48910 );
nand U88315 ( n42014, n41090, n76388 );
xor U88316 ( n40942, n40826, n41226 );
nor U88317 ( n41226, n41227, n40824 );
nor U88318 ( n41227, n759, n40825 );
buf U88319 ( n76382, n75705 );
nand U88320 ( n42015, n40913, n76388 );
nand U88321 ( n71275, n71276, n71277 );
nand U88322 ( n71277, n1243, n71278 );
not U88323 ( n1243, n71271 );
nand U88324 ( n71256, n71257, n1205 );
nor U88325 ( n71257, n1240, n71258 );
nor U88326 ( n71249, n71250, n71251 );
nor U88327 ( n71250, n1207, n71267 );
nand U88328 ( n71251, n71252, n71253 );
nand U88329 ( n71252, n71260, n71261 );
nand U88330 ( n71258, n71268, n71269 );
nand U88331 ( n71269, n71270, n71271 );
nand U88332 ( n71268, n71275, n71266 );
nand U88333 ( n71270, n71272, n71273 );
nand U88334 ( n67338, n68820, n68821 );
nor U88335 ( n68821, n68822, n68823 );
nor U88336 ( n68820, n68836, n68837 );
nand U88337 ( n68822, n68830, n68831 );
nand U88338 ( n25331, n26821, n26822 );
nor U88339 ( n26822, n26823, n26824 );
nor U88340 ( n26821, n26837, n26838 );
nand U88341 ( n26823, n26831, n26832 );
nand U88342 ( n58470, n59961, n59962 );
nor U88343 ( n59962, n59963, n59964 );
nor U88344 ( n59961, n59977, n59978 );
nand U88345 ( n59963, n59971, n59972 );
not U88346 ( n2169, n36532 );
nand U88347 ( n63698, n63699, n63700 );
nand U88348 ( n63699, n813, n41006 );
nand U88349 ( n63700, n837, n63686 );
xor U88350 ( n40841, n40826, n41302 );
nor U88351 ( n41302, n41303, n40824 );
nor U88352 ( n41303, n754, n40825 );
or U88353 ( n39729, n39554, n38866 );
nand U88354 ( n41573, n66442, n41989 );
nand U88355 ( n66442, n553, n42001 );
nand U88356 ( n41571, n41572, n41573 );
nor U88357 ( n41572, n662, n41574 );
not U88358 ( n662, n41560 );
nand U88359 ( n41870, n41906, n41632 );
nand U88360 ( n41906, n40834, n76378 );
nand U88361 ( n63658, n63659, n63660 );
nand U88362 ( n63660, n48570, n76076 );
nand U88363 ( n63659, n48567, n827 );
nand U88364 ( n41872, n41876, n41632 );
nand U88365 ( n41876, n40950, n76380 );
and U88366 ( n41869, n41905, n41635 );
nand U88367 ( n41905, n76010, n40834 );
nand U88368 ( n42026, n42064, n42065 );
nor U88369 ( n42064, n42068, n41598 );
nor U88370 ( n42065, n41504, n42066 );
nor U88371 ( n42068, n780, n76385 );
nand U88372 ( n41987, n42008, n769 );
nor U88373 ( n42008, n637, n41574 );
nor U88374 ( n41995, n42003, n42004 );
nand U88375 ( n42004, n42005, n749 );
nand U88376 ( n42003, n42007, n633 );
nor U88377 ( n42005, n649, n42006 );
not U88378 ( n2505, n19693 );
nand U88379 ( n37593, n1994, n36398 );
xor U88380 ( n41051, n41052, n41053 );
nand U88381 ( n41046, n41047, n41048 );
nand U88382 ( n41047, n584, n41054 );
nand U88383 ( n41048, n76851, n41049 );
xor U88384 ( n41049, n41050, n41051 );
nand U88385 ( n1916, n41043, n41044 );
nor U88386 ( n41043, n41055, n41056 );
nor U88387 ( n41044, n41045, n41046 );
nand U88388 ( n41056, n41057, n41058 );
xnor U88389 ( n11673, n11675, n11677 );
and U88390 ( n41871, n41875, n41635 );
nand U88391 ( n41875, n76383, n40950 );
nand U88392 ( n33798, n33884, n33885 );
nor U88393 ( n33885, n33886, n33887 );
nor U88394 ( n33884, n33900, n33901 );
nand U88395 ( n33886, n33894, n33895 );
not U88396 ( n1309, n52184 );
nand U88397 ( n71261, n71262, n71263 );
nand U88398 ( n71262, n1205, n71258 );
nand U88399 ( n71263, n71264, n1207 );
nor U88400 ( n71264, n1205, n1240 );
nand U88401 ( n40965, n40962, n40961 );
nor U88402 ( n41259, n592, n41005 );
nor U88403 ( n39706, n39711, n39712 );
and U88404 ( n39712, n37491, n37501 );
nor U88405 ( n39711, n39713, n39714 );
nand U88406 ( n39713, n39717, n39718 );
nor U88407 ( n39566, n38346, n38764 );
nand U88408 ( n49035, n64502, n64503 );
nor U88409 ( n64502, n64520, n64521 );
nor U88410 ( n64503, n64504, n64505 );
nor U88411 ( n64520, n684, n61441 );
not U88412 ( n3407, n34130 );
not U88413 ( n3405, n31138 );
nand U88414 ( n41590, n805, n40801 );
nor U88415 ( n71290, n71294, n71295 );
and U88416 ( n71294, n71293, n71292 );
nand U88417 ( n1506, n49020, n49021 );
nor U88418 ( n49021, n49022, n49023 );
nor U88419 ( n49020, n49030, n49031 );
nand U88420 ( n49022, n49027, n49028 );
nand U88421 ( n38401, n39775, n39776 );
nor U88422 ( n39775, n39793, n39794 );
nor U88423 ( n39776, n39777, n39778 );
nor U88424 ( n39793, n2170, n38822 );
nand U88425 ( n39788, n39747, n39838 );
nand U88426 ( n39838, n39742, n39738 );
nor U88427 ( n38746, n38833, n2145 );
nor U88428 ( n38898, n39031, n2128 );
nand U88429 ( n39922, n39965, n1937 );
nand U88430 ( n39821, n39866, n1947 );
nand U88431 ( n38737, n38745, n38746 );
nor U88432 ( n38745, n2148, n2149 );
nand U88433 ( n38616, n38732, n38733 );
nand U88434 ( n38733, n2152, n76409 );
nor U88435 ( n38732, n2075, n38734 );
nor U88436 ( n38734, n38601, n38110 );
nand U88437 ( n38833, n38899, n38898 );
nor U88438 ( n38899, n2138, n2133 );
nand U88439 ( n39031, n39086, n39084 );
nor U88440 ( n39086, n2122, n2117 );
and U88441 ( n39084, n39210, n39209 );
nor U88442 ( n39210, n2113, n2107 );
and U88443 ( n39694, n39765, n1959 );
nand U88444 ( n38110, n38735, n38736 );
nand U88445 ( n38736, n2152, n38737 );
or U88446 ( n38735, n38737, n2152 );
nand U88447 ( n63307, n707, n803 );
and U88448 ( n63305, n63307, n63308 );
nand U88449 ( n63308, n804, n714 );
nand U88450 ( n62832, n730, n807 );
nand U88451 ( n71630, n72499, n71302 );
nand U88452 ( n2731, n38387, n38388 );
nor U88453 ( n38388, n38389, n38390 );
nor U88454 ( n38387, n38396, n38397 );
nand U88455 ( n38389, n38393, n38394 );
or U88456 ( n64361, n63706, n41487 );
nor U88457 ( n32740, n32604, n31945 );
nand U88458 ( n63983, n63984, n63985 );
nand U88459 ( n63984, n784, n41178 );
nand U88460 ( n63985, n48676, n827 );
nand U88461 ( n39420, n2178, n1994 );
not U88462 ( n1350, n52343 );
or U88463 ( n64363, n63706, n61617 );
not U88464 ( n2170, n36730 );
not U88465 ( n709, n63312 );
buf U88466 ( n76415, n76413 );
nand U88467 ( n41983, n41984, n41985 );
nor U88468 ( n41984, n41986, n41987 );
nor U88469 ( n41986, n41988, n627 );
not U88470 ( n627, n41989 );
nor U88471 ( n71855, n1239, n71247 );
nand U88472 ( n62578, n745, n76388 );
and U88473 ( n72497, n72453, n71302 );
nand U88474 ( n39803, n39747, n39836 );
nand U88475 ( n39836, n39739, n39738 );
nand U88476 ( n39801, n1864, n39749 );
nand U88477 ( n63311, n804, n63312 );
or U88478 ( n40966, n40961, n40962 );
not U88479 ( n3408, n31130 );
nand U88480 ( n36570, n36567, n36566 );
nor U88481 ( n36873, n1984, n36612 );
nand U88482 ( n38624, n38741, n38742 );
nand U88483 ( n38742, n2149, n76409 );
nor U88484 ( n38741, n2075, n38743 );
nor U88485 ( n38743, n38601, n38117 );
nand U88486 ( n48563, n48564, n48565 );
nand U88487 ( n48565, n76335, n1774 );
nand U88488 ( n48564, n48567, n45754 );
not U88489 ( n684, n41114 );
buf U88490 ( n76249, n76247 );
nand U88491 ( n39292, n39319, n39320 );
nand U88492 ( n39320, n39321, n39322 );
nand U88493 ( n39321, n2102, n36512 );
nand U88494 ( n40742, n40829, n41237 );
nand U88495 ( n41237, n76848, n41134 );
and U88496 ( n41860, n41878, n41632 );
nand U88497 ( n41878, n41024, n76380 );
nand U88498 ( n41861, n41877, n41635 );
nand U88499 ( n41877, n76383, n41024 );
nor U88500 ( n39869, n38408, n76404 );
nand U88501 ( n41568, n41577, n41578 );
nand U88502 ( n71755, n71754, n71756 );
nand U88503 ( n41019, n40829, n41233 );
nand U88504 ( n41233, n76848, n40747 );
nor U88505 ( n45484, n76093, n76835 );
nand U88506 ( n39787, n1879, n39749 );
not U88507 ( n1879, n39788 );
and U88508 ( n40945, n40829, n41228 );
nand U88509 ( n41228, n76848, n41024 );
not U88510 ( n2172, n36322 );
nor U88511 ( n39128, n37402, n39129 );
nor U88512 ( n39129, n2112, n37457 );
nand U88513 ( n37542, n2183, n2113 );
nand U88514 ( n33744, n33806, n33807 );
nor U88515 ( n33807, n33808, n33809 );
nor U88516 ( n33806, n33822, n33823 );
nand U88517 ( n33808, n33816, n33817 );
nand U88518 ( n37554, n2054, n36702 );
or U88519 ( n36571, n36566, n36567 );
nand U88520 ( n61587, n76386, n40834 );
nand U88521 ( n38417, n39831, n39832 );
nor U88522 ( n39831, n39839, n39840 );
nor U88523 ( n39832, n39833, n39834 );
nor U88524 ( n39840, n2169, n38822 );
not U88525 ( n2428, n19116 );
and U88526 ( n41215, n40829, n41224 );
nand U88527 ( n41224, n76849, n40950 );
nand U88528 ( n39346, n2179, n2054 );
nand U88529 ( n39294, n39319, n39346 );
nor U88530 ( n71583, n71247, n1229 );
nor U88531 ( n65321, n49136, n76242 );
nand U88532 ( n64491, n64492, n64493 );
nand U88533 ( n64492, n784, n41329 );
nand U88534 ( n64493, n49026, n827 );
nand U88535 ( n46563, n76658, n45718 );
nand U88536 ( n2726, n38402, n38403 );
nor U88537 ( n38403, n38404, n38405 );
nor U88538 ( n38402, n38413, n38414 );
nand U88539 ( n38404, n38410, n38411 );
nand U88540 ( n67610, n76706, n66644 );
nand U88541 ( n25605, n76752, n24809 );
nand U88542 ( n58742, n76685, n57943 );
nand U88543 ( n49145, n64793, n64794 );
nand U88544 ( n64794, n813, n40930 );
nor U88545 ( n64793, n64795, n64796 );
nor U88546 ( n64796, n64784, n64797 );
not U88547 ( n1267, n51814 );
nand U88548 ( n1501, n49130, n49131 );
nor U88549 ( n49131, n49132, n49133 );
nor U88550 ( n49130, n49141, n49142 );
nand U88551 ( n49132, n49138, n49139 );
nand U88552 ( n62680, n720, n805 );
or U88553 ( n64512, n64513, n64514 );
nand U88554 ( n46510, n76659, n45695 );
nand U88555 ( n41586, n807, n41284 );
nand U88556 ( n67571, n76707, n66619 );
nand U88557 ( n25566, n76753, n24784 );
nand U88558 ( n58703, n76686, n57918 );
nor U88559 ( n71426, n71247, n1228 );
nor U88560 ( n38115, n38109, n38117 );
nand U88561 ( n36454, n36455, n36456 );
nand U88562 ( n36455, n76821, n36462 );
nand U88563 ( n36456, n76831, n36457 );
xnor U88564 ( n36457, n36458, n36459 );
xnor U88565 ( n36459, n36460, n36461 );
nand U88566 ( n3191, n36451, n36452 );
nor U88567 ( n36451, n36463, n36464 );
nor U88568 ( n36452, n36453, n36454 );
nand U88569 ( n36464, n36465, n36466 );
not U88570 ( n2173, n36961 );
nand U88571 ( n71737, n71276, n71738 );
nand U88572 ( n71738, n1239, n76044 );
nand U88573 ( n71061, n71731, n71732 );
nand U88574 ( n71731, n71519, n71516 );
nand U88575 ( n71732, n71518, n71733 );
or U88576 ( n71733, n71516, n71519 );
nand U88577 ( n33609, n33714, n33715 );
nor U88578 ( n33715, n33716, n33717 );
nor U88579 ( n33714, n33730, n33731 );
nand U88580 ( n33716, n33724, n33725 );
not U88581 ( n2175, n36613 );
not U88582 ( n700, n40967 );
nor U88583 ( n71719, n71247, n1222 );
nand U88584 ( n37557, n2180, n2102 );
xor U88585 ( n40832, n40826, n40835 );
nor U88586 ( n40835, n40836, n40824 );
nor U88587 ( n40836, n768, n40825 );
nand U88588 ( n72366, n71312, n71302 );
nand U88589 ( n40856, n40857, n40858 );
nand U88590 ( n40857, n584, n40864 );
nand U88591 ( n40858, n76851, n40859 );
xnor U88592 ( n40859, n40860, n40861 );
xnor U88593 ( n40861, n40862, n40863 );
nand U88594 ( n1966, n40853, n40854 );
nor U88595 ( n40853, n40865, n40866 );
nor U88596 ( n40854, n40855, n40856 );
nand U88597 ( n40866, n40867, n40868 );
nand U88598 ( n62474, n750, n76388 );
nand U88599 ( n38357, n38362, n38363 );
nand U88600 ( n38362, n76439, n36613 );
nand U88601 ( n38363, n38364, n76443 );
not U88602 ( n689, n40727 );
nand U88603 ( n39689, n39690, n39691 );
nand U88604 ( n39691, n38380, n76797 );
nand U88605 ( n39690, n2033, n38381 );
nand U88606 ( n62847, n62781, n41933 );
nor U88607 ( n39768, n38377, n76404 );
nand U88608 ( n37546, n2182, n2107 );
xnor U88609 ( n71058, n71741, n71742 );
xnor U88610 ( n71742, n71743, n71744 );
nor U88611 ( n39638, n38345, n76404 );
nor U88612 ( n37552, n2053, n37553 );
not U88613 ( n2053, n37554 );
and U88614 ( n37450, n37549, n37550 );
nand U88615 ( n37550, n37551, n1993 );
nor U88616 ( n37549, n2059, n37552 );
not U88617 ( n2059, n37555 );
not U88618 ( n707, n41006 );
nand U88619 ( n41553, n42079, n42080 );
or U88620 ( n42080, n42081, n668 );
not U88621 ( n609, n41004 );
nand U88622 ( n38433, n39875, n39876 );
nor U88623 ( n39875, n39903, n39904 );
nor U88624 ( n39876, n39877, n39878 );
nor U88625 ( n39904, n2168, n38822 );
nand U88626 ( n39882, n39883, n39884 );
nand U88627 ( n39884, n39885, n37422 );
or U88628 ( n39883, n39742, n2002 );
nand U88629 ( n39885, n39886, n39887 );
nand U88630 ( n42102, n40747, n76388 );
nand U88631 ( n42041, n42095, n42096 );
nor U88632 ( n42095, n42099, n42024 );
nor U88633 ( n42096, n41589, n42097 );
nand U88634 ( n42097, n42016, n42014 );
nor U88635 ( n42038, n42039, n42040 );
nor U88636 ( n42040, n42041, n42042 );
nor U88637 ( n42039, n42043, n42006 );
nor U88638 ( n42043, n42044, n688 );
or U88639 ( n42006, n75773, n42041 );
or U88640 ( n75773, n697, n42049 );
nor U88641 ( n39761, n39773, n38764 );
nand U88642 ( n38449, n39933, n39934 );
nor U88643 ( n39933, n39946, n39947 );
nor U88644 ( n39934, n39935, n39936 );
nor U88645 ( n39947, n2167, n38822 );
nand U88646 ( n39942, n39899, n39985 );
nand U88647 ( n39985, n39902, n39901 );
nand U88648 ( n1491, n49367, n49368 );
nor U88649 ( n49368, n49369, n49370 );
nor U88650 ( n49367, n49376, n49377 );
nand U88651 ( n49370, n49371, n49372 );
nand U88652 ( n38429, n38430, n38431 );
nand U88653 ( n38431, n76819, n38432 );
nand U88654 ( n38430, n76812, n38433 );
nand U88655 ( n2721, n38418, n38419 );
nor U88656 ( n38419, n38420, n38421 );
nor U88657 ( n38418, n38428, n38429 );
nand U88658 ( n38421, n38422, n38423 );
nand U88659 ( n65354, n42082, n65816 );
nand U88660 ( n65816, n64809, n42079 );
nand U88661 ( n49268, n65327, n65328 );
nor U88662 ( n65327, n65349, n65350 );
nor U88663 ( n65328, n65329, n65330 );
nor U88664 ( n65350, n672, n61441 );
nand U88665 ( n2716, n38434, n38435 );
nor U88666 ( n38435, n38436, n38437 );
nor U88667 ( n38434, n38445, n38446 );
nand U88668 ( n38436, n38442, n38443 );
nand U88669 ( n38964, n38187, n76797 );
nor U88670 ( n71519, n1218, n1205 );
nand U88671 ( n72417, n71308, n71302 );
nand U88672 ( n1496, n49253, n49254 );
nor U88673 ( n49254, n49255, n49256 );
nor U88674 ( n49253, n49264, n49265 );
nand U88675 ( n49256, n49257, n49258 );
nand U88676 ( n66640, n66641, n66642 );
nand U88677 ( n66642, n5660, n63168 );
nand U88678 ( n66641, n76711, n66644 );
nand U88679 ( n24805, n24806, n24807 );
nand U88680 ( n24807, n3903, n22086 );
nand U88681 ( n24806, n76759, n24809 );
nand U88682 ( n57939, n57940, n57941 );
nand U88683 ( n57941, n6535, n55196 );
nand U88684 ( n57940, n76692, n57943 );
nor U88685 ( n39817, n38409, n38764 );
not U88686 ( n2384, n18750 );
nor U88687 ( n64504, n64519, n61617 );
xor U88688 ( n64519, n64376, n64515 );
nand U88689 ( n72411, n71410, n71308 );
nand U88690 ( n71260, n71265, n71266 );
nor U88691 ( n64197, n48679, n76242 );
nand U88692 ( n65798, n65799, n65800 );
nand U88693 ( n65799, n784, n40930 );
nand U88694 ( n65800, n528, n827 );
nand U88695 ( n36269, n36270, n36271 );
nand U88696 ( n36270, n76821, n36286 );
nand U88697 ( n36271, n36272, n76830 );
nor U88698 ( n36272, n36273, n36274 );
nand U88699 ( n3231, n36266, n36267 );
nor U88700 ( n36266, n36288, n36289 );
nor U88701 ( n36267, n36268, n36269 );
nand U88702 ( n36289, n36290, n36291 );
nor U88703 ( n39839, n39841, n39842 );
nor U88704 ( n39841, n39849, n39850 );
xor U88705 ( n39842, n39798, n1955 );
nand U88706 ( n39849, n38956, n37513 );
nor U88707 ( n36273, n36282, n36283 );
xor U88708 ( n36282, n36284, n36285 );
xor U88709 ( n40816, n40821, n40822 );
nor U88710 ( n40822, n40823, n40824 );
xor U88711 ( n40821, n40826, n40827 );
nor U88712 ( n40823, n775, n40825 );
nand U88713 ( n72490, n71410, n72453 );
nand U88714 ( n45691, n45692, n45693 );
nand U88715 ( n45693, n7434, n7958 );
nand U88716 ( n45692, n45695, n76662 );
nand U88717 ( n33563, n33627, n33628 );
nor U88718 ( n33628, n33629, n33630 );
nor U88719 ( n33627, n33651, n33652 );
nand U88720 ( n33629, n33641, n33642 );
not U88721 ( n1989, n36611 );
nand U88722 ( n39256, n2107, n36747 );
nor U88723 ( n41807, n802, n76378 );
not U88724 ( n1393, n51162 );
not U88725 ( n695, n41329 );
and U88726 ( n71984, n71357, n71302 );
nand U88727 ( n39908, n37442, n39949 );
nand U88728 ( n39949, n39848, n37445 );
nand U88729 ( n64338, n64339, n64340 );
nand U88730 ( n64340, n48914, n76076 );
nand U88731 ( n64339, n48915, n827 );
nand U88732 ( n39081, n38215, n76797 );
nand U88733 ( n40673, n40674, n40675 );
nand U88734 ( n40674, n584, n40690 );
nand U88735 ( n40675, n40676, n76850 );
nor U88736 ( n40676, n40677, n40678 );
nand U88737 ( n2006, n40670, n40671 );
nor U88738 ( n40670, n40692, n40693 );
nor U88739 ( n40671, n40672, n40673 );
nand U88740 ( n40693, n40694, n40695 );
nand U88741 ( n49577, n65934, n65935 );
nand U88742 ( n65935, n813, n41054 );
nor U88743 ( n65934, n65936, n65937 );
nor U88744 ( n65937, n65938, n65939 );
nor U88745 ( n40677, n40686, n40687 );
xor U88746 ( n40686, n40688, n40689 );
nand U88747 ( n40707, n40829, n40833 );
nand U88748 ( n40833, n76849, n40834 );
not U88749 ( n1100, n71410 );
nand U88750 ( n38373, n38378, n38379 );
nand U88751 ( n38379, n38380, n76819 );
nand U88752 ( n38378, n38381, n76443 );
nand U88753 ( n1486, n49562, n49563 );
nor U88754 ( n49563, n49564, n49565 );
nor U88755 ( n49562, n49573, n49574 );
nand U88756 ( n49564, n49570, n49571 );
xor U88757 ( n53889, n51761, n51759 );
nor U88758 ( n48701, n48139, n48692 );
nor U88759 ( n48607, n48139, n48598 );
nor U88760 ( n49067, n48139, n49058 );
nor U88761 ( n48972, n48139, n48963 );
nor U88762 ( n49336, n48139, n49327 );
nor U88763 ( n49429, n48139, n49420 );
nand U88764 ( n71472, n71574, n71302 );
nor U88765 ( n39918, n38441, n38764 );
nand U88766 ( n14032, n14619, n5157 );
nand U88767 ( n11304, n14485, n14487 );
nor U88768 ( n14487, n14488, n14489 );
nor U88769 ( n14485, n14505, n14507 );
nand U88770 ( n14488, n14498, n14499 );
nand U88771 ( n14797, n5144, n5150 );
not U88772 ( n5142, n9327 );
nor U88773 ( n14619, n14610, n5142 );
nor U88774 ( n12684, n12688, n76596 );
nor U88775 ( n12688, n12690, n12692 );
nand U88776 ( n12690, n12720, n12722 );
nand U88777 ( n12692, n12693, n12694 );
nand U88778 ( n47682, n47831, n47832 );
nor U88779 ( n47832, n47833, n47834 );
nor U88780 ( n47831, n47850, n47851 );
nand U88781 ( n47833, n47842, n47843 );
nand U88782 ( n14044, n14628, n5157 );
nor U88783 ( n49249, n48139, n49180 );
nor U88784 ( n48880, n48139, n48811 );
nor U88785 ( n51669, n48139, n49648 );
nor U88786 ( n12925, n12969, n12970 );
and U88787 ( n12970, n12930, n76035 );
nand U88788 ( n14038, n14619, n5152 );
nand U88789 ( n36510, n36696, n36695 );
nor U88790 ( n64496, n48911, n76242 );
nand U88791 ( n36895, n2020, n36511 );
nand U88792 ( n14050, n14628, n5152 );
nand U88793 ( n26702, n26852, n26853 );
nor U88794 ( n26853, n26854, n26855 );
nor U88795 ( n26852, n26871, n26872 );
nand U88796 ( n26854, n26863, n26864 );
nand U88797 ( n59844, n59992, n59993 );
nor U88798 ( n59993, n59994, n59995 );
nor U88799 ( n59992, n60011, n60012 );
nand U88800 ( n59994, n60003, n60004 );
nand U88801 ( n68703, n68851, n68852 );
nor U88802 ( n68852, n68853, n68854 );
nor U88803 ( n68851, n68870, n68871 );
nand U88804 ( n68853, n68862, n68863 );
or U88805 ( n65822, n65823, n65824 );
nand U88806 ( n41809, n41815, n41819 );
nand U88807 ( n41819, n41814, n41813 );
not U88808 ( n2725, n16832 );
nand U88809 ( n41815, n41824, n41825 );
nor U88810 ( n42048, n42049, n42041 );
nand U88811 ( n38461, n38462, n38463 );
nand U88812 ( n38463, n76819, n38464 );
nand U88813 ( n38462, n76812, n38465 );
nand U88814 ( n2711, n38450, n38451 );
nor U88815 ( n38451, n38452, n38453 );
nor U88816 ( n38450, n38460, n38461 );
nand U88817 ( n38453, n38454, n38455 );
nand U88818 ( n14412, n14419, n14420 );
nor U88819 ( n14420, n14422, n14423 );
nor U88820 ( n14419, n14439, n14440 );
nand U88821 ( n14422, n14432, n14433 );
nand U88822 ( n32573, n34066, n34067 );
nor U88823 ( n34067, n34068, n34069 );
nor U88824 ( n34066, n34082, n34083 );
nand U88825 ( n34068, n34076, n34077 );
nand U88826 ( n39863, n39864, n39865 );
nand U88827 ( n39864, n76798, n38432 );
nand U88828 ( n39865, n2033, n38427 );
not U88829 ( n1424, n51347 );
nand U88830 ( n72265, n71371, n71302 );
nand U88831 ( n49369, n49374, n49375 );
nand U88832 ( n49374, n76338, n40930 );
nand U88833 ( n49375, n528, n45754 );
nand U88834 ( n42100, n41024, n76388 );
not U88835 ( n1573, n49993 );
not U88836 ( n710, n41811 );
nand U88837 ( n62253, n754, n76388 );
nand U88838 ( n41642, n41812, n717 );
not U88839 ( n717, n41813 );
nor U88840 ( n41812, n41814, n723 );
not U88841 ( n723, n41815 );
nand U88842 ( n71215, n71413, n71302 );
nand U88843 ( n14004, n14598, n5157 );
nor U88844 ( n14598, n5148, n9327 );
nand U88845 ( n36897, n36908, n36909 );
nand U88846 ( n36909, n76807, n36747 );
nand U88847 ( n36908, n2107, n76826 );
nand U88848 ( n3101, n36803, n36804 );
nor U88849 ( n36803, n36818, n36819 );
nor U88850 ( n36804, n36805, n36806 );
nand U88851 ( n36819, n36820, n36821 );
nand U88852 ( n36806, n36807, n36808 );
nand U88853 ( n36807, n76822, n36817 );
nand U88854 ( n36808, n76830, n36809 );
nand U88855 ( n36809, n36810, n36811 );
nand U88856 ( n36811, n36812, n1847 );
xor U88857 ( n36812, n36814, n36815 );
nand U88858 ( n48907, n48912, n48913 );
nand U88859 ( n48913, n48914, n568 );
nand U88860 ( n48912, n48915, n45754 );
nor U88861 ( n39903, n39905, n39906 );
nand U88862 ( n39905, n37337, n37466 );
nand U88863 ( n39906, n39907, n38792 );
nand U88864 ( n39907, n39908, n37422 );
nand U88865 ( n14017, n14607, n5157 );
nor U88866 ( n14607, n9327, n14610 );
nand U88867 ( n14010, n14598, n5152 );
nand U88868 ( n38214, n38215, n76818 );
and U88869 ( n71518, n71734, n71265 );
nor U88870 ( n71734, n1218, n1222 );
not U88871 ( n5148, n14610 );
nand U88872 ( n62325, n759, n76388 );
and U88873 ( n36696, n36910, n36911 );
nand U88874 ( n36911, n76807, n36512 );
nand U88875 ( n36910, n2102, n76826 );
nand U88876 ( n14023, n14607, n5152 );
nand U88877 ( n37594, n2184, n2117 );
nand U88878 ( n39962, n39963, n39964 );
nand U88879 ( n39963, n76798, n38464 );
nand U88880 ( n39964, n2033, n38459 );
not U88881 ( n549, n62786 );
nor U88882 ( n45361, n45406, n45407 );
nor U88883 ( n45407, n45408, n45363 );
nand U88884 ( n62331, n764, n76388 );
nor U88885 ( n37185, n2102, n76803 );
nand U88886 ( n41187, n41188, n41189 );
nand U88887 ( n41188, n584, n41198 );
nand U88888 ( n41189, n76851, n41190 );
nand U88889 ( n41190, n41191, n41192 );
nand U88890 ( n41192, n41193, n520 );
xor U88891 ( n41193, n41195, n41196 );
nand U88892 ( n1876, n41184, n41185 );
nor U88893 ( n41184, n41199, n41200 );
nor U88894 ( n41185, n41186, n41187 );
nand U88895 ( n41200, n41201, n41202 );
nor U88896 ( n65349, n65351, n65352 );
nand U88897 ( n65351, n42077, n41931 );
nand U88898 ( n65352, n61410, n65353 );
nand U88899 ( n65353, n65354, n64814 );
nand U88900 ( n36698, n36394, n36396 );
nand U88901 ( n41543, n42091, n797 );
nor U88902 ( n42091, n679, n683 );
not U88903 ( n683, n42045 );
nand U88904 ( n14207, n14314, n14315 );
nor U88905 ( n14315, n14317, n14318 );
nor U88906 ( n14314, n14334, n14335 );
nand U88907 ( n14317, n14327, n14328 );
nor U88908 ( n48204, n549, n62825 );
and U88909 ( n62825, n76386, n62826 );
nand U88910 ( n62826, n62827, n807 );
nand U88911 ( n72210, n71371, n71410 );
not U88912 ( n714, n41178 );
xnor U88913 ( n38479, n39902, n37352 );
not U88914 ( n2174, n36572 );
xor U88915 ( n36586, n36587, n36588 );
nand U88916 ( n36581, n36582, n36583 );
nand U88917 ( n36582, n76822, n36589 );
nand U88918 ( n36583, n76831, n36584 );
xor U88919 ( n36584, n36585, n36586 );
nand U88920 ( n3161, n36578, n36579 );
nor U88921 ( n36578, n36590, n36591 );
nor U88922 ( n36579, n36580, n36581 );
nand U88923 ( n36591, n36592, n36593 );
nand U88924 ( n2706, n38470, n38471 );
nor U88925 ( n38471, n38472, n38473 );
nor U88926 ( n38470, n38481, n38482 );
nand U88927 ( n38473, n38474, n38475 );
nand U88928 ( n39181, n2113, n36339 );
not U88929 ( n7535, n46770 );
nand U88930 ( n46757, n76658, n45855 );
not U88931 ( n5749, n67817 );
not U88932 ( n3992, n25814 );
not U88933 ( n6624, n58952 );
nand U88934 ( n67804, n76706, n66806 );
nand U88935 ( n25801, n76752, n24928 );
nand U88936 ( n58939, n76685, n58065 );
nand U88937 ( n38420, n38425, n38426 );
nand U88938 ( n38425, n76438, n36730 );
nand U88939 ( n38426, n38427, n76443 );
nor U88940 ( n36701, n36695, n36696 );
or U88941 ( n71636, n1223, n71196 );
nor U88942 ( n38279, n39209, n39332 );
and U88943 ( n39332, n2102, n39333 );
nand U88944 ( n39333, n39334, n2054 );
nand U88945 ( n41982, n41991, n76385 );
nor U88946 ( n41991, n41598, n41992 );
nor U88947 ( n41992, n779, n780 );
nand U88948 ( n65312, n65313, n65314 );
nand U88949 ( n65314, n49262, n76078 );
nand U88950 ( n65313, n49263, n827 );
nand U88951 ( n61296, n810, n62784 );
nand U88952 ( n62784, n62785, n62786 );
nor U88953 ( n62785, n834, n76385 );
not U88954 ( n5153, n10724 );
not U88955 ( n5154, n14629 );
nand U88956 ( n71977, n71357, n71410 );
nand U88957 ( n49565, n49566, n49567 );
nand U88958 ( n49567, n76335, n1794 );
or U88959 ( n49566, n49569, n573 );
nor U88960 ( n72381, n1234, n71196 );
nor U88961 ( n36700, n36396, n36394 );
nor U88962 ( n16109, n14954, n16098 );
nor U88963 ( n16010, n14954, n15990 );
nor U88964 ( n15903, n14954, n15892 );
nor U88965 ( n15588, n14954, n15577 );
nor U88966 ( n15490, n14954, n15470 );
nor U88967 ( n16320, n14954, n16309 );
nor U88968 ( n16423, n14954, n16412 );
nand U88969 ( n46611, n76658, n45730 );
nand U88970 ( n67658, n76706, n66656 );
nand U88971 ( n25653, n76752, n24821 );
nand U88972 ( n58793, n76685, n57955 );
not U88973 ( n5155, n10714 );
nand U88974 ( n36504, n2024, n36897 );
not U88975 ( n2024, n36511 );
nand U88976 ( n62273, n40950, n76388 );
nand U88977 ( n42067, n40834, n76388 );
not U88978 ( n2108, n37457 );
nor U88979 ( n15807, n14954, n15712 );
nor U88980 ( n16223, n14954, n16130 );
nand U88981 ( n38501, n40055, n40056 );
nor U88982 ( n40055, n40065, n40066 );
nor U88983 ( n40056, n40057, n40058 );
nor U88984 ( n40066, n2163, n38822 );
nand U88985 ( n40053, n40061, n1935 );
not U88986 ( n1935, n37359 );
nor U88987 ( n40061, n1929, n40062 );
nor U88988 ( n40062, n40029, n40028 );
nor U88989 ( n71060, n1218, n1173 );
not U88990 ( n2468, n19550 );
nand U88991 ( n38452, n38457, n38458 );
nand U88992 ( n38457, n76438, n36762 );
nand U88993 ( n38458, n38459, n76443 );
nor U88994 ( n39976, n39979, n39980 );
and U88995 ( n39979, n37442, n37445 );
nand U88996 ( n39980, n39848, n38792 );
xor U88997 ( n20933, n18803, n18805 );
nand U88998 ( n2701, n38486, n38487 );
nor U88999 ( n38487, n38488, n38489 );
nor U89000 ( n38486, n38496, n38497 );
nand U89001 ( n38488, n38493, n38494 );
not U89002 ( n719, n41594 );
nor U89003 ( n41829, n41830, n41831 );
nor U89004 ( n41828, n41824, n41825 );
nand U89005 ( n55523, n550, n45408 );
not U89006 ( n550, n61296 );
not U89007 ( n2427, n19228 );
nand U89008 ( n40976, n40977, n40978 );
nand U89009 ( n40977, n584, n40984 );
nand U89010 ( n40978, n76851, n40979 );
xnor U89011 ( n40979, n40980, n40981 );
xnor U89012 ( n40981, n40982, n40983 );
nand U89013 ( n1936, n40973, n40974 );
nor U89014 ( n40973, n40985, n40986 );
nor U89015 ( n40974, n40975, n40976 );
nand U89016 ( n40986, n40987, n40988 );
nand U89017 ( n32845, n76773, n32041 );
xor U89018 ( n38299, n2054, n39334 );
nand U89019 ( n37490, n37494, n37495 );
nor U89020 ( n37495, n37496, n37497 );
and U89021 ( n37494, n37456, n1993 );
nand U89022 ( n37497, n37457, n37498 );
nand U89023 ( n37307, n37375, n37376 );
nor U89024 ( n37376, n37377, n37378 );
nor U89025 ( n37375, n37423, n37424 );
nand U89026 ( n37377, n37391, n37392 );
nor U89027 ( n37458, n37461, n37382 );
nor U89028 ( n37461, n37469, n37274 );
nor U89029 ( n37469, n37273, n37470 );
nor U89030 ( n37470, n37471, n1914 );
not U89031 ( n688, n41542 );
not U89032 ( n1103, n71910 );
not U89033 ( n2177, n36797 );
nand U89034 ( n14139, n14217, n14218 );
nor U89035 ( n14218, n14219, n14220 );
nor U89036 ( n14217, n14237, n14238 );
nand U89037 ( n14219, n14229, n14230 );
nor U89038 ( n37181, n2107, n76803 );
xnor U89039 ( n54618, n65945, n41949 );
nand U89040 ( n54623, n66014, n66015 );
nor U89041 ( n66014, n66031, n66032 );
nor U89042 ( n66015, n66016, n66017 );
nor U89043 ( n66032, n654, n61441 );
not U89044 ( n1265, n51830 );
nor U89045 ( n42062, n40834, n76387 );
nand U89046 ( n39440, n38317, n76797 );
nand U89047 ( n55261, n61170, n45408 );
nand U89048 ( n61170, n61171, n61172 );
nand U89049 ( n61172, n76386, n76070 );
nor U89050 ( n61171, n549, n61174 );
nand U89051 ( n39132, n2117, n36633 );
nand U89052 ( n32806, n76773, n32016 );
not U89053 ( n2178, n36398 );
nand U89054 ( n37431, n37432, n37433 );
nand U89055 ( n37432, n37434, n37435 );
nor U89056 ( n37435, n37436, n37437 );
or U89057 ( n37437, n37421, n1944 );
nand U89058 ( n1481, n54608, n54609 );
nor U89059 ( n54609, n54610, n54611 );
nor U89060 ( n54608, n54619, n54620 );
nand U89061 ( n54610, n54615, n54616 );
nand U89062 ( n40052, n40063, n37359 );
nor U89063 ( n40063, n40029, n40064 );
and U89064 ( n40064, n40026, n40028 );
nor U89065 ( n33026, n33055, n33056 );
nor U89066 ( n33056, n33025, n76021 );
nand U89067 ( n37596, n2185, n2122 );
not U89068 ( n548, n63262 );
nor U89069 ( n48452, n62827, n63261 );
nor U89070 ( n63261, n805, n548 );
or U89071 ( n72272, n1235, n71196 );
nand U89072 ( n61590, n768, n76388 );
nand U89073 ( n12863, n12864, n4890 );
not U89074 ( n720, n40801 );
nand U89075 ( n49255, n49260, n49261 );
nand U89076 ( n49261, n49262, n568 );
nand U89077 ( n49260, n49263, n45754 );
xor U89078 ( n48336, n62827, n807 );
nor U89079 ( n61429, n76387, n775 );
nand U89080 ( n61412, n775, n76388 );
nand U89081 ( n38517, n40099, n40100 );
nand U89082 ( n40100, n2074, n36817 );
nor U89083 ( n40099, n40101, n40102 );
nor U89084 ( n40101, n2034, n40115 );
and U89085 ( n37406, n37509, n37510 );
nor U89086 ( n37510, n2134, n2123 );
nor U89087 ( n37509, n2129, n37511 );
nor U89088 ( n37511, n2120, n37512 );
nor U89089 ( n39514, n38313, n76404 );
nor U89090 ( n42056, n42059, n41577 );
nor U89091 ( n42050, n42052, n42053 );
nand U89092 ( n42052, n42057, n42058 );
nand U89093 ( n42053, n42054, n42055 );
nand U89094 ( n42057, n41567, n655 );
nor U89095 ( n45356, n289, n45391 );
nand U89096 ( n13964, n14102, n14103 );
nor U89097 ( n14103, n14104, n14105 );
nor U89098 ( n14102, n14122, n14123 );
nand U89099 ( n14104, n14114, n14115 );
nand U89100 ( n2696, n38502, n38503 );
nor U89101 ( n38503, n38504, n38505 );
nor U89102 ( n38502, n38513, n38514 );
nand U89103 ( n38504, n38510, n38511 );
xor U89104 ( n38337, n39443, n1987 );
nor U89105 ( n40041, n38492, n38764 );
nor U89106 ( n63673, n48449, n76242 );
nor U89107 ( n71478, n1224, n71196 );
nor U89108 ( n44926, n289, n44561 );
nor U89109 ( n44208, n289, n43799 );
nor U89110 ( n72170, n1237, n71196 );
nand U89111 ( n66091, n66112, n66113 );
nand U89112 ( n66112, n66117, n66105 );
nand U89113 ( n66113, n66114, n652 );
nor U89114 ( n66117, n66026, n66118 );
nor U89115 ( n66114, n66020, n66115 );
nor U89116 ( n66115, n66026, n543 );
nand U89117 ( n39569, n38349, n76797 );
not U89118 ( n3149, n32936 );
nand U89119 ( n32925, n76773, n32093 );
nand U89120 ( n33050, n76773, n32160 );
nor U89121 ( n33059, n3160, n33061 );
nor U89122 ( n33061, n33055, n3145 );
not U89123 ( n3145, n33025 );
nand U89124 ( n12803, n76726, n11829 );
nor U89125 ( n71913, n1239, n71196 );
nor U89126 ( n37436, n37438, n37439 );
nand U89127 ( n37439, n37440, n37441 );
nand U89128 ( n37438, n37444, n37445 );
nand U89129 ( n37441, n1939, n37442 );
nor U89130 ( n40010, n37352, n40015 );
nand U89131 ( n40015, n40016, n37260 );
nand U89132 ( n40016, n40017, n40018 );
nand U89133 ( n40018, n1932, n38792 );
nand U89134 ( n1476, n54624, n54625 );
nor U89135 ( n54625, n54626, n54627 );
nor U89136 ( n54624, n54633, n54634 );
nand U89137 ( n54627, n54628, n54629 );
nor U89138 ( n37174, n2113, n76803 );
nand U89139 ( n38316, n38317, n76818 );
nand U89140 ( n65999, n66000, n66001 );
nand U89141 ( n66001, n54617, n76077 );
nand U89142 ( n66000, n54618, n827 );
nand U89143 ( n41669, n40727, n76378 );
nor U89144 ( n72038, n1238, n71196 );
not U89145 ( n737, n41297 );
nand U89146 ( n38948, n2128, n36925 );
nand U89147 ( n38949, n2122, n36551 );
nor U89148 ( n40120, n37273, n40162 );
nor U89149 ( n40162, n1904, n37274 );
nor U89150 ( n40115, n40116, n40117 );
nor U89151 ( n40116, n37368, n40121 );
nor U89152 ( n40117, n40118, n40119 );
nand U89153 ( n40121, n40122, n37268 );
nand U89154 ( n32037, n32038, n32039 );
nand U89155 ( n32039, n3059, n29405 );
nand U89156 ( n32038, n76777, n32041 );
not U89157 ( n730, n41284 );
buf U89158 ( n76252, n76251 );
nor U89159 ( n42044, n692, n42045 );
nor U89160 ( n11714, n76788, n76160 );
and U89161 ( n71230, n71302, n71303 );
not U89162 ( n2383, n18858 );
nand U89163 ( n36641, n36642, n36643 );
nand U89164 ( n36642, n76822, n36649 );
nand U89165 ( n36643, n76831, n36644 );
xnor U89166 ( n36644, n36645, n36646 );
xnor U89167 ( n36646, n36647, n36648 );
nand U89168 ( n3146, n36638, n36639 );
nor U89169 ( n36638, n36650, n36651 );
nor U89170 ( n36639, n36640, n36641 );
nand U89171 ( n36651, n36652, n36653 );
or U89172 ( n37440, n37260, n37443 );
nor U89173 ( n66016, n41949, n66027 );
nand U89174 ( n66027, n66028, n41578 );
nand U89175 ( n66028, n66029, n66030 );
nand U89176 ( n66030, n657, n61410 );
nand U89177 ( n66088, n66089, n66090 );
nand U89178 ( n66089, n784, n41054 );
nand U89179 ( n66090, n527, n827 );
not U89180 ( n2183, n36339 );
nand U89181 ( n46639, n76658, n45788 );
nand U89182 ( n67686, n76706, n66696 );
nand U89183 ( n25681, n76752, n24861 );
nand U89184 ( n58821, n76685, n57995 );
not U89185 ( n283, n48113 );
nor U89186 ( n66118, n66020, n66116 );
nand U89187 ( n37408, n37463, n37464 );
nor U89188 ( n37464, n37265, n37465 );
nor U89189 ( n37463, n37421, n37443 );
nand U89190 ( n37465, n37263, n37466 );
nand U89191 ( n41028, n41029, n41030 );
nand U89192 ( n41029, n584, n41036 );
nand U89193 ( n41030, n76851, n41031 );
xnor U89194 ( n41031, n41032, n41033 );
xnor U89195 ( n41033, n41034, n41035 );
nand U89196 ( n1921, n41025, n41026 );
nor U89197 ( n41025, n41037, n41038 );
nor U89198 ( n41026, n41027, n41028 );
nand U89199 ( n41038, n41039, n41040 );
nand U89200 ( n38533, n40146, n40147 );
nand U89201 ( n40147, n2074, n36589 );
nor U89202 ( n40146, n40148, n40149 );
nor U89203 ( n40149, n2000, n38524 );
not U89204 ( n699, n42042 );
xor U89205 ( n38369, n1975, n39572 );
nand U89206 ( n37460, n2187, n2128 );
or U89207 ( n71190, n1232, n71196 );
xnor U89208 ( n41952, n76388, n779 );
nor U89209 ( n40058, n37359, n40059 );
or U89210 ( n40059, n2034, n40014 );
nand U89211 ( n41941, n41942, n41943 );
nor U89212 ( n41943, n41944, n41945 );
nor U89213 ( n41942, n41950, n41951 );
nand U89214 ( n41944, n41949, n665 );
nand U89215 ( n33947, n34097, n34098 );
nor U89216 ( n34098, n34099, n34100 );
nor U89217 ( n34097, n34116, n34117 );
nand U89218 ( n34099, n34108, n34109 );
nand U89219 ( n37485, n37486, n37487 );
nand U89220 ( n37486, n2100, n37457 );
nand U89221 ( n37487, n37468, n37488 );
nand U89222 ( n2691, n38518, n38519 );
nor U89223 ( n38519, n38520, n38521 );
nor U89224 ( n38518, n38528, n38529 );
nand U89225 ( n38520, n38525, n38526 );
not U89226 ( n729, n41595 );
not U89227 ( n2179, n36702 );
nand U89228 ( n13915, n13994, n13995 );
nor U89229 ( n13995, n13997, n13998 );
nor U89230 ( n13994, n14024, n14025 );
nand U89231 ( n13997, n14012, n14013 );
not U89232 ( n2134, n37532 );
not U89233 ( n547, n64194 );
nor U89234 ( n48797, n63663, n64193 );
nor U89235 ( n64193, n802, n547 );
nor U89236 ( n40083, n1855, n38764 );
nand U89237 ( n46797, n76658, n45878 );
nand U89238 ( n67844, n76706, n66829 );
nand U89239 ( n25841, n76752, n24953 );
nand U89240 ( n58979, n76685, n58088 );
xnor U89241 ( n36743, n36916, n2040 );
nand U89242 ( n36916, n36917, n36918 );
nand U89243 ( n36917, n76827, n36339 );
nand U89244 ( n36918, n2113, n2035 );
nand U89245 ( n38348, n38349, n76818 );
and U89246 ( n38903, n38994, n39000 );
nand U89247 ( n48569, n48570, n568 );
nand U89248 ( n45363, n579, n54996 );
nand U89249 ( n54996, n54997, n41477 );
nand U89250 ( n54997, n54998, n618 );
nor U89251 ( n54998, n41458, n41479 );
nand U89252 ( n41477, n827, n838 );
nand U89253 ( n54923, n41463, n76857 );
xor U89254 ( n48684, n63663, n803 );
nand U89255 ( n38945, n2133, n36305 );
nand U89256 ( n46935, n76335, n1783 );
nand U89257 ( n54611, n54612, n54613 );
nand U89258 ( n54613, n76338, n40760 );
nand U89259 ( n54612, n76335, n1793 );
nand U89260 ( n49257, n76335, n1797 );
nand U89261 ( n48792, n76335, n1790 );
nand U89262 ( n46547, n76335, n1784 );
nand U89263 ( n48200, n76335, n1778 );
nand U89264 ( n47956, n76335, n1780 );
nand U89265 ( n48329, n76335, n1777 );
nand U89266 ( n49027, n76335, n1799 );
nand U89267 ( n54626, n54630, n54631 );
nand U89268 ( n54631, n76338, n41054 );
nand U89269 ( n54630, n76335, n1792 );
nand U89270 ( n54665, n54670, n54671 );
nand U89271 ( n54671, n76338, n40690 );
nand U89272 ( n54670, n76335, n1812 );
nor U89273 ( n66102, n66105, n66106 );
or U89274 ( n66106, n823, n66035 );
not U89275 ( n2119, n38904 );
nand U89276 ( n37433, n2188, n2133 );
nand U89277 ( n37413, n37504, n37385 );
nor U89278 ( n37504, n2140, n37390 );
not U89279 ( n2140, n37507 );
nand U89280 ( n37476, n2194, n2152 );
nand U89281 ( n37383, n37409, n37410 );
nor U89282 ( n37410, n37273, n1908 );
nor U89283 ( n37409, n37412, n37413 );
not U89284 ( n1908, n37411 );
and U89285 ( n37385, n37505, n37480 );
nor U89286 ( n37505, n37506, n2150 );
not U89287 ( n2150, n37476 );
nand U89288 ( n66363, n66435, n66436 );
nand U89289 ( n66436, n66205, n66207 );
nand U89290 ( n54678, n66284, n66285 );
nor U89291 ( n66284, n66296, n66297 );
nor U89292 ( n66285, n66286, n66287 );
nor U89293 ( n66297, n639, n61441 );
nand U89294 ( n11825, n11827, n11828 );
nand U89295 ( n11827, n4790, n8478 );
nand U89296 ( n11828, n76730, n11829 );
nand U89297 ( n32089, n32090, n32091 );
nand U89298 ( n32091, n3059, n29456 );
nand U89299 ( n32090, n76777, n32093 );
nand U89300 ( n46218, n76335, n1785 );
nand U89301 ( n45746, n76335, n1788 );
nand U89302 ( n37418, n37419, n37420 );
or U89303 ( n37419, n37268, n37408 );
nand U89304 ( n37391, n37414, n37415 );
nor U89305 ( n37414, n37416, n37407 );
nor U89306 ( n37416, n37417, n37418 );
nor U89307 ( n37417, n37421, n37422 );
not U89308 ( n743, n41090 );
nor U89309 ( n37171, n2117, n76803 );
xor U89310 ( n38400, n39694, n1967 );
nand U89311 ( n72395, n71396, n71312 );
nor U89312 ( n37390, n2190, n2145 );
not U89313 ( n2180, n36512 );
nor U89314 ( n32982, n3149, n32947 );
nand U89315 ( n32978, n76773, n32100 );
nor U89316 ( n40155, n40106, n40157 );
nor U89317 ( n40157, n40107, n40154 );
nand U89318 ( n40154, n40111, n40191 );
nand U89319 ( n40191, n40112, n40114 );
not U89320 ( n2123, n37595 );
buf U89321 ( n76418, n76417 );
nor U89322 ( n37506, n2192, n2148 );
nor U89323 ( n37493, n37499, n37500 );
nor U89324 ( n37499, n1974, n37501 );
not U89325 ( n2129, n37535 );
nor U89326 ( n33160, n32604, n32224 );
nand U89327 ( n37389, n2189, n2138 );
nor U89328 ( n37471, n37412, n37472 );
nand U89329 ( n33088, n76773, n32183 );
not U89330 ( n2510, n18206 );
nand U89331 ( n66281, n66294, n66291 );
nor U89332 ( n66294, n638, n66295 );
and U89333 ( n66295, n66198, n66293 );
nor U89334 ( n11548, n36, n11594 );
nand U89335 ( n12660, n14549, n14550 );
nor U89336 ( n14550, n14552, n14553 );
nor U89337 ( n14549, n14569, n14570 );
nand U89338 ( n14552, n14562, n14563 );
nor U89339 ( n42061, n40713, n76387 );
nor U89340 ( n42025, n41589, n41596 );
nor U89341 ( n42020, n729, n42022 );
nor U89342 ( n42022, n42023, n42024 );
nor U89343 ( n42023, n42025, n713 );
not U89344 ( n713, n41593 );
buf U89345 ( n76244, n61295 );
nor U89346 ( n49227, n48113, n49180 );
nor U89347 ( n48858, n48113, n48811 );
nor U89348 ( n48393, n48113, n48346 );
nor U89349 ( n48296, n48113, n48249 );
nor U89350 ( n48213, n48113, n48151 );
nand U89351 ( n66692, n66693, n66694 );
nand U89352 ( n66694, n5660, n63219 );
nand U89353 ( n66693, n76711, n66696 );
nand U89354 ( n24857, n24858, n24859 );
nand U89355 ( n24859, n3903, n22137 );
nand U89356 ( n24858, n76759, n24861 );
nand U89357 ( n57991, n57992, n57993 );
nand U89358 ( n57993, n6535, n55247 );
nand U89359 ( n57992, n76692, n57995 );
nor U89360 ( n37381, n37383, n37384 );
not U89361 ( n2182, n36747 );
xnor U89362 ( n54646, n66116, n41958 );
nand U89363 ( n54654, n66189, n66190 );
nor U89364 ( n66189, n66215, n66216 );
nor U89365 ( n66190, n66191, n66192 );
nor U89366 ( n66216, n648, n61441 );
nand U89367 ( n36366, n36367, n36368 );
nand U89368 ( n36367, n76821, n36381 );
nand U89369 ( n36368, n36369, n76830 );
nor U89370 ( n36369, n36370, n36371 );
nand U89371 ( n3206, n36363, n36364 );
nor U89372 ( n36363, n36382, n36383 );
nor U89373 ( n36364, n36365, n36366 );
nand U89374 ( n36383, n36384, n36385 );
nor U89375 ( n11224, n36, n10785 );
nand U89376 ( n72284, n71396, n71371 );
nor U89377 ( n10355, n36, n9897 );
nand U89378 ( n54762, n66358, n66359 );
nand U89379 ( n66359, n813, n41036 );
nor U89380 ( n66358, n66360, n66361 );
nor U89381 ( n66360, n823, n66364 );
nor U89382 ( n41582, n41591, n41592 );
nand U89383 ( n41592, n41593, n41594 );
nand U89384 ( n41591, n41595, n41596 );
nand U89385 ( n14410, n14588, n14589 );
nor U89386 ( n14589, n14590, n14592 );
nor U89387 ( n14588, n14612, n14613 );
nand U89388 ( n14590, n14602, n14603 );
nand U89389 ( n46835, n76658, n45891 );
nand U89390 ( n67882, n76706, n66842 );
nand U89391 ( n25879, n76752, n24966 );
nand U89392 ( n59017, n76685, n58101 );
not U89393 ( n7547, n46657 );
nand U89394 ( n40769, n40770, n40771 );
nand U89395 ( n40770, n584, n40784 );
nand U89396 ( n40771, n40772, n76850 );
nor U89397 ( n40772, n40773, n40774 );
nand U89398 ( n1981, n40766, n40767 );
nor U89399 ( n40766, n40785, n40786 );
nor U89400 ( n40767, n40768, n40769 );
nand U89401 ( n40786, n40787, n40788 );
xor U89402 ( n38412, n1959, n39765 );
nor U89403 ( n37163, n2122, n76803 );
nand U89404 ( n54616, n54617, n568 );
nand U89405 ( n54641, n54647, n54648 );
nand U89406 ( n54647, n76338, n40864 );
nand U89407 ( n54648, n54649, n568 );
nand U89408 ( n54864, n54869, n54870 );
nand U89409 ( n54869, n76338, n41036 );
nand U89410 ( n54870, n54871, n568 );
nand U89411 ( n54750, n54755, n54756 );
nand U89412 ( n54755, n76338, n41198 );
nand U89413 ( n54756, n54757, n568 );
buf U89414 ( n76410, n38757 );
not U89415 ( n4890, n12809 );
nor U89416 ( n66191, n41958, n66211 );
nand U89417 ( n66211, n66212, n41562 );
nand U89418 ( n66212, n66213, n66214 );
nand U89419 ( n66214, n643, n61410 );
nor U89420 ( n71065, n1218, n71247 );
xnor U89421 ( n36335, n36919, n2040 );
nand U89422 ( n36919, n36920, n36921 );
nand U89423 ( n36920, n76827, n36633 );
nand U89424 ( n36921, n2117, n2035 );
nand U89425 ( n32935, n32903, n32936 );
not U89426 ( n5760, n67704 );
not U89427 ( n4003, n25699 );
not U89428 ( n6635, n58839 );
not U89429 ( n1079, n71396 );
nor U89430 ( n45352, n284, n45391 );
not U89431 ( n545, n64783 );
nor U89432 ( n49140, n64343, n64782 );
nor U89433 ( n64782, n798, n545 );
nor U89434 ( n12902, n12904, n76596 );
nor U89435 ( n12904, n12905, n12907 );
nand U89436 ( n12905, n12932, n12933 );
nand U89437 ( n12907, n12908, n12909 );
not U89438 ( n750, n41134 );
not U89439 ( n2545, n18391 );
nand U89440 ( n36746, n36859, n36860 );
nand U89441 ( n36860, n76808, n36339 );
nand U89442 ( n36859, n2113, n76826 );
nor U89443 ( n42078, n42083, n41578 );
not U89444 ( n31, n14914 );
nor U89445 ( n44937, n284, n44561 );
nor U89446 ( n44251, n284, n43799 );
nand U89447 ( n37395, n37399, n37400 );
nand U89448 ( n37400, n2072, n37401 );
nor U89449 ( n37399, n37402, n37403 );
xor U89450 ( n49034, n64343, n799 );
nand U89451 ( n32897, n76773, n32053 );
nor U89452 ( n40134, n38524, n38764 );
xor U89453 ( n36549, n36922, n2040 );
nand U89454 ( n36922, n36923, n36924 );
nand U89455 ( n36923, n76827, n36925 );
nand U89456 ( n36924, n2128, n2035 );
not U89457 ( n1074, n72093 );
nand U89458 ( n38548, n40187, n40188 );
nand U89459 ( n40188, n2074, n36649 );
nor U89460 ( n40187, n40189, n40190 );
nor U89461 ( n40189, n2034, n40192 );
not U89462 ( n523, n54988 );
nand U89463 ( n37302, n37316, n37317 );
nor U89464 ( n37316, n37345, n37346 );
nor U89465 ( n37317, n37318, n37319 );
nand U89466 ( n37346, n37347, n37348 );
nand U89467 ( n46860, n76658, n45927 );
nand U89468 ( n67907, n76706, n66879 );
nand U89469 ( n25904, n76752, n25003 );
nand U89470 ( n59042, n76685, n58138 );
nor U89471 ( n40192, n40193, n40194 );
nor U89472 ( n40194, n37336, n37591 );
nor U89473 ( n40193, n1904, n40195 );
nor U89474 ( n40195, n37273, n37274 );
nand U89475 ( n2686, n38534, n38535 );
nor U89476 ( n38535, n38536, n38537 );
nor U89477 ( n38534, n38544, n38545 );
nand U89478 ( n38536, n38541, n38542 );
nand U89479 ( n66174, n66175, n66176 );
nand U89480 ( n66176, n54649, n76076 );
nand U89481 ( n66175, n54646, n827 );
not U89482 ( n1983, n37453 );
not U89483 ( n2694, n17039 );
nor U89484 ( n71642, n1235, n71171 );
nand U89485 ( n36439, n2025, n36841 );
not U89486 ( n2025, n36630 );
nand U89487 ( n38835, n2138, n36442 );
not U89488 ( n277, n48102 );
xor U89489 ( n49616, n49617, n49618 );
nor U89490 ( n65938, n65348, n65824 );
nor U89491 ( n64515, n64382, n64386 );
nor U89492 ( n64784, n64387, n64514 );
nand U89493 ( n13013, n76725, n11982 );
nand U89494 ( n36776, n36777, n1848 );
xor U89495 ( n36777, n36779, n36780 );
nor U89496 ( n66364, n66365, n66366 );
nor U89497 ( n66365, n66367, n66368 );
nor U89498 ( n66366, n41938, n565 );
and U89499 ( n66368, n42087, n42084 );
not U89500 ( n645, n41562 );
nor U89501 ( n41939, n65343, n65347 );
nand U89502 ( n41159, n41160, n522 );
xor U89503 ( n41160, n41162, n41163 );
not U89504 ( n669, n64814 );
not U89505 ( n1852, n38602 );
nor U89506 ( n71780, n71196, n1222 );
not U89507 ( n694, n41535 );
xor U89508 ( n38444, n1947, n39866 );
nand U89509 ( n12963, n76726, n11952 );
nand U89510 ( n33126, n76773, n32196 );
nand U89511 ( n39938, n39891, n39893 );
nand U89512 ( n39829, n39749, n39792 );
nand U89513 ( n36840, n36926, n36927 );
nand U89514 ( n36927, n76807, n36925 );
nand U89515 ( n36926, n2128, n76826 );
nand U89516 ( n38563, n40222, n40223 );
nand U89517 ( n40223, n2074, n36381 );
nor U89518 ( n40222, n40224, n40225 );
nor U89519 ( n40224, n2034, n40232 );
not U89520 ( n745, n40913 );
nor U89521 ( n37160, n2128, n76803 );
or U89522 ( n41958, n66020, n66026 );
nand U89523 ( n40173, n40174, n40175 );
nand U89524 ( n40175, n38543, n76797 );
nand U89525 ( n40174, n2033, n38540 );
nand U89526 ( n36632, n2021, n36630 );
nor U89527 ( n36838, n36928, n36929 );
nand U89528 ( n2681, n38549, n38550 );
nor U89529 ( n38550, n38551, n38552 );
nor U89530 ( n38549, n38558, n38559 );
nand U89531 ( n38551, n38556, n38557 );
xor U89532 ( n36684, n37758, n36485 );
xor U89533 ( n37758, n36481, n1849 );
nand U89534 ( n41924, n63312, n63307 );
nand U89535 ( n54821, n66431, n66432 );
nand U89536 ( n66432, n813, n40784 );
nor U89537 ( n66431, n66433, n66434 );
nor U89538 ( n66433, n823, n66437 );
or U89539 ( n72176, n1237, n71171 );
nor U89540 ( n37369, n40106, n40103 );
nor U89541 ( n71484, n1234, n71171 );
nand U89542 ( n41932, n62781, n62832 );
nor U89543 ( n15779, n14914, n15712 );
nor U89544 ( n15248, n14914, n15180 );
nor U89545 ( n15138, n14914, n15073 );
nor U89546 ( n15028, n14914, n14969 );
nor U89547 ( n16195, n14914, n16130 );
nor U89548 ( n38834, n2143, n38773 );
not U89549 ( n2143, n38771 );
nor U89550 ( n39521, n37360, n39495 );
nand U89551 ( n37330, n40229, n40226 );
not U89552 ( n544, n65925 );
nor U89553 ( n49572, n65317, n65924 );
nor U89554 ( n65924, n794, n544 );
nand U89555 ( n37329, n40114, n40111 );
nand U89556 ( n36338, n36854, n36855 );
nand U89557 ( n36855, n76808, n36633 );
nand U89558 ( n36854, n2117, n76826 );
nand U89559 ( n37352, n39901, n39899 );
nand U89560 ( n45924, n45925, n45926 );
nand U89561 ( n45925, n42863, n45841 );
nand U89562 ( n45926, n45927, n76662 );
xor U89563 ( n40878, n40879, n40880 );
nand U89564 ( n37338, n39322, n39346 );
nand U89565 ( n37447, n37456, n37457 );
nand U89566 ( n36435, n36929, n36928 );
nand U89567 ( n36841, n36849, n36850 );
nand U89568 ( n36850, n76808, n36551 );
nand U89569 ( n36849, n2122, n76826 );
nand U89570 ( n66875, n66876, n66877 );
nand U89571 ( n66877, n63515, n66792 );
nand U89572 ( n66876, n66879, n76710 );
nand U89573 ( n24999, n25000, n25001 );
nand U89574 ( n25001, n22295, n24914 );
nand U89575 ( n25000, n25003, n76758 );
nand U89576 ( n58134, n58135, n58136 );
nand U89577 ( n58136, n55407, n58051 );
nand U89578 ( n58135, n58138, n76691 );
nand U89579 ( n41923, n66207, n66435 );
nand U89580 ( n54876, n66735, n66736 );
nor U89581 ( n66735, n66748, n66749 );
nor U89582 ( n66736, n66737, n66738 );
nor U89583 ( n66749, n623, n61441 );
nor U89584 ( n61175, n76066, n76387 );
nor U89585 ( n13249, n13284, n13285 );
nor U89586 ( n13285, n13248, n76603 );
nand U89587 ( n41925, n62680, n62687 );
nor U89588 ( n71195, n71196, n1230 );
nor U89589 ( n37152, n2133, n76803 );
nor U89590 ( n40232, n40233, n40234 );
nor U89591 ( n40233, n37329, n40236 );
nor U89592 ( n40234, n40198, n40235 );
nand U89593 ( n40236, n40237, n37472 );
nand U89594 ( n37374, n39612, n39609 );
nand U89595 ( n38578, n40265, n40266 );
nor U89596 ( n40265, n40280, n40281 );
nor U89597 ( n40266, n40267, n40268 );
nor U89598 ( n40281, n2157, n38822 );
and U89599 ( n40275, n40230, n40231 );
xor U89600 ( n49380, n65317, n795 );
not U89601 ( n2184, n36633 );
nor U89602 ( n72054, n1238, n71171 );
nand U89603 ( n37356, n39744, n39748 );
or U89604 ( n37368, n1929, n40029 );
not U89605 ( n4889, n13127 );
nand U89606 ( n13113, n76725, n12047 );
nand U89607 ( n39791, n39749, n37356 );
nand U89608 ( n37337, n39738, n39747 );
nand U89609 ( n37372, n40230, n40283 );
nor U89610 ( n41988, n629, n41990 );
nand U89611 ( n41957, n64025, n64022 );
nor U89612 ( n49219, n48102, n49180 );
nor U89613 ( n48850, n48102, n48811 );
nor U89614 ( n48385, n48102, n48346 );
nor U89615 ( n48288, n48102, n48249 );
nor U89616 ( n48190, n48102, n48151 );
nand U89617 ( n37324, n39255, n39256 );
not U89618 ( n640, n66198 );
nand U89619 ( n37367, n39420, n39417 );
nand U89620 ( n36928, n36930, n36931 );
nand U89621 ( n36931, n76807, n36305 );
nand U89622 ( n36930, n2133, n76826 );
nand U89623 ( n37343, n39000, n38945 );
nand U89624 ( n38985, n38992, n38993 );
nand U89625 ( n38993, n2127, n2125 );
or U89626 ( n38992, n38994, n2130 );
nand U89627 ( n37355, n39896, n39943 );
nor U89628 ( n11543, n32, n11594 );
nand U89629 ( n37397, n1893, n37288 );
not U89630 ( n652, n66105 );
nand U89631 ( n41962, n66750, n66753 );
nand U89632 ( n41963, n64233, n64230 );
not U89633 ( n647, n66291 );
nand U89634 ( n37342, n38994, n38948 );
nand U89635 ( n37373, n39669, n39666 );
not U89636 ( n1929, n40026 );
nor U89637 ( n13289, n4898, n13292 );
nor U89638 ( n13292, n13284, n4886 );
not U89639 ( n4886, n13248 );
nand U89640 ( n13278, n76725, n12135 );
nor U89641 ( n11238, n32, n10785 );
nor U89642 ( n10409, n32, n9897 );
nand U89643 ( n37341, n38904, n38949 );
not U89644 ( n2382, n18874 );
nand U89645 ( n37331, n38838, n38835 );
nand U89646 ( n37326, n39135, n39132 );
not U89647 ( n712, n63695 );
and U89648 ( n39786, n39737, n39748 );
nand U89649 ( n36480, n36485, n1849 );
nand U89650 ( n36476, n2009, n36477 );
not U89651 ( n2009, n36482 );
nand U89652 ( n36477, n36478, n36479 );
nand U89653 ( n36479, n36480, n36481 );
nor U89654 ( n45348, n278, n45391 );
xor U89655 ( n38480, n1937, n39965 );
or U89656 ( n36478, n36485, n1849 );
nand U89657 ( n39347, n39322, n37344 );
nand U89658 ( n37344, n39319, n39321 );
nand U89659 ( n39524, n37360, n39491 );
not U89660 ( n754, n40747 );
buf U89661 ( n76250, n76247 );
nand U89662 ( n37325, n39184, n39181 );
nor U89663 ( n37521, n2152, n2194 );
nor U89664 ( n37528, n37599, n37479 );
or U89665 ( n37599, n37520, n37521 );
nor U89666 ( n40211, n38555, n38764 );
or U89667 ( n71167, n1223, n71171 );
xor U89668 ( n38500, n1889, n1933 );
not U89669 ( n1889, n39999 );
nor U89670 ( n44946, n278, n44561 );
nor U89671 ( n44295, n278, n43799 );
nor U89672 ( n42201, n41968, n45272 );
and U89673 ( n45272, n45273, n76389 );
nand U89674 ( n45273, n830, n818 );
nand U89675 ( n45202, n45268, n45269 );
or U89676 ( n45268, n41490, n42201 );
nand U89677 ( n45269, n579, n587 );
not U89678 ( n26, n14900 );
xor U89679 ( n16637, n16638, n16639 );
nor U89680 ( n71068, n1218, n1100 );
nand U89681 ( n46909, n76658, n45935 );
nand U89682 ( n67956, n76706, n66886 );
nand U89683 ( n25953, n76752, n25010 );
nand U89684 ( n59091, n76685, n58145 );
nor U89685 ( n37133, n2148, n76804 );
nor U89686 ( n37141, n37134, n37294 );
nor U89687 ( n37294, n37295, n37133 );
nor U89688 ( n37289, n37143, n37293 );
nand U89689 ( n37293, n37141, n36429 );
nand U89690 ( n42193, n812, n45202 );
nand U89691 ( n63668, n712, n63312 );
nand U89692 ( n40086, n38512, n76797 );
nor U89693 ( n64001, n42049, n702 );
nand U89694 ( n37134, n37296, n37138 );
nand U89695 ( n37296, n37137, n37136 );
nand U89696 ( n37292, n2152, n37297 );
not U89697 ( n2057, n39322 );
nand U89698 ( n63670, n63695, n63307 );
nand U89699 ( n37387, n2190, n2145 );
nand U89700 ( n37129, n37130, n37131 );
nand U89701 ( n37130, n37135, n2067 );
nand U89702 ( n37131, n37132, n37133 );
not U89703 ( n2067, n37136 );
nand U89704 ( n66738, n66739, n66740 );
nand U89705 ( n66740, n66741, n66742 );
nand U89706 ( n66739, n66743, n524 );
nand U89707 ( n66742, n42001, n41989 );
nand U89708 ( n3136, n36673, n36674 );
nor U89709 ( n36674, n36675, n36676 );
nor U89710 ( n36673, n36682, n36683 );
nor U89711 ( n36676, n2157, n76454 );
nand U89712 ( n40252, n40253, n40254 );
nand U89713 ( n40254, n38573, n76797 );
nand U89714 ( n40253, n2033, n38570 );
xor U89715 ( n36608, n36611, n36612 );
xor U89716 ( n36376, n36379, n36380 );
nand U89717 ( n40268, n40269, n40270 );
nand U89718 ( n40270, n40271, n40272 );
nand U89719 ( n40269, n40274, n40275 );
nand U89720 ( n40272, n37411, n37472 );
nor U89721 ( n36415, n36301, n36303 );
not U89722 ( n2185, n36551 );
buf U89723 ( n76416, n76413 );
not U89724 ( n270, n48091 );
not U89725 ( n1942, n39896 );
nor U89726 ( n37135, n37137, n2068 );
not U89727 ( n2068, n37138 );
nand U89728 ( n37478, n37479, n37480 );
nand U89729 ( n37694, n2197, n38039 );
nand U89730 ( n37745, n37603, n38101 );
nand U89731 ( n38101, n38102, n76457 );
nand U89732 ( n38102, n2082, n2198 );
nand U89733 ( n54924, n67006, n67007 );
nand U89734 ( n67007, n813, n42184 );
nor U89735 ( n67006, n67008, n67009 );
nor U89736 ( n67009, n823, n67010 );
xor U89737 ( n54637, n66004, n792 );
and U89738 ( n36417, n36301, n36303 );
nor U89739 ( n71929, n1239, n71171 );
nand U89740 ( n38593, n40306, n40307 );
nand U89741 ( n40307, n2074, n37288 );
nor U89742 ( n40306, n40308, n40309 );
nor U89743 ( n40308, n2034, n40310 );
nand U89744 ( n38719, n40293, n40294 );
nor U89745 ( n40294, n40295, n40296 );
nor U89746 ( n40293, n40305, n38593 );
and U89747 ( n40295, n38592, n76797 );
not U89748 ( n2093, n40402 );
nand U89749 ( n38109, n37094, n76811 );
nand U89750 ( n40444, n2094, n2199 );
not U89751 ( n2092, n38729 );
nand U89752 ( n38511, n38512, n76819 );
nand U89753 ( n38542, n38543, n76819 );
not U89754 ( n2030, n38119 );
not U89755 ( n732, n62781 );
nand U89756 ( n38566, n38571, n38572 );
nand U89757 ( n38571, n76438, n36649 );
nand U89758 ( n38572, n38573, n76818 );
nor U89759 ( n37148, n2138, n76803 );
nand U89760 ( n38589, n38590, n38591 );
nand U89761 ( n38590, n76814, n38593 );
nand U89762 ( n38591, n76819, n38592 );
nor U89763 ( n13193, n4889, n13140 );
nand U89764 ( n13188, n76725, n12055 );
nand U89765 ( n38225, n76815, n2117 );
nand U89766 ( n38257, n76815, n2107 );
xor U89767 ( n41001, n41004, n41005 );
nand U89768 ( n37477, n2193, n2149 );
xnor U89769 ( n40310, n37372, n37401 );
not U89770 ( n2147, n37361 );
nand U89771 ( n38766, n38820, n38821 );
nand U89772 ( n38821, n38773, n37361 );
nand U89773 ( n38820, n2143, n2147 );
xor U89774 ( n38532, n1925, n40089 );
nand U89775 ( n42194, n814, n45202 );
nand U89776 ( n45066, n45067, n45068 );
nand U89777 ( n45068, n45069, n577 );
nand U89778 ( n45067, n45078, n575 );
nor U89779 ( n45069, n45070, n45071 );
nand U89780 ( n42667, n42668, n42669 );
nand U89781 ( n42669, n42670, n577 );
nand U89782 ( n42668, n42679, n575 );
nor U89783 ( n42670, n42671, n42672 );
nand U89784 ( n42328, n42329, n42330 );
nand U89785 ( n42330, n42331, n577 );
nand U89786 ( n42329, n42345, n575 );
nor U89787 ( n42331, n42332, n42333 );
nand U89788 ( n37518, n37519, n37506 );
nor U89789 ( n37519, n37520, n37521 );
nand U89790 ( n45135, n45136, n45137 );
nand U89791 ( n45137, n577, n45138 );
nand U89792 ( n45136, n575, n45203 );
xor U89793 ( n45138, n45139, n45140 );
nand U89794 ( n44386, n44387, n44388 );
nand U89795 ( n44388, n577, n44389 );
nand U89796 ( n44387, n575, n44392 );
xor U89797 ( n44389, n44390, n44391 );
nand U89798 ( n42415, n42416, n42417 );
nand U89799 ( n42417, n577, n42418 );
nand U89800 ( n42416, n575, n42426 );
nand U89801 ( n42418, n42419, n42420 );
nand U89802 ( n42240, n42241, n42242 );
nand U89803 ( n42242, n577, n42243 );
nand U89804 ( n42241, n575, n42253 );
nand U89805 ( n42243, n42244, n42245 );
and U89806 ( n41070, n41071, n76850 );
nor U89807 ( n13414, n12887, n12215 );
xor U89808 ( n40779, n40782, n40783 );
not U89809 ( n759, n41024 );
xor U89810 ( n36414, n36419, n36420 );
nor U89811 ( n36420, n36421, n36422 );
xor U89812 ( n36419, n36426, n2040 );
nor U89813 ( n36422, n2190, n36423 );
nand U89814 ( n36426, n36427, n36428 );
nand U89815 ( n36428, n76808, n36429 );
nand U89816 ( n36427, n2145, n76826 );
xor U89817 ( n54677, n789, n66179 );
nand U89818 ( n13324, n76725, n12164 );
nor U89819 ( n16185, n14900, n16130 );
nor U89820 ( n15769, n14900, n15712 );
nor U89821 ( n15238, n14900, n15180 );
nor U89822 ( n15128, n14900, n15073 );
nor U89823 ( n15018, n14900, n14969 );
nand U89824 ( n45932, n45933, n45934 );
nand U89825 ( n45933, n7434, n7950 );
nand U89826 ( n45934, n76662, n45935 );
nand U89827 ( n66883, n66884, n66885 );
nand U89828 ( n66884, n5660, n6163 );
nand U89829 ( n66885, n76710, n66886 );
nand U89830 ( n25007, n25008, n25009 );
nand U89831 ( n25008, n3903, n4385 );
nand U89832 ( n25009, n76758, n25010 );
nand U89833 ( n58142, n58143, n58144 );
nand U89834 ( n58143, n6535, n7018 );
nand U89835 ( n58144, n76691, n58145 );
nand U89836 ( n36303, n36440, n36441 );
nand U89837 ( n36441, n76808, n36442 );
nand U89838 ( n36440, n2138, n76826 );
nand U89839 ( n49258, n76338, n41114 );
nand U89840 ( n46936, n76339, n41024 );
nand U89841 ( n48793, n76339, n41006 );
nand U89842 ( n48448, n76339, n41284 );
nand U89843 ( n47957, n76339, n41134 );
nand U89844 ( n46548, n76339, n40950 );
nand U89845 ( n48201, n76339, n41090 );
or U89846 ( n38772, n37361, n38773 );
nand U89847 ( n49028, n76339, n41329 );
nand U89848 ( n48910, n76339, n40967 );
xnor U89849 ( n67010, n41962, n42011 );
nand U89850 ( n48330, n76339, n41297 );
nand U89851 ( n48678, n76339, n41178 );
nand U89852 ( n66346, n54757, n76075 );
nand U89853 ( n48568, n76339, n40801 );
nand U89854 ( n49570, n76338, n41145 );
nand U89855 ( n49138, n76338, n40727 );
not U89856 ( n1052, n72189 );
nor U89857 ( n43849, n865, n42193 );
nor U89858 ( n43659, n864, n42193 );
nor U89859 ( n43552, n882, n42193 );
nor U89860 ( n45134, n847, n42193 );
nor U89861 ( n44999, n849, n42193 );
nor U89862 ( n44385, n859, n42193 );
nor U89863 ( n43424, n880, n42193 );
nor U89864 ( n43223, n888, n42193 );
nor U89865 ( n42950, n887, n42193 );
nor U89866 ( n42414, n893, n42193 );
nor U89867 ( n42239, n915, n42193 );
nor U89868 ( n42204, n917, n42193 );
nand U89869 ( n47077, n76657, n46050 );
nand U89870 ( n68108, n76705, n66990 );
nand U89871 ( n26105, n76751, n25114 );
nand U89872 ( n59246, n76684, n58252 );
nand U89873 ( n46219, n76340, n40834 );
xor U89874 ( n36482, n36486, n36487 );
nand U89875 ( n45747, n76340, n40852 );
not U89876 ( n2070, n38601 );
nand U89877 ( n40296, n40297, n40298 );
nand U89878 ( n40297, n2073, n36381 );
nand U89879 ( n40298, n2033, n38585 );
nand U89880 ( n37700, n37701, n37702 );
nand U89881 ( n37702, n37703, n2079 );
nand U89882 ( n37701, n37707, n2078 );
xnor U89883 ( n37703, n37704, n37705 );
not U89884 ( n2188, n36305 );
not U89885 ( n7529, n46958 );
nand U89886 ( n45824, n46745, n7907 );
nand U89887 ( n45910, n46894, n7900 );
nand U89888 ( n45617, n45688, n7917 );
not U89889 ( n7594, n47445 );
not U89890 ( n7528, n46597 );
not U89891 ( n7527, n46540 );
nor U89892 ( n46399, n46411, n46412 );
nor U89893 ( n46411, n46415, n46416 );
nor U89894 ( n46412, n46413, n46414 );
or U89895 ( n46416, n45597, n45596 );
or U89896 ( n46414, n45600, n45599 );
not U89897 ( n2187, n36925 );
nor U89898 ( n11538, n27, n11594 );
nand U89899 ( n37689, n2153, n38039 );
xor U89900 ( n38562, n40178, n1913 );
nor U89901 ( n40328, n1852, n38764 );
nand U89902 ( n38726, n40318, n40319 );
nor U89903 ( n40319, n38609, n40320 );
nor U89904 ( n40318, n40328, n40329 );
nor U89905 ( n40320, n1893, n40321 );
nor U89906 ( n49211, n48091, n49180 );
nor U89907 ( n48842, n48091, n48811 );
nor U89908 ( n48377, n48091, n48346 );
nor U89909 ( n48280, n48091, n48249 );
nor U89910 ( n48182, n48091, n48151 );
nand U89911 ( n39005, n37433, n37532 );
xor U89912 ( n54820, n66349, n787 );
nor U89913 ( n11255, n27, n10785 );
nor U89914 ( n10464, n27, n9897 );
nand U89915 ( n13125, n13085, n13127 );
nand U89916 ( n12052, n12053, n12054 );
nand U89917 ( n12053, n4790, n5300 );
nand U89918 ( n12054, n76729, n12055 );
buf U89919 ( n76383, n75705 );
nor U89920 ( n71828, n1239, n1057 );
nand U89921 ( n41631, n41297, n76379 );
nand U89922 ( n71957, n71307, n71357 );
nand U89923 ( n13078, n76725, n11997 );
nand U89924 ( n66724, n54871, n76074 );
nand U89925 ( n54995, n67219, n67220 );
nand U89926 ( n67220, n67221, n61410 );
nand U89927 ( n67219, n54988, n61439 );
nand U89928 ( n67221, n42011, n67225 );
and U89929 ( n38609, n38602, n40323 );
nand U89930 ( n40323, n2034, n2000 );
nor U89931 ( n71506, n1218, n71196 );
nor U89932 ( n45344, n272, n45391 );
nor U89933 ( n42265, n42304, n42194 );
nor U89934 ( n42304, n42305, n42306 );
nor U89935 ( n42305, n42310, n42311 );
nor U89936 ( n42306, n910, n42307 );
not U89937 ( n764, n40950 );
not U89938 ( n1057, n71307 );
nor U89939 ( n71796, n71171, n1222 );
nor U89940 ( n44309, n272, n43799 );
nor U89941 ( n44956, n272, n44561 );
not U89942 ( n3142, n33238 );
nand U89943 ( n32129, n33037, n3503 );
nand U89944 ( n32218, n33185, n3497 );
nand U89945 ( n31939, n32009, n3514 );
nand U89946 ( n32024, n32882, n3509 );
not U89947 ( n3208, n33710 );
nor U89948 ( n32698, n32710, n32711 );
nor U89949 ( n32710, n32714, n32715 );
nor U89950 ( n32711, n32712, n32713 );
or U89951 ( n32715, n31899, n31898 );
or U89952 ( n32713, n31902, n31901 );
not U89953 ( n21, n14887 );
nand U89954 ( n46046, n46047, n46048 );
nand U89955 ( n46048, n7434, n43031 );
nand U89956 ( n46047, n76662, n46050 );
nand U89957 ( n66986, n66987, n66988 );
nand U89958 ( n66988, n5660, n63730 );
nand U89959 ( n66987, n76710, n66990 );
nand U89960 ( n25110, n25111, n25112 );
nand U89961 ( n25112, n3903, n22449 );
nand U89962 ( n25111, n76758, n25114 );
nand U89963 ( n58248, n58249, n58250 );
nand U89964 ( n58250, n6535, n55564 );
nand U89965 ( n58249, n76691, n58252 );
not U89966 ( n5743, n67993 );
not U89967 ( n3985, n25990 );
not U89968 ( n6618, n59128 );
nand U89969 ( n66775, n67792, n6118 );
nand U89970 ( n24897, n25789, n4340 );
nand U89971 ( n58034, n58927, n6973 );
nand U89972 ( n66861, n67941, n6112 );
nand U89973 ( n24985, n25938, n4334 );
nand U89974 ( n58120, n59076, n6967 );
nand U89975 ( n66542, n66612, n6129 );
nand U89976 ( n66627, n67643, n6124 );
nand U89977 ( n24707, n24777, n4352 );
nand U89978 ( n24792, n25638, n4347 );
nand U89979 ( n57841, n57911, n6984 );
nand U89980 ( n57926, n58775, n6979 );
not U89981 ( n5807, n68466 );
not U89982 ( n4040, n26465 );
not U89983 ( n6673, n59604 );
nor U89984 ( n67463, n67475, n67476 );
nor U89985 ( n67475, n67479, n67480 );
nor U89986 ( n67476, n67477, n67478 );
or U89987 ( n67480, n66522, n66521 );
nor U89988 ( n25458, n25470, n25471 );
nor U89989 ( n25470, n25474, n25475 );
nor U89990 ( n25471, n25472, n25473 );
or U89991 ( n25475, n24687, n24686 );
nor U89992 ( n58595, n58607, n58608 );
nor U89993 ( n58607, n58611, n58612 );
nor U89994 ( n58608, n58609, n58610 );
or U89995 ( n58612, n57821, n57820 );
or U89996 ( n67478, n66525, n66524 );
or U89997 ( n25473, n24690, n24689 );
or U89998 ( n58610, n57824, n57823 );
not U89999 ( n2192, n37295 );
not U90000 ( n619, n67261 );
nand U90001 ( n70967, n620, n817 );
xor U90002 ( n54922, n785, n552 );
not U90003 ( n2190, n36429 );
not U90004 ( n2189, n36442 );
not U90005 ( n775, n40713 );
not U90006 ( n3153, n33320 );
nand U90007 ( n33351, n76772, n32351 );
nand U90008 ( n67225, n552, n42184 );
not U90009 ( n7559, n46955 );
nand U90010 ( n45921, n7900, n46897 );
nand U90011 ( n45821, n7907, n46748 );
nand U90012 ( n45614, n7917, n45685 );
not U90013 ( n7557, n46542 );
not U90014 ( n7558, n46600 );
not U90015 ( n7560, n47108 );
nand U90016 ( n47540, n47596, n47617 );
nor U90017 ( n37920, n1972, n37689 );
nor U90018 ( n37862, n1950, n37689 );
nor U90019 ( n37806, n1930, n37689 );
nand U90020 ( n33240, n76773, n32272 );
not U90021 ( n2045, n38866 );
nand U90022 ( n36843, n37075, n2087 );
nor U90023 ( n37075, n37076, n36943 );
nor U90024 ( n71072, n1218, n1079 );
nand U90025 ( n37108, n40446, n2198 );
nor U90026 ( n40446, n76039, n2088 );
not U90027 ( n264, n48066 );
xor U90028 ( n49541, n49543, n49544 );
not U90029 ( n4884, n13512 );
nand U90030 ( n12208, n13445, n5247 );
nand U90031 ( n12092, n13263, n5253 );
not U90032 ( n4940, n14097 );
not U90033 ( n4883, n13059 );
not U90034 ( n4882, n12800 );
nand U90035 ( n12694, n76727, n11780 );
nor U90036 ( n47340, n47336, n47337 );
nand U90037 ( n45578, n45593, n45594 );
nand U90038 ( n45594, n45595, n76346 );
nand U90039 ( n45593, n45598, n76670 );
nor U90040 ( n45595, n45596, n45597 );
nor U90041 ( n45598, n45599, n45600 );
xor U90042 ( MUL_1411_U13, n71508, n71509 );
xor U90043 ( n71508, n71510, n71511 );
nor U90044 ( n16175, n14887, n16130 );
nor U90045 ( n15759, n14887, n15712 );
nor U90046 ( n15228, n14887, n15180 );
nor U90047 ( n15118, n14887, n15073 );
nor U90048 ( n15008, n14887, n14969 );
nor U90049 ( n39525, n1987, n76407 );
nor U90050 ( n67214, n552, n67216 );
and U90051 ( n67216, n76071, n834 );
nor U90052 ( n39643, n1975, n76407 );
not U90053 ( n4881, n12859 );
nor U90054 ( n39394, n2054, n76406 );
nor U90055 ( n40264, n1909, n76407 );
nor U90056 ( n40145, n1925, n76406 );
nor U90057 ( n40305, n2098, n76407 );
nor U90058 ( n40186, n1919, n76406 );
nor U90059 ( n40221, n1913, n76407 );
nor U90060 ( n39774, n1967, n76407 );
not U90061 ( n768, n40834 );
nor U90062 ( n39582, n1982, n76407 );
nor U90063 ( n39830, n1959, n76407 );
nor U90064 ( n40007, n1937, n76407 );
nor U90065 ( n39932, n1947, n76407 );
nand U90066 ( n32347, n32348, n32349 );
nand U90067 ( n32349, n3059, n29770 );
nand U90068 ( n32348, n76776, n32351 );
nand U90069 ( n71654, n71357, n71313 );
nor U90070 ( n39452, n1994, n76406 );
not U90071 ( n779, n40852 );
not U90072 ( n3173, n33235 );
nand U90073 ( n32126, n3503, n33040 );
nand U90074 ( n32215, n3497, n33188 );
nand U90075 ( n31936, n3514, n32006 );
nand U90076 ( n32034, n3509, n32885 );
not U90077 ( n3174, n33387 );
nand U90078 ( n33805, n33861, n33882 );
nor U90079 ( n39874, n1953, n76407 );
nor U90080 ( n40054, n1933, n76407 );
not U90081 ( n7592, n47539 );
not U90082 ( n5772, n67990 );
not U90083 ( n4013, n25987 );
not U90084 ( n6645, n59125 );
nand U90085 ( n66872, n6112, n67944 );
nand U90086 ( n24996, n4334, n25941 );
nand U90087 ( n58131, n6967, n59079 );
nand U90088 ( n66772, n6118, n67795 );
nand U90089 ( n24894, n4340, n25792 );
nand U90090 ( n58031, n6973, n58930 );
nand U90091 ( n24704, n4352, n24774 );
nand U90092 ( n66539, n6129, n66609 );
nand U90093 ( n57838, n6984, n57908 );
nand U90094 ( n66637, n6124, n67646 );
nand U90095 ( n24802, n4347, n25641 );
nand U90096 ( n57936, n6979, n58778 );
not U90097 ( n5773, n68139 );
not U90098 ( n4014, n26136 );
not U90099 ( n6647, n59277 );
nand U90100 ( n68561, n68617, n68638 );
nand U90101 ( n26560, n26616, n26637 );
nand U90102 ( n59702, n59758, n59779 );
nor U90103 ( n39973, n1940, n76407 );
nor U90104 ( n39703, n1969, n76407 );
nor U90105 ( n66099, n792, n76072 );
nor U90106 ( n40098, n1928, n76407 );
nor U90107 ( n32826, n32834, n32835 );
nor U90108 ( n32834, n32714, n32837 );
nor U90109 ( n32835, n32712, n32836 );
or U90110 ( n32837, n32007, n32006 );
or U90111 ( n32836, n32010, n32009 );
nor U90112 ( n64501, n799, n76068 );
nor U90113 ( n65809, n795, n76073 );
nor U90114 ( n67591, n67599, n67600 );
nor U90115 ( n67599, n67479, n67602 );
nor U90116 ( n67600, n67477, n67601 );
or U90117 ( n67602, n66610, n66609 );
nor U90118 ( n25586, n25594, n25595 );
nor U90119 ( n25594, n25474, n25597 );
nor U90120 ( n25595, n25472, n25596 );
or U90121 ( n25597, n24775, n24774 );
nor U90122 ( n58723, n58731, n58732 );
nor U90123 ( n58731, n58611, n58734 );
nor U90124 ( n58732, n58609, n58733 );
or U90125 ( n58734, n57909, n57908 );
or U90126 ( n67601, n66613, n66612 );
or U90127 ( n25596, n24778, n24777 );
or U90128 ( n58733, n57912, n57911 );
nor U90129 ( n11533, n22, n11594 );
nor U90130 ( n64792, n798, n76068 );
nor U90131 ( n65326, n797, n76066 );
nor U90132 ( n65933, n794, n76072 );
nor U90133 ( n64202, n802, n76073 );
nor U90134 ( n66283, n789, n76066 );
nor U90135 ( n62948, n807, n76069 );
nor U90136 ( n63678, n804, n76067 );
nor U90137 ( n63270, n805, n76068 );
nor U90138 ( n66188, n790, n76067 );
nor U90139 ( n66013, n793, n76070 );
nor U90140 ( n63993, n803, n76071 );
nor U90141 ( n66430, n787, n76071 );
nor U90142 ( n10482, n22, n9897 );
nor U90143 ( n67005, n785, n76069 );
nor U90144 ( n64352, n800, n76069 );
nor U90145 ( n66734, n786, n76070 );
nor U90146 ( n36682, n1893, n36492 );
nor U90147 ( n11268, n22, n10785 );
nor U90148 ( n48834, n48066, n48811 );
nor U90149 ( n48369, n48066, n48346 );
nor U90150 ( n48272, n48066, n48249 );
nor U90151 ( n48174, n48066, n48151 );
nor U90152 ( n49203, n48066, n49180 );
nand U90153 ( n31880, n31895, n31896 );
nand U90154 ( n31896, n31897, n76480 );
nand U90155 ( n31895, n31900, n76784 );
nor U90156 ( n31897, n31898, n31899 );
nor U90157 ( n31900, n31901, n31902 );
nor U90158 ( n33616, n33612, n33613 );
nand U90159 ( n66503, n66518, n66519 );
nand U90160 ( n66519, n66520, n76202 );
nand U90161 ( n66518, n66523, n76718 );
nor U90162 ( n66520, n66521, n66522 );
nand U90163 ( n24668, n24683, n24684 );
nand U90164 ( n24684, n24685, n76526 );
nand U90165 ( n24683, n24688, n76766 );
nor U90166 ( n24685, n24686, n24687 );
nand U90167 ( n57802, n57817, n57818 );
nand U90168 ( n57818, n57819, n76268 );
nand U90169 ( n57817, n57822, n76699 );
nor U90170 ( n57819, n57820, n57821 );
nor U90171 ( n66523, n66524, n66525 );
nor U90172 ( n24688, n24689, n24690 );
nor U90173 ( n57822, n57823, n57824 );
nor U90174 ( n26371, n26367, n26368 );
nor U90175 ( n59510, n59506, n59507 );
nor U90176 ( n68372, n68368, n68369 );
nand U90177 ( n41445, n70969, n818 );
nor U90178 ( n70969, n76041, n604 );
nor U90179 ( n36783, n1909, n36492 );
nor U90180 ( n41069, n552, n40884 );
nor U90181 ( n36491, n2098, n36492 );
nor U90182 ( n66357, n788, n76067 );
nand U90183 ( n36448, n36449, n36450 );
nand U90184 ( n36450, n2904, n36310 );
nand U90185 ( n36449, n2145, n76805 );
nor U90186 ( n71937, n71311, n1239 );
not U90187 ( n4910, n13508 );
nand U90188 ( n12088, n5253, n13267 );
nand U90189 ( n12204, n5247, n13449 );
not U90190 ( n4907, n12854 );
not U90191 ( n4909, n13064 );
not U90192 ( n4911, n13700 );
nand U90193 ( n14215, n14285, n14312 );
nand U90194 ( n71315, n71371, n71313 );
nand U90195 ( n12850, n11889, n76727 );
nand U90196 ( n36514, n36515, n36516 );
nand U90197 ( n36516, n2895, n36310 );
nand U90198 ( n36515, n2107, n76805 );
nand U90199 ( n36937, n36938, n36939 );
nand U90200 ( n36939, n2902, n36310 );
nand U90201 ( n36938, n2133, n76805 );
nand U90202 ( n36341, n36342, n36343 );
nand U90203 ( n36343, n2898, n36310 );
nand U90204 ( n36342, n2117, n76805 );
nand U90205 ( n36553, n36554, n36555 );
nand U90206 ( n36555, n2900, n36310 );
nand U90207 ( n36554, n2128, n76805 );
nand U90208 ( n36307, n36308, n36309 );
nand U90209 ( n36309, n2903, n36310 );
nand U90210 ( n36308, n2138, n76805 );
nand U90211 ( n36635, n36636, n36637 );
nand U90212 ( n36637, n2899, n36310 );
nand U90213 ( n36636, n2122, n76805 );
nand U90214 ( n36704, n36705, n36706 );
nand U90215 ( n36706, n2894, n36310 );
nand U90216 ( n36705, n2102, n76805 );
nand U90217 ( n36749, n36750, n36751 );
nand U90218 ( n36751, n2897, n36310 );
nand U90219 ( n36750, n2113, n76805 );
not U90220 ( n76377, n42109 );
nand U90221 ( n42109, n42293, n818 );
nor U90222 ( n42293, n76041, n40665 );
not U90223 ( n4908, n12799 );
nor U90224 ( n45340, n265, n45391 );
nor U90225 ( n40883, n785, n40884 );
nand U90226 ( n12722, n4848, n11763 );
nor U90227 ( n41166, n786, n40884 );
not U90228 ( n16, n14873 );
xor U90229 ( n16562, n16564, n16565 );
nor U90230 ( n37598, n2194, n2193 );
not U90231 ( n3205, n33804 );
nor U90232 ( n44967, n265, n44561 );
nor U90233 ( n44380, n265, n43799 );
not U90234 ( n5804, n68560 );
not U90235 ( n4038, n26559 );
not U90236 ( n6670, n59701 );
nor U90237 ( n71036, n1218, n71171 );
nand U90238 ( n46671, n45782, n7528 );
nor U90239 ( n46658, n46669, n46670 );
nor U90240 ( n46669, n46415, n46673 );
nor U90241 ( n46670, n46413, n46671 );
nand U90242 ( n46673, n45780, n7558 );
nand U90243 ( n32964, n32087, n3140 );
nor U90244 ( n32951, n32962, n32963 );
nor U90245 ( n32962, n32714, n32966 );
nor U90246 ( n32963, n32712, n32964 );
nand U90247 ( n32966, n32085, n3172 );
not U90248 ( n3140, n32882 );
nand U90249 ( n13162, n12039, n4883 );
nor U90250 ( n13145, n13159, n13160 );
nor U90251 ( n13159, n13060, n13164 );
nor U90252 ( n13160, n13055, n13162 );
nand U90253 ( n13164, n12037, n4909 );
nand U90254 ( n67718, n66690, n5742 );
nand U90255 ( n25713, n24855, n3984 );
nand U90256 ( n58853, n57989, n6617 );
nor U90257 ( n67705, n67716, n67717 );
nor U90258 ( n67716, n67479, n67720 );
nor U90259 ( n67717, n67477, n67718 );
nand U90260 ( n67720, n66688, n5770 );
nor U90261 ( n25700, n25711, n25712 );
nor U90262 ( n25711, n25474, n25715 );
nor U90263 ( n25712, n25472, n25713 );
nand U90264 ( n25715, n24853, n4012 );
nor U90265 ( n58840, n58851, n58852 );
nor U90266 ( n58851, n58611, n58855 );
nor U90267 ( n58852, n58609, n58853 );
nand U90268 ( n58855, n57987, n6644 );
not U90269 ( n5742, n67643 );
not U90270 ( n3984, n25638 );
not U90271 ( n6617, n58775 );
nor U90272 ( n13973, n13968, n13969 );
nand U90273 ( n36292, n37085, n37086 );
and U90274 ( n37085, n36681, n36680 );
nand U90275 ( n37086, n36944, n76920 );
not U90276 ( n258, n48055 );
nor U90277 ( n71310, n1235, n71311 );
not U90278 ( n2003, n36944 );
nand U90279 ( n36310, n36680, n36940 );
nand U90280 ( n36940, n36941, n76920 );
nand U90281 ( n36941, n2003, n36942 );
nand U90282 ( n36942, n76409, n36943 );
nand U90283 ( n33431, n76772, n32380 );
nor U90284 ( n71536, n71311, n1238 );
not U90285 ( n76291, n55262 );
nand U90286 ( n55262, n61071, n61072 );
nor U90287 ( n61071, n618, n41445 );
not U90288 ( n76452, n37612 );
nand U90289 ( n37612, n37778, n2198 );
nor U90290 ( n37778, n76039, n36265 );
nor U90291 ( n37089, n2032, n36264 );
nand U90292 ( n11884, n11885, n11887 );
nand U90293 ( n11887, n11888, n76607 );
nand U90294 ( n11885, n11889, n76737 );
not U90295 ( n4938, n14214 );
nand U90296 ( n36617, n2890, n36292 );
nand U90297 ( n37084, n2908, n36292 );
nand U90298 ( n36734, n2917, n36292 );
nand U90299 ( n36766, n2914, n36292 );
nand U90300 ( n36291, n2909, n36292 );
nand U90301 ( n36593, n2929, n36292 );
nand U90302 ( n36671, n2912, n36292 );
nand U90303 ( n13662, n76724, n12377 );
nand U90304 ( n31988, n32003, n32004 );
nand U90305 ( n32004, n32005, n76480 );
nand U90306 ( n32003, n32008, n76784 );
nor U90307 ( n32005, n32006, n32007 );
nor U90308 ( n32008, n32009, n32010 );
nand U90309 ( n66591, n66606, n66607 );
nand U90310 ( n66607, n66608, n76202 );
nand U90311 ( n66606, n66611, n76718 );
nor U90312 ( n66608, n66609, n66610 );
nand U90313 ( n24756, n24771, n24772 );
nand U90314 ( n24772, n24773, n76526 );
nand U90315 ( n24771, n24776, n76766 );
nor U90316 ( n24773, n24774, n24775 );
nand U90317 ( n57890, n57905, n57906 );
nand U90318 ( n57906, n57907, n76268 );
nand U90319 ( n57905, n57910, n76699 );
nor U90320 ( n57907, n57908, n57909 );
nor U90321 ( n66611, n66612, n66613 );
nor U90322 ( n24776, n24777, n24778 );
nor U90323 ( n57910, n57911, n57912 );
nand U90324 ( n37291, n2194, n37297 );
nand U90325 ( n12852, n4848, n11888 );
nand U90326 ( n37100, n38872, n38875 );
and U90327 ( n75774, n38728, n38613 );
nor U90328 ( n16165, n14873, n16130 );
nor U90329 ( n15749, n14873, n15712 );
nor U90330 ( n15218, n14873, n15180 );
nor U90331 ( n15108, n14873, n15073 );
nor U90332 ( n14998, n14873, n14969 );
nor U90333 ( n71040, n1218, n1057 );
nand U90334 ( n33476, n76773, n32414 );
nor U90335 ( n71366, n71311, n1237 );
nor U90336 ( n49195, n48055, n49180 );
nor U90337 ( n48826, n48055, n48811 );
nor U90338 ( n48361, n48055, n48346 );
nor U90339 ( n48264, n48055, n48249 );
nor U90340 ( n48166, n48055, n48151 );
not U90341 ( n252, n48044 );
nor U90342 ( n11528, n17, n11594 );
nand U90343 ( n32975, n76774, n32113 );
nand U90344 ( n13184, n76727, n12072 );
nand U90345 ( n46682, n76660, n45808 );
nand U90346 ( n67729, n76708, n66716 );
nand U90347 ( n25724, n76754, n24881 );
nand U90348 ( n58864, n76687, n58018 );
nor U90349 ( n11282, n17, n10785 );
nor U90350 ( n10570, n17, n9897 );
and U90351 ( n75775, n579, n67261 );
nand U90352 ( n33112, n32169, n3139 );
nor U90353 ( n33100, n33110, n33111 );
nor U90354 ( n33110, n32714, n33114 );
nor U90355 ( n33111, n32712, n33112 );
nand U90356 ( n33114, n32178, n3170 );
not U90357 ( n3139, n33037 );
nand U90358 ( n71147, n71307, n71308 );
nand U90359 ( n46821, n45864, n7525 );
nor U90360 ( n46809, n46819, n46820 );
nor U90361 ( n46819, n46415, n46823 );
nor U90362 ( n46820, n46413, n46821 );
nand U90363 ( n46823, n45873, n7555 );
not U90364 ( n7525, n46745 );
nand U90365 ( n67868, n66815, n5740 );
nand U90366 ( n25865, n24939, n3983 );
nand U90367 ( n59003, n58074, n6615 );
nor U90368 ( n67856, n67866, n67867 );
nor U90369 ( n67866, n67479, n67870 );
nor U90370 ( n67867, n67477, n67868 );
nand U90371 ( n67870, n66824, n5769 );
nor U90372 ( n25853, n25863, n25864 );
nor U90373 ( n25863, n25474, n25867 );
nor U90374 ( n25864, n25472, n25865 );
nand U90375 ( n25867, n24948, n4010 );
nor U90376 ( n58991, n59001, n59002 );
nor U90377 ( n59001, n58611, n59005 );
nor U90378 ( n59002, n58609, n59003 );
nand U90379 ( n59005, n58083, n6643 );
not U90380 ( n5740, n67792 );
not U90381 ( n3983, n25789 );
not U90382 ( n6615, n58927 );
nand U90383 ( n13354, n12147, n4880 );
nor U90384 ( n13339, n13352, n13353 );
nor U90385 ( n13352, n13060, n13357 );
nor U90386 ( n13353, n13055, n13354 );
nand U90387 ( n13357, n12158, n4906 );
not U90388 ( n4880, n13263 );
nand U90389 ( n13514, n76725, n12278 );
nand U90390 ( n12372, n12373, n12374 );
nand U90391 ( n12374, n4790, n9024 );
nand U90392 ( n12373, n76729, n12377 );
nor U90393 ( n71810, n71311, n1222 );
nor U90394 ( n45336, n259, n45391 );
not U90395 ( n3172, n32885 );
not U90396 ( n5770, n67646 );
not U90397 ( n4012, n25641 );
not U90398 ( n6644, n58778 );
nor U90399 ( n44975, n259, n44561 );
nor U90400 ( n44438, n259, n43799 );
nand U90401 ( n12014, n12033, n12034 );
nand U90402 ( n12034, n12035, n76607 );
nand U90403 ( n12033, n12038, n76738 );
and U90404 ( n12035, n4909, n12037 );
and U90405 ( n12038, n4883, n12039 );
nand U90406 ( n45762, n45777, n45778 );
nand U90407 ( n45778, n45779, n76346 );
nand U90408 ( n45777, n45781, n76671 );
and U90409 ( n45779, n7558, n45780 );
and U90410 ( n45781, n7528, n45782 );
nand U90411 ( n32067, n32082, n32083 );
nand U90412 ( n32083, n32084, n76480 );
nand U90413 ( n32082, n32086, n76785 );
and U90414 ( n32084, n3172, n32085 );
and U90415 ( n32086, n3140, n32087 );
not U90416 ( n11, n14859 );
nand U90417 ( n3241, n36260, n76920 );
nand U90418 ( n36260, n36261, n76457 );
nand U90419 ( n36261, n2198, n36263 );
nand U90420 ( n36263, n36264, n36265 );
nand U90421 ( n24835, n24850, n24851 );
nand U90422 ( n24851, n24852, n76526 );
nand U90423 ( n24850, n24854, n76767 );
and U90424 ( n24852, n4012, n24853 );
nand U90425 ( n57969, n57984, n57985 );
nand U90426 ( n57985, n57986, n76268 );
nand U90427 ( n57984, n57988, n76700 );
and U90428 ( n57986, n6644, n57987 );
nand U90429 ( n66670, n66685, n66686 );
nand U90430 ( n66686, n66687, n76202 );
nand U90431 ( n66685, n66689, n76719 );
and U90432 ( n66687, n5770, n66688 );
and U90433 ( n66689, n5742, n66690 );
and U90434 ( n24854, n3984, n24855 );
and U90435 ( n57988, n6617, n57989 );
nand U90436 ( n23826, n28728, n28729 );
nor U90437 ( n28728, n28744, n28745 );
nor U90438 ( n28729, n28730, n28731 );
nand U90439 ( n28744, n28752, n28753 );
nand U90440 ( n56950, n62033, n62034 );
nor U90441 ( n62033, n62049, n62050 );
nor U90442 ( n62034, n62035, n62036 );
nand U90443 ( n62049, n62057, n62058 );
nand U90444 ( n24322, n28624, n28625 );
nand U90445 ( n28624, n25408, n4224 );
or U90446 ( n28625, n22781, n167 );
nand U90447 ( n55895, n57739, n60030 );
nand U90448 ( n22781, n24607, n26890 );
and U90449 ( n56380, n6553, n57442 );
nand U90450 ( n57442, n438, n57443 );
nand U90451 ( n57443, n57444, n6640 );
not U90452 ( n438, n57445 );
and U90453 ( n23256, n3920, n24319 );
nand U90454 ( n24319, n165, n24320 );
nand U90455 ( n24320, n24321, n4008 );
not U90456 ( n165, n24322 );
nand U90457 ( n57445, n61929, n61930 );
nand U90458 ( n61929, n58545, n6857 );
or U90459 ( n61930, n55895, n439 );
nand U90460 ( n64119, n66415, n68889 );
nand U90461 ( n65424, n70633, n70634 );
nor U90462 ( n70633, n70649, n70650 );
nor U90463 ( n70634, n70635, n70636 );
nand U90464 ( n70649, n70657, n70658 );
and U90465 ( n64736, n5678, n65901 );
nand U90466 ( n65901, n470, n65902 );
nand U90467 ( n65902, n65903, n5767 );
not U90468 ( n470, n65904 );
nand U90469 ( n65904, n70529, n70530 );
nand U90470 ( n70529, n67413, n6002 );
or U90471 ( n70530, n64119, n472 );
nand U90472 ( n31618, n35803, n35804 );
nand U90473 ( n35803, n32648, n3387 );
or U90474 ( n35804, n30102, n200 );
nand U90475 ( n30102, n31823, n34135 );
nand U90476 ( n31170, n35907, n35908 );
nor U90477 ( n35907, n35923, n35924 );
nor U90478 ( n35908, n35909, n35910 );
nand U90479 ( n35923, n35931, n35932 );
and U90480 ( n30577, n3077, n31615 );
nand U90481 ( n31615, n199, n31616 );
nand U90482 ( n31616, n31617, n3168 );
not U90483 ( n199, n31618 );
nand U90484 ( n26918, n28758, n28759 );
nor U90485 ( n28758, n28774, n28775 );
nor U90486 ( n28759, n28760, n28761 );
nand U90487 ( n28774, n28782, n28783 );
nand U90488 ( n60058, n62063, n62064 );
nor U90489 ( n62063, n62079, n62080 );
nor U90490 ( n62064, n62065, n62066 );
nand U90491 ( n62079, n62087, n62088 );
nand U90492 ( n68917, n70663, n70664 );
nor U90493 ( n70663, n70679, n70680 );
nor U90494 ( n70664, n70665, n70666 );
nand U90495 ( n70679, n70687, n70688 );
nand U90496 ( n34163, n35937, n35938 );
nor U90497 ( n35937, n35953, n35954 );
nor U90498 ( n35938, n35939, n35940 );
nand U90499 ( n35953, n35961, n35962 );
not U90500 ( n1357, n49719 );
nand U90501 ( n28664, n4229, n4252 );
nand U90502 ( n61969, n6862, n6884 );
nand U90503 ( n24601, n28696, n28697 );
nor U90504 ( n28696, n28712, n28713 );
nor U90505 ( n28697, n28698, n28699 );
nand U90506 ( n28712, n28720, n28721 );
nand U90507 ( n57733, n62001, n62002 );
nor U90508 ( n62001, n62017, n62018 );
nor U90509 ( n62002, n62003, n62004 );
nand U90510 ( n62017, n62025, n62026 );
not U90511 ( n4252, n24210 );
not U90512 ( n6884, n57332 );
nand U90513 ( n70569, n6007, n6029 );
nand U90514 ( n66409, n70601, n70602 );
nor U90515 ( n70601, n70617, n70618 );
nor U90516 ( n70602, n70603, n70604 );
nand U90517 ( n70617, n70625, n70626 );
not U90518 ( n6029, n65754 );
nand U90519 ( n35843, n3392, n3414 );
nand U90520 ( n31817, n35875, n35876 );
nor U90521 ( n35875, n35891, n35892 );
nor U90522 ( n35876, n35877, n35878 );
nand U90523 ( n35891, n35899, n35900 );
not U90524 ( n3414, n31504 );
nand U90525 ( n28694, n4234, n4252 );
nand U90526 ( n61999, n6867, n6884 );
nand U90527 ( n70599, n6012, n6029 );
nand U90528 ( n23077, n28788, n28789 );
nor U90529 ( n28788, n28804, n28805 );
nor U90530 ( n28789, n28790, n28791 );
nand U90531 ( n28804, n28812, n28813 );
nand U90532 ( n56198, n62093, n62094 );
nor U90533 ( n62093, n62109, n62110 );
nor U90534 ( n62094, n62095, n62096 );
nand U90535 ( n62109, n62117, n62118 );
nand U90536 ( n35873, n3397, n3414 );
nand U90537 ( n64567, n70693, n70694 );
nor U90538 ( n70693, n70709, n70710 );
nor U90539 ( n70694, n70695, n70696 );
nand U90540 ( n70709, n70717, n70718 );
nand U90541 ( n30408, n35967, n35968 );
nor U90542 ( n35967, n35983, n35984 );
nor U90543 ( n35968, n35969, n35970 );
nand U90544 ( n35983, n35991, n35992 );
nand U90545 ( n61512, n61957, n61958 );
nor U90546 ( n61957, n61980, n61981 );
nor U90547 ( n61958, n61959, n61960 );
nand U90548 ( n61980, n61992, n61993 );
nand U90549 ( n28290, n28652, n28653 );
nor U90550 ( n28652, n28675, n28676 );
nor U90551 ( n28653, n28654, n28655 );
nand U90552 ( n28675, n28687, n28688 );
nand U90553 ( n70246, n70557, n70558 );
nor U90554 ( n70557, n70580, n70581 );
nor U90555 ( n70558, n70559, n70560 );
nand U90556 ( n70580, n70592, n70593 );
nand U90557 ( n35518, n35831, n35832 );
nor U90558 ( n35831, n35854, n35855 );
nor U90559 ( n35832, n35833, n35834 );
nand U90560 ( n35854, n35866, n35867 );
nand U90561 ( n28691, n4234, n4248 );
nand U90562 ( n61996, n6867, n6880 );
nand U90563 ( n70596, n6012, n6025 );
nand U90564 ( n35870, n3397, n3410 );
nor U90565 ( n41458, n40664, n840 );
nand U90566 ( n2016, n40660, n76925 );
nand U90567 ( n40660, n40661, n76389 );
nand U90568 ( n40661, n818, n40663 );
nand U90569 ( n40663, n40664, n40665 );
nand U90570 ( n47232, n76658, n46122 );
nand U90571 ( n28660, n4229, n4248 );
nand U90572 ( n28695, n4234, n4250 );
nand U90573 ( n61965, n6862, n6880 );
nand U90574 ( n62000, n6867, n6883 );
nand U90575 ( n68263, n76706, n67086 );
nand U90576 ( n26262, n76752, n25188 );
nand U90577 ( n59401, n76685, n58324 );
nand U90578 ( n70565, n6007, n6025 );
nand U90579 ( n35839, n3392, n3410 );
nand U90580 ( n70600, n6012, n6028 );
nor U90581 ( n49187, n48044, n49180 );
nor U90582 ( n48818, n48044, n48811 );
nor U90583 ( n48353, n48044, n48346 );
nor U90584 ( n48256, n48044, n48249 );
nor U90585 ( n48158, n48044, n48151 );
nand U90586 ( n35874, n3397, n3413 );
not U90587 ( n1272, n50605 );
nand U90588 ( n28336, n28818, n28819 );
nor U90589 ( n28818, n28834, n28835 );
nor U90590 ( n28819, n28820, n28821 );
nand U90591 ( n28834, n28842, n28843 );
nand U90592 ( n61558, n62123, n62124 );
nor U90593 ( n62123, n62139, n62140 );
nor U90594 ( n62124, n62125, n62126 );
nand U90595 ( n62139, n62147, n62148 );
nand U90596 ( n70274, n70723, n70724 );
nor U90597 ( n70723, n70739, n70740 );
nor U90598 ( n70724, n70725, n70726 );
nand U90599 ( n70739, n70747, n70748 );
nand U90600 ( n35546, n35997, n35998 );
nor U90601 ( n35997, n36013, n36014 );
nor U90602 ( n35998, n35999, n36000 );
nand U90603 ( n36013, n36021, n36022 );
and U90604 ( n75776, n2087, n40402 );
nand U90605 ( n36492, n2087, n37109 );
nand U90606 ( n37109, n37110, n37111 );
nand U90607 ( n37111, n76409, n2090 );
not U90608 ( n2090, n36943 );
nand U90609 ( n28665, n4229, n4250 );
nand U90610 ( n61970, n6862, n6883 );
nand U90611 ( n70570, n6007, n6028 );
nand U90612 ( n32109, n32110, n32111 );
nand U90613 ( n32111, n76481, n32112 );
nand U90614 ( n32110, n76785, n32113 );
nand U90615 ( n35844, n3392, n3413 );
nand U90616 ( n12067, n12068, n12069 );
nand U90617 ( n12069, n76607, n12070 );
nand U90618 ( n12068, n76738, n12072 );
nand U90619 ( n45804, n45805, n45806 );
nand U90620 ( n45806, n76347, n45807 );
nand U90621 ( n45805, n76671, n45808 );
nand U90622 ( n66712, n66713, n66714 );
nand U90623 ( n66714, n76203, n66715 );
nand U90624 ( n66713, n76719, n66716 );
nand U90625 ( n24877, n24878, n24879 );
nand U90626 ( n24879, n76527, n24880 );
nand U90627 ( n24878, n76767, n24881 );
nand U90628 ( n58014, n58015, n58016 );
nand U90629 ( n58016, n76269, n58017 );
nand U90630 ( n58015, n76700, n58018 );
nand U90631 ( n26903, n28848, n28849 );
nor U90632 ( n28848, n28864, n28865 );
nor U90633 ( n28849, n28850, n28851 );
nand U90634 ( n28864, n28872, n28873 );
nand U90635 ( n60043, n62153, n62154 );
nor U90636 ( n62153, n62169, n62170 );
nor U90637 ( n62154, n62155, n62156 );
nand U90638 ( n62169, n62177, n62178 );
nand U90639 ( n68902, n70753, n70754 );
nor U90640 ( n70753, n70769, n70770 );
nor U90641 ( n70754, n70755, n70756 );
nand U90642 ( n70769, n70777, n70778 );
nand U90643 ( n34148, n36027, n36028 );
nor U90644 ( n36027, n36043, n36044 );
nor U90645 ( n36028, n36029, n36030 );
nand U90646 ( n36043, n36051, n36052 );
nor U90647 ( n67222, n829, n845 );
nand U90648 ( n41229, n41442, n41443 );
nor U90649 ( n41442, n41444, n41445 );
nand U90650 ( n33508, n76773, n32430 );
nand U90651 ( n8659, n8438, n8660 );
nand U90652 ( n8660, n76744, n5273 );
not U90653 ( n5310, n12328 );
not U90654 ( n5309, n12167 );
nor U90655 ( n45332, n253, n45391 );
nand U90656 ( n9114, n8438, n9115 );
nand U90657 ( n9115, n76744, n5282 );
nand U90658 ( n9109, n9110, n9112 );
nand U90659 ( n9112, n9113, n76743 );
nand U90660 ( n9110, n9080, n9114 );
nor U90661 ( n9113, n5282, n9080 );
nand U90662 ( n8725, n8438, n8727 );
nand U90663 ( n8727, n76744, n5274 );
nand U90664 ( n8597, n8438, n8598 );
nand U90665 ( n8598, n76744, n5272 );
nand U90666 ( n8933, n8438, n8934 );
nand U90667 ( n8934, n76744, n5278 );
nand U90668 ( n9194, n8438, n9195 );
nand U90669 ( n9195, n76744, n5283 );
nand U90670 ( n8999, n8438, n9000 );
nand U90671 ( n9000, n76744, n5279 );
nand U90672 ( n8805, n8438, n8807 );
nand U90673 ( n8807, n76744, n5275 );
nand U90674 ( n38376, n76439, n36572 );
nor U90675 ( n38146, n38604, n38119 );
nand U90676 ( n38475, n76438, n36355 );
nand U90677 ( n38331, n76439, n36398 );
nand U90678 ( n38557, n76438, n36589 );
nand U90679 ( n38194, n76439, n36305 );
nand U90680 ( n38394, n76439, n36961 );
nand U90681 ( n38242, n76439, n36633 );
nand U90682 ( n38293, n76439, n36512 );
nand U90683 ( n38587, n76438, n36381 );
nand U90684 ( n38494, n76438, n36667 );
nand U90685 ( n38526, n76438, n36286 );
nand U90686 ( n42721, n42512, n42722 );
nand U90687 ( n42722, n76677, n7928 );
not U90688 ( n7965, n46011 );
not U90689 ( n7964, n45880 );
nand U90690 ( n38510, n76438, n36462 );
nand U90691 ( n38213, n76439, n36925 );
nand U90692 ( n38541, n76438, n36817 );
nand U90693 ( n38315, n76439, n36702 );
not U90694 ( n6, n14845 );
nand U90695 ( n38410, n76438, n36322 );
nand U90696 ( n38442, n76438, n36532 );
not U90697 ( n2047, n38875 );
nand U90698 ( n38277, n76439, n36747 );
nand U90699 ( n33123, n76774, n32207 );
nand U90700 ( n38347, n76439, n36797 );
nor U90701 ( n16155, n14859, n16130 );
nor U90702 ( n15730, n14859, n15712 );
nor U90703 ( n15199, n14859, n15180 );
nor U90704 ( n15098, n14859, n15073 );
nor U90705 ( n14988, n14859, n14969 );
nand U90706 ( n43103, n42512, n43104 );
nand U90707 ( n43104, n76677, n7937 );
nand U90708 ( n43099, n43100, n43101 );
nand U90709 ( n43101, n43102, n76677 );
nand U90710 ( n43100, n43076, n43103 );
nor U90711 ( n43102, n7937, n43076 );
nand U90712 ( n13368, n76727, n12194 );
nand U90713 ( n42944, n42512, n42945 );
nand U90714 ( n42945, n76677, n7933 );
nand U90715 ( n46832, n76660, n45902 );
nand U90716 ( n43167, n42512, n43168 );
nand U90717 ( n43168, n76677, n7938 );
nand U90718 ( n43011, n42512, n43012 );
nand U90719 ( n43012, n76677, n7934 );
nand U90720 ( n42842, n42512, n42843 );
nand U90721 ( n42843, n76677, n7930 );
nand U90722 ( n67879, n76708, n66853 );
nand U90723 ( n25876, n76754, n24977 );
nand U90724 ( n59014, n76687, n58112 );
nor U90725 ( n38129, n38119, n37103 );
nor U90726 ( n65818, n667, n61441 );
nor U90727 ( n44983, n253, n44561 );
nor U90728 ( n44480, n253, n43799 );
nand U90729 ( n71125, n71357, n71144 );
nor U90730 ( n38127, n38119, n37110 );
nand U90731 ( n38145, n76440, n37295 );
nand U90732 ( n38181, n76440, n36442 );
nand U90733 ( n38162, n76440, n36429 );
nand U90734 ( n38423, n76446, n2914 );
nand U90735 ( n38455, n76446, n2912 );
nand U90736 ( n38360, n76447, n2908 );
nand U90737 ( n38258, n76447, n2895 );
nand U90738 ( n38226, n76447, n2898 );
nand U90739 ( n32976, n3103, n32112 );
nand U90740 ( n13185, n4848, n12070 );
nor U90741 ( n62332, n759, n61441 );
nand U90742 ( n38241, n76447, n2897 );
nand U90743 ( n33523, n3103, n32429 );
nand U90744 ( n46683, n7490, n45807 );
nand U90745 ( n38330, n76447, n2890 );
nand U90746 ( n38292, n76447, n2893 );
nand U90747 ( n38393, n76447, n2917 );
nand U90748 ( n38525, n76446, n2929 );
nand U90749 ( n38493, n76446, n2909 );
nand U90750 ( n67730, n5704, n66715 );
nand U90751 ( n25725, n3947, n24880 );
nand U90752 ( n58865, n6579, n58017 );
nor U90753 ( n66111, n650, n61441 );
nor U90754 ( n39305, n2180, n38822 );
nand U90755 ( n38193, n76448, n2900 );
nand U90756 ( n38161, n76448, n2903 );
nand U90757 ( n38144, n76448, n2904 );
nand U90758 ( n38180, n76448, n2902 );
not U90759 ( n3063, n31969 );
nand U90760 ( n32172, n32154, n32192 );
nand U90761 ( n32192, n3055, n3560 );
and U90762 ( n32154, n31969, n32193 );
nand U90763 ( n32193, n76779, n32152 );
buf U90764 ( n76779, n3058 );
and U90765 ( n31891, n31969, n31970 );
nand U90766 ( n31970, n76779, n31888 );
not U90767 ( n3053, n31960 );
nand U90768 ( n54341, n7794, n7817 );
not U90769 ( n3907, n24737 );
not U90770 ( n7438, n45648 );
not U90771 ( n5664, n66572 );
not U90772 ( n6539, n57871 );
nand U90773 ( n45509, n54373, n54374 );
nor U90774 ( n54373, n54389, n54390 );
nor U90775 ( n54374, n54375, n54376 );
nand U90776 ( n54389, n54397, n54398 );
not U90777 ( n7817, n44889 );
nand U90778 ( n45867, n45849, n45887 );
nand U90779 ( n45887, n7430, n7964 );
nand U90780 ( n66818, n66800, n66838 );
nand U90781 ( n66838, n5657, n6175 );
nand U90782 ( n24942, n24922, n24962 );
nand U90783 ( n24962, n3899, n4398 );
nand U90784 ( n58077, n58059, n58097 );
nand U90785 ( n58097, n6532, n7030 );
nor U90786 ( n39720, n2172, n38822 );
and U90787 ( n66800, n66572, n66839 );
nand U90788 ( n66839, n76713, n66798 );
and U90789 ( n45849, n45648, n45888 );
nand U90790 ( n45888, n76665, n45847 );
and U90791 ( n24922, n24737, n24963 );
nand U90792 ( n24963, n76761, n24920 );
and U90793 ( n58059, n57871, n58098 );
nand U90794 ( n58098, n76694, n58057 );
buf U90795 ( n76665, n7433 );
buf U90796 ( n76761, n3902 );
buf U90797 ( n76694, n6534 );
buf U90798 ( n76713, n5659 );
and U90799 ( n24679, n24737, n24738 );
nand U90800 ( n24738, n76761, n24676 );
and U90801 ( n66514, n66572, n66573 );
nand U90802 ( n66573, n76713, n66511 );
and U90803 ( n57813, n57871, n57872 );
nand U90804 ( n57872, n76694, n57810 );
not U90805 ( n3897, n24728 );
not U90806 ( n5654, n66563 );
not U90807 ( n6529, n57862 );
nand U90808 ( n68278, n5704, n67085 );
nand U90809 ( n47247, n7490, n46121 );
nand U90810 ( n26277, n3947, n25187 );
nand U90811 ( n59416, n6579, n58323 );
and U90812 ( n32078, n31969, n32136 );
nand U90813 ( n32136, n76779, n32075 );
and U90814 ( n45678, n45648, n45726 );
nand U90815 ( n45726, n76665, n45675 );
not U90816 ( n7428, n45706 );
and U90817 ( n45589, n45648, n45649 );
nand U90818 ( n45649, n76665, n45586 );
not U90819 ( n7429, n45639 );
and U90820 ( n66681, n66572, n66782 );
nand U90821 ( n66782, n76713, n66678 );
and U90822 ( n24846, n24737, n24904 );
nand U90823 ( n24904, n76761, n24843 );
and U90824 ( n57980, n57871, n58041 );
nand U90825 ( n58041, n76694, n57977 );
and U90826 ( n31999, n31969, n32049 );
nand U90827 ( n32049, n76779, n31996 );
not U90828 ( n3052, n32028 );
nand U90829 ( n26905, n28878, n28879 );
nor U90830 ( n28878, n28894, n28895 );
nor U90831 ( n28879, n28880, n28881 );
nand U90832 ( n28894, n28902, n28903 );
nand U90833 ( n60045, n62183, n62184 );
nor U90834 ( n62183, n62199, n62200 );
nor U90835 ( n62184, n62185, n62186 );
nand U90836 ( n62199, n62207, n62208 );
nand U90837 ( n32320, n32297, n32335 );
nand U90838 ( n32335, n3055, n3562 );
and U90839 ( n32297, n31969, n32336 );
nand U90840 ( n32336, n76780, n32295 );
buf U90841 ( n76780, n3058 );
not U90842 ( n824, n61617 );
nor U90843 ( n40020, n2164, n38822 );
and U90844 ( n45773, n45648, n45831 );
nand U90845 ( n45831, n76665, n45770 );
nand U90846 ( n68904, n70783, n70784 );
nor U90847 ( n70783, n70799, n70800 );
nor U90848 ( n70784, n70785, n70786 );
nand U90849 ( n70799, n70807, n70808 );
and U90850 ( n66602, n66572, n66652 );
nand U90851 ( n66652, n76713, n66599 );
and U90852 ( n24767, n24737, n24817 );
nand U90853 ( n24817, n76761, n24764 );
and U90854 ( n57901, n57871, n57951 );
nand U90855 ( n57951, n76694, n57898 );
not U90856 ( n5653, n66631 );
not U90857 ( n3895, n24796 );
not U90858 ( n6528, n57930 );
nand U90859 ( n34150, n36057, n36058 );
nor U90860 ( n36057, n36073, n36074 );
nor U90861 ( n36058, n36059, n36060 );
nand U90862 ( n36073, n36081, n36082 );
nand U90863 ( n46019, n45985, n46034 );
nand U90864 ( n46034, n7430, n7965 );
nand U90865 ( n66959, n66936, n66974 );
nand U90866 ( n66974, n5657, n6177 );
nand U90867 ( n25083, n25060, n25098 );
nand U90868 ( n25098, n3899, n4399 );
nand U90869 ( n58218, n58195, n58236 );
nand U90870 ( n58236, n6532, n7032 );
and U90871 ( n66936, n66572, n66975 );
nand U90872 ( n66975, n76714, n66934 );
and U90873 ( n45985, n45648, n46035 );
nand U90874 ( n46035, n76666, n45983 );
and U90875 ( n25060, n24737, n25099 );
nand U90876 ( n25099, n76762, n25058 );
and U90877 ( n58195, n57871, n58237 );
nand U90878 ( n58237, n76695, n58193 );
buf U90879 ( n76714, n5659 );
buf U90880 ( n76762, n3902 );
buf U90881 ( n76695, n6534 );
buf U90882 ( n76666, n7433 );
nand U90883 ( n32514, n31969, n32532 );
nand U90884 ( n67170, n66572, n67188 );
nand U90885 ( n25272, n24737, n25290 );
nand U90886 ( n58408, n57871, n58426 );
nand U90887 ( n46206, n45648, n46236 );
nand U90888 ( n43725, n54465, n54466 );
nor U90889 ( n54465, n54481, n54482 );
nor U90890 ( n54466, n54467, n54468 );
nand U90891 ( n54481, n54489, n54490 );
and U90892 ( n12145, n4880, n12147 );
nand U90893 ( n68310, n76705, n67106 );
nand U90894 ( n26309, n76751, n25208 );
nand U90895 ( n59448, n76684, n58344 );
nor U90896 ( n39984, n2165, n38822 );
nand U90897 ( n33554, n76772, n32450 );
nand U90898 ( n47279, n76657, n46142 );
nand U90899 ( n36489, n37077, n37078 );
nor U90900 ( n37077, n2153, n36943 );
nand U90901 ( n47884, n54555, n54556 );
nor U90902 ( n54555, n54571, n54572 );
nor U90903 ( n54556, n54557, n54558 );
nand U90904 ( n54571, n54579, n54580 );
not U90905 ( n4895, n13035 );
nand U90906 ( n54371, n7799, n7817 );
nor U90907 ( n41443, n41479, n618 );
nor U90908 ( n39001, n2187, n38822 );
nand U90909 ( n9312, n8438, n9313 );
nand U90910 ( n9313, n76745, n5285 );
buf U90911 ( n76745, n76741 );
buf U90912 ( n76741, n4760 );
nand U90913 ( n32460, n31969, n32474 );
nand U90914 ( n32474, n76780, n32409 );
nand U90915 ( n67116, n66572, n67130 );
nand U90916 ( n67130, n76714, n67072 );
nand U90917 ( n32392, n31969, n32406 );
nand U90918 ( n32406, n76780, n32339 );
nand U90919 ( n46152, n45648, n46166 );
nand U90920 ( n46166, n76666, n46108 );
nand U90921 ( n25218, n24737, n25232 );
nand U90922 ( n25232, n76762, n25174 );
nand U90923 ( n58354, n57871, n58368 );
nand U90924 ( n58368, n76695, n58310 );
nand U90925 ( n67055, n66572, n67069 );
nand U90926 ( n67069, n76714, n66978 );
nand U90927 ( n46091, n45648, n46105 );
nand U90928 ( n46105, n76666, n46038 );
nand U90929 ( n25155, n24737, n25171 );
nand U90930 ( n25171, n76762, n25102 );
nand U90931 ( n58293, n57871, n58307 );
nand U90932 ( n58307, n76695, n58240 );
nand U90933 ( n54337, n7794, n7813 );
nand U90934 ( n21358, n5139, n5162 );
not U90935 ( n4794, n11899 );
nand U90936 ( n11733, n21390, n21391 );
nor U90937 ( n21390, n21406, n21407 );
nor U90938 ( n21391, n21392, n21393 );
nand U90939 ( n21406, n21414, n21415 );
not U90940 ( n5162, n11178 );
not U90941 ( n4906, n13267 );
and U90942 ( n11842, n11899, n11900 );
nand U90943 ( n11900, n76732, n11838 );
not U90944 ( n4785, n11864 );
buf U90945 ( n76732, n4789 );
xor U90946 ( MUL_1411_U12, n71512, n71513 );
xor U90947 ( n71513, n71514, n71515 );
nand U90948 ( n8533, n8438, n8534 );
nand U90949 ( n8534, n76745, n5270 );
not U90950 ( n3170, n33040 );
nand U90951 ( n49545, n54495, n54496 );
nor U90952 ( n54495, n54511, n54512 );
nor U90953 ( n54496, n54497, n54498 );
nand U90954 ( n54511, n54519, n54520 );
nand U90955 ( n9063, n8438, n9064 );
nand U90956 ( n9064, n76745, n5280 );
nand U90957 ( n9257, n8438, n9258 );
nand U90958 ( n9258, n76745, n5284 );
nand U90959 ( n32176, n32197, n32198 );
nand U90960 ( n32198, n3055, n32185 );
nand U90961 ( n32197, n76779, n3569 );
not U90962 ( n4224, n26901 );
not U90963 ( n6857, n60041 );
nand U90964 ( n66822, n66843, n66844 );
nand U90965 ( n66844, n5657, n66831 );
nand U90966 ( n66843, n76713, n6184 );
nand U90967 ( n24946, n24967, n24968 );
nand U90968 ( n24968, n3899, n24955 );
nand U90969 ( n24967, n76761, n4407 );
nand U90970 ( n58081, n58102, n58103 );
nand U90971 ( n58103, n6532, n58090 );
nand U90972 ( n58102, n76694, n7039 );
nand U90973 ( n43275, n42512, n43276 );
nand U90974 ( n43276, n76678, n7940 );
nand U90975 ( n12150, n12128, n12175 );
nand U90976 ( n12175, n4787, n5309 );
not U90977 ( n7555, n46748 );
and U90978 ( n12128, n11899, n12177 );
nand U90979 ( n12177, n76732, n12125 );
buf U90980 ( n76678, n76674 );
buf U90981 ( n76674, n7405 );
not U90982 ( n6002, n68900 );
not U90983 ( n3387, n34146 );
nand U90984 ( n45871, n45892, n45893 );
nand U90985 ( n45893, n7430, n45880 );
nand U90986 ( n45892, n76665, n7973 );
not U90987 ( n4893, n13522 );
not U90988 ( n5769, n67795 );
and U90989 ( n11942, n11899, n11992 );
nand U90990 ( n11992, n76732, n11938 );
nand U90991 ( n32252, n32273, n32274 );
nand U90992 ( n32274, n3055, n3549 );
nand U90993 ( n32273, n76780, n3570 );
not U90994 ( n4010, n25792 );
not U90995 ( n6643, n58930 );
nand U90996 ( n45940, n45961, n45962 );
nand U90997 ( n45962, n7430, n7952 );
nand U90998 ( n45961, n76666, n7974 );
nand U90999 ( n66891, n66912, n66913 );
nand U91000 ( n66913, n5657, n6164 );
nand U91001 ( n66912, n76714, n6185 );
nand U91002 ( n32317, n32333, n32334 );
nand U91003 ( n32334, n3055, n32312 );
nand U91004 ( n32333, n76780, n3572 );
nand U91005 ( n25015, n25036, n25037 );
nand U91006 ( n25037, n3899, n4387 );
nand U91007 ( n25036, n76762, n4408 );
nand U91008 ( n58150, n58171, n58172 );
nand U91009 ( n58172, n6532, n7019 );
nand U91010 ( n58171, n76695, n7040 );
nand U91011 ( n46118, n46119, n46120 );
nand U91012 ( n46120, n76347, n46121 );
nand U91013 ( n46119, n46122, n76662 );
nand U91014 ( n67082, n67083, n67084 );
nand U91015 ( n67084, n76203, n67085 );
nand U91016 ( n67083, n67086, n76710 );
nand U91017 ( n25184, n25185, n25186 );
nand U91018 ( n25186, n76527, n25187 );
nand U91019 ( n25185, n25188, n76758 );
nand U91020 ( n58320, n58321, n58322 );
nand U91021 ( n58322, n76269, n58323 );
nand U91022 ( n58321, n58324, n76691 );
nand U91023 ( n46016, n46032, n46033 );
nand U91024 ( n46033, n7430, n46011 );
nand U91025 ( n46032, n76666, n7975 );
nand U91026 ( n66956, n66972, n66973 );
nand U91027 ( n66973, n5657, n66951 );
nand U91028 ( n66972, n76714, n6187 );
nand U91029 ( n25080, n25096, n25097 );
nand U91030 ( n25097, n3899, n25075 );
nand U91031 ( n25096, n76762, n4409 );
nand U91032 ( n58215, n58234, n58235 );
nand U91033 ( n58235, n6532, n58210 );
nand U91034 ( n58234, n76695, n7042 );
and U91035 ( n12028, n11899, n12100 );
nand U91036 ( n12100, n76732, n12024 );
nand U91037 ( n12338, n12309, n12357 );
nand U91038 ( n12357, n4787, n5310 );
and U91039 ( n12309, n11899, n12358 );
nand U91040 ( n12358, n76733, n12307 );
buf U91041 ( n76733, n4789 );
nand U91042 ( n4501, n32444, n32445 );
nor U91043 ( n32445, n32446, n32447 );
nor U91044 ( n32444, n32456, n32457 );
nand U91045 ( n32446, n32452, n32453 );
nand U91046 ( n42778, n42512, n42779 );
nand U91047 ( n42779, n76678, n7929 );
nand U91048 ( n42647, n42512, n42648 );
nand U91049 ( n42648, n76678, n7927 );
nand U91050 ( n42596, n42512, n42597 );
nand U91051 ( n42597, n76678, n7925 );
nand U91052 ( n11236, n67100, n67101 );
nor U91053 ( n67101, n67102, n67103 );
nor U91054 ( n67100, n67112, n67113 );
nand U91055 ( n67102, n67108, n67109 );
nand U91056 ( n15726, n46136, n46137 );
nor U91057 ( n46137, n46138, n46139 );
nor U91058 ( n46136, n46148, n46149 );
nand U91059 ( n46138, n46144, n46145 );
nand U91060 ( n6746, n25202, n25203 );
nor U91061 ( n25203, n25204, n25205 );
nor U91062 ( n25202, n25214, n25215 );
nand U91063 ( n25204, n25210, n25211 );
nand U91064 ( n13481, n58338, n58339 );
nor U91065 ( n58339, n58340, n58341 );
nor U91066 ( n58338, n58350, n58351 );
nand U91067 ( n58340, n58346, n58347 );
nand U91068 ( n43062, n42512, n43063 );
nand U91069 ( n43063, n76678, n7935 );
nand U91070 ( n43217, n42512, n43218 );
nand U91071 ( n43218, n76678, n7939 );
nand U91072 ( n8437, n8438, n8439 );
nand U91073 ( n8439, n76745, n8400 );
nand U91074 ( n42507, n42508, n42509 );
nand U91075 ( n42509, n42510, n76675 );
nand U91076 ( n42508, n42490, n42511 );
nor U91077 ( n42510, n7924, n42490 );
nand U91078 ( n42511, n42512, n42513 );
nand U91079 ( n42513, n76678, n7924 );
nand U91080 ( n9804, n21482, n21483 );
nor U91081 ( n21482, n21498, n21499 );
nor U91082 ( n21483, n21484, n21485 );
nand U91083 ( n21498, n21506, n21507 );
nor U91084 ( n11523, n12, n11594 );
nor U91085 ( n71324, n1238, n71325 );
nand U91086 ( n12578, n11899, n12600 );
nand U91087 ( n14654, n21572, n21573 );
nor U91088 ( n21572, n21588, n21589 );
nor U91089 ( n21573, n21574, n21575 );
nand U91090 ( n21588, n21596, n21597 );
and U91091 ( n75777, n2064, n2083 );
nand U91092 ( n21388, n5144, n5162 );
not U91093 ( n835, n41487 );
nor U91094 ( n67224, n838, n842 );
nand U91095 ( n21354, n5139, n5158 );
nand U91096 ( n47897, n54435, n54436 );
nor U91097 ( n54435, n54451, n54452 );
nor U91098 ( n54436, n54437, n54438 );
nand U91099 ( n54451, n54459, n54460 );
nand U91100 ( n12510, n11899, n12528 );
nand U91101 ( n12528, n76733, n12455 );
not U91102 ( n2044, n38865 );
nand U91103 ( n54368, n7799, n7813 );
nand U91104 ( n12434, n11899, n12452 );
nand U91105 ( n12452, n76733, n12362 );
nand U91106 ( n16567, n21512, n21513 );
nor U91107 ( n21512, n21528, n21529 );
nor U91108 ( n21513, n21514, n21515 );
nand U91109 ( n21528, n21536, n21537 );
nand U91110 ( n44495, n54405, n54406 );
nor U91111 ( n54405, n54421, n54422 );
nor U91112 ( n54406, n54407, n54408 );
nand U91113 ( n54421, n54429, n54430 );
nand U91114 ( n54372, n7799, n7815 );
nand U91115 ( n12155, n12182, n12183 );
nand U91116 ( n12183, n4787, n12167 );
nand U91117 ( n12182, n76732, n5318 );
nand U91118 ( n9202, n9214, n8789 );
nand U91119 ( n9214, n9215, n76744 );
nor U91120 ( n9215, n5283, n9217 );
nor U91121 ( n9217, n9218, n9219 );
nand U91122 ( n12253, n12279, n12280 );
nand U91123 ( n12280, n4787, n5297 );
nand U91124 ( n12279, n76733, n5319 );
nand U91125 ( n12334, n12354, n12355 );
nand U91126 ( n12355, n4787, n12328 );
nand U91127 ( n12354, n76733, n5320 );
nand U91128 ( n8940, n8952, n8789 );
nand U91129 ( n8952, n8953, n76743 );
nor U91130 ( n8953, n5278, n8954 );
nor U91131 ( n8954, n8955, n5294 );
nand U91132 ( n9007, n9019, n8789 );
nand U91133 ( n9019, n9020, n76743 );
nor U91134 ( n9020, n5279, n9022 );
nor U91135 ( n9022, n9023, n5293 );
nand U91136 ( n8813, n8825, n8789 );
nand U91137 ( n8825, n8827, n76742 );
nor U91138 ( n8827, n5275, n8828 );
nor U91139 ( n8828, n8829, n5298 );
nand U91140 ( n9006, n12410, n12412 );
nor U91141 ( n12412, n12413, n12414 );
nor U91142 ( n12410, n12429, n12430 );
nand U91143 ( n12413, n12420, n12422 );
nand U91144 ( n8991, n12490, n12492 );
nor U91145 ( n12492, n12493, n12494 );
nor U91146 ( n12490, n12505, n12507 );
nand U91147 ( n12494, n12495, n12497 );
nand U91148 ( n47882, n54525, n54526 );
nor U91149 ( n54525, n54541, n54542 );
nor U91150 ( n54526, n54527, n54528 );
nand U91151 ( n54541, n54549, n54550 );
nand U91152 ( n13714, n76724, n12385 );
nand U91153 ( n32426, n32427, n32428 );
nand U91154 ( n32428, n32429, n76480 );
nand U91155 ( n32427, n76776, n32430 );
nor U91156 ( n11292, n12, n10785 );
nor U91157 ( n10625, n12, n9897 );
buf U91158 ( n76778, n3058 );
buf U91159 ( n76712, n5659 );
buf U91160 ( n76760, n3902 );
buf U91161 ( n76693, n6534 );
buf U91162 ( n76664, n7433 );
nand U91163 ( n54342, n7794, n7815 );
nand U91164 ( n14670, n21452, n21453 );
nor U91165 ( n21452, n21468, n21469 );
nor U91166 ( n21453, n21454, n21455 );
nand U91167 ( n21468, n21476, n21477 );
nand U91168 ( n21385, n5144, n5158 );
nand U91169 ( n10697, n21422, n21423 );
nor U91170 ( n21422, n21438, n21439 );
nor U91171 ( n21423, n21424, n21425 );
nand U91172 ( n21438, n21446, n21447 );
nand U91173 ( n42964, n42973, n42829 );
nand U91174 ( n42973, n42974, n76676 );
nor U91175 ( n42974, n7933, n42975 );
nor U91176 ( n42975, n42976, n7949 );
nand U91177 ( n43017, n43027, n42829 );
nand U91178 ( n43027, n43028, n76676 );
nor U91179 ( n43028, n7934, n43029 );
nor U91180 ( n43029, n43030, n7948 );
nand U91181 ( n42848, n42858, n42829 );
nand U91182 ( n42858, n42859, n76676 );
nor U91183 ( n42859, n7930, n42860 );
nor U91184 ( n42860, n42861, n7953 );
nand U91185 ( n43173, n43183, n42829 );
nand U91186 ( n43183, n43184, n76676 );
nor U91187 ( n43184, n7938, n43185 );
nor U91188 ( n43185, n43186, n43187 );
nand U91189 ( n42531, n42546, n42547 );
nand U91190 ( n42547, n42548, n76862 );
nand U91191 ( n42546, n42551, n76675 );
nor U91192 ( n42548, n42497, n42549 );
nand U91193 ( n21389, n5144, n5160 );
not U91194 ( n3155, n32864 );
buf U91195 ( n76456, n76453 );
nand U91196 ( n14652, n21542, n21543 );
nor U91197 ( n21542, n21558, n21559 );
nor U91198 ( n21543, n21544, n21545 );
nand U91199 ( n21558, n21566, n21567 );
nand U91200 ( n45799, n45816, n45817 );
nand U91201 ( n45817, n7430, n7962 );
nand U91202 ( n45816, n76665, n7972 );
nand U91203 ( n67301, n67302, n67226 );
nand U91204 ( n67302, n829, n67217 );
not U91205 ( n3062, n31848 );
buf U91206 ( n76731, n4789 );
nand U91207 ( n21359, n5139, n5160 );
nand U91208 ( n33230, n32283, n76774 );
nor U91209 ( n71354, n1239, n71325 );
nor U91210 ( n71044, n1218, n71311 );
nand U91211 ( n13502, n12292, n76727 );
nand U91212 ( n46950, n45971, n76660 );
nand U91213 ( n67985, n66922, n76708 );
nand U91214 ( n25982, n25046, n76754 );
nand U91215 ( n59120, n58181, n76687 );
nor U91216 ( n16145, n14845, n16130 );
nor U91217 ( n15720, n14845, n15712 );
nor U91218 ( n15189, n14845, n15180 );
nor U91219 ( n15088, n14845, n15073 );
nor U91220 ( n14978, n14845, n14969 );
not U91221 ( n3905, n24634 );
not U91222 ( n5663, n66471 );
not U91223 ( n6538, n57766 );
nand U91224 ( n32203, n32204, n32205 );
nand U91225 ( n32205, n76480, n32206 );
nand U91226 ( n32204, n76785, n32207 );
nand U91227 ( n12189, n12190, n12192 );
nand U91228 ( n12192, n76607, n12193 );
nand U91229 ( n12190, n76738, n12194 );
nand U91230 ( n45898, n45899, n45900 );
nand U91231 ( n45900, n76346, n45901 );
nand U91232 ( n45899, n76671, n45902 );
nand U91233 ( n12060, n12082, n12083 );
nand U91234 ( n12083, n4787, n5307 );
nand U91235 ( n12082, n76732, n5317 );
nand U91236 ( n67217, n838, n842 );
nand U91237 ( n66849, n66850, n66851 );
nand U91238 ( n66851, n76202, n66852 );
nand U91239 ( n66850, n76719, n66853 );
nand U91240 ( n24973, n24974, n24975 );
nand U91241 ( n24975, n76526, n24976 );
nand U91242 ( n24974, n76767, n24977 );
nand U91243 ( n58108, n58109, n58110 );
nand U91244 ( n58110, n76268, n58111 );
nand U91245 ( n58109, n76700, n58112 );
not U91246 ( n7437, n45629 );
nand U91247 ( n40696, n41454, n41455 );
and U91248 ( n41454, n41068, n41067 );
nand U91249 ( n41455, n41312, n76925 );
not U91250 ( n4793, n12223 );
nor U91251 ( n32570, n32562, n32571 );
nand U91252 ( n4466, n32567, n32568 );
nor U91253 ( n32567, n32580, n32581 );
nor U91254 ( n32568, n32569, n32570 );
nor U91255 ( n32580, n3243, n32566 );
nand U91256 ( n67103, n67104, n67105 );
nand U91257 ( n67104, n76719, n67107 );
nand U91258 ( n67105, n67106, n76710 );
nand U91259 ( n25205, n25206, n25207 );
nand U91260 ( n25206, n76767, n25209 );
nand U91261 ( n25207, n25208, n76758 );
nand U91262 ( n58341, n58342, n58343 );
nand U91263 ( n58342, n76700, n58345 );
nand U91264 ( n58343, n58344, n76691 );
nand U91265 ( n46139, n46140, n46141 );
nand U91266 ( n46140, n76671, n46143 );
nand U91267 ( n46141, n46142, n76662 );
nand U91268 ( n32447, n32448, n32449 );
nand U91269 ( n32448, n76785, n32451 );
nand U91270 ( n32449, n32450, n76776 );
nand U91271 ( n49449, n54329, n54330 );
nor U91272 ( n54329, n54352, n54353 );
nor U91273 ( n54330, n54331, n54332 );
nand U91274 ( n54352, n54364, n54365 );
nor U91275 ( n25328, n25320, n25329 );
nor U91276 ( n67335, n67327, n67336 );
nor U91277 ( n58467, n58459, n58468 );
nand U91278 ( n6711, n25325, n25326 );
nor U91279 ( n25325, n25338, n25339 );
nor U91280 ( n25326, n25327, n25328 );
nor U91281 ( n25338, n4068, n25324 );
nand U91282 ( n11201, n67332, n67333 );
nor U91283 ( n67332, n67345, n67346 );
nor U91284 ( n67333, n67334, n67335 );
nor U91285 ( n67345, n5843, n67331 );
nand U91286 ( n13446, n58464, n58465 );
nor U91287 ( n58464, n58477, n58478 );
nor U91288 ( n58465, n58466, n58467 );
nor U91289 ( n58477, n6700, n58463 );
not U91290 ( n3138, n32386 );
and U91291 ( n32494, n32476, n76778 );
not U91292 ( n7524, n46085 );
nand U91293 ( n40849, n40850, n40851 );
nand U91294 ( n40851, n583, n40852 );
nand U91295 ( n40850, n1788, n40714 );
nand U91296 ( n41305, n41306, n41307 );
nand U91297 ( n41307, n583, n40834 );
nand U91298 ( n41306, n1785, n40714 );
nand U91299 ( n40947, n40948, n40949 );
nand U91300 ( n40949, n583, n40950 );
nand U91301 ( n40948, n1784, n40714 );
nand U91302 ( n41021, n41022, n41023 );
nand U91303 ( n41023, n583, n41024 );
nand U91304 ( n41022, n1783, n40714 );
nand U91305 ( n41131, n41132, n41133 );
nand U91306 ( n41133, n583, n41134 );
nand U91307 ( n41132, n1780, n40714 );
nand U91308 ( n41087, n41088, n41089 );
nand U91309 ( n41089, n583, n41090 );
nand U91310 ( n41088, n1778, n40714 );
not U91311 ( n603, n41312 );
and U91312 ( n67150, n67132, n76712 );
and U91313 ( n25252, n25234, n76760 );
and U91314 ( n58388, n58370, n76693 );
and U91315 ( n46186, n46168, n76664 );
not U91316 ( n5739, n67049 );
not U91317 ( n4879, n12427 );
not U91318 ( n3982, n25149 );
not U91319 ( n6614, n58287 );
nor U91320 ( n46274, n46266, n46275 );
nand U91321 ( n15691, n46271, n46272 );
nor U91322 ( n46271, n46284, n46285 );
nor U91323 ( n46272, n46273, n46274 );
nor U91324 ( n46284, n7630, n46270 );
nor U91325 ( n11513, n7, n11594 );
nand U91326 ( n16448, n21346, n21347 );
nor U91327 ( n21346, n21369, n21370 );
nor U91328 ( n21347, n21348, n21349 );
nand U91329 ( n21369, n21381, n21382 );
nand U91330 ( n66997, n784, n40784 );
nand U91331 ( n66345, n784, n41198 );
nand U91332 ( n12382, n12383, n12384 );
nand U91333 ( n12383, n9025, n12118 );
nand U91334 ( n12384, n76729, n12385 );
and U91335 ( n12553, n12530, n76731 );
nand U91336 ( n66422, n784, n40984 );
nand U91337 ( n13749, n76724, n12419 );
nor U91338 ( n11302, n7, n10785 );
nor U91339 ( n10678, n7, n9897 );
nand U91340 ( n66723, n784, n41036 );
nand U91341 ( n66272, n784, n40690 );
nand U91342 ( n33124, n3103, n32206 );
nor U91343 ( n12657, n12638, n12658 );
nand U91344 ( n13369, n4848, n12193 );
nand U91345 ( n8956, n12653, n12654 );
nor U91346 ( n12653, n12669, n12670 );
nor U91347 ( n12654, n12655, n12657 );
nor U91348 ( n12669, n4977, n12643 );
nand U91349 ( n65922, n784, n41145 );
nand U91350 ( n46833, n7490, n45901 );
nand U91351 ( n39568, n2073, n36797 );
nand U91352 ( n67880, n5704, n66852 );
nand U91353 ( n25877, n3947, n24976 );
nand U91354 ( n59015, n6579, n58111 );
nand U91355 ( n40085, n2073, n36462 );
nand U91356 ( n40213, n2073, n36589 );
nand U91357 ( n39080, n2073, n36925 );
nand U91358 ( n40136, n2073, n36286 );
nand U91359 ( n40043, n2073, n36667 );
nand U91360 ( n39510, n2073, n36398 );
nand U91361 ( n38963, n2073, n36442 );
nand U91362 ( n39439, n2073, n36702 );
nand U91363 ( n39763, n2073, n36961 );
nand U91364 ( n39819, n2073, n36322 );
nand U91365 ( n39920, n2073, n36532 );
nand U91366 ( n41010, n1774, n40696 );
nand U91367 ( n41453, n1790, n40696 );
nand U91368 ( n41118, n1799, n40696 );
nand U91369 ( n41149, n1797, n40696 );
nand U91370 ( n41058, n1794, n40696 );
nand U91371 ( n40695, n1792, n40696 );
nand U91372 ( n40988, n1812, n40696 );
nand U91373 ( n39330, n2073, n36747 );
nand U91374 ( n39385, n2073, n36512 );
nand U91375 ( n32486, n32487, n32488 );
nand U91376 ( n32488, n76481, n32489 );
nand U91377 ( n32487, n32490, n76776 );
nand U91378 ( n39850, n38866, n38865 );
nand U91379 ( n32542, n32532, n32543 );
nand U91380 ( n32543, n76776, n32544 );
nor U91381 ( n41446, n812, n617 );
nand U91382 ( n67198, n67188, n67199 );
nand U91383 ( n67199, n76710, n67200 );
nand U91384 ( n46246, n46236, n46247 );
nand U91385 ( n46247, n76662, n46248 );
nand U91386 ( n25300, n25290, n25301 );
nand U91387 ( n25301, n76758, n25302 );
nand U91388 ( n58439, n58426, n58440 );
nand U91389 ( n58440, n76691, n58441 );
nand U91390 ( n32517, n32518, n32519 );
nand U91391 ( n32518, n76786, n32521 );
nand U91392 ( n32519, n76776, n32520 );
nand U91393 ( n32466, n32467, n32468 );
nand U91394 ( n32468, n76481, n32469 );
nand U91395 ( n32467, n76776, n32470 );
nand U91396 ( n32279, n32280, n32281 );
nand U91397 ( n32281, n32282, n76480 );
nand U91398 ( n32280, n32283, n76784 );
nand U91399 ( n32534, n32535, n32536 );
nand U91400 ( n32535, n32538, n76784 );
nand U91401 ( n32536, n76776, n32537 );
nand U91402 ( n12287, n12288, n12289 );
nand U91403 ( n12289, n12290, n76607 );
nand U91404 ( n12288, n12292, n76737 );
nand U91405 ( n45967, n45968, n45969 );
nand U91406 ( n45969, n45970, n76346 );
nand U91407 ( n45968, n45971, n76670 );
nand U91408 ( n66918, n66919, n66920 );
nand U91409 ( n66920, n66921, n76202 );
nand U91410 ( n66919, n66922, n76718 );
nand U91411 ( n25042, n25043, n25044 );
nand U91412 ( n25044, n25045, n76526 );
nand U91413 ( n25043, n25046, n76766 );
nand U91414 ( n58177, n58178, n58179 );
nand U91415 ( n58179, n58180, n76268 );
nand U91416 ( n58178, n58181, n76699 );
nand U91417 ( n67142, n67143, n67144 );
nand U91418 ( n67144, n76203, n67145 );
nand U91419 ( n67143, n67146, n76710 );
nand U91420 ( n25244, n25245, n25246 );
nand U91421 ( n25246, n76527, n25247 );
nand U91422 ( n25245, n25248, n76758 );
nand U91423 ( n58380, n58381, n58382 );
nand U91424 ( n58382, n76269, n58383 );
nand U91425 ( n58381, n58384, n76691 );
nand U91426 ( n32173, n32177, n76480 );
and U91427 ( n32177, n3170, n32178 );
nand U91428 ( n12152, n12157, n76607 );
and U91429 ( n12157, n4906, n12158 );
nand U91430 ( n67173, n67174, n67175 );
nand U91431 ( n67174, n76720, n67177 );
nand U91432 ( n67175, n76710, n67176 );
nand U91433 ( n25275, n25276, n25277 );
nand U91434 ( n25276, n76768, n25279 );
nand U91435 ( n25277, n76758, n25278 );
nand U91436 ( n58411, n58412, n58413 );
nand U91437 ( n58412, n76701, n58415 );
nand U91438 ( n58413, n76691, n58414 );
nand U91439 ( n67122, n67123, n67124 );
nand U91440 ( n67124, n76203, n67125 );
nand U91441 ( n67123, n76710, n67126 );
nand U91442 ( n25224, n25225, n25226 );
nand U91443 ( n25226, n76527, n25227 );
nand U91444 ( n25225, n76758, n25228 );
nand U91445 ( n58360, n58361, n58362 );
nand U91446 ( n58362, n76269, n58363 );
nand U91447 ( n58361, n76691, n58364 );
nand U91448 ( n45868, n45872, n76346 );
and U91449 ( n45872, n7555, n45873 );
nand U91450 ( n46178, n46179, n46180 );
nand U91451 ( n46180, n76347, n46181 );
nand U91452 ( n46179, n46182, n76662 );
nand U91453 ( n67190, n67191, n67192 );
nand U91454 ( n67191, n67194, n76718 );
nand U91455 ( n67192, n76710, n67193 );
nand U91456 ( n25292, n25293, n25294 );
nand U91457 ( n25293, n25296, n76766 );
nand U91458 ( n25294, n76758, n25295 );
nand U91459 ( n58428, n58429, n58430 );
nand U91460 ( n58429, n58432, n76699 );
nand U91461 ( n58430, n76691, n58431 );
nand U91462 ( n66819, n66823, n76202 );
and U91463 ( n66823, n5769, n66824 );
nand U91464 ( n24943, n24947, n76526 );
and U91465 ( n24947, n4010, n24948 );
nand U91466 ( n58078, n58082, n76268 );
and U91467 ( n58082, n6643, n58083 );
not U91468 ( n872, n43880 );
nand U91469 ( n42686, n42431, n42433 );
not U91470 ( n890, n42959 );
nand U91471 ( n46158, n46159, n46160 );
nand U91472 ( n46160, n76347, n46161 );
nand U91473 ( n46159, n76662, n46162 );
nand U91474 ( n46209, n46210, n46211 );
nand U91475 ( n46210, n76672, n46213 );
nand U91476 ( n46211, n76662, n46212 );
nand U91477 ( n12613, n12600, n12614 );
nand U91478 ( n12614, n76730, n12615 );
nand U91479 ( n46238, n46239, n46240 );
nand U91480 ( n46239, n46242, n76670 );
nand U91481 ( n46240, n76662, n46241 );
nand U91482 ( n40409, n37304, n40325 );
and U91483 ( n37078, n37105, n2087 );
nor U91484 ( n37105, n2083, n37106 );
nand U91485 ( n12497, n12498, n76729 );
nand U91486 ( n41968, n45274, n76925 );
nand U91487 ( n45274, n818, n604 );
nand U91488 ( n12543, n12544, n12545 );
nand U91489 ( n12545, n76608, n12547 );
nand U91490 ( n12544, n12548, n76729 );
not U91491 ( n1274, n50359 );
nand U91492 ( n42677, n42423, n42425 );
not U91493 ( n892, n42955 );
not U91494 ( n875, n43557 );
nand U91495 ( n45199, n42247, n42227 );
nor U91496 ( n33441, n33452, n33453 );
nor U91497 ( n33452, n32714, n33457 );
nor U91498 ( n33453, n32712, n33454 );
nand U91499 ( n33457, n32384, n3174 );
nor U91500 ( n13767, n13780, n13782 );
nor U91501 ( n13780, n13060, n13787 );
nor U91502 ( n13782, n13055, n13783 );
nand U91503 ( n13787, n12424, n4911 );
nor U91504 ( n47161, n47172, n47173 );
nor U91505 ( n47172, n46415, n47177 );
nor U91506 ( n47173, n46413, n47174 );
nand U91507 ( n47177, n46083, n7560 );
not U91508 ( n839, n42287 );
nor U91509 ( n68192, n68203, n68204 );
nor U91510 ( n68203, n67479, n68208 );
nor U91511 ( n68204, n67477, n68205 );
nand U91512 ( n68208, n67047, n5773 );
nor U91513 ( n26191, n26202, n26203 );
nor U91514 ( n26202, n25474, n26207 );
nor U91515 ( n26203, n25472, n26204 );
nand U91516 ( n26207, n25147, n4014 );
nor U91517 ( n59330, n59341, n59342 );
nor U91518 ( n59341, n58611, n59346 );
nor U91519 ( n59342, n58609, n59343 );
nand U91520 ( n59346, n58285, n6647 );
nor U91521 ( n71523, n1222, n71325 );
nand U91522 ( n12468, n12469, n12470 );
nand U91523 ( n12470, n12472, n76607 );
nand U91524 ( n12469, n76730, n12473 );
nand U91525 ( n12582, n12583, n12584 );
nand U91526 ( n12583, n76739, n12587 );
nand U91527 ( n12584, n76730, n12585 );
nand U91528 ( n12603, n12604, n12605 );
nand U91529 ( n12604, n12608, n76737 );
nand U91530 ( n12605, n76730, n12607 );
nand U91531 ( n13847, n76725, n12473 );
nand U91532 ( n12533, n12534, n12535 );
nand U91533 ( n12535, n5289, n12118 );
nand U91534 ( n12534, n76730, n12538 );
not U91535 ( n3040, n32566 );
not U91536 ( n3884, n25324 );
not U91537 ( n7417, n46270 );
not U91538 ( n5642, n67331 );
not U91539 ( n6517, n58463 );
not U91540 ( n2007, n37106 );
nand U91541 ( n33231, n3103, n32282 );
nand U91542 ( n13503, n4848, n12290 );
nand U91543 ( n46951, n7490, n45970 );
nand U91544 ( n67986, n5704, n66921 );
nand U91545 ( n25983, n3947, n25045 );
nand U91546 ( n59121, n6579, n58180 );
nand U91547 ( n32439, n32440, n32441 );
nand U91548 ( n32440, n3543, n32146 );
nand U91549 ( n32441, n32442, n76784 );
buf U91550 ( n76039, n76921 );
nand U91551 ( n67095, n67096, n67097 );
nand U91552 ( n67096, n6158, n66792 );
nand U91553 ( n67097, n67098, n76718 );
nand U91554 ( n46131, n46132, n46133 );
nand U91555 ( n46132, n7945, n45841 );
nand U91556 ( n46133, n46134, n76670 );
nand U91557 ( n25197, n25198, n25199 );
nand U91558 ( n25198, n4380, n24914 );
nand U91559 ( n25199, n25200, n76766 );
nand U91560 ( n58333, n58334, n58335 );
nand U91561 ( n58334, n7013, n58051 );
nand U91562 ( n58335, n58336, n76699 );
nand U91563 ( n32375, n32381, n32382 );
nand U91564 ( n32382, n32383, n76480 );
nand U91565 ( n32381, n32385, n76784 );
and U91566 ( n32383, n3174, n32384 );
nand U91567 ( n67038, n67044, n67045 );
nand U91568 ( n67045, n67046, n76202 );
nand U91569 ( n67044, n67048, n76718 );
and U91570 ( n67046, n5773, n67047 );
nand U91571 ( n46074, n46080, n46081 );
nand U91572 ( n46081, n46082, n76346 );
nand U91573 ( n46080, n46084, n76670 );
and U91574 ( n46082, n7560, n46083 );
nand U91575 ( n25138, n25144, n25145 );
nand U91576 ( n25145, n25146, n76526 );
nand U91577 ( n25144, n25148, n76766 );
and U91578 ( n25146, n4014, n25147 );
nand U91579 ( n58276, n58282, n58283 );
nand U91580 ( n58283, n58284, n76268 );
nand U91581 ( n58282, n58286, n76699 );
and U91582 ( n58284, n6647, n58285 );
nand U91583 ( n32499, n32500, n32501 );
nand U91584 ( n32501, n29931, n32146 );
nand U91585 ( n32500, n32503, n76784 );
nand U91586 ( n67155, n67156, n67157 );
nand U91587 ( n67157, n63887, n66792 );
nand U91588 ( n67156, n67159, n76718 );
nand U91589 ( n25257, n25258, n25259 );
nand U91590 ( n25259, n22608, n24914 );
nand U91591 ( n25258, n25261, n76766 );
nand U91592 ( n58393, n58394, n58395 );
nand U91593 ( n58395, n55721, n58051 );
nand U91594 ( n58394, n58397, n76699 );
nand U91595 ( n46191, n46192, n46193 );
nand U91596 ( n46193, n43188, n45841 );
nand U91597 ( n46192, n46195, n76670 );
not U91598 ( n834, n61176 );
nand U91599 ( n32478, n32479, n32480 );
nand U91600 ( n32479, n3542, n32146 );
nand U91601 ( n32480, n76786, n32481 );
nand U91602 ( n67134, n67135, n67136 );
nand U91603 ( n67135, n6157, n66792 );
nand U91604 ( n67136, n76720, n67137 );
nand U91605 ( n46170, n46171, n46172 );
nand U91606 ( n46171, n7944, n45841 );
nand U91607 ( n46172, n76672, n46173 );
nand U91608 ( n25236, n25237, n25238 );
nand U91609 ( n25237, n4379, n24914 );
nand U91610 ( n25238, n76768, n25239 );
nand U91611 ( n58372, n58373, n58374 );
nand U91612 ( n58373, n7012, n58051 );
nand U91613 ( n58374, n76701, n58375 );
not U91614 ( n4773, n12643 );
nand U91615 ( n40691, n41448, n41447 );
nand U91616 ( n12484, n12485, n12487 );
nand U91617 ( n12485, n5290, n12118 );
nand U91618 ( n12487, n12488, n76737 );
buf U91619 ( n76516, n76513 );
buf U91620 ( n76512, n76509 );
not U91621 ( n76476, n76477 );
nand U91622 ( n12495, n76738, n12499 );
buf U91623 ( n76511, n76509 );
buf U91624 ( n76510, n76509 );
not U91625 ( n4762, n8559 );
nand U91626 ( n9437, n11749, n4845 );
and U91627 ( n8263, n4819, n9434 );
nand U91628 ( n9434, n9435, n9437 );
nand U91629 ( n12559, n12560, n12562 );
nand U91630 ( n12562, n9220, n12118 );
nand U91631 ( n12560, n12564, n76737 );
and U91632 ( n32563, n32565, n76784 );
and U91633 ( n67328, n67330, n76718 );
and U91634 ( n46267, n46269, n76670 );
and U91635 ( n25321, n25323, n76766 );
and U91636 ( n58460, n58462, n76699 );
not U91637 ( n7407, n42617 );
nand U91638 ( n43376, n45522, n7488 );
and U91639 ( n42323, n7463, n43374 );
nand U91640 ( n43374, n43375, n43376 );
nand U91641 ( n21195, n14767, n21202 );
nand U91642 ( n12518, n12519, n12520 );
nand U91643 ( n12520, n76608, n12522 );
nand U91644 ( n12519, n76739, n12523 );
nor U91645 ( n32553, n29162, n3063 );
nor U91646 ( n25311, n21849, n3907 );
nor U91647 ( n67209, n62884, n5664 );
nor U91648 ( n58450, n54940, n6539 );
nor U91649 ( n46257, n42375, n7438 );
and U91650 ( n12639, n12642, n76737 );
nand U91651 ( n30405, n3077, n30409 );
nand U91652 ( n30409, n30410, n30411 );
nand U91653 ( n30411, n30412, n3168 );
nand U91654 ( n30410, n3387, n30414 );
nand U91655 ( n64564, n5678, n64568 );
nand U91656 ( n64568, n64569, n64570 );
nand U91657 ( n64570, n64571, n5767 );
nand U91658 ( n64569, n6002, n64573 );
nand U91659 ( n43722, n7463, n43726 );
nand U91660 ( n43726, n43727, n43728 );
nand U91661 ( n43728, n43729, n7553 );
nand U91662 ( n43727, n7789, n43731 );
nand U91663 ( n9800, n4819, n9805 );
nand U91664 ( n9805, n9807, n9808 );
nand U91665 ( n9808, n9809, n4904 );
nand U91666 ( n9807, n5134, n9812 );
nand U91667 ( n23074, n3920, n23078 );
nand U91668 ( n23078, n23079, n23080 );
nand U91669 ( n23080, n23081, n4008 );
nand U91670 ( n23079, n4224, n23083 );
nand U91671 ( n56195, n6553, n56199 );
nand U91672 ( n56199, n56200, n56201 );
nand U91673 ( n56201, n56202, n6640 );
nand U91674 ( n56200, n6857, n56204 );
nand U91675 ( n36680, n37078, n36943 );
nand U91676 ( n13865, n4848, n12472 );
nor U91677 ( n12627, n8285, n4794 );
nand U91678 ( n76104, n41448, n41447 );
nand U91679 ( n76103, n41448, n41447 );
nor U91680 ( n17401, n76929, n76788 );
not U91681 ( n5134, n14649 );
and U91682 ( n41447, n41474, n839 );
nor U91683 ( n41474, n829, n41445 );
xnor U91684 ( n16525, n16528, n16529 );
nand U91685 ( n9435, n11749, n14635 );
nand U91686 ( n13904, n76724, n12498 );
nand U91687 ( n54990, n830, n812 );
nand U91688 ( n43375, n45522, n47869 );
nor U91689 ( n71048, n1218, n71325 );
and U91690 ( n37603, n38103, n76920 );
nand U91691 ( n38103, n2198, n2088 );
not U91692 ( n7789, n47880 );
not U91693 ( n3032, n29274 );
not U91694 ( n3875, n21957 );
not U91695 ( n5633, n63041 );
not U91696 ( n6508, n55069 );
nand U91697 ( n30103, n31823, n3100 );
nand U91698 ( n22782, n24607, n3944 );
nand U91699 ( n64120, n66415, n5702 );
nand U91700 ( n55896, n57739, n6577 );
and U91701 ( n29144, n3077, n30101 );
nand U91702 ( n30101, n30102, n30103 );
and U91703 ( n62811, n5678, n64118 );
nand U91704 ( n64118, n64119, n64120 );
and U91705 ( n21829, n3920, n22780 );
nand U91706 ( n22780, n22781, n22782 );
and U91707 ( n54905, n6553, n55894 );
nand U91708 ( n55894, n55895, n55896 );
nand U91709 ( n63199, n63064, n63200 );
nand U91710 ( n63200, n76875, n6324 );
nand U91711 ( n29436, n29297, n29437 );
nand U91712 ( n29437, n76901, n3690 );
nand U91713 ( n22117, n21982, n22118 );
nand U91714 ( n22118, n76910, n4584 );
nand U91715 ( n55227, n55092, n55228 );
nand U91716 ( n55228, n76884, n7217 );
nand U91717 ( n63367, n76875, n6327 );
nand U91718 ( n29538, n76901, n3693 );
nand U91719 ( n22219, n76910, n4587 );
nand U91720 ( n55333, n76884, n7219 );
buf U91721 ( n76910, n170 );
buf U91722 ( n76901, n204 );
buf U91723 ( n76875, n475 );
buf U91724 ( n76884, n443 );
nand U91725 ( n63533, n63064, n63534 );
nand U91726 ( n63534, n76875, n6329 );
nand U91727 ( n29634, n29297, n29635 );
nand U91728 ( n29635, n76901, n3695 );
nand U91729 ( n22313, n21982, n22314 );
nand U91730 ( n22314, n76910, n4589 );
nand U91731 ( n55425, n55092, n55426 );
nand U91732 ( n55426, n76884, n7222 );
nand U91733 ( n63239, n63064, n63240 );
nand U91734 ( n63240, n76875, n6325 );
nand U91735 ( n29476, n29297, n29477 );
nand U91736 ( n29477, n76901, n3692 );
nand U91737 ( n22157, n21982, n22158 );
nand U91738 ( n22158, n76910, n4585 );
nand U91739 ( n55271, n55092, n55272 );
nand U91740 ( n55272, n76884, n7218 );
nand U91741 ( n63815, n76875, n6334 );
nand U91742 ( n29859, n76901, n3700 );
nand U91743 ( n22536, n76910, n4594 );
nand U91744 ( n55649, n76884, n7227 );
nand U91745 ( n63148, n76875, n6323 );
nand U91746 ( n29385, n76901, n3689 );
nand U91747 ( n22066, n76910, n4583 );
nand U91748 ( n55176, n76884, n7215 );
nand U91749 ( n63496, n63064, n63497 );
nand U91750 ( n63497, n76875, n6328 );
nand U91751 ( n63598, n63064, n63599 );
nand U91752 ( n63599, n76875, n6330 );
nand U91753 ( n63651, n63064, n63652 );
nand U91754 ( n63652, n76875, n6332 );
nand U91755 ( n63763, n63064, n63764 );
nand U91756 ( n63764, n76875, n6333 );
nand U91757 ( n63868, n63064, n63869 );
nand U91758 ( n63869, n76875, n6335 );
nand U91759 ( n63918, n63064, n63919 );
nand U91760 ( n63919, n76875, n6337 );
nand U91761 ( n29597, n29297, n29598 );
nand U91762 ( n29598, n76901, n3694 );
nand U91763 ( n29699, n29297, n29700 );
nand U91764 ( n29700, n76901, n3697 );
nand U91765 ( n29752, n29297, n29753 );
nand U91766 ( n29753, n76901, n3698 );
nand U91767 ( n29803, n29297, n29804 );
nand U91768 ( n29804, n76901, n3699 );
nand U91769 ( n29912, n29297, n29913 );
nand U91770 ( n29913, n76901, n3702 );
nand U91771 ( n29962, n29297, n29963 );
nand U91772 ( n29963, n76901, n3703 );
nand U91773 ( n22431, n21982, n22432 );
nand U91774 ( n22432, n76910, n4592 );
nand U91775 ( n22589, n21982, n22590 );
nand U91776 ( n22590, n76910, n4595 );
nand U91777 ( n22276, n21982, n22277 );
nand U91778 ( n22277, n76910, n4588 );
nand U91779 ( n22378, n21982, n22379 );
nand U91780 ( n22379, n76910, n4590 );
nand U91781 ( n22482, n21982, n22483 );
nand U91782 ( n22483, n76910, n4593 );
nand U91783 ( n22639, n21982, n22640 );
nand U91784 ( n22640, n76910, n4597 );
nand U91785 ( n55546, n55092, n55547 );
nand U91786 ( n55547, n76884, n7224 );
nand U91787 ( n55702, n55092, n55703 );
nand U91788 ( n55703, n76884, n7228 );
nand U91789 ( n55388, n55092, n55389 );
nand U91790 ( n55389, n76884, n7220 );
nand U91791 ( n55490, n55092, n55491 );
nand U91792 ( n55491, n76884, n7223 );
nand U91793 ( n55597, n55092, n55598 );
nand U91794 ( n55598, n76884, n7225 );
nand U91795 ( n55752, n55092, n55753 );
nand U91796 ( n55753, n76884, n7229 );
buf U91797 ( n76900, n204 );
nor U91798 ( n26896, n26909, n26910 );
nor U91799 ( n26909, n26911, n24605 );
nor U91800 ( n26911, n26912, n26913 );
nor U91801 ( n26912, n26916, n24601 );
nor U91802 ( n60036, n60049, n60050 );
nor U91803 ( n60049, n60051, n57737 );
nor U91804 ( n60051, n60052, n60053 );
nor U91805 ( n60052, n60056, n57733 );
buf U91806 ( n76519, n25360 );
buf U91807 ( n76261, n58497 );
buf U91808 ( n76907, n179 );
buf U91809 ( n76881, n450 );
buf U91810 ( n76909, n170 );
buf U91811 ( n76874, n475 );
buf U91812 ( n76883, n443 );
nor U91813 ( n34141, n34154, n34155 );
nor U91814 ( n34154, n34156, n31821 );
nor U91815 ( n34156, n34157, n34158 );
nor U91816 ( n34157, n34161, n31817 );
buf U91817 ( n76468, n32600 );
buf U91818 ( n76898, n213 );
nor U91819 ( n68895, n68908, n68909 );
nor U91820 ( n68908, n68910, n66413 );
nor U91821 ( n68910, n68911, n68912 );
nor U91822 ( n68911, n68915, n66409 );
buf U91823 ( n76195, n67365 );
buf U91824 ( n76872, n484 );
buf U91825 ( n76897, n213 );
buf U91826 ( n76871, n484 );
buf U91827 ( n76906, n179 );
buf U91828 ( n76880, n450 );
not U91829 ( n215, n32592 );
not U91830 ( n487, n67357 );
not U91831 ( n182, n25352 );
not U91832 ( n453, n58489 );
buf U91833 ( n76908, n179 );
buf U91834 ( n76882, n450 );
buf U91835 ( n76899, n213 );
nor U91836 ( n35734, n35699, n35735 );
nor U91837 ( n35735, n35736, n35737 );
nand U91838 ( n35736, n34136, n31822 );
nand U91839 ( n35737, n34061, n34134 );
nor U91840 ( n28555, n28520, n28556 );
nor U91841 ( n28556, n28557, n28558 );
nand U91842 ( n28557, n26891, n24606 );
nand U91843 ( n28558, n26816, n26889 );
nor U91844 ( n70460, n70425, n70461 );
nor U91845 ( n70461, n70462, n70463 );
nand U91846 ( n70462, n68890, n66414 );
nand U91847 ( n70463, n68815, n68888 );
nor U91848 ( n61860, n61825, n61861 );
nor U91849 ( n61861, n61862, n61863 );
nand U91850 ( n61862, n60031, n57738 );
nand U91851 ( n61863, n59956, n60029 );
buf U91852 ( n76873, n484 );
nor U91853 ( n54232, n54197, n54233 );
nor U91854 ( n54233, n54234, n54235 );
nand U91855 ( n54234, n47870, n45521 );
nand U91856 ( n54235, n47795, n47868 );
not U91857 ( n5132, n14658 );
buf U91858 ( n76911, n170 );
buf U91859 ( n76902, n204 );
buf U91860 ( n76876, n475 );
buf U91861 ( n76885, n443 );
nand U91862 ( n10478, n9965, n10529 );
nand U91863 ( n10529, n76892, n10475 );
nand U91864 ( n44306, n43889, n44347 );
nand U91865 ( n44347, n76866, n44304 );
and U91866 ( n9965, n4819, n11314 );
nand U91867 ( n11314, n225, n11315 );
nand U91868 ( n11315, n11317, n4904 );
not U91869 ( n225, n11318 );
and U91870 ( n43889, n7463, n44993 );
nand U91871 ( n44993, n497, n44994 );
nand U91872 ( n44994, n44995, n7553 );
not U91873 ( n497, n44996 );
nand U91874 ( n11318, n21318, n21319 );
nand U91875 ( n21318, n12777, n5134 );
or U91876 ( n21319, n9435, n227 );
nand U91877 ( n44996, n54301, n54302 );
nand U91878 ( n54301, n46349, n7789 );
or U91879 ( n54302, n43375, n498 );
nand U91880 ( n63962, n63064, n63963 );
nand U91881 ( n63963, n76876, n6338 );
nand U91882 ( n30006, n29297, n30007 );
nand U91883 ( n30007, n76902, n3704 );
nand U91884 ( n22683, n21982, n22684 );
nand U91885 ( n22684, n76911, n4598 );
nand U91886 ( n55799, n55092, n55800 );
nand U91887 ( n55800, n76885, n7230 );
nand U91888 ( n10247, n9965, n10368 );
nand U91889 ( n10368, n76892, n10245 );
nand U91890 ( n44121, n43889, n44218 );
nand U91891 ( n44218, n76866, n44120 );
nand U91892 ( n44448, n43889, n44490 );
nand U91893 ( n44490, n76866, n44447 );
nand U91894 ( n10638, n9965, n10690 );
nand U91895 ( n10690, n76892, n10637 );
nand U91896 ( n9909, n9965, n9967 );
nand U91897 ( n9967, n76893, n9907 );
nand U91898 ( n10069, n9965, n10130 );
nand U91899 ( n10130, n76893, n10068 );
nand U91900 ( n43809, n43889, n43890 );
nand U91901 ( n43890, n76867, n43807 );
nand U91902 ( n43983, n43889, n44028 );
nand U91903 ( n44028, n76867, n43982 );
nand U91904 ( n29296, n29297, n29298 );
nand U91905 ( n29298, n76902, n29269 );
nand U91906 ( n63063, n63064, n63065 );
nand U91907 ( n63065, n76876, n63036 );
nand U91908 ( n55091, n55092, n55093 );
nand U91909 ( n55093, n76885, n55064 );
nand U91910 ( n21981, n21982, n21983 );
nand U91911 ( n21983, n76911, n21952 );
not U91912 ( n3384, n34153 );
not U91913 ( n4222, n26908 );
not U91914 ( n5999, n68907 );
not U91915 ( n6854, n60048 );
and U91916 ( n10999, n9965, n11048 );
nand U91917 ( n11048, n76892, n11002 );
and U91918 ( n44732, n43889, n44771 );
nand U91919 ( n44771, n76866, n44734 );
and U91920 ( n10849, n9965, n10898 );
nand U91921 ( n10898, n76892, n10852 );
and U91922 ( n44612, n43889, n44651 );
nand U91923 ( n44651, n76866, n44614 );
and U91924 ( n11149, n9965, n11219 );
nand U91925 ( n11219, n76893, n11152 );
and U91926 ( n11252, n9965, n11263 );
nand U91927 ( n11263, n76893, n11254 );
and U91928 ( n44866, n43889, n44922 );
nand U91929 ( n44922, n76867, n44868 );
and U91930 ( n44943, n43889, n44952 );
nand U91931 ( n44952, n76867, n44945 );
nand U91932 ( n32525, n32526, n32527 );
nand U91933 ( n32526, n29984, n32146 );
nand U91934 ( n32527, n32528, n76480 );
nand U91935 ( n67181, n67182, n67183 );
nand U91936 ( n67182, n63940, n66792 );
nand U91937 ( n67183, n67184, n76202 );
nand U91938 ( n25283, n25284, n25285 );
nand U91939 ( n25284, n22661, n24914 );
nand U91940 ( n25285, n25286, n76526 );
nand U91941 ( n58419, n58420, n58421 );
nand U91942 ( n58420, n55774, n58051 );
nand U91943 ( n58421, n58422, n76268 );
nand U91944 ( n46229, n46230, n46231 );
nand U91945 ( n46230, n43255, n45841 );
nand U91946 ( n46231, n46232, n76346 );
nand U91947 ( n32399, n32402, n76480 );
nand U91948 ( n67062, n67065, n76202 );
nand U91949 ( n46098, n46101, n76346 );
nand U91950 ( n25164, n25167, n76526 );
nand U91951 ( n58300, n58303, n76268 );
nand U91952 ( n35678, n35782, n35783 );
nor U91953 ( n35783, n35784, n35785 );
nor U91954 ( n35782, n31618, n34155 );
nor U91955 ( n35785, n3130, n34146 );
nand U91956 ( n28499, n28603, n28604 );
nor U91957 ( n28604, n28605, n28606 );
nor U91958 ( n28603, n24322, n26910 );
nor U91959 ( n28606, n3974, n26901 );
nand U91960 ( n70404, n70508, n70509 );
nor U91961 ( n70509, n70510, n70511 );
nor U91962 ( n70508, n65904, n68909 );
nor U91963 ( n70511, n5732, n68900 );
nand U91964 ( n61804, n61908, n61909 );
nor U91965 ( n61909, n61910, n61911 );
nor U91966 ( n61908, n57445, n60050 );
nor U91967 ( n61911, n6607, n60041 );
nand U91968 ( n32507, n32508, n32509 );
nand U91969 ( n32509, n3540, n32146 );
nand U91970 ( n32508, n32511, n76480 );
not U91971 ( n2474, n16763 );
nand U91972 ( n67163, n67164, n67165 );
nand U91973 ( n67165, n6155, n66792 );
nand U91974 ( n67164, n67167, n76202 );
nand U91975 ( n25265, n25266, n25267 );
nand U91976 ( n25267, n4378, n24914 );
nand U91977 ( n25266, n25269, n76526 );
nand U91978 ( n58401, n58402, n58403 );
nand U91979 ( n58403, n7010, n58051 );
nand U91980 ( n58402, n58405, n76268 );
nand U91981 ( n46199, n46200, n46201 );
nand U91982 ( n46201, n7943, n45841 );
nand U91983 ( n46200, n46203, n76346 );
not U91984 ( n7787, n47887 );
and U91985 ( n30142, n3075, n30150 );
nand U91986 ( n30150, n76023, n30144 );
and U91987 ( n43411, n7462, n43419 );
nand U91988 ( n43419, n76007, n43413 );
and U91989 ( n64155, n5677, n64163 );
nand U91990 ( n64163, n75991, n64157 );
and U91991 ( n22817, n3919, n22825 );
nand U91992 ( n22825, n76028, n22819 );
and U91993 ( n55931, n6552, n55939 );
nand U91994 ( n55939, n75999, n55933 );
nand U91995 ( n54176, n54280, n54281 );
nor U91996 ( n54281, n54282, n54283 );
nor U91997 ( n54280, n44996, n47889 );
nor U91998 ( n54283, n7517, n47880 );
and U91999 ( n9480, n4818, n9490 );
nand U92000 ( n9490, n76036, n9483 );
buf U92001 ( n76436, n76433 );
buf U92002 ( n76432, n76429 );
not U92003 ( n76611, n76612 );
nand U92004 ( n12592, n12593, n12594 );
nand U92005 ( n12593, n9287, n12118 );
nand U92006 ( n12594, n12595, n76607 );
buf U92007 ( n76431, n76429 );
buf U92008 ( n76430, n76429 );
nand U92009 ( n12442, n12443, n12444 );
nand U92010 ( n12444, n9080, n12118 );
nand U92011 ( n12443, n12447, n76607 );
nand U92012 ( n12422, n12423, n76607 );
and U92013 ( n12423, n4911, n12424 );
nand U92014 ( n21202, n21297, n21298 );
nor U92015 ( n21298, n21299, n21300 );
nor U92016 ( n21297, n11318, n14660 );
nor U92017 ( n21300, n4872, n14649 );
nand U92018 ( n12569, n12570, n12572 );
nand U92019 ( n12572, n5288, n12118 );
nand U92020 ( n12570, n12574, n76607 );
buf U92021 ( n76481, n31833 );
buf U92022 ( n76527, n24619 );
buf U92023 ( n76347, n45532 );
buf U92024 ( n76203, n66456 );
buf U92025 ( n76269, n57751 );
nand U92026 ( n32452, n76481, n32455 );
nand U92027 ( n67108, n76203, n67111 );
nand U92028 ( n46144, n76347, n46147 );
nand U92029 ( n25210, n76527, n25213 );
nand U92030 ( n58346, n76269, n58349 );
nand U92031 ( n21991, n22005, n22006 );
nand U92032 ( n22005, n22010, n76547 );
nand U92033 ( n22006, n22007, n76909 );
nor U92034 ( n22010, n4359, n22011 );
nand U92035 ( n29310, n29324, n29325 );
nand U92036 ( n29324, n29329, n76494 );
nand U92037 ( n29325, n29326, n76900 );
nor U92038 ( n29329, n3522, n29330 );
nand U92039 ( n63073, n63087, n63088 );
nand U92040 ( n63087, n63092, n76227 );
nand U92041 ( n63088, n63089, n76874 );
nor U92042 ( n63092, n6137, n63093 );
nand U92043 ( n55101, n55115, n55116 );
nand U92044 ( n55115, n55120, n76293 );
nand U92045 ( n55116, n55117, n76883 );
nor U92046 ( n55120, n6992, n55121 );
nor U92047 ( n30110, n30112, n76489 );
nor U92048 ( n43379, n43381, n76363 );
nor U92049 ( n64123, n64125, n76222 );
nor U92050 ( n22785, n22787, n76542 );
nor U92051 ( n55899, n55901, n76284 );
nor U92052 ( n9440, n9443, n76633 );
not U92053 ( n6175, n66831 );
not U92054 ( n3560, n32185 );
not U92055 ( n4398, n24955 );
not U92056 ( n7030, n58090 );
not U92057 ( n6177, n66951 );
not U92058 ( n3562, n32312 );
not U92059 ( n4399, n25075 );
not U92060 ( n7032, n58210 );
nand U92061 ( n63238, n76227, n6140 );
nand U92062 ( n29475, n76494, n3525 );
nand U92063 ( n22156, n76547, n4363 );
nand U92064 ( n55270, n76293, n6995 );
buf U92065 ( n76608, n11762 );
nand U92066 ( n63799, n63775, n63802 );
nand U92067 ( n63802, n63052, n63803 );
nand U92068 ( n63803, n76227, n6149 );
nand U92069 ( n29843, n29815, n29846 );
nand U92070 ( n29846, n29285, n29847 );
nand U92071 ( n29847, n76494, n3534 );
nand U92072 ( n22520, n22496, n22523 );
nand U92073 ( n22523, n21970, n22524 );
nand U92074 ( n22524, n76547, n4372 );
nand U92075 ( n55633, n55609, n55636 );
nand U92076 ( n55636, n55080, n55637 );
nand U92077 ( n55637, n76293, n7004 );
nand U92078 ( n63184, n63168, n63187 );
nand U92079 ( n63187, n63052, n63188 );
nand U92080 ( n63188, n76227, n6139 );
nand U92081 ( n63353, n63342, n63356 );
nand U92082 ( n63356, n63052, n63357 );
nand U92083 ( n63357, n76227, n6142 );
nand U92084 ( n29421, n29405, n29424 );
nand U92085 ( n29424, n29285, n29425 );
nand U92086 ( n29425, n76494, n3524 );
nand U92087 ( n29524, n29513, n29527 );
nand U92088 ( n29527, n29285, n29528 );
nand U92089 ( n29528, n76494, n3527 );
nand U92090 ( n22205, n22194, n22208 );
nand U92091 ( n22208, n21970, n22209 );
nand U92092 ( n22209, n76547, n4364 );
nand U92093 ( n22102, n22086, n22105 );
nand U92094 ( n22105, n21970, n22106 );
nand U92095 ( n22106, n76547, n4362 );
nand U92096 ( n55319, n55308, n55322 );
nand U92097 ( n55322, n55080, n55323 );
nand U92098 ( n55323, n76293, n6997 );
nand U92099 ( n55212, n55196, n55215 );
nand U92100 ( n55215, n55080, n55216 );
nand U92101 ( n55216, n76293, n6994 );
nand U92102 ( n63597, n76227, n6145 );
nand U92103 ( n63762, n76227, n6148 );
nand U92104 ( n63867, n76227, n6150 );
nand U92105 ( n63917, n76227, n6152 );
nand U92106 ( n29698, n76494, n3530 );
nand U92107 ( n29802, n76494, n3533 );
nand U92108 ( n29911, n76494, n3535 );
nand U92109 ( n29961, n76494, n3537 );
nand U92110 ( n22588, n76547, n4373 );
nand U92111 ( n22377, n76547, n4368 );
nand U92112 ( n22481, n76547, n4370 );
nand U92113 ( n22638, n76547, n4374 );
nand U92114 ( n55701, n76293, n7005 );
nand U92115 ( n55489, n76293, n7000 );
nand U92116 ( n55596, n76293, n7003 );
nand U92117 ( n55751, n76293, n7007 );
nand U92118 ( n63495, n76227, n6143 );
nand U92119 ( n63650, n76227, n6147 );
nand U92120 ( n29596, n76494, n3528 );
nand U92121 ( n29751, n76494, n3532 );
nand U92122 ( n22430, n76547, n4369 );
nand U92123 ( n22275, n76547, n4365 );
nand U92124 ( n55545, n76293, n7002 );
nand U92125 ( n55387, n76293, n6998 );
not U92126 ( n245, n48033 );
not U92127 ( n830, n40664 );
nand U92128 ( n42789, n76863, n8108 );
nand U92129 ( n42659, n42524, n42660 );
nand U92130 ( n42660, n76863, n8105 );
not U92131 ( n502, n42495 );
nand U92132 ( n42882, n76863, n8110 );
nand U92133 ( n42724, n76863, n8107 );
nand U92134 ( n43116, n76863, n8115 );
nand U92135 ( n42607, n76863, n8104 );
nand U92136 ( n30160, n3075, n30168 );
nand U92137 ( n30168, n76024, n30169 );
nand U92138 ( n30179, n3075, n30187 );
nand U92139 ( n30187, n76024, n30188 );
nand U92140 ( n30198, n3075, n30210 );
nand U92141 ( n30210, n76024, n30211 );
nand U92142 ( n30221, n3075, n30229 );
nand U92143 ( n30229, n76024, n30230 );
nand U92144 ( n30240, n3075, n30248 );
nand U92145 ( n30248, n76023, n30249 );
nand U92146 ( n30259, n3075, n30267 );
nand U92147 ( n30267, n76023, n30268 );
nand U92148 ( n30278, n3075, n30286 );
nand U92149 ( n30286, n76023, n30287 );
nand U92150 ( n30356, n3075, n30363 );
nand U92151 ( n30363, n76024, n30364 );
not U92152 ( n76620, n11504 );
nand U92153 ( n11504, n4819, n11743 );
nand U92154 ( n11743, n11744, n11745 );
nand U92155 ( n11744, n4878, n11749 );
or U92156 ( n11745, n11747, n11748 );
nand U92157 ( n43462, n7462, n43470 );
nand U92158 ( n43470, n76008, n43471 );
nand U92159 ( n43481, n7462, n43489 );
nand U92160 ( n43489, n76008, n43490 );
nand U92161 ( n43500, n7462, n43508 );
nand U92162 ( n43508, n76008, n43509 );
nand U92163 ( n43519, n7462, n43527 );
nand U92164 ( n43527, n76008, n43528 );
nand U92165 ( n43538, n7462, n43546 );
nand U92166 ( n43546, n76007, n43547 );
nand U92167 ( n43570, n7462, n43578 );
nand U92168 ( n43578, n76007, n43579 );
nand U92169 ( n64173, n5677, n64181 );
nand U92170 ( n64181, n75992, n64182 );
nand U92171 ( n64245, n5677, n64253 );
nand U92172 ( n64253, n75992, n64254 );
nand U92173 ( n64264, n5677, n64272 );
nand U92174 ( n64272, n75992, n64273 );
nand U92175 ( n64283, n5677, n64291 );
nand U92176 ( n64291, n75992, n64292 );
nand U92177 ( n64302, n5677, n64310 );
nand U92178 ( n64310, n75991, n64311 );
nand U92179 ( n64321, n5677, n64329 );
nand U92180 ( n64329, n75991, n64330 );
nand U92181 ( n64401, n5677, n64409 );
nand U92182 ( n64409, n75991, n64410 );
nand U92183 ( n22835, n3919, n22843 );
nand U92184 ( n22843, n76029, n22844 );
nand U92185 ( n22854, n3919, n22862 );
nand U92186 ( n22862, n76029, n22863 );
nand U92187 ( n22875, n3919, n22883 );
nand U92188 ( n22883, n76029, n22884 );
nand U92189 ( n22894, n3919, n22902 );
nand U92190 ( n22902, n76029, n22903 );
nand U92191 ( n22913, n3919, n22921 );
nand U92192 ( n22921, n76028, n22922 );
nand U92193 ( n22932, n3919, n22940 );
nand U92194 ( n22940, n76028, n22941 );
nand U92195 ( n22951, n3919, n22959 );
nand U92196 ( n22959, n76028, n22960 );
nand U92197 ( n23027, n3919, n23034 );
nand U92198 ( n23034, n76029, n23035 );
nand U92199 ( n9503, n4818, n9513 );
nand U92200 ( n9513, n76037, n9514 );
nand U92201 ( n9527, n4818, n9537 );
nand U92202 ( n9537, n76037, n9538 );
nand U92203 ( n9550, n4818, n9560 );
nand U92204 ( n9560, n76037, n9562 );
nand U92205 ( n9574, n4818, n9584 );
nand U92206 ( n9584, n76037, n9585 );
nand U92207 ( n9597, n4818, n9607 );
nand U92208 ( n9607, n76036, n9608 );
nand U92209 ( n9644, n4818, n9658 );
nand U92210 ( n9658, n76036, n9659 );
nand U92211 ( n9740, n4818, n9749 );
nand U92212 ( n9749, n76037, n9750 );
nand U92213 ( n64475, n5677, n64482 );
nand U92214 ( n64482, n75992, n64483 );
nand U92215 ( n55949, n6552, n55960 );
nand U92216 ( n55960, n76000, n55961 );
nand U92217 ( n55971, n6552, n55979 );
nand U92218 ( n55979, n76000, n55980 );
nand U92219 ( n55990, n6552, n55998 );
nand U92220 ( n55998, n76000, n55999 );
nand U92221 ( n56009, n6552, n56017 );
nand U92222 ( n56017, n76000, n56018 );
nand U92223 ( n56028, n6552, n56036 );
nand U92224 ( n56036, n75999, n56037 );
nand U92225 ( n56047, n6552, n56058 );
nand U92226 ( n56058, n75999, n56059 );
nand U92227 ( n56069, n6552, n56077 );
nand U92228 ( n56077, n75999, n56078 );
nand U92229 ( n56143, n6552, n56153 );
nand U92230 ( n56153, n76000, n56154 );
nand U92231 ( n43589, n7462, n43597 );
nand U92232 ( n43597, n76007, n43598 );
nand U92233 ( n43677, n7462, n43684 );
nand U92234 ( n43684, n76008, n43685 );
nand U92235 ( n9620, n4818, n9630 );
nand U92236 ( n9630, n76036, n9632 );
nor U92237 ( n21234, n21214, n21235 );
nor U92238 ( n21235, n21236, n21237 );
nand U92239 ( n21236, n14637, n11748 );
nand U92240 ( n21237, n14543, n14634 );
nand U92241 ( n42947, n76863, n8112 );
nand U92242 ( n43014, n76863, n8113 );
nand U92243 ( n43065, n76863, n8114 );
nand U92244 ( n43170, n76863, n8117 );
nand U92245 ( n42845, n76863, n8109 );
nand U92246 ( n43220, n76863, n8118 );
not U92247 ( n76534, n24463 );
nand U92248 ( n24463, n3920, n24602 );
nand U92249 ( n24602, n24603, n24604 );
nand U92250 ( n24603, n3980, n24607 );
not U92251 ( n76276, n57592 );
nand U92252 ( n57592, n6553, n57734 );
nand U92253 ( n57734, n57735, n57736 );
nand U92254 ( n57735, n6613, n57739 );
or U92255 ( n24604, n24605, n24606 );
or U92256 ( n57736, n57737, n57738 );
nand U92257 ( n30297, n3075, n30309 );
nand U92258 ( n30309, n76025, n30310 );
nand U92259 ( n30320, n3075, n30328 );
nand U92260 ( n30328, n76025, n30329 );
nand U92261 ( n30339, n3075, n30346 );
nand U92262 ( n30346, n76025, n30347 );
nand U92263 ( n64420, n5677, n64428 );
nand U92264 ( n64428, n75993, n64429 );
nand U92265 ( n22972, n3919, n22980 );
nand U92266 ( n22980, n76030, n22981 );
nand U92267 ( n22991, n3919, n22999 );
nand U92268 ( n22999, n76030, n23000 );
nand U92269 ( n23010, n3919, n23017 );
nand U92270 ( n23017, n76030, n23018 );
nand U92271 ( n9672, n4818, n9682 );
nand U92272 ( n9682, n76038, n9683 );
nand U92273 ( n9695, n4818, n9705 );
nand U92274 ( n9705, n76038, n9707 );
nand U92275 ( n9719, n4818, n9728 );
nand U92276 ( n9728, n76038, n9729 );
nand U92277 ( n64439, n5677, n64447 );
nand U92278 ( n64447, n75993, n64448 );
nand U92279 ( n64458, n5677, n64465 );
nand U92280 ( n64465, n75993, n64466 );
nand U92281 ( n56088, n6552, n56096 );
nand U92282 ( n56096, n76001, n56097 );
nand U92283 ( n56107, n6552, n56115 );
nand U92284 ( n56115, n76001, n56116 );
nand U92285 ( n56126, n6552, n56133 );
nand U92286 ( n56133, n76001, n56134 );
nand U92287 ( n43608, n7462, n43616 );
nand U92288 ( n43616, n76009, n43617 );
nand U92289 ( n43627, n7462, n43635 );
nand U92290 ( n43635, n76009, n43636 );
nand U92291 ( n43646, n7462, n43653 );
nand U92292 ( n43653, n76009, n43654 );
not U92293 ( n76210, n66165 );
nand U92294 ( n66165, n5678, n66410 );
nand U92295 ( n66410, n66411, n66412 );
nand U92296 ( n66411, n5738, n66415 );
or U92297 ( n66412, n66413, n66414 );
nand U92298 ( n29190, n35805, n35806 );
nand U92299 ( n35806, n32588, n34153 );
nor U92300 ( n35805, n35810, n35811 );
nor U92301 ( n35810, n31823, n35825 );
nand U92302 ( n21873, n28626, n28627 );
nand U92303 ( n28627, n25346, n26908 );
nor U92304 ( n28626, n28631, n28632 );
nor U92305 ( n28631, n24607, n28646 );
nand U92306 ( n62908, n70531, n70532 );
nand U92307 ( n70532, n67353, n68907 );
nor U92308 ( n70531, n70536, n70537 );
nor U92309 ( n70536, n66415, n70551 );
nand U92310 ( n54964, n61931, n61932 );
nand U92311 ( n61932, n58485, n60048 );
nor U92312 ( n61931, n61936, n61937 );
nor U92313 ( n61936, n57739, n61951 );
nand U92314 ( n42399, n54303, n54304 );
nand U92315 ( n54304, n46292, n47887 );
nor U92316 ( n54303, n54308, n54309 );
nor U92317 ( n54308, n45522, n54323 );
not U92318 ( n230, n8408 );
nand U92319 ( n8612, n8428, n8613 );
nand U92320 ( n8613, n76890, n5452 );
nand U92321 ( n8739, n76890, n5454 );
nand U92322 ( n8855, n76890, n5457 );
nand U92323 ( n9315, n76890, n5465 );
nand U92324 ( n8663, n76890, n5453 );
nand U92325 ( n9130, n76890, n5462 );
nand U92326 ( n8547, n76890, n5450 );
nand U92327 ( n63961, n76228, n6153 );
nand U92328 ( n30005, n76495, n3538 );
nand U92329 ( n22682, n76548, n4375 );
nand U92330 ( n55798, n76294, n7008 );
nand U92331 ( n47231, n46134, n76660 );
nand U92332 ( n13845, n12488, n76727 );
nand U92333 ( n68262, n67098, n76708 );
nand U92334 ( n26261, n25200, n76754 );
nand U92335 ( n59400, n58336, n76687 );
nand U92336 ( n8937, n76890, n5458 );
nand U92337 ( n9003, n76890, n5459 );
nand U92338 ( n9067, n76890, n5460 );
nand U92339 ( n9198, n76890, n5463 );
nand U92340 ( n8809, n76890, n5455 );
nand U92341 ( n9260, n76890, n5464 );
nand U92342 ( n63134, n63123, n63137 );
nand U92343 ( n63137, n63052, n63138 );
nand U92344 ( n63138, n76228, n6138 );
nand U92345 ( n29371, n29360, n29374 );
nand U92346 ( n29374, n29285, n29375 );
nand U92347 ( n29375, n76495, n3523 );
nand U92348 ( n22052, n22041, n22055 );
nand U92349 ( n22055, n21970, n22056 );
nand U92350 ( n22056, n76548, n4360 );
nand U92351 ( n55162, n55151, n55165 );
nand U92352 ( n55165, n55080, n55166 );
nand U92353 ( n55166, n76294, n6993 );
nand U92354 ( n33507, n32442, n76774 );
not U92355 ( n76354, n45325 );
nand U92356 ( n45325, n7463, n45517 );
nand U92357 ( n45517, n45518, n45519 );
nand U92358 ( n45518, n7523, n45522 );
or U92359 ( n45519, n45520, n45521 );
xor U92360 ( MUL_1411_U11, n71516, n71517 );
xor U92361 ( n71517, n71518, n71519 );
nand U92362 ( n21966, n21958, n21969 );
nand U92363 ( n21969, n21970, n21971 );
nand U92364 ( n21971, n76548, n4359 );
nand U92365 ( n29281, n29275, n29284 );
nand U92366 ( n29284, n29285, n29286 );
nand U92367 ( n29286, n76495, n3522 );
nand U92368 ( n63048, n63042, n63051 );
nand U92369 ( n63051, n63052, n63053 );
nand U92370 ( n63053, n76228, n6137 );
nand U92371 ( n55076, n55070, n55079 );
nand U92372 ( n55079, n55080, n55081 );
nand U92373 ( n55081, n76294, n6992 );
nor U92374 ( n26897, n26898, n26899 );
nor U92375 ( n26899, n26900, n26901 );
nor U92376 ( n26898, n26906, n26907 );
nor U92377 ( n26900, n26902, n26903 );
nor U92378 ( n60037, n60038, n60039 );
nor U92379 ( n60039, n60040, n60041 );
nor U92380 ( n60038, n60046, n60047 );
nor U92381 ( n60040, n60042, n60043 );
nor U92382 ( n34142, n34143, n34144 );
nor U92383 ( n34144, n34145, n34146 );
nor U92384 ( n34143, n34151, n34152 );
nor U92385 ( n34145, n34147, n34148 );
nor U92386 ( n68896, n68897, n68898 );
nor U92387 ( n68898, n68899, n68900 );
nor U92388 ( n68897, n68905, n68906 );
nor U92389 ( n68899, n68901, n68902 );
nand U92390 ( n22002, n22751, n22752 );
nor U92391 ( n22752, n21864, n22753 );
and U92392 ( n22751, n22754, n3822 );
nand U92393 ( n29321, n30072, n30073 );
nor U92394 ( n30073, n29177, n30074 );
and U92395 ( n30072, n30075, n2978 );
nand U92396 ( n55112, n55865, n55866 );
nor U92397 ( n55866, n54955, n55867 );
and U92398 ( n55865, n55868, n6454 );
nand U92399 ( n63084, n64089, n64090 );
nor U92400 ( n64090, n62899, n64091 );
and U92401 ( n64089, n64092, n5579 );
not U92402 ( n4759, n8438 );
nand U92403 ( n43278, n76864, n8119 );
not U92404 ( n7404, n42512 );
nand U92405 ( n8315, n21320, n21321 );
nand U92406 ( n21321, n12679, n14658 );
nor U92407 ( n21320, n21325, n21326 );
nor U92408 ( n21325, n11749, n21340 );
not U92409 ( n154, n23640 );
not U92410 ( n153, n23729 );
not U92411 ( n155, n23551 );
nand U92412 ( n42525, n76864, n42497 );
not U92413 ( n427, n56762 );
not U92414 ( n428, n56673 );
not U92415 ( n425, n56851 );
not U92416 ( n464, n65062 );
not U92417 ( n463, n65147 );
not U92418 ( n462, n65232 );
not U92419 ( n190, n31030 );
not U92420 ( n193, n30860 );
not U92421 ( n192, n30945 );
not U92422 ( n158, n23307 );
not U92423 ( n430, n56431 );
not U92424 ( n429, n56526 );
not U92425 ( n157, n23404 );
not U92426 ( n467, n64831 );
not U92427 ( n465, n64920 );
not U92428 ( n195, n30625 );
not U92429 ( n194, n30714 );
and U92430 ( n10020, n9969, n76891 );
and U92431 ( n10422, n10370, n76891 );
and U92432 ( n10188, n10133, n76891 );
and U92433 ( n43936, n43892, n76865 );
and U92434 ( n44261, n44220, n76865 );
and U92435 ( n44074, n44030, n76865 );
and U92436 ( n44404, n44349, n76865 );
and U92437 ( n10583, n10532, n76891 );
nand U92438 ( n11834, n4787, n11809 );
nand U92439 ( n21997, n22755, n22754 );
nor U92440 ( n22755, n22756, n22753 );
nand U92441 ( n29316, n30076, n30075 );
nor U92442 ( n30076, n30077, n30074 );
nand U92443 ( n63079, n64093, n64092 );
nor U92444 ( n64093, n64094, n64091 );
nand U92445 ( n55107, n55869, n55868 );
nor U92446 ( n55869, n55870, n55867 );
nand U92447 ( n11102, n11052, n76892 );
nand U92448 ( n11279, n11267, n76892 );
nand U92449 ( n44814, n44774, n76866 );
nand U92450 ( n44965, n44955, n76866 );
nand U92451 ( n10952, n10902, n76891 );
nand U92452 ( n44694, n44654, n76865 );
nand U92453 ( n44935, n44925, n76865 );
nand U92454 ( n10779, n10693, n76891 );
nand U92455 ( n11235, n11223, n76891 );
nand U92456 ( n44556, n44492, n76865 );
nand U92457 ( n63135, n63136, n76227 );
nor U92458 ( n63136, n6138, n63123 );
nand U92459 ( n63185, n63186, n76227 );
nor U92460 ( n63186, n6139, n63168 );
nand U92461 ( n63354, n63355, n76227 );
nor U92462 ( n63355, n6142, n63342 );
nand U92463 ( n29372, n29373, n76494 );
nor U92464 ( n29373, n3523, n29360 );
nand U92465 ( n29422, n29423, n76494 );
nor U92466 ( n29423, n3524, n29405 );
nand U92467 ( n29525, n29526, n76494 );
nor U92468 ( n29526, n3527, n29513 );
nand U92469 ( n22053, n22054, n76547 );
nor U92470 ( n22054, n4360, n22041 );
nand U92471 ( n22206, n22207, n76547 );
nor U92472 ( n22207, n4364, n22194 );
nand U92473 ( n22103, n22104, n76547 );
nor U92474 ( n22104, n4362, n22086 );
nand U92475 ( n55163, n55164, n76293 );
nor U92476 ( n55164, n6993, n55151 );
nand U92477 ( n55320, n55321, n76293 );
nor U92478 ( n55321, n6997, n55308 );
nand U92479 ( n55213, n55214, n76293 );
nor U92480 ( n55214, n6994, n55196 );
nand U92481 ( n68309, n76708, n67107 );
nand U92482 ( n26308, n76754, n25209 );
nand U92483 ( n59447, n76687, n58345 );
nand U92484 ( n63800, n63801, n76226 );
nor U92485 ( n63801, n6149, n63775 );
nand U92486 ( n29844, n29845, n76493 );
nor U92487 ( n29845, n3534, n29815 );
nand U92488 ( n22521, n22522, n76546 );
nor U92489 ( n22522, n4372, n22496 );
nand U92490 ( n55634, n55635, n76292 );
nor U92491 ( n55635, n7004, n55609 );
nand U92492 ( n33553, n76774, n32451 );
nand U92493 ( n47278, n76660, n46143 );
nand U92494 ( n21967, n21968, n76546 );
nor U92495 ( n21968, n4359, n21958 );
nand U92496 ( n29282, n29283, n76493 );
nor U92497 ( n29283, n3522, n29275 );
nand U92498 ( n63049, n63050, n76226 );
nor U92499 ( n63050, n6137, n63042 );
nand U92500 ( n55077, n55078, n76292 );
nor U92501 ( n55078, n6992, n55070 );
nand U92502 ( n13903, n76727, n12499 );
nand U92503 ( n63500, n63510, n63481 );
nand U92504 ( n63510, n63511, n76227 );
nor U92505 ( n63511, n6143, n63512 );
nor U92506 ( n63512, n63513, n6165 );
nand U92507 ( n29601, n29611, n29582 );
nand U92508 ( n29611, n29612, n76494 );
nor U92509 ( n29612, n3528, n29613 );
nor U92510 ( n29613, n29614, n3550 );
nand U92511 ( n22280, n22290, n22261 );
nand U92512 ( n22290, n22291, n76547 );
nor U92513 ( n22291, n4365, n22292 );
nor U92514 ( n22292, n22293, n4388 );
nand U92515 ( n55392, n55402, n55373 );
nand U92516 ( n55402, n55403, n76293 );
nor U92517 ( n55403, n6998, n55404 );
nor U92518 ( n55404, n55405, n7020 );
nand U92519 ( n63602, n63611, n63481 );
nand U92520 ( n63611, n63612, n76226 );
nor U92521 ( n63612, n6145, n63613 );
nor U92522 ( n63613, n63614, n6162 );
nand U92523 ( n63716, n63726, n63481 );
nand U92524 ( n63726, n63727, n76226 );
nor U92525 ( n63727, n6147, n63728 );
nor U92526 ( n63728, n63729, n6160 );
nand U92527 ( n63872, n63882, n63481 );
nand U92528 ( n63882, n63883, n76226 );
nor U92529 ( n63883, n6150, n63884 );
nor U92530 ( n63884, n63885, n63886 );
nand U92531 ( n29703, n29712, n29582 );
nand U92532 ( n29712, n29713, n76493 );
nor U92533 ( n29713, n3530, n29714 );
nor U92534 ( n29714, n29715, n3547 );
nand U92535 ( n29756, n29766, n29582 );
nand U92536 ( n29766, n29767, n76493 );
nor U92537 ( n29767, n3532, n29768 );
nor U92538 ( n29768, n29769, n3545 );
nand U92539 ( n29916, n29926, n29582 );
nand U92540 ( n29926, n29927, n76493 );
nor U92541 ( n29927, n3535, n29928 );
nor U92542 ( n29928, n29929, n29930 );
nand U92543 ( n22382, n22391, n22261 );
nand U92544 ( n22391, n22392, n76546 );
nor U92545 ( n22392, n4368, n22393 );
nor U92546 ( n22393, n22394, n4384 );
nand U92547 ( n22435, n22445, n22261 );
nand U92548 ( n22445, n22446, n76546 );
nor U92549 ( n22446, n4369, n22447 );
nor U92550 ( n22447, n22448, n4383 );
nand U92551 ( n22593, n22603, n22261 );
nand U92552 ( n22603, n22604, n76546 );
nor U92553 ( n22604, n4373, n22605 );
nor U92554 ( n22605, n22606, n22607 );
nand U92555 ( n55494, n55503, n55373 );
nand U92556 ( n55503, n55504, n76292 );
nor U92557 ( n55504, n7000, n55505 );
nor U92558 ( n55505, n55506, n7017 );
nand U92559 ( n55550, n55560, n55373 );
nand U92560 ( n55560, n55561, n76292 );
nor U92561 ( n55561, n7002, n55562 );
nor U92562 ( n55562, n55563, n7015 );
nand U92563 ( n55706, n55716, n55373 );
nand U92564 ( n55716, n55717, n76292 );
nor U92565 ( n55717, n7005, n55718 );
nor U92566 ( n55718, n55719, n55720 );
nand U92567 ( n30116, n3075, n30119 );
nand U92568 ( n30119, n76023, n30112 );
nand U92569 ( n64129, n5677, n64132 );
nand U92570 ( n64132, n75991, n64125 );
nand U92571 ( n22791, n3919, n22794 );
nand U92572 ( n22794, n76028, n22787 );
nand U92573 ( n55905, n6552, n55908 );
nand U92574 ( n55908, n75999, n55901 );
nand U92575 ( n43385, n7462, n43388 );
nand U92576 ( n43388, n76007, n43381 );
nand U92577 ( n9448, n4818, n9452 );
nand U92578 ( n9452, n76036, n9443 );
nand U92579 ( n30135, n30125, n76023 );
nand U92580 ( n32400, n29815, n32146 );
nand U92581 ( n67063, n63775, n66792 );
nand U92582 ( n25165, n22496, n24914 );
nand U92583 ( n58301, n55609, n58051 );
nand U92584 ( n43404, n43394, n76007 );
nand U92585 ( n64148, n64138, n75991 );
nand U92586 ( n22810, n22800, n76028 );
nand U92587 ( n55924, n55914, n75999 );
nand U92588 ( n9472, n9459, n76036 );
nand U92589 ( n46099, n43076, n45841 );
not U92590 ( n2082, n36264 );
nor U92591 ( n12151, n63017, n63018 );
nor U92592 ( n63017, n63021, n63020 );
nor U92593 ( n63018, n76226, n63020 );
nor U92594 ( n63021, n63042, n63043 );
nor U92595 ( n5416, n29250, n29251 );
nor U92596 ( n29250, n29254, n29253 );
nor U92597 ( n29251, n76493, n29253 );
nor U92598 ( n29254, n29275, n29276 );
nor U92599 ( n7661, n21933, n21934 );
nor U92600 ( n21933, n21937, n21936 );
nor U92601 ( n21934, n76546, n21936 );
nor U92602 ( n21937, n21958, n21959 );
nor U92603 ( n14396, n55045, n55046 );
nor U92604 ( n55045, n55049, n55048 );
nor U92605 ( n55046, n76292, n55048 );
nor U92606 ( n55049, n55070, n55071 );
nor U92607 ( n63193, n63161, n478 );
nor U92608 ( n63337, n63252, n478 );
nor U92609 ( n63484, n63453, n478 );
nor U92610 ( n63568, n63546, n478 );
nor U92611 ( n29430, n29398, n207 );
nor U92612 ( n29508, n29489, n207 );
nor U92613 ( n29585, n29550, n207 );
nor U92614 ( n29669, n29647, n207 );
nor U92615 ( n22189, n22170, n173 );
nor U92616 ( n22111, n22079, n173 );
nor U92617 ( n22264, n22233, n173 );
nor U92618 ( n22348, n22326, n173 );
nor U92619 ( n55303, n55284, n445 );
nor U92620 ( n55221, n55189, n445 );
nor U92621 ( n55376, n55345, n445 );
nor U92622 ( n55460, n55438, n445 );
nand U92623 ( n30375, n76024, n3688 );
nand U92624 ( n9764, n76037, n5448 );
nand U92625 ( n64538, n75992, n6322 );
nand U92626 ( n43696, n76008, n8103 );
nand U92627 ( n23046, n76029, n4582 );
nand U92628 ( n56165, n76000, n7214 );
nand U92629 ( n42527, n42538, n42539 );
nand U92630 ( n42538, n43349, n7409 );
nor U92631 ( n43349, n43350, n43346 );
nor U92632 ( n49175, n48033, n49180 );
nor U92633 ( n48806, n48033, n48811 );
nor U92634 ( n48340, n48033, n48346 );
nor U92635 ( n48243, n48033, n48249 );
nor U92636 ( n48145, n48033, n48151 );
not U92637 ( n2074, n38822 );
nand U92638 ( n8448, n8462, n8463 );
nand U92639 ( n8462, n9403, n4764 );
nor U92640 ( n9403, n9404, n9399 );
and U92641 ( n35609, n35610, n3077 );
and U92642 ( n54109, n54110, n7463 );
and U92643 ( n28432, n28433, n3920 );
and U92644 ( n70337, n70338, n5678 );
and U92645 ( n61737, n61738, n6553 );
not U92646 ( n2060, n37110 );
not U92647 ( n76925, n72968 );
not U92648 ( n813, n61441 );
nand U92649 ( n33468, n3103, n32402 );
nand U92650 ( n47188, n7490, n46101 );
nand U92651 ( n68219, n5704, n67065 );
nand U92652 ( n26218, n3947, n25167 );
nand U92653 ( n59357, n6579, n58303 );
nor U92654 ( n45327, n247, n45391 );
nand U92655 ( n13815, n4848, n12447 );
nor U92656 ( n42294, n812, n814 );
nor U92657 ( n44988, n247, n44561 );
nor U92658 ( n42759, n42736, n504 );
nor U92659 ( n42916, n42894, n504 );
nor U92660 ( n42653, n42621, n504 );
nor U92661 ( n42832, n42801, n504 );
nor U92662 ( n44496, n247, n43799 );
and U92663 ( n21126, n21127, n4819 );
nor U92664 ( n54214, n7802, n46408 );
nor U92665 ( n35716, n3399, n32707 );
nor U92666 ( n28537, n4237, n25467 );
nor U92667 ( n70442, n6014, n67472 );
nor U92668 ( n61842, n6869, n58604 );
buf U92669 ( n76041, n76926 );
nor U92670 ( n8702, n8678, n233 );
nor U92671 ( n8898, n8870, n233 );
nor U92672 ( n8604, n8564, n233 );
nor U92673 ( n8793, n8754, n233 );
nand U92674 ( n71502, n71276, n71503 );
nand U92675 ( n71503, n1222, n76043 );
not U92676 ( n169, n21982 );
not U92677 ( n203, n29297 );
not U92678 ( n474, n63064 );
not U92679 ( n442, n55092 );
nand U92680 ( n13960, n76727, n12523 );
nand U92681 ( n68355, n76708, n67137 );
nand U92682 ( n47323, n76660, n46173 );
nand U92683 ( n26354, n76754, n25239 );
nand U92684 ( n59493, n76687, n58375 );
nand U92685 ( n33599, n76774, n32481 );
nand U92686 ( n42489, n42553, n42554 );
nand U92687 ( n26913, n26914, n26915 );
nand U92688 ( n26915, n3822, n26905 );
nand U92689 ( n26914, n4045, n4020 );
nand U92690 ( n60053, n60054, n60055 );
nand U92691 ( n60055, n6454, n60045 );
nand U92692 ( n60054, n6678, n6653 );
nand U92693 ( n34158, n34159, n34160 );
nand U92694 ( n34160, n2978, n34150 );
nand U92695 ( n34159, n3215, n3183 );
nand U92696 ( n68912, n68913, n68914 );
nand U92697 ( n68914, n5579, n68904 );
nand U92698 ( n68913, n5814, n5782 );
not U92699 ( n1022, n71055 );
nor U92700 ( n37779, n2153, n2197 );
nand U92701 ( n12729, n12768, n12769 );
nor U92702 ( n12768, n12779, n12780 );
nor U92703 ( n12769, n12770, n12772 );
nor U92704 ( n12779, n12755, n4872 );
nand U92705 ( n63976, n63041, n64049 );
nand U92706 ( n30020, n29274, n30032 );
nand U92707 ( n55813, n55069, n55825 );
nand U92708 ( n22697, n21957, n22709 );
nand U92709 ( n46329, n46359, n46360 );
nor U92710 ( n46359, n46367, n46368 );
nor U92711 ( n46360, n46361, n46362 );
nor U92712 ( n46367, n46348, n7518 );
nand U92713 ( n63149, n63041, n63158 );
nand U92714 ( n63158, n63068, n63157 );
nand U92715 ( n29386, n29274, n29395 );
nand U92716 ( n29395, n29301, n29394 );
nand U92717 ( n22067, n21957, n22076 );
nand U92718 ( n22076, n21986, n22075 );
nand U92719 ( n55177, n55069, n55186 );
nand U92720 ( n55186, n55096, n55185 );
nand U92721 ( n63524, n63041, n63541 );
nand U92722 ( n63541, n63068, n63453 );
nand U92723 ( n63740, n63041, n63755 );
nand U92724 ( n63755, n63068, n63628 );
nand U92725 ( n63896, n63041, n63911 );
nand U92726 ( n63911, n63068, n63845 );
nand U92727 ( n29625, n29274, n29642 );
nand U92728 ( n29642, n29301, n29550 );
nand U92729 ( n29780, n29274, n29795 );
nand U92730 ( n29795, n29301, n29729 );
nand U92731 ( n29940, n29274, n29955 );
nand U92732 ( n29955, n29301, n29889 );
nand U92733 ( n22459, n21957, n22474 );
nand U92734 ( n22474, n21986, n22408 );
nand U92735 ( n22617, n21957, n22632 );
nand U92736 ( n22632, n21986, n22566 );
nand U92737 ( n22304, n21957, n22321 );
nand U92738 ( n22321, n21986, n22233 );
nand U92739 ( n55574, n55069, n55589 );
nand U92740 ( n55589, n55096, n55520 );
nand U92741 ( n55730, n55069, n55745 );
nand U92742 ( n55745, n55096, n55679 );
nand U92743 ( n55416, n55069, n55433 );
nand U92744 ( n55433, n55096, n55345 );
nand U92745 ( n63368, n63041, n63450 );
nand U92746 ( n63450, n63068, n63252 );
nand U92747 ( n29539, n29274, n29547 );
nand U92748 ( n29547, n29301, n29489 );
nand U92749 ( n22220, n21957, n22230 );
nand U92750 ( n22230, n21986, n22170 );
nand U92751 ( n55334, n55069, n55342 );
nand U92752 ( n55342, n55096, n55284 );
nand U92753 ( n63592, n63041, n63625 );
nand U92754 ( n63625, n63068, n63546 );
nand U92755 ( n63810, n63041, n63842 );
nand U92756 ( n63842, n63068, n63758 );
nand U92757 ( n29693, n29274, n29726 );
nand U92758 ( n29726, n29301, n29647 );
nand U92759 ( n29854, n29274, n29886 );
nand U92760 ( n29886, n29301, n29798 );
nand U92761 ( n22531, n21957, n22563 );
nand U92762 ( n22563, n21986, n22477 );
nand U92763 ( n22372, n21957, n22405 );
nand U92764 ( n22405, n21986, n22326 );
nand U92765 ( n55644, n55069, n55676 );
nand U92766 ( n55676, n55096, n55592 );
nand U92767 ( n55484, n55069, n55517 );
nand U92768 ( n55517, n55096, n55438 );
nand U92769 ( n63211, n63041, n63249 );
nand U92770 ( n63249, n63068, n63161 );
nand U92771 ( n29448, n29274, n29486 );
nand U92772 ( n29486, n29301, n29398 );
nand U92773 ( n22129, n21957, n22167 );
nand U92774 ( n22167, n21986, n22079 );
nand U92775 ( n55239, n55069, n55281 );
nand U92776 ( n55281, n55096, n55189 );
not U92777 ( n7925, n42583 );
not U92778 ( n2389, n17404 );
nor U92779 ( n8400, n8479, n8478 );
nor U92780 ( n42551, n7924, n42552 );
nor U92781 ( n42552, n42553, n42554 );
nor U92782 ( n11507, n2, n11594 );
not U92783 ( n7927, n42629 );
nor U92784 ( n24488, n29, n24530 );
nor U92785 ( n24474, n14, n24530 );
nor U92786 ( n24480, n19, n24530 );
nor U92787 ( n57619, n287, n57658 );
nor U92788 ( n57615, n280, n57658 );
nor U92789 ( n57607, n268, n57658 );
nor U92790 ( n57603, n262, n57658 );
nor U92791 ( n57623, n292, n57658 );
nor U92792 ( n57611, n274, n57658 );
nor U92793 ( n57594, n249, n57658 );
nor U92794 ( n24496, n38, n24530 );
nor U92795 ( n24492, n34, n24530 );
nor U92796 ( n24484, n24, n24530 );
nor U92797 ( n24465, n4, n24530 );
nor U92798 ( n24470, n9, n24530 );
nor U92799 ( n57599, n255, n57658 );
not U92800 ( n3873, n21970 );
not U92801 ( n3029, n29285 );
not U92802 ( n5630, n63052 );
not U92803 ( n6505, n55080 );
nand U92804 ( n63572, n5630, n6163 );
nand U92805 ( n63737, n5630, n63730 );
nand U92806 ( n29673, n3029, n3548 );
nand U92807 ( n29777, n3029, n29770 );
nand U92808 ( n22352, n3873, n4385 );
nand U92809 ( n22456, n3873, n22449 );
nand U92810 ( n55464, n6505, n7018 );
nand U92811 ( n55571, n6505, n55564 );
nor U92812 ( n40482, n40359, n76399 );
nor U92813 ( n40644, n40242, n76399 );
nor U92814 ( n40503, n40464, n76399 );
nor U92815 ( n40521, n2084, n76399 );
not U92816 ( n2084, n40461 );
nor U92817 ( n40486, n2097, n76399 );
not U92818 ( n2097, n40342 );
not U92819 ( n76920, n72969 );
nor U92820 ( n40585, n39808, n76398 );
nor U92821 ( n40596, n39913, n76398 );
nor U92822 ( n40607, n39990, n76398 );
nor U92823 ( n40618, n40078, n76398 );
nor U92824 ( n40633, n40167, n76398 );
nor U92825 ( n40533, n40421, n76398 );
nor U92826 ( n40550, n40412, n76398 );
nor U92827 ( n40559, n39561, n76398 );
nor U92828 ( n40574, n39683, n76398 );
not U92829 ( n7928, n42704 );
nor U92830 ( n13648, n76626, n13652 );
nor U92831 ( n14775, n76625, n14778 );
nor U92832 ( n15082, n76625, n15084 );
nor U92833 ( n15345, n76625, n15348 );
nor U92834 ( n15617, n76625, n15619 );
nor U92835 ( n15870, n76625, n15873 );
nor U92836 ( n16139, n76625, n16142 );
nor U92837 ( n40554, n76397, n40556 );
nand U92838 ( n40556, n1990, n40547 );
not U92839 ( n1990, n39502 );
nor U92840 ( n40492, n76397, n40494 );
or U92841 ( n40494, n2154, n40347 );
nor U92842 ( n40527, n76397, n40529 );
or U92843 ( n40529, n2095, n40451 );
not U92844 ( n5270, n8517 );
not U92845 ( n7929, n42765 );
nand U92846 ( n42809, n42865, n7932 );
nor U92847 ( n42865, n42863, n42862 );
not U92848 ( n7932, n42864 );
buf U92849 ( n76515, n76513 );
buf U92850 ( n76514, n76513 );
nor U92851 ( n16390, n76626, n16393 );
nor U92852 ( n42488, n42489, n42490 );
nand U92853 ( n25388, n25418, n25419 );
nor U92854 ( n25418, n25426, n25427 );
nor U92855 ( n25419, n25420, n25421 );
nor U92856 ( n25426, n25407, n3975 );
nand U92857 ( n58525, n58555, n58556 );
nor U92858 ( n58555, n58563, n58564 );
nor U92859 ( n58556, n58557, n58558 );
nor U92860 ( n58563, n58544, n6608 );
nand U92861 ( n32628, n32658, n32659 );
nor U92862 ( n32658, n32666, n32667 );
nor U92863 ( n32659, n32660, n32661 );
nor U92864 ( n32666, n32647, n3132 );
nand U92865 ( n67393, n67423, n67424 );
nor U92866 ( n67423, n67431, n67432 );
nor U92867 ( n67424, n67425, n67426 );
nor U92868 ( n67431, n67412, n5733 );
nor U92869 ( n47875, n47888, n47889 );
nor U92870 ( n47888, n47890, n45520 );
nor U92871 ( n47890, n47891, n47892 );
nor U92872 ( n47891, n47895, n45509 );
nor U92873 ( n14643, n14659, n14660 );
nor U92874 ( n14659, n14662, n11747 );
nor U92875 ( n14662, n14663, n14664 );
nor U92876 ( n14663, n14668, n11733 );
buf U92877 ( n76334, n76331 );
buf U92878 ( n76600, n76597 );
buf U92879 ( n76333, n76331 );
buf U92880 ( n76599, n76597 );
buf U92881 ( n76332, n76331 );
buf U92882 ( n76598, n76597 );
not U92883 ( n5272, n8574 );
nor U92884 ( n32932, n3113, n32877 );
nor U92885 ( n67693, n5714, n67638 );
nor U92886 ( n25688, n3957, n25633 );
nor U92887 ( n58828, n6589, n58770 );
nor U92888 ( n33278, n33218, n3113 );
nor U92889 ( n68037, n67973, n5714 );
nor U92890 ( n26034, n25970, n3957 );
nor U92891 ( n59175, n59108, n6589 );
nor U92892 ( n13218, n4832, n13157 );
not U92893 ( n7933, n42906 );
not U92894 ( n7947, n43075 );
nand U92895 ( n42979, n43034, n7935 );
nor U92896 ( n43034, n43031, n43032 );
nand U92897 ( n43033, n43078, n7937 );
nor U92898 ( n43078, n7947, n43076 );
nor U92899 ( n67596, n67514, n5714 );
nor U92900 ( n32831, n32749, n3113 );
nor U92901 ( n25591, n25509, n3957 );
nor U92902 ( n58728, n58646, n6589 );
or U92903 ( n13492, n13432, n4832 );
or U92904 ( n46502, n46450, n7500 );
not U92905 ( n5273, n8638 );
nand U92906 ( n21987, n21999, n22000 );
nand U92907 ( n22000, n178, n21998 );
nor U92908 ( n21999, n3875, n22003 );
nor U92909 ( n22003, n21946, n21997 );
nand U92910 ( n29302, n29318, n29319 );
nand U92911 ( n29319, n212, n29317 );
nor U92912 ( n29318, n3032, n29322 );
nor U92913 ( n29322, n29263, n29316 );
nand U92914 ( n63069, n63081, n63082 );
nand U92915 ( n63082, n483, n63080 );
nor U92916 ( n63081, n5633, n63085 );
nor U92917 ( n63085, n63030, n63079 );
nand U92918 ( n55097, n55109, n55110 );
nand U92919 ( n55110, n449, n55108 );
nor U92920 ( n55109, n6508, n55113 );
nor U92921 ( n55113, n55058, n55107 );
or U92922 ( n12998, n12898, n4855 );
nor U92923 ( n13122, n4855, n13050 );
nor U92924 ( n46646, n7500, n46591 );
nor U92925 ( n13567, n13487, n4855 );
not U92926 ( n5274, n8709 );
nand U92927 ( n8764, n8834, n5277 );
nor U92928 ( n8834, n8832, n8830 );
not U92929 ( n5277, n8833 );
not U92930 ( n7945, n43127 );
nand U92931 ( n43077, n43130, n7938 );
nor U92932 ( n43130, n7945, n43128 );
nor U92933 ( n47002, n46926, n7500 );
nand U92934 ( n21988, P1_P2_STATE2_REG_3_, n21957 );
nand U92935 ( n29303, P1_P3_STATE2_REG_3_, n29274 );
nand U92936 ( n63070, P2_P3_STATE2_REG_3_, n63041 );
nand U92937 ( n55098, P2_P2_STATE2_REG_3_, n55069 );
nand U92938 ( n76102, n42538, n42539 );
nand U92939 ( n43291, n42617, n43303 );
and U92940 ( n41311, n54987, n829 );
nor U92941 ( n42544, n42537, n42538 );
nand U92942 ( n42528, n42541, n42542 );
nand U92943 ( n42542, n510, n42540 );
nor U92944 ( n42541, n7407, n42544 );
not U92945 ( n510, n42539 );
nand U92946 ( n42608, n42617, n42618 );
nand U92947 ( n42618, n42527, n42616 );
nand U92948 ( n43041, n42617, n43056 );
nand U92949 ( n43056, n42527, n42990 );
nand U92950 ( n43197, n42617, n43212 );
nand U92951 ( n43212, n42527, n43146 );
nand U92952 ( n42872, n42617, n42889 );
nand U92953 ( n42889, n42527, n42801 );
not U92954 ( n6138, n63124 );
not U92955 ( n3523, n29361 );
not U92956 ( n4360, n22042 );
not U92957 ( n6993, n55152 );
not U92958 ( n6139, n63169 );
not U92959 ( n6140, n63220 );
not U92960 ( n6142, n63343 );
not U92961 ( n6143, n63461 );
not U92962 ( n3524, n29406 );
not U92963 ( n3525, n29457 );
not U92964 ( n3527, n29514 );
not U92965 ( n3528, n29558 );
not U92966 ( n4364, n22195 );
not U92967 ( n4362, n22087 );
not U92968 ( n4363, n22138 );
not U92969 ( n4365, n22241 );
not U92970 ( n6997, n55309 );
not U92971 ( n6994, n55197 );
not U92972 ( n6995, n55248 );
not U92973 ( n6998, n55353 );
not U92974 ( n4359, n21959 );
not U92975 ( n3522, n29276 );
not U92976 ( n6137, n63043 );
not U92977 ( n6992, n55071 );
nand U92978 ( n42790, n42617, n42798 );
nand U92979 ( n42798, n42527, n42736 );
not U92980 ( n6144, n63516 );
not U92981 ( n3529, n29617 );
not U92982 ( n4367, n22296 );
not U92983 ( n6999, n55408 );
nand U92984 ( n43111, n42617, n43143 );
nand U92985 ( n43143, n42527, n43059 );
nand U92986 ( n42940, n42617, n42987 );
nand U92987 ( n42987, n42527, n42894 );
nand U92988 ( n76172, n8462, n8463 );
nand U92989 ( n9332, n8559, n9347 );
nand U92990 ( n42695, n42617, n42733 );
nand U92991 ( n42733, n42527, n42621 );
nor U92992 ( n8469, n8460, n8462 );
nand U92993 ( n8449, n8465, n8467 );
nand U92994 ( n8467, n239, n8464 );
nor U92995 ( n8465, n4762, n8469 );
not U92996 ( n239, n8463 );
nor U92997 ( n37117, n76039, n2198 );
nand U92998 ( n8548, n8559, n8560 );
nand U92999 ( n8560, n8448, n8558 );
nand U93000 ( n9037, n8559, n9055 );
nand U93001 ( n9055, n8448, n8973 );
nand U93002 ( n9232, n8559, n9250 );
nand U93003 ( n9250, n8448, n9168 );
nand U93004 ( n8843, n8559, n8864 );
nand U93005 ( n8864, n8448, n8754 );
nand U93006 ( n8740, n8559, n8750 );
nand U93007 ( n8750, n8448, n8678 );
nand U93008 ( n9124, n8559, n9164 );
nand U93009 ( n9164, n8448, n9059 );
nand U93010 ( n8928, n8559, n8969 );
nand U93011 ( n8969, n8448, n8870 );
nor U93012 ( n68286, n68287, n68288 );
nand U93013 ( n68287, n68246, n68249 );
nand U93014 ( n68288, n68289, n68290 );
nand U93015 ( n68290, n6078, n67395 );
nor U93016 ( n26285, n26286, n26287 );
nand U93017 ( n26286, n26245, n26248 );
nand U93018 ( n26287, n26288, n26289 );
nand U93019 ( n26289, n4300, n25390 );
nor U93020 ( n59424, n59425, n59426 );
nand U93021 ( n59425, n59384, n59387 );
nand U93022 ( n59426, n59427, n59428 );
nand U93023 ( n59428, n6933, n58527 );
nand U93024 ( n8627, n8559, n8674 );
nand U93025 ( n8674, n8448, n8564 );
nor U93026 ( n68158, n68159, n68160 );
nand U93027 ( n68159, n68116, n5709 );
nand U93028 ( n68160, n68161, n68162 );
not U93029 ( n5709, n68113 );
nor U93030 ( n26157, n26158, n26159 );
nand U93031 ( n26158, n26113, n3952 );
nand U93032 ( n26159, n26160, n26161 );
not U93033 ( n3952, n26110 );
nor U93034 ( n59296, n59297, n59298 );
nand U93035 ( n59297, n59254, n6584 );
nand U93036 ( n59298, n59299, n59300 );
not U93037 ( n6584, n59251 );
not U93038 ( n7944, n43187 );
nand U93039 ( n43129, n43190, n7939 );
nor U93040 ( n43190, n7944, n43188 );
nor U93041 ( n33530, n33531, n33532 );
nand U93042 ( n33531, n33491, n33494 );
nand U93043 ( n33532, n33533, n33534 );
nand U93044 ( n33534, n3463, n32630 );
nor U93045 ( n33408, n33409, n33410 );
nand U93046 ( n33409, n33359, n3108 );
nand U93047 ( n33410, n33411, n33412 );
not U93048 ( n3108, n33356 );
nor U93049 ( n13347, n13312, n4832 );
nand U93050 ( n21975, n21995, n21996 );
nand U93051 ( n21996, n177, n21946 );
nand U93052 ( n21995, n178, n21946 );
nand U93053 ( n55085, n55105, n55106 );
nand U93054 ( n55106, n448, n55058 );
nand U93055 ( n55105, n449, n55058 );
nand U93056 ( n29290, n29314, n29315 );
nand U93057 ( n29315, n210, n29263 );
nand U93058 ( n29314, n212, n29263 );
nand U93059 ( n63057, n63077, n63078 );
nand U93060 ( n63078, n482, n63030 );
nand U93061 ( n63077, n483, n63030 );
nor U93062 ( n13048, n13002, n4832 );
not U93063 ( n6145, n63558 );
not U93064 ( n3530, n29659 );
not U93065 ( n4368, n22338 );
not U93066 ( n7000, n55450 );
not U93067 ( n6155, n63939 );
not U93068 ( n3540, n29983 );
not U93069 ( n4378, n22660 );
not U93070 ( n7010, n55773 );
nand U93071 ( n63617, n63733, n6148 );
nor U93072 ( n63733, n63730, n63731 );
nand U93073 ( n63732, n63777, n6149 );
nor U93074 ( n63777, n6159, n63775 );
nand U93075 ( n63776, n63829, n6150 );
nor U93076 ( n63829, n6158, n63827 );
nand U93077 ( n63828, n63889, n6152 );
nor U93078 ( n63889, n6157, n63887 );
nand U93079 ( n63888, n63942, n6153 );
nor U93080 ( n63942, n6155, n63940 );
nand U93081 ( n29718, n29773, n3533 );
nor U93082 ( n29773, n29770, n29771 );
nand U93083 ( n29772, n29817, n3534 );
nor U93084 ( n29817, n3544, n29815 );
nand U93085 ( n29816, n29873, n3535 );
nor U93086 ( n29873, n3543, n29871 );
nand U93087 ( n29872, n29933, n3537 );
nor U93088 ( n29933, n3542, n29931 );
nand U93089 ( n29932, n29986, n3538 );
nor U93090 ( n29986, n3540, n29984 );
nand U93091 ( n22397, n22452, n4370 );
nor U93092 ( n22452, n22449, n22450 );
nand U93093 ( n22497, n22550, n4373 );
nor U93094 ( n22550, n4380, n22548 );
nand U93095 ( n22549, n22610, n4374 );
nor U93096 ( n22610, n4379, n22608 );
nand U93097 ( n22451, n22498, n4372 );
nor U93098 ( n22498, n4382, n22496 );
nand U93099 ( n22609, n22663, n4375 );
nor U93100 ( n22663, n4378, n22661 );
nand U93101 ( n55509, n55567, n7003 );
nor U93102 ( n55567, n55564, n55565 );
nand U93103 ( n55610, n55663, n7005 );
nor U93104 ( n55663, n7013, n55661 );
nand U93105 ( n55662, n55723, n7007 );
nor U93106 ( n55723, n7012, n55721 );
nand U93107 ( n55566, n55611, n7004 );
nor U93108 ( n55611, n7014, n55609 );
nand U93109 ( n55722, n55776, n7008 );
nor U93110 ( n55776, n7010, n55774 );
not U93111 ( n6158, n63826 );
not U93112 ( n3543, n29870 );
not U93113 ( n4380, n22547 );
not U93114 ( n7013, n55660 );
not U93115 ( n6157, n63886 );
not U93116 ( n3542, n29930 );
not U93117 ( n4379, n22607 );
not U93118 ( n7012, n55720 );
not U93119 ( n6159, n63774 );
not U93120 ( n3544, n29814 );
not U93121 ( n4382, n22495 );
not U93122 ( n7014, n55608 );
nand U93123 ( n33499, n33538, n33539 );
nand U93124 ( n33538, n3474, n76128 );
nand U93125 ( n33539, n33540, n3469 );
not U93126 ( n3469, n33451 );
not U93127 ( n5278, n8885 );
not U93128 ( n5292, n9079 );
nand U93129 ( n8959, n9028, n5280 );
nor U93130 ( n9028, n9024, n9025 );
nand U93131 ( n9027, n9083, n5282 );
nor U93132 ( n9083, n5292, n9080 );
nand U93133 ( n68254, n68294, n68295 );
nand U93134 ( n68294, n6089, n76058 );
nand U93135 ( n68295, n68296, n6084 );
not U93136 ( n6084, n68202 );
nand U93137 ( n26253, n26293, n26294 );
nand U93138 ( n26293, n4312, n76156 );
nand U93139 ( n26294, n26295, n4307 );
not U93140 ( n4307, n26201 );
nand U93141 ( n59392, n59432, n59433 );
nand U93142 ( n59432, n6944, n76084 );
nand U93143 ( n59433, n59434, n6939 );
not U93144 ( n6939, n59340 );
not U93145 ( n1, n14832 );
nor U93146 ( n13874, n13875, n13877 );
nand U93147 ( n13875, n13825, n13829 );
nand U93148 ( n13877, n13878, n13879 );
nand U93149 ( n13879, n5214, n12732 );
nor U93150 ( n13724, n13725, n13727 );
nand U93151 ( n13725, n13672, n4852 );
nand U93152 ( n13727, n13728, n13729 );
not U93153 ( n4852, n13668 );
buf U93154 ( n76682, n7319 );
nor U93155 ( MUL_1411_U5, n1218, n1209 );
not U93156 ( n7943, n43254 );
nand U93157 ( n43189, n43257, n7940 );
nor U93158 ( n43257, n7943, n43255 );
or U93159 ( n33164, n3113, n33108 );
or U93160 ( n67915, n5714, n67864 );
or U93161 ( n25912, n3957, n25861 );
or U93162 ( n59050, n6589, n58999 );
nor U93163 ( n47255, n47256, n47257 );
nand U93164 ( n47256, n47215, n47218 );
nand U93165 ( n47257, n47258, n47259 );
nand U93166 ( n47259, n7868, n46331 );
not U93167 ( n500, n42524 );
nor U93168 ( n47127, n47128, n47129 );
nand U93169 ( n47128, n47085, n7495 );
nand U93170 ( n47129, n47130, n47131 );
not U93171 ( n7495, n47082 );
nand U93172 ( n8477, n8478, n8479 );
nor U93173 ( n14644, n14645, n14647 );
nor U93174 ( n14647, n14648, n14649 );
nor U93175 ( n14645, n14655, n14657 );
nor U93176 ( n14648, n14650, n14652 );
or U93177 ( n12879, n4832, n12838 );
not U93178 ( n229, n8428 );
nand U93179 ( n12735, n12753, n12754 );
nand U93180 ( n12754, n12755, n9812 );
nor U93181 ( n12753, n12757, n12758 );
nor U93182 ( n12758, n4873, n12759 );
nand U93183 ( n46356, n7874, n46365 );
not U93184 ( n7874, n46432 );
nor U93185 ( n12813, n12814, n12815 );
nand U93186 ( n12815, n12817, n4843 );
nand U93187 ( n12814, n12825, n12827 );
not U93188 ( n4843, n12780 );
nand U93189 ( n46334, n46346, n46347 );
nand U93190 ( n46347, n46348, n46349 );
nor U93191 ( n46346, n46350, n46351 );
nor U93192 ( n46351, n7517, n46352 );
not U93193 ( n5290, n9144 );
nand U93194 ( n9082, n9148, n5283 );
nor U93195 ( n9148, n5290, n9145 );
nand U93196 ( n13924, n4848, n12504 );
nand U93197 ( n68326, n5704, n67111 );
nand U93198 ( n47295, n7490, n46147 );
nand U93199 ( n26325, n3947, n25213 );
nand U93200 ( n59464, n6579, n58349 );
nand U93201 ( n33570, n3103, n32455 );
nor U93202 ( n67832, n67758, n5714 );
nor U93203 ( n33076, n33002, n3113 );
nor U93204 ( n25829, n25753, n3957 );
nor U93205 ( n58967, n58893, n6589 );
or U93206 ( n13419, n4855, n13349 );
or U93207 ( n46868, n7500, n46817 );
nor U93208 ( n67757, n5689, n67714 );
nor U93209 ( n46710, n7474, n46667 );
nor U93210 ( n25752, n3932, n25709 );
nor U93211 ( n58892, n6564, n58849 );
nor U93212 ( n33001, n3088, n32960 );
nor U93213 ( n68113, n5714, n68095 );
nor U93214 ( n26110, n3957, n26092 );
nor U93215 ( n59251, n6589, n59233 );
nor U93216 ( n33356, n3113, n33338 );
nand U93217 ( n61173, n54987, n829 );
not U93218 ( n5289, n9219 );
nand U93219 ( n9147, n9223, n5284 );
nor U93220 ( n9223, n5289, n9220 );
or U93221 ( n33222, n33174, n3088 );
nor U93222 ( n33341, n33288, n3123 );
nor U93223 ( n68098, n68047, n5723 );
nor U93224 ( n47067, n47012, n7509 );
nor U93225 ( n26095, n26044, n3965 );
nor U93226 ( n59236, n59185, n6598 );
nor U93227 ( n13309, n13219, n4855 );
or U93228 ( n67977, n67937, n5689 );
or U93229 ( n46930, n46890, n7474 );
or U93230 ( n25974, n25934, n3932 );
or U93231 ( n59112, n59072, n6564 );
nor U93232 ( n47314, n7509, n47270 );
nor U93233 ( n46785, n46711, n7500 );
nor U93234 ( n47876, n47877, n47878 );
nor U93235 ( n47878, n47879, n47880 );
nor U93236 ( n47877, n47885, n47886 );
nor U93237 ( n47879, n47881, n47882 );
nor U93238 ( n68346, n5723, n68301 );
nor U93239 ( n33590, n3123, n33545 );
nor U93240 ( n26345, n3965, n26300 );
nor U93241 ( n59484, n6598, n59439 );
nand U93242 ( n42517, n42535, n42536 );
or U93243 ( n42535, n42539, n42540 );
nand U93244 ( n42536, n509, n42537 );
not U93245 ( n509, n42538 );
not U93246 ( n5288, n9285 );
nand U93247 ( n9222, n9289, n5285 );
nor U93248 ( n9289, n5288, n9287 );
nor U93249 ( n13668, n4855, n13638 );
nor U93250 ( n47082, n7500, n47064 );
nand U93251 ( n14064, n14158, n14159 );
nand U93252 ( n14158, n13944, n12775 );
or U93253 ( n14159, n13889, n4832 );
nand U93254 ( n8435, n8458, n8459 );
or U93255 ( n8458, n8463, n8464 );
nand U93256 ( n8459, n238, n8460 );
not U93257 ( n238, n8462 );
not U93258 ( n512, n47786 );
not U93259 ( n240, n14532 );
buf U93260 ( n76683, n7319 );
and U93261 ( n67159, n68458, n68459 );
nand U93262 ( n68458, n68463, n5783 );
nand U93263 ( n68459, n68460, n68461 );
not U93264 ( n5783, n68461 );
and U93265 ( n46195, n47437, n47438 );
nand U93266 ( n47437, n47442, n7570 );
nand U93267 ( n47438, n47439, n47440 );
not U93268 ( n7570, n47440 );
and U93269 ( n25261, n26457, n26458 );
nand U93270 ( n26457, n26462, n4022 );
nand U93271 ( n26458, n26459, n26460 );
not U93272 ( n4022, n26460 );
and U93273 ( n58397, n59596, n59597 );
nand U93274 ( n59596, n59601, n6654 );
nand U93275 ( n59597, n59598, n59599 );
not U93276 ( n6654, n59599 );
nor U93277 ( n13642, n13579, n4864 );
and U93278 ( n32503, n33702, n33703 );
nand U93279 ( n33702, n33707, n3184 );
nand U93280 ( n33703, n33704, n33705 );
not U93281 ( n3184, n33705 );
and U93282 ( n12564, n14087, n14088 );
nand U93283 ( n14087, n14093, n4919 );
nand U93284 ( n14088, n14089, n14090 );
not U93285 ( n4919, n14090 );
nor U93286 ( n13948, n4864, n13893 );
nor U93287 ( n33448, n33413, n3123 );
nor U93288 ( n68199, n68163, n5723 );
nor U93289 ( n47168, n47132, n7509 );
nor U93290 ( n26198, n26162, n3965 );
nor U93291 ( n59337, n59301, n6598 );
nor U93292 ( n46587, n46536, n7474 );
nor U93293 ( n67636, n67598, n5689 );
nor U93294 ( n25631, n25593, n3932 );
nor U93295 ( n58768, n58730, n6564 );
nor U93296 ( n32875, n32833, n3088 );
nor U93297 ( n33106, n33078, n3088 );
nor U93298 ( n67862, n67834, n5689 );
nor U93299 ( n46815, n46787, n7474 );
nor U93300 ( n25859, n25831, n3932 );
nor U93301 ( n58997, n58969, n6564 );
not U93302 ( n7940, n43256 );
not U93303 ( n6153, n63941 );
not U93304 ( n3538, n29985 );
not U93305 ( n4375, n22662 );
not U93306 ( n7008, n55775 );
not U93307 ( n3122, n33093 );
not U93308 ( n5722, n67849 );
not U93309 ( n7508, n46802 );
not U93310 ( n3964, n25846 );
not U93311 ( n6597, n58984 );
not U93312 ( n7960, n42554 );
nor U93313 ( n13775, n13730, n4864 );
nand U93314 ( n67551, n67578, n67495 );
nand U93315 ( n32786, n32813, n32730 );
nand U93316 ( n25546, n25573, n25490 );
nand U93317 ( n58683, n58710, n58627 );
or U93318 ( n46431, n7474, n46410 );
not U93319 ( n4863, n13330 );
not U93320 ( n877, n45174 );
not U93321 ( n873, n45239 );
buf U93322 ( n76469, n32600 );
buf U93323 ( n76520, n25360 );
buf U93324 ( n76196, n67365 );
buf U93325 ( n76262, n58497 );
nand U93326 ( n67712, n67638, n67429 );
nand U93327 ( n32958, n32877, n32664 );
nand U93328 ( n46665, n46591, n46365 );
nand U93329 ( n25707, n25633, n25424 );
nand U93330 ( n58847, n58770, n58561 );
nand U93331 ( n13154, n13050, n12775 );
and U93332 ( n13428, n13349, n12775 );
and U93333 ( n33171, n33108, n32664 );
and U93334 ( n67934, n67864, n67429 );
and U93335 ( n46887, n46817, n46365 );
and U93336 ( n25931, n25861, n25424 );
and U93337 ( n59069, n58999, n58561 );
nand U93338 ( n32655, n3470, n32664 );
not U93339 ( n3470, n32731 );
nand U93340 ( n25415, n4308, n25424 );
not U93341 ( n4308, n25491 );
nand U93342 ( n67420, n6085, n67429 );
not U93343 ( n6085, n67496 );
nand U93344 ( n58552, n6940, n58561 );
not U93345 ( n6940, n58628 );
nand U93346 ( n32633, n32645, n32646 );
nand U93347 ( n32646, n32647, n32648 );
nor U93348 ( n32645, n32649, n32650 );
nor U93349 ( n32650, n3130, n32651 );
nand U93350 ( n25393, n25405, n25406 );
nand U93351 ( n25406, n25407, n25408 );
nor U93352 ( n25405, n25409, n25410 );
nor U93353 ( n25410, n3974, n25411 );
nand U93354 ( n67398, n67410, n67411 );
nand U93355 ( n67411, n67412, n67413 );
nor U93356 ( n67410, n67414, n67415 );
nor U93357 ( n67415, n5732, n67416 );
nand U93358 ( n58530, n58542, n58543 );
nand U93359 ( n58543, n58544, n58545 );
nor U93360 ( n58542, n58546, n58547 );
nor U93361 ( n58547, n6607, n58548 );
buf U93362 ( n76213, n76211 );
buf U93363 ( n76279, n76277 );
not U93364 ( n5285, n9288 );
buf U93365 ( n76537, n76535 );
buf U93366 ( n76214, n76211 );
buf U93367 ( n76280, n76277 );
nor U93368 ( n16124, n14832, n16130 );
nor U93369 ( n15705, n14832, n15712 );
nor U93370 ( n15173, n14832, n15180 );
nor U93371 ( n15065, n14832, n15073 );
nor U93372 ( n14962, n14832, n14969 );
buf U93373 ( n76538, n76535 );
nand U93374 ( n68356, n76705, n67126 );
nand U93375 ( n47324, n76657, n46162 );
nand U93376 ( n26355, n76751, n25228 );
nand U93377 ( n59494, n76684, n58364 );
nand U93378 ( n68439, n68515, n68516 );
nand U93379 ( n68515, n68343, n67429 );
or U93380 ( n68516, n68299, n5689 );
nand U93381 ( n33683, n33759, n33760 );
nand U93382 ( n33759, n33587, n32664 );
or U93383 ( n33760, n33543, n3088 );
nand U93384 ( n47407, n47494, n47495 );
nand U93385 ( n47494, n47311, n46365 );
or U93386 ( n47495, n47267, n7474 );
nand U93387 ( n26438, n26514, n26515 );
nand U93388 ( n26514, n26342, n25424 );
or U93389 ( n26515, n26298, n3932 );
nand U93390 ( n59577, n59653, n59654 );
nand U93391 ( n59653, n59481, n58561 );
or U93392 ( n59654, n59437, n6564 );
nand U93393 ( n33600, n76772, n32470 );
buf U93394 ( n76278, n76277 );
buf U93395 ( n76212, n76211 );
buf U93396 ( n76536, n76535 );
nand U93397 ( n42500, n76180, n42617 );
nor U93398 ( n68603, n5714, n68518 );
nor U93399 ( n33847, n3113, n33762 );
nor U93400 ( n26602, n3957, n26517 );
nor U93401 ( n59744, n6589, n59656 );
buf U93402 ( n76357, n76355 );
nand U93403 ( n13959, n76724, n12538 );
buf U93404 ( n76358, n76355 );
nand U93405 ( n13987, n4848, n12522 );
nand U93406 ( n47345, n7490, n46161 );
nand U93407 ( n8414, n76190, n8559 );
buf U93408 ( n76356, n76355 );
nand U93409 ( n46368, n46389, n46390 );
nand U93410 ( n46390, n46391, n46392 );
nand U93411 ( n46391, n46393, n46394 );
nand U93412 ( n46389, n46365, n46432 );
buf U93413 ( n76434, n76433 );
buf U93414 ( n76435, n76433 );
buf U93415 ( n76623, n76621 );
nand U93416 ( n12780, n12818, n12819 );
nand U93417 ( n12819, n12820, n12822 );
nand U93418 ( n12820, n12823, n12824 );
or U93419 ( n68162, n68132, n5723 );
or U93420 ( n47131, n47101, n7509 );
or U93421 ( n26161, n26129, n3965 );
or U93422 ( n59300, n59270, n6598 );
or U93423 ( n33412, n33380, n3123 );
buf U93424 ( n76624, n76621 );
nor U93425 ( n14268, n4855, n14162 );
nor U93426 ( n47582, n7500, n47497 );
nand U93427 ( n14734, n21109, n21110 );
or U93428 ( n21110, n5183, n15278 );
nor U93429 ( n21109, n15809, n5184 );
nor U93430 ( n15395, n14728, n18715 );
nand U93431 ( n14728, n21111, n21112 );
nand U93432 ( n21112, n15272, n20929 );
nor U93433 ( n21111, n15698, n15804 );
nor U93434 ( n15698, n15390, n20929 );
nor U93435 ( n18701, n14733, n5178 );
nor U93436 ( n18710, n18712, n14947 );
and U93437 ( n18712, n16449, n5168 );
not U93438 ( n5193, n15272 );
buf U93439 ( n76622, n76621 );
nand U93440 ( n48240, n54094, n54095 );
or U93441 ( n54095, n7838, n48417 );
nor U93442 ( n54094, n48882, n7839 );
not U93443 ( n7863, n48130 );
nor U93444 ( n48522, n48418, n51671 );
nand U93445 ( n48418, n54096, n54097 );
nand U93446 ( n54097, n48412, n53885 );
nor U93447 ( n54096, n48784, n48878 );
nor U93448 ( n48784, n48518, n53885 );
nor U93449 ( n48783, n48785, n48133 );
nor U93450 ( n48785, n7839, n7832 );
or U93451 ( n13729, n13692, n4864 );
nand U93452 ( n23162, n3797, n23819 );
nand U93453 ( n56283, n56944, n6429 );
buf U93454 ( n76074, n61176 );
nand U93455 ( n15925, n16013, n76591 );
nor U93456 ( n16013, n16014, n16015 );
and U93457 ( n16015, n15927, n76189 );
nor U93458 ( n16014, n16017, n16012 );
nand U93459 ( n16340, n16425, n76591 );
nor U93460 ( n16425, n16427, n16428 );
and U93461 ( n16428, n16342, n76191 );
nor U93462 ( n16427, n16429, n16424 );
nand U93463 ( n15932, n16024, n14958 );
nand U93464 ( n16347, n16024, n15397 );
nor U93465 ( n16024, n14692, n5178 );
nor U93466 ( n16429, n16432, n14947 );
and U93467 ( n16432, n16345, n16347 );
nor U93468 ( n16017, n16019, n14947 );
and U93469 ( n16019, n15930, n15932 );
nor U93470 ( n33283, n33284, n33252 );
nor U93471 ( n33284, n3123, n33256 );
nor U93472 ( n47007, n47008, n46976 );
nor U93473 ( n47008, n7509, n46980 );
nand U93474 ( n22738, n22754, n22767 );
nand U93475 ( n22767, n22768, n22769 );
nand U93476 ( n55854, n55868, n55881 );
nand U93477 ( n55881, n55882, n55883 );
nand U93478 ( n30061, n30075, n30088 );
nand U93479 ( n30088, n30089, n30090 );
nand U93480 ( n64078, n64092, n64105 );
nand U93481 ( n64105, n64106, n64107 );
nor U93482 ( n68042, n68043, n68011 );
nor U93483 ( n68043, n5723, n68015 );
nor U93484 ( n26039, n26040, n26008 );
nor U93485 ( n26040, n3965, n26012 );
nor U93486 ( n59180, n59181, n59146 );
nor U93487 ( n59181, n6598, n59150 );
nand U93488 ( n63971, n5632, n63972 );
nand U93489 ( n30015, n3030, n30016 );
nand U93490 ( n22692, n3874, n22693 );
nand U93491 ( n55808, n6507, n55809 );
nand U93492 ( n21172, n21173, n11749 );
nor U93493 ( n21173, n21174, n21175 );
nor U93494 ( n21174, n4965, n4963 );
and U93495 ( n8270, n21170, n21171 );
nand U93496 ( n21170, n14654, n21176 );
nand U93497 ( n21171, n4949, n21172 );
nand U93498 ( n21176, n21177, n11749 );
nand U93499 ( n14099, n4848, n12547 );
nand U93500 ( n68468, n5704, n67145 );
nand U93501 ( n47447, n7490, n46181 );
nand U93502 ( n26467, n3947, n25247 );
nand U93503 ( n59606, n6579, n58383 );
nand U93504 ( n33712, n3103, n32489 );
nand U93505 ( n46457, n46410, n46438 );
nor U93506 ( n49341, n49343, n48133 );
and U93507 ( n49343, n49279, n49280 );
nand U93508 ( n49275, n49338, n76325 );
nor U93509 ( n49338, n49339, n49340 );
and U93510 ( n49340, n49276, n76182 );
nor U93511 ( n49339, n49341, n49337 );
nand U93512 ( n15820, n15905, n76591 );
nor U93513 ( n15905, n15907, n15908 );
and U93514 ( n15908, n15822, n76190 );
nor U93515 ( n15907, n15909, n15904 );
nor U93516 ( n15909, n15912, n14947 );
and U93517 ( n15912, n15825, n15827 );
nand U93518 ( n16033, n16112, n76591 );
nor U93519 ( n16112, n16113, n16114 );
and U93520 ( n16114, n16034, n76187 );
nor U93521 ( n16113, n16115, n16110 );
nor U93522 ( n16115, n16118, n14947 );
and U93523 ( n16118, n16038, n16039 );
nand U93524 ( n68528, n76708, n67177 );
nand U93525 ( n47507, n76660, n46213 );
nand U93526 ( n26527, n76754, n25279 );
nand U93527 ( n59669, n76687, n58415 );
nand U93528 ( n48990, n49069, n76325 );
nor U93529 ( n49069, n49070, n49071 );
and U93530 ( n49071, n48991, n76179 );
nor U93531 ( n49070, n49072, n49068 );
nand U93532 ( n48995, n49078, n48142 );
nand U93533 ( n49358, n49078, n48523 );
nor U93534 ( n49078, n47921, n7833 );
nor U93535 ( n49072, n49074, n48133 );
and U93536 ( n49074, n48994, n48995 );
nor U93537 ( n49434, n49436, n48133 );
and U93538 ( n49436, n49357, n49358 );
nand U93539 ( n49353, n49431, n76325 );
nor U93540 ( n49431, n49432, n49433 );
and U93541 ( n49433, n49354, n76181 );
nor U93542 ( n49432, n49434, n49430 );
nand U93543 ( n33772, n76774, n32521 );
nand U93544 ( n14174, n76727, n12587 );
nand U93545 ( n16235, n16322, n76591 );
nor U93546 ( n16322, n16323, n16324 );
and U93547 ( n16324, n16237, n76192 );
nor U93548 ( n16323, n16325, n16321 );
nor U93549 ( n16325, n16328, n14947 );
and U93550 ( n16328, n16240, n16242 );
nand U93551 ( n68044, n67429, n67973 );
nand U93552 ( n47009, n46365, n46926 );
nand U93553 ( n26041, n25424, n25970 );
nand U93554 ( n59182, n58561, n59108 );
nand U93555 ( n28478, n28479, n24607 );
nor U93556 ( n28479, n28480, n28481 );
nor U93557 ( n28480, n4060, n4058 );
nand U93558 ( n61783, n61784, n57739 );
nor U93559 ( n61784, n61785, n61786 );
nor U93560 ( n61785, n6693, n6690 );
nand U93561 ( n35657, n35658, n31823 );
nor U93562 ( n35658, n35659, n35660 );
nor U93563 ( n35659, n3233, n3230 );
nand U93564 ( n70383, n70384, n66415 );
nor U93565 ( n70384, n70385, n70386 );
nor U93566 ( n70385, n5832, n5829 );
and U93567 ( n21835, n28476, n28477 );
nand U93568 ( n28476, n26905, n28482 );
nand U93569 ( n28477, n4047, n28478 );
nand U93570 ( n28482, n28483, n24607 );
and U93571 ( n54928, n61781, n61782 );
nand U93572 ( n61781, n60045, n61787 );
nand U93573 ( n61782, n6679, n61783 );
nand U93574 ( n61787, n61788, n57739 );
and U93575 ( n29150, n35655, n35656 );
nand U93576 ( n35655, n34150, n35661 );
nand U93577 ( n35656, n3217, n35657 );
nand U93578 ( n35661, n35662, n31823 );
and U93579 ( n62817, n70381, n70382 );
nand U93580 ( n70381, n68904, n70387 );
nand U93581 ( n70382, n5815, n70383 );
nand U93582 ( n70387, n70388, n66415 );
nand U93583 ( n33285, n32664, n33218 );
nand U93584 ( n13575, n12775, n13487 );
nand U93585 ( n67827, n67429, n67758 );
nand U93586 ( n46780, n46365, n46711 );
nand U93587 ( n25824, n25424, n25753 );
nand U93588 ( n58962, n58561, n58893 );
nand U93589 ( n33071, n32664, n33002 );
nand U93590 ( n12990, n12775, n12898 );
nand U93591 ( n13303, n12775, n13219 );
nand U93592 ( n68170, n68095, n67429 );
nand U93593 ( n33420, n33338, n32664 );
nand U93594 ( n13739, n13638, n12775 );
nand U93595 ( n47139, n47064, n46365 );
nand U93596 ( n26169, n26092, n25424 );
nand U93597 ( n59308, n59233, n58561 );
nand U93598 ( n15717, n15812, n14958 );
nand U93599 ( n16135, n15812, n15397 );
nor U93600 ( n15802, n15805, n14947 );
and U93601 ( n15805, n15717, n15715 );
nor U93602 ( n16218, n16222, n14947 );
and U93603 ( n16222, n16135, n16134 );
nand U93604 ( n48815, n48884, n48142 );
nand U93605 ( n49184, n48884, n48523 );
nor U93606 ( n49245, n49248, n48133 );
and U93607 ( n49248, n49184, n49183 );
nor U93608 ( n48876, n48879, n48133 );
and U93609 ( n48879, n48815, n48814 );
nand U93610 ( n13020, n12999, n13002 );
nand U93611 ( n13483, n12999, n13432 );
nand U93612 ( n13333, n12999, n13312 );
nor U93613 ( n13573, n13574, n13534 );
nor U93614 ( n13574, n4864, n13539 );
nor U93615 ( n27695, n85, n4269 );
buf U93616 ( n76077, n61176 );
buf U93617 ( n76517, n26979 );
and U93618 ( n28395, n76517, n3910 );
nand U93619 ( n13672, n12999, n13643 );
nand U93620 ( n13632, n13672, n13673 );
nand U93621 ( n13673, n13579, n12732 );
buf U93622 ( n76079, n61176 );
buf U93623 ( n76078, n61176 );
buf U93624 ( n76075, n61176 );
buf U93625 ( n76076, n61176 );
nor U93626 ( n28195, n85, n28127 );
nor U93627 ( n28276, n85, n28208 );
nor U93628 ( n28114, n85, n28045 );
nor U93629 ( n28033, n85, n27969 );
nor U93630 ( n27951, n85, n27887 );
nor U93631 ( n27873, n85, n27805 );
nor U93632 ( n27791, n85, n27720 );
nor U93633 ( n27630, n85, n27566 );
nor U93634 ( n27551, n85, n27480 );
nand U93635 ( n13758, n13825, n13827 );
nand U93636 ( n13827, n13730, n12732 );
nand U93637 ( n33858, n76772, n32537 );
nand U93638 ( n13825, n12999, n13880 );
nor U93639 ( n48977, n48979, n48133 );
and U93640 ( n48979, n48895, n48896 );
nand U93641 ( n48891, n48974, n76325 );
nor U93642 ( n48974, n48975, n48976 );
and U93643 ( n48976, n48892, n76180 );
nor U93644 ( n48975, n48977, n48973 );
nor U93645 ( n11308, n2, n10785 );
and U93646 ( n28287, n28395, n3797 );
nand U93647 ( n46517, n46365, n46450 );
nand U93648 ( n67578, n67429, n67514 );
nand U93649 ( n32813, n32664, n32749 );
nand U93650 ( n25573, n25424, n25509 );
nand U93651 ( n58710, n58561, n58646 );
nand U93652 ( n13939, n14059, n14060 );
nand U93653 ( n14060, n13893, n12732 );
nand U93654 ( n14059, n12999, n13889 );
nor U93655 ( n27645, n68, n4269 );
nor U93656 ( n27687, n83, n4269 );
nor U93657 ( n27634, n65, n4269 );
nor U93658 ( n27679, n80, n4269 );
nor U93659 ( n27663, n74, n4269 );
nor U93660 ( n27671, n77, n4269 );
nor U93661 ( n27655, n71, n4269 );
nand U93662 ( n54159, n54160, n45522 );
nor U93663 ( n54160, n54161, n54162 );
nor U93664 ( n54161, n7620, n7615 );
and U93665 ( n42363, n54153, n54154 );
nand U93666 ( n54154, n7603, n54155 );
nand U93667 ( n54153, n47884, n54159 );
nand U93668 ( n54155, n54156, n45522 );
nor U93669 ( n60830, n344, n6902 );
nor U93670 ( n60814, n337, n6902 );
nor U93671 ( n60838, n348, n6902 );
nor U93672 ( n60798, n329, n6902 );
nor U93673 ( n60787, n325, n6902 );
nor U93674 ( n60806, n333, n6902 );
nor U93675 ( n60822, n340, n6902 );
nor U93676 ( n60846, n350, n6902 );
buf U93677 ( n76259, n60119 );
and U93678 ( n61676, n76259, n6543 );
nor U93679 ( n28136, n68, n28127 );
nor U93680 ( n28172, n80, n28127 );
nor U93681 ( n28152, n74, n28127 );
nor U93682 ( n28164, n77, n28127 );
nor U93683 ( n28144, n71, n28127 );
nor U93684 ( n27978, n68, n27969 );
nor U93685 ( n27896, n68, n27887 );
nor U93686 ( n27814, n68, n27805 );
nor U93687 ( n27575, n68, n27566 );
nor U93688 ( n27490, n68, n27480 );
nor U93689 ( n28098, n83, n28045 );
nor U93690 ( n27775, n83, n27720 );
nor U93691 ( n28044, n65, n28045 );
nor U93692 ( n27719, n65, n27720 );
nor U93693 ( n28090, n80, n28045 );
nor U93694 ( n28010, n80, n27969 );
nor U93695 ( n27928, n80, n27887 );
nor U93696 ( n27846, n80, n27805 );
nor U93697 ( n27767, n80, n27720 );
nor U93698 ( n27607, n80, n27566 );
nor U93699 ( n27526, n80, n27480 );
nor U93700 ( n28233, n74, n28208 );
nor U93701 ( n27994, n74, n27969 );
nor U93702 ( n27912, n74, n27887 );
nor U93703 ( n27830, n74, n27805 );
nor U93704 ( n27591, n74, n27566 );
nor U93705 ( n27508, n74, n27480 );
nor U93706 ( n28241, n77, n28208 );
nor U93707 ( n28002, n77, n27969 );
nor U93708 ( n27920, n77, n27887 );
nor U93709 ( n27838, n77, n27805 );
nor U93710 ( n27599, n77, n27566 );
nor U93711 ( n27517, n77, n27480 );
nor U93712 ( n28225, n71, n28208 );
nor U93713 ( n27986, n71, n27969 );
nor U93714 ( n27904, n71, n27887 );
nor U93715 ( n27822, n71, n27805 );
nor U93716 ( n27583, n71, n27566 );
nor U93717 ( n27499, n71, n27480 );
nor U93718 ( n28249, n80, n28208 );
nand U93719 ( n14153, n14263, n14264 );
nand U93720 ( n14263, n12775, n14162 );
nand U93721 ( n68511, n68599, n68600 );
nand U93722 ( n68599, n67429, n68518 );
nand U93723 ( n33755, n33843, n33844 );
nand U93724 ( n33843, n32664, n33762 );
nand U93725 ( n47490, n47578, n47579 );
nand U93726 ( n47578, n46365, n47497 );
nand U93727 ( n26510, n26598, n26599 );
nand U93728 ( n26598, n25424, n26517 );
nand U93729 ( n59649, n59740, n59741 );
nand U93730 ( n59740, n58561, n59656 );
nor U93731 ( n28217, n68, n28208 );
nor U93732 ( n28180, n83, n28127 );
nor U93733 ( n28126, n65, n28127 );
nor U93734 ( n61336, n344, n61282 );
nor U93735 ( n61320, n337, n61282 );
nor U93736 ( n61304, n329, n61282 );
nor U93737 ( n61312, n333, n61282 );
nor U93738 ( n61328, n340, n61282 );
nor U93739 ( n61359, n350, n61282 );
nor U93740 ( n28054, n68, n28045 );
nor U93741 ( n27729, n68, n27720 );
nor U93742 ( n28018, n83, n27969 );
nor U93743 ( n27936, n83, n27887 );
nor U93744 ( n27858, n83, n27805 );
nor U93745 ( n27615, n83, n27566 );
nor U93746 ( n27535, n83, n27480 );
nor U93747 ( n28207, n65, n28208 );
nor U93748 ( n27968, n65, n27969 );
nor U93749 ( n27886, n65, n27887 );
nor U93750 ( n27804, n65, n27805 );
nor U93751 ( n27565, n65, n27566 );
nor U93752 ( n27479, n65, n27480 );
nor U93753 ( n28074, n74, n28045 );
nor U93754 ( n27745, n74, n27720 );
nor U93755 ( n28082, n77, n28045 );
nor U93756 ( n27759, n77, n27720 );
nor U93757 ( n28066, n71, n28045 );
nor U93758 ( n27737, n71, n27720 );
nor U93759 ( n61475, n344, n61372 );
nor U93760 ( n61245, n344, n61204 );
nor U93761 ( n61159, n344, n61118 );
nor U93762 ( n61081, n344, n61034 );
nor U93763 ( n60997, n344, n60953 );
nor U93764 ( n60915, n344, n60871 );
nor U93765 ( n60757, n344, n60716 );
nor U93766 ( n60678, n344, n60629 );
nor U93767 ( n61143, n337, n61118 );
nor U93768 ( n61059, n337, n61034 );
nor U93769 ( n60981, n337, n60953 );
nor U93770 ( n60741, n337, n60716 );
nor U93771 ( n60657, n337, n60629 );
nor U93772 ( n61253, n348, n61204 );
nor U93773 ( n60923, n348, n60871 );
nor U93774 ( n61381, n329, n61372 );
nor U93775 ( n61127, n329, n61118 );
nor U93776 ( n61043, n329, n61034 );
nor U93777 ( n60962, n329, n60953 );
nor U93778 ( n60725, n329, n60716 );
nor U93779 ( n60639, n329, n60629 );
nor U93780 ( n61203, n325, n61204 );
nor U93781 ( n60870, n325, n60871 );
nor U93782 ( n61389, n333, n61372 );
nor U93783 ( n61135, n333, n61118 );
nor U93784 ( n61051, n333, n61034 );
nor U93785 ( n60970, n333, n60953 );
nor U93786 ( n60733, n333, n60716 );
nor U93787 ( n60648, n333, n60629 );
nor U93788 ( n61467, n340, n61372 );
nor U93789 ( n61151, n340, n61118 );
nor U93790 ( n61067, n340, n61034 );
nor U93791 ( n60989, n340, n60953 );
nor U93792 ( n60749, n340, n60716 );
nor U93793 ( n60666, n340, n60629 );
nor U93794 ( n61459, n337, n61372 );
nor U93795 ( n61269, n350, n61204 );
nor U93796 ( n61192, n350, n61118 );
nor U93797 ( n61104, n350, n61034 );
nor U93798 ( n61020, n350, n60953 );
nor U93799 ( n60939, n350, n60871 );
nor U93800 ( n60783, n350, n60716 );
nor U93801 ( n60703, n350, n60629 );
nor U93802 ( n28261, n83, n28208 );
nor U93803 ( n61498, n350, n61372 );
nor U93804 ( n61344, n348, n61282 );
nor U93805 ( n61281, n325, n61282 );
nor U93806 ( n61229, n337, n61204 );
nor U93807 ( n60899, n337, n60871 );
nor U93808 ( n61483, n348, n61372 );
nor U93809 ( n61167, n348, n61118 );
nor U93810 ( n61089, n348, n61034 );
nor U93811 ( n61005, n348, n60953 );
nor U93812 ( n60765, n348, n60716 );
nor U93813 ( n60687, n348, n60629 );
nor U93814 ( n61213, n329, n61204 );
nor U93815 ( n60883, n329, n60871 );
nor U93816 ( n61371, n325, n61372 );
nor U93817 ( n61117, n325, n61118 );
nor U93818 ( n61033, n325, n61034 );
nor U93819 ( n60952, n325, n60953 );
nor U93820 ( n60715, n325, n60716 );
nor U93821 ( n60628, n325, n60629 );
nor U93822 ( n61221, n333, n61204 );
nor U93823 ( n60891, n333, n60871 );
nor U93824 ( n61237, n340, n61204 );
nor U93825 ( n60907, n340, n60871 );
and U93826 ( n12893, n12838, n12999 );
and U93827 ( n61509, n61676, n6429 );
not U93828 ( n7848, n48412 );
nand U93829 ( n67494, n67453, n67495 );
nand U93830 ( n32729, n32688, n32730 );
nand U93831 ( n25489, n25448, n25490 );
nand U93832 ( n58626, n58585, n58627 );
nor U93833 ( n28316, n52, n28291 );
nor U93834 ( n28359, n58, n28291 );
nor U93835 ( n28330, n54, n28291 );
nor U93836 ( n28302, n50, n28291 );
nor U93837 ( n28345, n56, n28291 );
nor U93838 ( n28279, n48, n28291 );
nor U93839 ( n28373, n60, n28291 );
nor U93840 ( n28387, n62, n28291 );
nand U93841 ( n5871, n28357, n28358 );
nor U93842 ( n28357, n28367, n28368 );
nor U93843 ( n28358, n28359, n28360 );
nor U93844 ( n28367, n27099, n28297 );
nand U93845 ( n5896, n28277, n28278 );
nor U93846 ( n28277, n28294, n28295 );
nor U93847 ( n28278, n28279, n28280 );
nor U93848 ( n28294, n27043, n28297 );
nand U93849 ( n5866, n28371, n28372 );
nor U93850 ( n28371, n28381, n28382 );
nor U93851 ( n28372, n28373, n28374 );
nor U93852 ( n28381, n27110, n28297 );
nand U93853 ( n5861, n28385, n28386 );
nor U93854 ( n28385, n28396, n28397 );
nor U93855 ( n28386, n28387, n28388 );
nor U93856 ( n28397, n27133, n28297 );
nand U93857 ( n68614, n76705, n67193 );
nand U93858 ( n26613, n76751, n25295 );
nand U93859 ( n59755, n76684, n58431 );
nand U93860 ( n5886, n28314, n28315 );
nor U93861 ( n28314, n28324, n28325 );
nor U93862 ( n28315, n28316, n28317 );
nor U93863 ( n28324, n27066, n28297 );
nand U93864 ( n5881, n28328, n28329 );
nor U93865 ( n28328, n28339, n28340 );
nor U93866 ( n28329, n28330, n28331 );
nor U93867 ( n28339, n27077, n28297 );
nand U93868 ( n5891, n28300, n28301 );
nor U93869 ( n28300, n28310, n28311 );
nor U93870 ( n28301, n28302, n28303 );
nor U93871 ( n28310, n27055, n28297 );
nand U93872 ( n5876, n28343, n28344 );
nor U93873 ( n28343, n28353, n28354 );
nor U93874 ( n28344, n28345, n28346 );
nor U93875 ( n28353, n27088, n28297 );
nor U93876 ( n61552, n312, n61513 );
nor U93877 ( n61636, n317, n61513 );
nor U93878 ( n61538, n309, n61513 );
nor U93879 ( n61524, n307, n61513 );
nor U93880 ( n61567, n314, n61513 );
nor U93881 ( n61650, n319, n61513 );
nor U93882 ( n61668, n322, n61513 );
nor U93883 ( n61501, n304, n61513 );
nor U93884 ( n27318, n50, n27311 );
nor U93885 ( n27236, n50, n27229 );
nor U93886 ( n27154, n50, n27147 );
nor U93887 ( n27368, n62, n27311 );
nor U93888 ( n27286, n62, n27229 );
nor U93889 ( n27202, n62, n27147 );
nor U93890 ( n27360, n60, n27311 );
nor U93891 ( n27278, n60, n27229 );
nor U93892 ( n27194, n60, n27147 );
nor U93893 ( n27305, n48, n27311 );
nor U93894 ( n27223, n48, n27229 );
nor U93895 ( n27141, n48, n27147 );
nor U93896 ( n27352, n58, n27311 );
nor U93897 ( n27270, n58, n27229 );
nor U93898 ( n27186, n58, n27147 );
nor U93899 ( n27334, n54, n27311 );
nor U93900 ( n27254, n54, n27229 );
nor U93901 ( n27170, n54, n27147 );
nor U93902 ( n27344, n56, n27311 );
nor U93903 ( n27262, n56, n27229 );
nor U93904 ( n27178, n56, n27147 );
nor U93905 ( n27326, n52, n27311 );
nor U93906 ( n27246, n52, n27229 );
nor U93907 ( n27162, n52, n27147 );
nand U93908 ( n12606, n61634, n61635 );
nor U93909 ( n61634, n61644, n61645 );
nor U93910 ( n61635, n61636, n61637 );
nor U93911 ( n61644, n60243, n61519 );
nand U93912 ( n12601, n61648, n61649 );
nor U93913 ( n61648, n61658, n61659 );
nor U93914 ( n61649, n61650, n61651 );
nor U93915 ( n61658, n60254, n61519 );
nand U93916 ( n12596, n61666, n61667 );
nor U93917 ( n61666, n61677, n61678 );
nor U93918 ( n61667, n61668, n61669 );
nor U93919 ( n61678, n60277, n61519 );
nand U93920 ( n12631, n61499, n61500 );
nor U93921 ( n61499, n61516, n61517 );
nor U93922 ( n61500, n61501, n61502 );
nor U93923 ( n61516, n60184, n61519 );
nand U93924 ( n12616, n61550, n61551 );
nor U93925 ( n61550, n61561, n61562 );
nor U93926 ( n61551, n61552, n61553 );
nor U93927 ( n61561, n60218, n61519 );
nand U93928 ( n12621, n61536, n61537 );
nor U93929 ( n61536, n61546, n61547 );
nor U93930 ( n61537, n61538, n61539 );
nor U93931 ( n61546, n60207, n61519 );
nand U93932 ( n12626, n61522, n61523 );
nor U93933 ( n61522, n61532, n61533 );
nor U93934 ( n61523, n61524, n61525 );
nor U93935 ( n61532, n60196, n61519 );
nand U93936 ( n12611, n61565, n61566 );
nor U93937 ( n61565, n61575, n61576 );
nor U93938 ( n61566, n61567, n61568 );
nor U93939 ( n61575, n60229, n61519 );
nor U93940 ( n12763, n12822, n12832 );
and U93941 ( n12832, n12823, n12824 );
nor U93942 ( n60500, n317, n60454 );
nor U93943 ( n60413, n317, n60374 );
nor U93944 ( n60328, n317, n60289 );
nor U93945 ( n60484, n312, n60454 );
nor U93946 ( n60397, n312, n60374 );
nor U93947 ( n60312, n312, n60289 );
nor U93948 ( n60508, n319, n60454 );
nor U93949 ( n60421, n319, n60374 );
nor U93950 ( n60336, n319, n60289 );
nor U93951 ( n60464, n307, n60454 );
nor U93952 ( n60381, n307, n60374 );
nor U93953 ( n60296, n307, n60289 );
nor U93954 ( n60448, n304, n60454 );
nor U93955 ( n60368, n304, n60374 );
nor U93956 ( n60283, n304, n60289 );
nor U93957 ( n60472, n309, n60454 );
nor U93958 ( n60389, n309, n60374 );
nor U93959 ( n60304, n309, n60289 );
nor U93960 ( n60492, n314, n60454 );
nor U93961 ( n60405, n314, n60374 );
nor U93962 ( n60320, n314, n60289 );
nor U93963 ( n60516, n322, n60454 );
nor U93964 ( n60429, n322, n60374 );
nor U93965 ( n60347, n322, n60289 );
buf U93966 ( n76081, n61176 );
nor U93967 ( n27650, n50, n27642 );
nor U93968 ( n27708, n62, n27642 );
nor U93969 ( n27692, n60, n27642 );
nor U93970 ( n27641, n48, n27642 );
nor U93971 ( n27684, n58, n27642 );
nor U93972 ( n27668, n54, n27642 );
nor U93973 ( n27676, n56, n27642 );
nor U93974 ( n27660, n52, n27642 );
nor U93975 ( n60835, n317, n60795 );
nor U93976 ( n60819, n312, n60795 );
nor U93977 ( n60843, n319, n60795 );
nor U93978 ( n60803, n307, n60795 );
nor U93979 ( n60794, n304, n60795 );
nor U93980 ( n60811, n309, n60795 );
nor U93981 ( n60827, n314, n60795 );
nor U93982 ( n60859, n322, n60795 );
nor U93983 ( n27465, n62, n27397 );
nor U93984 ( n27394, n48, n27397 );
nor U93985 ( n27436, n58, n27397 );
nor U93986 ( n27446, n60, n27397 );
nor U93987 ( n27131, n62, n27044 );
nor U93988 ( n27108, n60, n27044 );
nor U93989 ( n27040, n48, n27044 );
nor U93990 ( n27097, n58, n27044 );
nor U93991 ( n60587, n317, n60545 );
nor U93992 ( n60542, n304, n60545 );
nor U93993 ( n60595, n319, n60545 );
nor U93994 ( n60614, n322, n60545 );
nor U93995 ( n27404, n50, n27397 );
nor U93996 ( n27053, n50, n27044 );
nor U93997 ( n27420, n54, n27397 );
nor U93998 ( n27075, n54, n27044 );
nor U93999 ( n27086, n56, n27044 );
nor U94000 ( n27428, n56, n27397 );
nor U94001 ( n27412, n52, n27397 );
nor U94002 ( n27064, n52, n27044 );
nor U94003 ( n60241, n317, n60185 );
nor U94004 ( n60252, n319, n60185 );
nor U94005 ( n60181, n304, n60185 );
nor U94006 ( n60275, n322, n60185 );
nor U94007 ( n46355, n46392, n46404 );
and U94008 ( n46404, n46393, n46394 );
nor U94009 ( n60571, n312, n60545 );
nor U94010 ( n60216, n312, n60185 );
nor U94011 ( n60194, n307, n60185 );
nor U94012 ( n60560, n309, n60545 );
nor U94013 ( n60205, n309, n60185 );
nor U94014 ( n60579, n314, n60545 );
nor U94015 ( n60227, n314, n60185 );
nor U94016 ( n60552, n307, n60545 );
nand U94017 ( n14282, n76724, n12607 );
nand U94018 ( n14387, n76725, n12615 );
not U94019 ( n162, n23209 );
buf U94020 ( n76749, n4687 );
buf U94021 ( n76080, n61176 );
nand U94022 ( n47593, n76657, n46241 );
nand U94023 ( n67432, n67453, n67454 );
nand U94024 ( n67454, n67455, n67456 );
nand U94025 ( n67455, n67457, n67458 );
nand U94026 ( n32667, n32688, n32689 );
nand U94027 ( n32689, n32690, n32691 );
nand U94028 ( n32690, n32692, n32693 );
nand U94029 ( n25427, n25448, n25449 );
nand U94030 ( n25449, n25450, n25451 );
nand U94031 ( n25450, n25452, n25453 );
nand U94032 ( n58564, n58585, n58586 );
nand U94033 ( n58586, n58587, n58588 );
nand U94034 ( n58587, n58589, n58590 );
nand U94035 ( n67453, n67429, n67496 );
nand U94036 ( n32688, n32664, n32731 );
nand U94037 ( n25448, n25424, n25491 );
nand U94038 ( n58585, n58561, n58628 );
not U94039 ( n3823, n24323 );
not U94040 ( n434, n56330 );
not U94041 ( n5580, n65905 );
not U94042 ( n6455, n57446 );
nand U94043 ( n13207, n13157, n12999 );
nand U94044 ( n32851, n32737, n32833 );
nand U94045 ( n46569, n46438, n46536 );
nand U94046 ( n67616, n67502, n67598 );
nand U94047 ( n25611, n25497, n25593 );
nand U94048 ( n58748, n58634, n58730 );
nand U94049 ( n33333, n33359, n33360 );
nand U94050 ( n33360, n33288, n32630 );
nand U94051 ( n33359, n32737, n33342 );
nand U94052 ( n68090, n68116, n68117 );
nand U94053 ( n68117, n68047, n67395 );
nand U94054 ( n47059, n47085, n47086 );
nand U94055 ( n47086, n47012, n46331 );
nand U94056 ( n26087, n26113, n26114 );
nand U94057 ( n26114, n26044, n25390 );
nand U94058 ( n59228, n59254, n59255 );
nand U94059 ( n59255, n59185, n58527 );
nand U94060 ( n68116, n67502, n68099 );
nand U94061 ( n47085, n46438, n47068 );
nand U94062 ( n26113, n25497, n26096 );
nand U94063 ( n59254, n58634, n59237 );
nand U94064 ( n67970, n76058, n67937 );
nand U94065 ( n46923, n76101, n46890 );
nand U94066 ( n25967, n76156, n25934 );
nand U94067 ( n59105, n76084, n59072 );
nand U94068 ( n33215, n76128, n33174 );
nand U94069 ( n33095, n76127, n33078 );
nand U94070 ( n67851, n76057, n67834 );
nand U94071 ( n46804, n76100, n46787 );
nand U94072 ( n25848, n76155, n25831 );
nand U94073 ( n58986, n76083, n58969 );
nand U94074 ( n68185, n68246, n68247 );
nand U94075 ( n68247, n68163, n67395 );
nand U94076 ( n47154, n47215, n47216 );
nand U94077 ( n47216, n47132, n46331 );
nand U94078 ( n26184, n26245, n26246 );
nand U94079 ( n26246, n26162, n25390 );
nand U94080 ( n59323, n59384, n59385 );
nand U94081 ( n59385, n59301, n58527 );
nand U94082 ( n68246, n76058, n68291 );
nand U94083 ( n47215, n76101, n47260 );
nand U94084 ( n26245, n76156, n26290 );
nand U94085 ( n59384, n76084, n59429 );
nand U94086 ( n33438, n33491, n33492 );
nand U94087 ( n33492, n33413, n32630 );
nand U94088 ( n33491, n76128, n33535 );
not U94089 ( n7344, n45317 );
nand U94090 ( n8322, n21210, n21211 );
nor U94091 ( n21211, n4975, n21212 );
nor U94092 ( n21210, n4858, n14658 );
nor U94093 ( n21212, n5134, n11733 );
nand U94094 ( n68338, n68435, n68436 );
nand U94095 ( n68436, n68301, n67395 );
nand U94096 ( n33582, n33679, n33680 );
nand U94097 ( n33680, n33545, n32630 );
nand U94098 ( n26337, n26434, n26435 );
nand U94099 ( n26435, n26300, n25390 );
nand U94100 ( n59476, n59573, n59574 );
nand U94101 ( n59574, n59439, n58527 );
nand U94102 ( n68435, n76058, n68299 );
nand U94103 ( n33679, n76128, n33543 );
nand U94104 ( n26434, n76156, n26298 );
nand U94105 ( n59573, n76084, n59437 );
nand U94106 ( n47307, n47403, n47404 );
nand U94107 ( n47404, n47270, n46331 );
nand U94108 ( n47403, n76101, n47267 );
nand U94109 ( n14264, n5219, n12732 );
nand U94110 ( n26969, n28410, n28411 );
or U94111 ( n28411, n4273, n27379 );
nor U94112 ( n28410, n27788, n4274 );
nand U94113 ( n60109, n61719, n61720 );
or U94114 ( n61720, n6905, n60527 );
nor U94115 ( n61719, n60936, n6907 );
nand U94116 ( n60104, n61723, n61724 );
nand U94117 ( n61724, n60531, n61717 );
nor U94118 ( n61723, n60857, n60941 );
nand U94119 ( n26964, n28414, n28415 );
nand U94120 ( n28415, n27383, n28408 );
nor U94121 ( n28414, n27706, n27793 );
nor U94122 ( n27467, n26964, n28412 );
nor U94123 ( n60616, n60104, n61721 );
nor U94124 ( n27952, n26935, n4268 );
nor U94125 ( n61105, n60075, n6900 );
nor U94126 ( n27706, n27460, n28408 );
nor U94127 ( n60857, n60609, n61717 );
nand U94128 ( n28204, n28268, n76517 );
nor U94129 ( n28268, n28269, n28270 );
and U94130 ( n28270, n28209, P1_P2_STATE2_REG_3_ );
nor U94131 ( n28269, n28271, n28272 );
nand U94132 ( n61368, n61490, n76259 );
nor U94133 ( n61490, n61491, n61492 );
and U94134 ( n61492, n61373, P2_P2_STATE2_REG_3_ );
nor U94135 ( n61491, n61493, n61494 );
not U94136 ( n4283, n27383 );
not U94137 ( n6915, n60531 );
nand U94138 ( n69629, n69456, n69370 );
nand U94139 ( n34214, n35591, n35592 );
or U94140 ( n35592, n3435, n34624 );
nor U94141 ( n35591, n35029, n3437 );
nand U94142 ( n68968, n70319, n70320 );
or U94143 ( n70320, n6050, n69370 );
nor U94144 ( n70319, n69767, n6052 );
nand U94145 ( n70171, n69927, n69451 );
nand U94146 ( n35441, n35191, n34707 );
nand U94147 ( n68963, n70323, n70324 );
nand U94148 ( n70324, n69374, n70317 );
nor U94149 ( n70323, n69691, n69772 );
nor U94150 ( n34712, n34209, n35593 );
nor U94151 ( n69456, n68963, n70321 );
nor U94152 ( n69927, n68934, n6045 );
nor U94153 ( n35191, n34180, n3430 );
nand U94154 ( n27883, n27943, n76517 );
nor U94155 ( n27943, n27944, n27945 );
and U94156 ( n27945, n27888, P1_P2_STATE2_REG_3_ );
nor U94157 ( n27944, n27946, n27947 );
nand U94158 ( n61030, n61096, n76259 );
nor U94159 ( n61096, n61097, n61098 );
and U94160 ( n61098, n61035, P2_P2_STATE2_REG_3_ );
nor U94161 ( n61097, n61099, n61100 );
nor U94162 ( n27946, n27948, n27124 );
nor U94163 ( n27948, n27882, n4260 );
not U94164 ( n4260, n27887 );
nor U94165 ( n61099, n61101, n60268 );
nor U94166 ( n61101, n61029, n6893 );
not U94167 ( n6893, n61034 );
nor U94168 ( n28271, n28273, n27124 );
nor U94169 ( n28273, n28203, n4259 );
not U94170 ( n4259, n28208 );
nor U94171 ( n61493, n61495, n60268 );
nor U94172 ( n61495, n61367, n6892 );
not U94173 ( n6892, n61372 );
nand U94174 ( n34887, n34712, n34624 );
nand U94175 ( n34209, n35595, n35596 );
nand U94176 ( n35596, n34628, n35589 );
nor U94177 ( n35595, n34951, n35034 );
nor U94178 ( n34951, n34705, n35589 );
nor U94179 ( n69691, n69449, n70317 );
nand U94180 ( n70167, n70227, n76193 );
nor U94181 ( n70227, n70228, n70229 );
and U94182 ( n70229, n70172, P2_P3_STATE2_REG_3_ );
nor U94183 ( n70228, n70230, n70231 );
nand U94184 ( n35437, n35499, n76461 );
nor U94185 ( n35499, n35500, n35501 );
and U94186 ( n35501, n35442, P1_P3_STATE2_REG_3_ );
nor U94187 ( n35500, n35502, n35503 );
not U94188 ( n3445, n34628 );
not U94189 ( n6060, n69374 );
nor U94190 ( n70230, n70232, n69121 );
nor U94191 ( n70232, n70166, n6037 );
not U94192 ( n6037, n70171 );
nor U94193 ( n35502, n35504, n34369 );
nor U94194 ( n35504, n35436, n3422 );
not U94195 ( n3422, n35441 );
nand U94196 ( n48344, n48407, n76325 );
nor U94197 ( n48407, n48408, n48409 );
and U94198 ( n48409, n48350, n76179 );
nor U94199 ( n48408, n48410, n48406 );
nand U94200 ( n35126, n35191, n34371 );
nand U94201 ( n69862, n69927, n69123 );
and U94202 ( n48345, n48419, n7833 );
nor U94203 ( n48419, n47934, n47935 );
nand U94204 ( n35122, n35182, n76461 );
nor U94205 ( n35182, n35183, n35184 );
and U94206 ( n35184, n35127, P1_P3_STATE2_REG_3_ );
nor U94207 ( n35183, n35185, n35186 );
nand U94208 ( n69858, n69918, n76193 );
nor U94209 ( n69918, n69919, n69920 );
and U94210 ( n69920, n69863, P2_P3_STATE2_REG_3_ );
nor U94211 ( n69919, n69921, n69922 );
nor U94212 ( n35185, n35187, n34369 );
nor U94213 ( n35187, n35121, n3423 );
not U94214 ( n3423, n35126 );
nor U94215 ( n69921, n69923, n69121 );
nor U94216 ( n69923, n69857, n6038 );
not U94217 ( n6038, n69862 );
nor U94218 ( n48410, n48414, n48133 );
nor U94219 ( n48414, n7842, n48345 );
not U94220 ( n7842, n48349 );
nand U94221 ( n14270, n14364, n14163 );
nand U94222 ( n14364, n5225, n12999 );
not U94223 ( n4712, n11494 );
nand U94224 ( n29195, n35695, n35696 );
nor U94225 ( n35696, n3242, n35697 );
nor U94226 ( n35695, n3117, n34153 );
nor U94227 ( n35697, n3387, n31817 );
nand U94228 ( n21878, n28516, n28517 );
nor U94229 ( n28517, n4067, n28518 );
nor U94230 ( n28516, n3960, n26908 );
nor U94231 ( n28518, n4224, n24601 );
nand U94232 ( n62913, n70421, n70422 );
nor U94233 ( n70422, n5842, n70423 );
nor U94234 ( n70421, n5718, n68907 );
nor U94235 ( n70423, n6002, n66409 );
nand U94236 ( n54969, n61821, n61822 );
nor U94237 ( n61822, n6699, n61823 );
nor U94238 ( n61821, n6593, n60048 );
nor U94239 ( n61823, n6857, n57733 );
and U94240 ( n35515, n76461, n3067 );
and U94241 ( n70243, n76193, n5668 );
buf U94242 ( n76461, n34224 );
buf U94243 ( n76193, n68978 );
nand U94244 ( n43332, n7409, n43361 );
nand U94245 ( n43361, n43362, n43363 );
nand U94246 ( n43286, n7408, n43287 );
nand U94247 ( n35552, n35553, n35554 );
or U94248 ( n35553, n35516, n34329 );
nand U94249 ( n35554, n35514, n140 );
nand U94250 ( n70280, n70281, n70282 );
or U94251 ( n70281, n70244, n69081 );
nand U94252 ( n70282, n70242, n413 );
nand U94253 ( n35576, n35577, n35578 );
or U94254 ( n35577, n35516, n34372 );
nand U94255 ( n35578, n35514, n147 );
nand U94256 ( n70304, n70305, n70306 );
or U94257 ( n70305, n70244, n69124 );
nand U94258 ( n70306, n70242, n419 );
nand U94259 ( n35560, n35561, n35562 );
or U94260 ( n35561, n35516, n34340 );
nand U94261 ( n35562, n35514, n143 );
nand U94262 ( n35568, n35569, n35570 );
or U94263 ( n35569, n35516, n34351 );
nand U94264 ( n35570, n35514, n145 );
nand U94265 ( n35543, n35544, n35545 );
or U94266 ( n35544, n35516, n34318 );
nand U94267 ( n35545, n35514, n138 );
nand U94268 ( n35535, n35536, n35537 );
or U94269 ( n35536, n35516, n34307 );
nand U94270 ( n35537, n35514, n135 );
nand U94271 ( n70263, n70264, n70265 );
or U94272 ( n70264, n70244, n69059 );
nand U94273 ( n70265, n70242, n408 );
nand U94274 ( n70271, n70272, n70273 );
or U94275 ( n70272, n70244, n69070 );
nand U94276 ( n70273, n70242, n410 );
nand U94277 ( n70296, n70297, n70298 );
or U94278 ( n70297, n70244, n69103 );
nand U94279 ( n70298, n70242, n418 );
nand U94280 ( n70288, n70289, n70290 );
or U94281 ( n70289, n70244, n69092 );
nand U94282 ( n70290, n70242, n415 );
nand U94283 ( n35511, n35512, n35513 );
or U94284 ( n35512, n35516, n34283 );
nand U94285 ( n35513, n35514, n130 );
nand U94286 ( n70239, n70240, n70241 );
or U94287 ( n70240, n70244, n69035 );
nand U94288 ( n70241, n70242, n403 );
nand U94289 ( n35527, n35528, n35529 );
or U94290 ( n35528, n35516, n34296 );
nand U94291 ( n35529, n35514, n133 );
nand U94292 ( n70255, n70256, n70257 );
or U94293 ( n70256, n70244, n69048 );
nand U94294 ( n70257, n70242, n405 );
nand U94295 ( n47579, n7873, n46331 );
nand U94296 ( n68600, n6083, n67395 );
nand U94297 ( n33844, n3468, n32630 );
nand U94298 ( n26599, n4305, n25390 );
nand U94299 ( n59741, n6938, n58527 );
nand U94300 ( n47892, n47893, n47894 );
nand U94301 ( n47894, n7343, n47884 );
nand U94302 ( n47893, n7602, n7569 );
nand U94303 ( n14664, n14665, n14667 );
nand U94304 ( n14667, n4711, n14654 );
nand U94305 ( n14665, n4948, n4918 );
nand U94306 ( n28041, n28105, n76517 );
nor U94307 ( n28105, n28106, n28107 );
and U94308 ( n28107, n28042, P1_P2_STATE2_REG_3_ );
nor U94309 ( n28106, n28108, n28109 );
nand U94310 ( n61200, n61260, n76259 );
nor U94311 ( n61260, n61261, n61262 );
and U94312 ( n61262, n61201, P2_P2_STATE2_REG_3_ );
nor U94313 ( n61261, n61263, n61264 );
nand U94314 ( n58486, n54947, n60034 );
nand U94315 ( n25347, n21856, n26894 );
nand U94316 ( n32589, n29169, n34139 );
nand U94317 ( n67354, n62891, n68893 );
nor U94318 ( n28109, n28110, n27124 );
nor U94319 ( n28110, n28040, n4263 );
not U94320 ( n4263, n28045 );
nor U94321 ( n61264, n61265, n60268 );
nor U94322 ( n61265, n61199, n6895 );
not U94323 ( n6895, n61204 );
nand U94324 ( n35278, n35340, n76461 );
nor U94325 ( n35340, n35341, n35342 );
and U94326 ( n35342, n35279, P1_P3_STATE2_REG_3_ );
nor U94327 ( n35341, n35343, n35344 );
nand U94328 ( n70012, n70072, n76193 );
nor U94329 ( n70072, n70073, n70074 );
and U94330 ( n70074, n70013, P2_P3_STATE2_REG_3_ );
nor U94331 ( n70073, n70075, n70076 );
nor U94332 ( n27786, n27787, n27124 );
nor U94333 ( n27787, n27715, n4264 );
not U94334 ( n4264, n27720 );
nand U94335 ( n35282, n35033, n34707 );
nand U94336 ( n70016, n69771, n69451 );
nand U94337 ( n69705, n69771, n69123 );
nor U94338 ( n60934, n60935, n60268 );
nor U94339 ( n60935, n60866, n6897 );
not U94340 ( n6897, n60871 );
nand U94341 ( n34965, n35033, n34371 );
nor U94342 ( n35027, n35028, n34369 );
nor U94343 ( n35028, n34960, n3427 );
not U94344 ( n3427, n34965 );
nor U94345 ( n69765, n69766, n69121 );
nor U94346 ( n69766, n69700, n6042 );
not U94347 ( n6042, n69705 );
nor U94348 ( n35344, n35345, n34369 );
nor U94349 ( n35345, n35277, n3425 );
not U94350 ( n3425, n35282 );
nor U94351 ( n70076, n70077, n69121 );
nor U94352 ( n70077, n70011, n6040 );
not U94353 ( n6040, n70016 );
nand U94354 ( n9383, n4764, n9418 );
nand U94355 ( n9418, n9419, n9420 );
nand U94356 ( n9325, n4763, n9327 );
not U94357 ( n863, n45161 );
nand U94358 ( n27801, n27865, n76517 );
nor U94359 ( n27865, n27866, n27867 );
and U94360 ( n27867, n27806, P1_P2_STATE2_REG_3_ );
nor U94361 ( n27866, n27868, n27869 );
nand U94362 ( n60949, n61012, n76259 );
nor U94363 ( n61012, n61013, n61014 );
and U94364 ( n61014, n60954, P2_P2_STATE2_REG_3_ );
nor U94365 ( n61013, n61015, n61016 );
nor U94366 ( n27868, n27870, n27124 );
nor U94367 ( n27870, n27800, n4267 );
not U94368 ( n4267, n27805 );
nor U94369 ( n61015, n61017, n60268 );
nor U94370 ( n61017, n60948, n6899 );
not U94371 ( n6899, n60953 );
nor U94372 ( n28028, n28030, n27124 );
nor U94373 ( n28030, n27964, n4265 );
not U94374 ( n4265, n27969 );
nor U94375 ( n61187, n61189, n60268 );
nor U94376 ( n61189, n61113, n6898 );
not U94377 ( n6898, n61118 );
nand U94378 ( n27965, n28025, n76517 );
nor U94379 ( n28025, n28026, n28027 );
and U94380 ( n28027, n27970, P1_P2_STATE2_REG_3_ );
nor U94381 ( n28026, n28028, n28029 );
nand U94382 ( n35042, n35104, n76461 );
nor U94383 ( n35104, n35105, n35106 );
and U94384 ( n35106, n35047, P1_P3_STATE2_REG_3_ );
nor U94385 ( n35105, n35107, n35108 );
nand U94386 ( n69780, n69840, n76193 );
nor U94387 ( n69840, n69841, n69842 );
and U94388 ( n69842, n69785, P2_P3_STATE2_REG_3_ );
nor U94389 ( n69841, n69843, n69844 );
nand U94390 ( n61114, n61184, n76259 );
nor U94391 ( n61184, n61185, n61186 );
and U94392 ( n61186, n61119, P2_P2_STATE2_REG_3_ );
nor U94393 ( n61185, n61187, n61188 );
nor U94394 ( n35107, n35109, n34369 );
nor U94395 ( n35109, n35041, n3429 );
not U94396 ( n3429, n35046 );
nor U94397 ( n69843, n69845, n69121 );
nor U94398 ( n69845, n69779, n6044 );
not U94399 ( n6044, n69784 );
nand U94400 ( n35200, n35262, n76461 );
nor U94401 ( n35262, n35263, n35264 );
and U94402 ( n35264, n35205, P1_P3_STATE2_REG_3_ );
nor U94403 ( n35263, n35265, n35266 );
nand U94404 ( n69936, n69996, n76193 );
nor U94405 ( n69996, n69997, n69998 );
and U94406 ( n69998, n69941, P2_P3_STATE2_REG_3_ );
nor U94407 ( n69997, n69999, n70000 );
nor U94408 ( n35265, n35267, n34369 );
nor U94409 ( n35267, n35199, n3428 );
not U94410 ( n3428, n35204 );
nor U94411 ( n69999, n70001, n69121 );
nor U94412 ( n70001, n69935, n6043 );
not U94413 ( n6043, n69940 );
nand U94414 ( n28123, n28187, n76517 );
nor U94415 ( n28187, n28188, n28189 );
and U94416 ( n28189, n28128, P1_P2_STATE2_REG_3_ );
nor U94417 ( n28188, n28190, n28191 );
nand U94418 ( n61278, n61351, n76259 );
nor U94419 ( n61351, n61352, n61353 );
and U94420 ( n61353, n61283, P2_P2_STATE2_REG_3_ );
nor U94421 ( n61352, n61354, n61355 );
nor U94422 ( n28190, n28192, n27124 );
nor U94423 ( n28192, n28122, n4262 );
not U94424 ( n4262, n28127 );
nor U94425 ( n61354, n61356, n60268 );
nor U94426 ( n61356, n61277, n6894 );
not U94427 ( n6894, n61282 );
nand U94428 ( n35358, n35420, n76461 );
nor U94429 ( n35420, n35421, n35422 );
and U94430 ( n35422, n35363, P1_P3_STATE2_REG_3_ );
nor U94431 ( n35421, n35423, n35424 );
nand U94432 ( n70090, n70150, n76193 );
nor U94433 ( n70150, n70151, n70152 );
and U94434 ( n70152, n70095, P2_P3_STATE2_REG_3_ );
nor U94435 ( n70151, n70153, n70154 );
nor U94436 ( n35423, n35425, n34369 );
nor U94437 ( n35425, n35357, n3424 );
not U94438 ( n3424, n35362 );
nor U94439 ( n70153, n70155, n69121 );
nor U94440 ( n70155, n70089, n6039 );
not U94441 ( n6039, n70094 );
not U94442 ( n862, n45226 );
nand U94443 ( n49085, n49164, n76325 );
nor U94444 ( n49164, n49165, n49166 );
and U94445 ( n49166, n49086, n76177 );
nor U94446 ( n49165, n49167, n49163 );
nor U94447 ( n49158, n49172, n47934 );
nand U94448 ( n49172, n48240, n7855 );
nor U94449 ( n49167, n49169, n48133 );
and U94450 ( n49169, n49089, n7834 );
nand U94451 ( n42404, n54193, n54194 );
nor U94452 ( n54194, n7629, n54195 );
nor U94453 ( n54193, n7504, n47887 );
nor U94454 ( n54195, n7789, n45509 );
buf U94455 ( n76750, n4687 );
and U94456 ( n48248, n48321, n48142 );
nor U94457 ( n48321, n47921, n48240 );
nor U94458 ( n48313, n48316, n48133 );
nor U94459 ( n48316, n7843, n48248 );
not U94460 ( n7843, n48252 );
nand U94461 ( n67749, n67714, n76058 );
nand U94462 ( n46702, n46667, n76101 );
nand U94463 ( n25744, n25709, n76156 );
nand U94464 ( n58884, n58849, n76084 );
nand U94465 ( n32993, n32960, n76128 );
not U94466 ( U39, n70997 );
nand U94467 ( n48624, n48703, n76325 );
nor U94468 ( n48703, n48704, n48705 );
and U94469 ( n48705, n48625, n76181 );
nor U94470 ( n48704, n48706, n48702 );
nand U94471 ( n48629, n48321, n48523 );
nor U94472 ( n48706, n48708, n48133 );
and U94473 ( n48708, n48628, n48629 );
and U94474 ( n48025, n48141, n48142 );
nor U94475 ( n48128, n48132, n48133 );
nor U94476 ( n48132, n48025, n7845 );
not U94477 ( n7845, n48030 );
and U94478 ( n48427, n48141, n48523 );
nand U94479 ( n48426, n48511, n76325 );
nor U94480 ( n48511, n48512, n48513 );
and U94481 ( n48513, n48429, n76181 );
nor U94482 ( n48512, n48516, n48517 );
nor U94483 ( n48516, n48519, n48133 );
nor U94484 ( n48519, n48427, n7840 );
not U94485 ( n7840, n48432 );
not U94486 ( n5634, n63481 );
not U94487 ( n3033, n29582 );
not U94488 ( n3877, n22261 );
not U94489 ( n6509, n55373 );
nand U94490 ( n15178, n15265, n76591 );
nor U94491 ( n15265, n15267, n15268 );
and U94492 ( n15268, n15185, n76189 );
nor U94493 ( n15267, n15269, n15264 );
nor U94494 ( n15269, n15274, n14947 );
nor U94495 ( n15274, n5187, n15179 );
not U94496 ( n5187, n15184 );
and U94497 ( n28289, n76517, P1_P2_STATE2_REG_3_ );
and U94498 ( n61511, n76259, P2_P2_STATE2_REG_3_ );
nor U94499 ( n57437, n249, n57007 );
nor U94500 ( n24314, n4, n23883 );
or U94501 ( n23822, n23152, n4 );
or U94502 ( n56947, n56273, n249 );
and U94503 ( n35517, n76461, P1_P3_STATE2_REG_3_ );
and U94504 ( n70245, n76193, P2_P3_STATE2_REG_3_ );
nand U94505 ( n34058, n76774, n32571 );
nand U94506 ( n26813, n76754, n25329 );
nand U94507 ( n59953, n76687, n58468 );
nand U94508 ( n47792, n76660, n46275 );
nand U94509 ( n68812, n76708, n67336 );
nor U94510 ( n57372, n292, n57007 );
nor U94511 ( n57383, n287, n57007 );
nor U94512 ( n57393, n280, n57007 );
nor U94513 ( n57404, n274, n57007 );
nor U94514 ( n57413, n268, n57007 );
nor U94515 ( n57424, n262, n57007 );
nor U94516 ( n24247, n38, n23883 );
nor U94517 ( n24258, n34, n23883 );
nor U94518 ( n24268, n29, n23883 );
nor U94519 ( n24281, n24, n23883 );
nor U94520 ( n24290, n19, n23883 );
nor U94521 ( n24301, n14, n23883 );
nand U94522 ( n68605, n68680, n68519 );
nand U94523 ( n68680, n6090, n67502 );
nand U94524 ( n33849, n33924, n33763 );
nand U94525 ( n33924, n3475, n32737 );
nand U94526 ( n26604, n26679, n26518 );
nand U94527 ( n26679, n4313, n25497 );
nand U94528 ( n59746, n59821, n59657 );
nand U94529 ( n59821, n6945, n58634 );
nand U94530 ( n47584, n47659, n47498 );
nand U94531 ( n47659, n7879, n46438 );
nand U94532 ( n68765, n76708, n67330 );
nand U94533 ( n34009, n76774, n32565 );
nand U94534 ( n26766, n76754, n25323 );
nand U94535 ( n59906, n76687, n58462 );
nand U94536 ( n47744, n76660, n46269 );
nand U94537 ( n48530, n48609, n76325 );
nor U94538 ( n48609, n48610, n48611 );
and U94539 ( n48611, n48531, n76182 );
nor U94540 ( n48610, n48612, n48608 );
nor U94541 ( n48612, n48614, n48133 );
and U94542 ( n48614, n48534, n48535 );
and U94543 ( n15072, n15169, n14958 );
nor U94544 ( n15169, n14692, n14734 );
nor U94545 ( n15159, n15163, n14947 );
nor U94546 ( n15163, n5188, n15072 );
not U94547 ( n5188, n15077 );
nand U94548 ( n15518, n15169, n15397 );
nand U94549 ( n15512, n15590, n76591 );
nor U94550 ( n15590, n15592, n15593 );
and U94551 ( n15593, n15513, n76191 );
nor U94552 ( n15592, n15594, n15589 );
nor U94553 ( n15594, n15597, n14947 );
and U94554 ( n15597, n15517, n15518 );
nor U94555 ( n48231, n48234, n48133 );
nor U94556 ( n48234, n7844, n48150 );
not U94557 ( n7844, n48154 );
nand U94558 ( n48149, n48228, n76325 );
nor U94559 ( n48228, n48229, n48230 );
and U94560 ( n48230, n48155, n76177 );
nor U94561 ( n48229, n48231, n48226 );
and U94562 ( n14822, n14957, n14958 );
nor U94563 ( n14942, n14945, n14947 );
nor U94564 ( n14945, n14822, n5190 );
not U94565 ( n5190, n14828 );
nand U94566 ( n15288, n15380, n76591 );
nor U94567 ( n15380, n15382, n15383 );
and U94568 ( n15383, n15292, n76191 );
nor U94569 ( n15382, n15387, n15388 );
and U94570 ( n15289, n14957, n15397 );
nor U94571 ( n15387, n15392, n14947 );
nor U94572 ( n15392, n15289, n5185 );
not U94573 ( n5185, n15295 );
nor U94574 ( n60103, n6513, n6515 );
nor U94575 ( n26963, n3880, n3883 );
nor U94576 ( n34208, n3037, n3039 );
nor U94577 ( n68962, n5638, n5640 );
nor U94578 ( n14213, n4937, n14214 );
and U94579 ( n12574, n14210, n14212 );
nand U94580 ( n14210, n4926, n14143 );
nand U94581 ( n14212, n14213, n14177 );
not U94582 ( n4926, n14177 );
nor U94583 ( n68559, n5803, n68560 );
nor U94584 ( n47538, n7590, n47539 );
nor U94585 ( n26558, n4037, n26559 );
nor U94586 ( n59700, n6669, n59701 );
and U94587 ( n67167, n68557, n68558 );
nand U94588 ( n68557, n5792, n68503 );
nand U94589 ( n68558, n68559, n68530 );
not U94590 ( n5792, n68530 );
and U94591 ( n46203, n47536, n47537 );
nand U94592 ( n47536, n7579, n47482 );
nand U94593 ( n47537, n47538, n47509 );
not U94594 ( n7579, n47509 );
and U94595 ( n25269, n26556, n26557 );
nand U94596 ( n26556, n4028, n26502 );
nand U94597 ( n26557, n26558, n26529 );
not U94598 ( n4028, n26529 );
and U94599 ( n58405, n59698, n59699 );
nand U94600 ( n59698, n6660, n59641 );
nand U94601 ( n59699, n59700, n59671 );
not U94602 ( n6660, n59671 );
nor U94603 ( n33803, n3204, n33804 );
and U94604 ( n32511, n33801, n33802 );
nand U94605 ( n33801, n3193, n33747 );
nand U94606 ( n33802, n33803, n33774 );
not U94607 ( n3193, n33774 );
nor U94608 ( n15497, n15499, n14947 );
and U94609 ( n15499, n15410, n15412 );
nand U94610 ( n15405, n15493, n76591 );
nor U94611 ( n15493, n15494, n15495 );
and U94612 ( n15495, n15407, n76192 );
nor U94613 ( n15494, n15497, n15492 );
not U94614 ( n7859, n47921 );
nor U94615 ( n47948, n47934, n7855 );
not U94616 ( n7860, n47916 );
nand U94617 ( n14479, n76727, n12642 );
nand U94618 ( n14539, n76727, n12658 );
nor U94619 ( n67419, n67456, n67468 );
and U94620 ( n67468, n67457, n67458 );
nor U94621 ( n32654, n32691, n32703 );
and U94622 ( n32703, n32692, n32693 );
nor U94623 ( n25414, n25451, n25463 );
and U94624 ( n25463, n25452, n25453 );
nor U94625 ( n58551, n58588, n58600 );
and U94626 ( n58600, n58589, n58590 );
nor U94627 ( n34894, n34215, n34296 );
nor U94628 ( n34928, n34215, n34340 );
nor U94629 ( n34936, n34215, n34351 );
nor U94630 ( n34952, n34215, n34372 );
nor U94631 ( n34912, n34215, n34318 );
nor U94632 ( n34920, n34215, n34329 );
nor U94633 ( n34902, n34215, n34307 );
nor U94634 ( n69636, n68969, n69048 );
nor U94635 ( n69644, n68969, n69059 );
nor U94636 ( n69652, n68969, n69070 );
nor U94637 ( n69676, n68969, n69103 );
nor U94638 ( n69692, n68969, n69124 );
nor U94639 ( n69668, n68969, n69092 );
nor U94640 ( n69660, n68969, n69081 );
nand U94641 ( n14967, n15047, n76591 );
nor U94642 ( n15047, n15048, n15049 );
and U94643 ( n15049, n14974, n76187 );
nor U94644 ( n15048, n15050, n15044 );
nor U94645 ( n15050, n15054, n14947 );
nor U94646 ( n15054, n5189, n14968 );
not U94647 ( n5189, n14973 );
nor U94648 ( n27349, n27085, n27314 );
nor U94649 ( n27183, n27085, n27150 );
nor U94650 ( n60497, n60226, n60457 );
nor U94651 ( n60325, n60226, n60292 );
nor U94652 ( n27323, n27052, n27314 );
nor U94653 ( n27159, n27052, n27150 );
nor U94654 ( n27381, n27128, n27314 );
nor U94655 ( n27216, n27128, n27150 );
nor U94656 ( n27357, n27096, n27314 );
nor U94657 ( n27191, n27096, n27150 );
nor U94658 ( n60505, n60240, n60457 );
nor U94659 ( n60333, n60240, n60292 );
nor U94660 ( n60469, n60193, n60457 );
nor U94661 ( n60301, n60193, n60292 );
nor U94662 ( n60529, n60272, n60457 );
nor U94663 ( n60361, n60272, n60292 );
nor U94664 ( n27339, n27074, n27314 );
nor U94665 ( n27175, n27074, n27150 );
nor U94666 ( n27331, n27063, n27314 );
nor U94667 ( n27167, n27063, n27150 );
nor U94668 ( n60489, n60215, n60457 );
nor U94669 ( n60317, n60215, n60292 );
nor U94670 ( n60477, n60204, n60457 );
nor U94671 ( n60309, n60204, n60292 );
nor U94672 ( n35312, n34329, n35279 );
nor U94673 ( n34669, n34329, n34638 );
nor U94674 ( n70044, n69081, n70013 );
nor U94675 ( n35286, n34296, n35279 );
nor U94676 ( n34645, n34296, n34638 );
nor U94677 ( n35320, n34340, n35279 );
nor U94678 ( n34677, n34340, n34638 );
nor U94679 ( n35328, n34351, n35279 );
nor U94680 ( n34685, n34351, n34638 );
nor U94681 ( n34695, n34372, n34638 );
nor U94682 ( n35336, n34372, n35279 );
nor U94683 ( n70020, n69048, n70013 );
nor U94684 ( n69391, n69048, n69384 );
nor U94685 ( n70060, n69103, n70013 );
nor U94686 ( n69431, n69103, n69384 );
nor U94687 ( n69439, n69124, n69384 );
nor U94688 ( n70068, n69124, n70013 );
nor U94689 ( n70052, n69092, n70013 );
nor U94690 ( n69423, n69092, n69384 );
nor U94691 ( n34661, n34318, n34638 );
nor U94692 ( n35304, n34318, n35279 );
nor U94693 ( n34653, n34307, n34638 );
nor U94694 ( n35294, n34307, n35279 );
nor U94695 ( n70028, n69059, n70013 );
nor U94696 ( n69399, n69059, n69384 );
nor U94697 ( n69407, n69070, n69384 );
nor U94698 ( n70036, n69070, n70013 );
nor U94699 ( n69415, n69081, n69384 );
nor U94700 ( n28240, n27085, n28209 );
nor U94701 ( n28001, n27085, n27970 );
nor U94702 ( n27919, n27085, n27888 );
nor U94703 ( n27837, n27085, n27806 );
nor U94704 ( n27598, n27085, n27567 );
nor U94705 ( n27516, n27085, n27481 );
nor U94706 ( n61466, n60226, n61373 );
nor U94707 ( n61150, n60226, n61119 );
nor U94708 ( n61066, n60226, n61035 );
nor U94709 ( n60988, n60226, n60954 );
nor U94710 ( n60748, n60226, n60717 );
nor U94711 ( n60665, n60226, n60630 );
nor U94712 ( n27977, n27052, n27970 );
nor U94713 ( n27895, n27052, n27888 );
nor U94714 ( n27813, n27052, n27806 );
nor U94715 ( n27574, n27052, n27567 );
nor U94716 ( n27489, n27052, n27481 );
nor U94717 ( n28275, n27128, n28209 );
nor U94718 ( n28032, n27128, n27970 );
nor U94719 ( n27950, n27128, n27888 );
nor U94720 ( n27872, n27128, n27806 );
nor U94721 ( n27629, n27128, n27567 );
nor U94722 ( n27550, n27128, n27481 );
nor U94723 ( n28009, n27096, n27970 );
nor U94724 ( n27927, n27096, n27888 );
nor U94725 ( n27845, n27096, n27806 );
nor U94726 ( n27606, n27096, n27567 );
nor U94727 ( n27525, n27096, n27481 );
nor U94728 ( n28248, n27096, n28209 );
nor U94729 ( n61474, n60240, n61373 );
nor U94730 ( n61158, n60240, n61119 );
nor U94731 ( n61080, n60240, n61035 );
nor U94732 ( n60996, n60240, n60954 );
nor U94733 ( n60756, n60240, n60717 );
nor U94734 ( n60677, n60240, n60630 );
nor U94735 ( n61380, n60193, n61373 );
nor U94736 ( n61126, n60193, n61119 );
nor U94737 ( n61042, n60193, n61035 );
nor U94738 ( n60961, n60193, n60954 );
nor U94739 ( n60724, n60193, n60717 );
nor U94740 ( n60638, n60193, n60630 );
nor U94741 ( n61191, n60272, n61119 );
nor U94742 ( n61103, n60272, n61035 );
nor U94743 ( n61019, n60272, n60954 );
nor U94744 ( n60782, n60272, n60717 );
nor U94745 ( n60702, n60272, n60630 );
nor U94746 ( n28216, n27052, n28209 );
nor U94747 ( n61497, n60272, n61373 );
nor U94748 ( n28232, n27074, n28209 );
nor U94749 ( n27993, n27074, n27970 );
nor U94750 ( n27911, n27074, n27888 );
nor U94751 ( n27829, n27074, n27806 );
nor U94752 ( n27590, n27074, n27567 );
nor U94753 ( n27507, n27074, n27481 );
nor U94754 ( n28224, n27063, n28209 );
nor U94755 ( n27985, n27063, n27970 );
nor U94756 ( n27903, n27063, n27888 );
nor U94757 ( n27821, n27063, n27806 );
nor U94758 ( n27582, n27063, n27567 );
nor U94759 ( n27498, n27063, n27481 );
nor U94760 ( n61142, n60215, n61119 );
nor U94761 ( n61058, n60215, n61035 );
nor U94762 ( n60980, n60215, n60954 );
nor U94763 ( n60740, n60215, n60717 );
nor U94764 ( n60656, n60215, n60630 );
nor U94765 ( n61388, n60204, n61373 );
nor U94766 ( n61134, n60204, n61119 );
nor U94767 ( n61050, n60204, n61035 );
nor U94768 ( n60969, n60204, n60954 );
nor U94769 ( n60732, n60204, n60717 );
nor U94770 ( n60647, n60204, n60630 );
nor U94771 ( n61458, n60215, n61373 );
nor U94772 ( n34592, n34329, n34559 );
nor U94773 ( n34428, n34329, n34393 );
nor U94774 ( n69340, n69081, n69307 );
nor U94775 ( n69178, n69081, n69145 );
nor U94776 ( n34568, n34296, n34559 );
nor U94777 ( n34404, n34296, n34393 );
nor U94778 ( n34602, n34340, n34559 );
nor U94779 ( n34436, n34340, n34393 );
nor U94780 ( n34610, n34351, n34559 );
nor U94781 ( n34444, n34351, n34393 );
nor U94782 ( n34626, n34372, n34559 );
nor U94783 ( n34461, n34372, n34393 );
nor U94784 ( n69316, n69048, n69307 );
nor U94785 ( n69154, n69048, n69145 );
nor U94786 ( n69356, n69103, n69307 );
nor U94787 ( n69194, n69103, n69145 );
nor U94788 ( n69372, n69124, n69307 );
nor U94789 ( n69211, n69124, n69145 );
nor U94790 ( n69348, n69092, n69307 );
nor U94791 ( n69186, n69092, n69145 );
nor U94792 ( n34584, n34318, n34559 );
nor U94793 ( n34420, n34318, n34393 );
nor U94794 ( n34576, n34307, n34559 );
nor U94795 ( n34412, n34307, n34393 );
nor U94796 ( n69324, n69059, n69307 );
nor U94797 ( n69162, n69059, n69145 );
nor U94798 ( n69332, n69070, n69307 );
nor U94799 ( n69170, n69070, n69145 );
nor U94800 ( n51666, n51668, n48133 );
and U94801 ( n51668, n49450, n49462 );
nor U94802 ( n35473, n34329, n35442 );
nor U94803 ( n35238, n34329, n35205 );
nor U94804 ( n35158, n34329, n35127 );
nor U94805 ( n35078, n34329, n35047 );
nor U94806 ( n34843, n34329, n34810 );
nor U94807 ( n34760, n34329, n34726 );
nor U94808 ( n70203, n69081, n70172 );
nor U94809 ( n69972, n69081, n69941 );
nor U94810 ( n69894, n69081, n69863 );
nor U94811 ( n69816, n69081, n69785 );
nor U94812 ( n69585, n69081, n69554 );
nor U94813 ( n69504, n69081, n69470 );
nor U94814 ( n35449, n34296, n35442 );
nor U94815 ( n35214, n34296, n35205 );
nor U94816 ( n35134, n34296, n35127 );
nor U94817 ( n35054, n34296, n35047 );
nor U94818 ( n34819, n34296, n34810 );
nor U94819 ( n34733, n34296, n34726 );
nor U94820 ( n35246, n34340, n35205 );
nor U94821 ( n35166, n34340, n35127 );
nor U94822 ( n35086, n34340, n35047 );
nor U94823 ( n34851, n34340, n34810 );
nor U94824 ( n34769, n34340, n34726 );
nor U94825 ( n35481, n34340, n35442 );
nor U94826 ( n35254, n34351, n35205 );
nor U94827 ( n35174, n34351, n35127 );
nor U94828 ( n35094, n34351, n35047 );
nor U94829 ( n34859, n34351, n34810 );
nor U94830 ( n34778, n34351, n34726 );
nor U94831 ( n35489, n34351, n35442 );
nor U94832 ( n35506, n34372, n35442 );
nor U94833 ( n35269, n34372, n35205 );
nor U94834 ( n35189, n34372, n35127 );
nor U94835 ( n35111, n34372, n35047 );
nor U94836 ( n34874, n34372, n34810 );
nor U94837 ( n34794, n34372, n34726 );
nor U94838 ( n70179, n69048, n70172 );
nor U94839 ( n69948, n69048, n69941 );
nor U94840 ( n69870, n69048, n69863 );
nor U94841 ( n69792, n69048, n69785 );
nor U94842 ( n69561, n69048, n69554 );
nor U94843 ( n69477, n69048, n69470 );
nor U94844 ( n69988, n69103, n69941 );
nor U94845 ( n69910, n69103, n69863 );
nor U94846 ( n69832, n69103, n69785 );
nor U94847 ( n69601, n69103, n69554 );
nor U94848 ( n69522, n69103, n69470 );
nor U94849 ( n70219, n69103, n70172 );
nor U94850 ( n70234, n69124, n70172 );
nor U94851 ( n70003, n69124, n69941 );
nor U94852 ( n69925, n69124, n69863 );
nor U94853 ( n69847, n69124, n69785 );
nor U94854 ( n69616, n69124, n69554 );
nor U94855 ( n69538, n69124, n69470 );
nor U94856 ( n69980, n69092, n69941 );
nor U94857 ( n69902, n69092, n69863 );
nor U94858 ( n69824, n69092, n69785 );
nor U94859 ( n69593, n69092, n69554 );
nor U94860 ( n69513, n69092, n69470 );
nor U94861 ( n70211, n69092, n70172 );
nor U94862 ( n35465, n34318, n35442 );
nor U94863 ( n35230, n34318, n35205 );
nor U94864 ( n35150, n34318, n35127 );
nor U94865 ( n35070, n34318, n35047 );
nor U94866 ( n34835, n34318, n34810 );
nor U94867 ( n34751, n34318, n34726 );
nor U94868 ( n35222, n34307, n35205 );
nor U94869 ( n35142, n34307, n35127 );
nor U94870 ( n35062, n34307, n35047 );
nor U94871 ( n34827, n34307, n34810 );
nor U94872 ( n34742, n34307, n34726 );
nor U94873 ( n69956, n69059, n69941 );
nor U94874 ( n69878, n69059, n69863 );
nor U94875 ( n69800, n69059, n69785 );
nor U94876 ( n69569, n69059, n69554 );
nor U94877 ( n69486, n69059, n69470 );
nor U94878 ( n70195, n69070, n70172 );
nor U94879 ( n69964, n69070, n69941 );
nor U94880 ( n69886, n69070, n69863 );
nor U94881 ( n69808, n69070, n69785 );
nor U94882 ( n69577, n69070, n69554 );
nor U94883 ( n69495, n69070, n69470 );
nor U94884 ( n70187, n69059, n70172 );
nor U94885 ( n35457, n34307, n35442 );
not U94886 ( n900, n42431 );
not U94887 ( n188, n34228 );
not U94888 ( n150, n26983 );
not U94889 ( n459, n68982 );
not U94890 ( n423, n60126 );
not U94891 ( n493, n47974 );
not U94892 ( n222, n14752 );
not U94893 ( n4865, n13314 );
not U94894 ( n76234, n76235 );
not U94895 ( n76233, n76235 );
nand U94896 ( n12993, n12732, n13098 );
nor U94897 ( n28283, n26968, n4268 );
nor U94898 ( n61505, n60108, n6900 );
nor U94899 ( n35587, n35590, n34369 );
nor U94900 ( n35590, n3420, n35514 );
not U94901 ( n3420, n35519 );
nor U94902 ( n28406, n28409, n27124 );
nor U94903 ( n28409, n4258, n28283 );
not U94904 ( n4258, n28291 );
nor U94905 ( n70315, n70318, n69121 );
nor U94906 ( n70318, n6035, n70242 );
not U94907 ( n6035, n70247 );
nor U94908 ( n61715, n61718, n60268 );
nor U94909 ( n61718, n6890, n61505 );
not U94910 ( n6890, n61513 );
and U94911 ( n35522, n35582, n76461 );
nor U94912 ( n35582, n35585, n35586 );
and U94913 ( n35586, n35516, P1_P3_STATE2_REG_3_ );
nor U94914 ( n35585, n35587, n35581 );
and U94915 ( n28296, n28401, n76517 );
nor U94916 ( n28401, n28404, n28405 );
and U94917 ( n28405, n28288, P1_P2_STATE2_REG_3_ );
nor U94918 ( n28404, n28406, n28398 );
and U94919 ( n70250, n70310, n76193 );
nor U94920 ( n70310, n70313, n70314 );
and U94921 ( n70314, n70244, P2_P3_STATE2_REG_3_ );
nor U94922 ( n70313, n70315, n70309 );
and U94923 ( n61518, n61710, n76259 );
nor U94924 ( n61710, n61713, n61714 );
and U94925 ( n61714, n61510, P2_P2_STATE2_REG_3_ );
nor U94926 ( n61713, n61715, n61679 );
not U94927 ( n6512, n60072 );
not U94928 ( n3879, n26932 );
not U94929 ( n3035, n34177 );
not U94930 ( n5637, n68931 );
not U94931 ( n76503, n76504 );
not U94932 ( n76502, n76504 );
not U94933 ( n7512, n46789 );
not U94934 ( n5725, n67836 );
not U94935 ( n3968, n25833 );
not U94936 ( n6600, n58971 );
not U94937 ( n76302, n76304 );
not U94938 ( n76303, n76304 );
not U94939 ( n3124, n33080 );
not U94940 ( n902, n42423 );
nor U94941 ( n34885, n34215, n34283 );
nor U94942 ( n69627, n68969, n69035 );
xor U94943 ( n47935, n48417, n7857 );
nand U94944 ( n13217, n13237, n12732 );
nor U94945 ( n27365, n27107, n27314 );
nor U94946 ( n27199, n27107, n27150 );
nor U94947 ( n27313, n27039, n27314 );
nor U94948 ( n27149, n27039, n27150 );
nor U94949 ( n60513, n60251, n60457 );
nor U94950 ( n60341, n60251, n60292 );
nor U94951 ( n60456, n60180, n60457 );
nor U94952 ( n60291, n60180, n60292 );
nor U94953 ( n35273, n34283, n35279 );
nor U94954 ( n34632, n34283, n34638 );
nor U94955 ( n70007, n69035, n70013 );
nor U94956 ( n69378, n69035, n69384 );
not U94957 ( n76561, n76563 );
not U94958 ( n76562, n76563 );
nor U94959 ( n28017, n27107, n27970 );
nor U94960 ( n27935, n27107, n27888 );
nor U94961 ( n27857, n27107, n27806 );
nor U94962 ( n27614, n27107, n27567 );
nor U94963 ( n28206, n27039, n28209 );
nor U94964 ( n27885, n27039, n27888 );
nor U94965 ( n27803, n27039, n27806 );
nor U94966 ( n27564, n27039, n27567 );
nor U94967 ( n27478, n27039, n27481 );
nor U94968 ( n61166, n60251, n61119 );
nor U94969 ( n61088, n60251, n61035 );
nor U94970 ( n61004, n60251, n60954 );
nor U94971 ( n60686, n60251, n60630 );
nor U94972 ( n61370, n60180, n61373 );
nor U94973 ( n61032, n60180, n61035 );
nor U94974 ( n28260, n27107, n28209 );
nand U94975 ( n46570, n46331, n46627 );
nor U94976 ( n27534, n27107, n27481 );
nor U94977 ( n27967, n27039, n27970 );
nor U94978 ( n61482, n60251, n61373 );
nor U94979 ( n60764, n60251, n60717 );
nor U94980 ( n61116, n60180, n61119 );
nor U94981 ( n60951, n60180, n60954 );
nor U94982 ( n60714, n60180, n60717 );
nor U94983 ( n60627, n60180, n60630 );
nand U94984 ( n32852, n32630, n32913 );
nor U94985 ( n34558, n34283, n34559 );
nor U94986 ( n34392, n34283, n34393 );
nor U94987 ( n69306, n69035, n69307 );
nor U94988 ( n69144, n69035, n69145 );
nand U94989 ( n67617, n67395, n67674 );
nand U94990 ( n25612, n25390, n25669 );
nand U94991 ( n58749, n58527, n58809 );
and U94992 ( n25296, n26623, n26624 );
nand U94993 ( n26623, n26629, n4039 );
nand U94994 ( n26624, n26625, n26626 );
not U94995 ( n4039, n26626 );
and U94996 ( n58432, n59765, n59766 );
nand U94997 ( n59765, n59771, n6672 );
nand U94998 ( n59766, n59767, n59768 );
not U94999 ( n6672, n59768 );
and U95000 ( n67194, n68624, n68625 );
nand U95001 ( n68624, n68630, n5805 );
nand U95002 ( n68625, n68626, n68627 );
not U95003 ( n5805, n68627 );
and U95004 ( n46242, n47603, n47604 );
nand U95005 ( n47603, n47609, n7593 );
nand U95006 ( n47604, n47605, n47606 );
not U95007 ( n7593, n47606 );
nand U95008 ( n27562, n27622, n76517 );
nor U95009 ( n27622, n27623, n27624 );
and U95010 ( n27624, n27567, P1_P2_STATE2_REG_3_ );
nor U95011 ( n27623, n27625, n27626 );
nand U95012 ( n34805, n34867, n76461 );
nor U95013 ( n34867, n34868, n34869 );
and U95014 ( n34869, n34810, P1_P3_STATE2_REG_3_ );
nor U95015 ( n34868, n34870, n34871 );
nand U95016 ( n69549, n69609, n76193 );
nor U95017 ( n69609, n69610, n69611 );
and U95018 ( n69611, n69554, P2_P3_STATE2_REG_3_ );
nor U95019 ( n69610, n69612, n69613 );
nand U95020 ( n60712, n60775, n76259 );
nor U95021 ( n60775, n60776, n60777 );
and U95022 ( n60777, n60717, P2_P2_STATE2_REG_3_ );
nor U95023 ( n60776, n60778, n60779 );
nand U95024 ( n34809, n34541, n34707 );
nand U95025 ( n69553, n69289, n69451 );
nor U95026 ( n27296, n26935, n26969 );
nor U95027 ( n34541, n34180, n34214 );
nor U95028 ( n60439, n60075, n60109 );
nor U95029 ( n69289, n68934, n68968 );
nor U95030 ( n27625, n27627, n27124 );
nor U95031 ( n27627, n27561, n4270 );
not U95032 ( n4270, n27566 );
nor U95033 ( n34870, n34872, n34369 );
nor U95034 ( n34872, n34804, n3433 );
not U95035 ( n3433, n34809 );
nor U95036 ( n69612, n69614, n69121 );
nor U95037 ( n69614, n69548, n6048 );
not U95038 ( n6048, n69553 );
nor U95039 ( n60778, n60780, n60268 );
nor U95040 ( n60780, n60711, n6903 );
not U95041 ( n6903, n60716 );
and U95042 ( n32538, n33868, n33869 );
nand U95043 ( n33868, n33874, n3207 );
nand U95044 ( n33869, n33870, n33871 );
not U95045 ( n3207, n33871 );
and U95046 ( n12608, n14294, n14295 );
nand U95047 ( n14294, n14302, n4939 );
nand U95048 ( n14295, n14297, n14298 );
not U95049 ( n4939, n14298 );
nand U95050 ( n33000, n33016, n32630 );
nand U95051 ( n46709, n46725, n46331 );
nand U95052 ( n67756, n67772, n67395 );
nand U95053 ( n25751, n25769, n25390 );
nand U95054 ( n58891, n58907, n58527 );
not U95055 ( n7857, n51671 );
nor U95056 ( n27546, n27548, n27124 );
nor U95057 ( n27548, n27474, n4272 );
not U95058 ( n4272, n27480 );
nor U95059 ( n34790, n34792, n34369 );
nor U95060 ( n34792, n34719, n3434 );
not U95061 ( n3434, n34725 );
nor U95062 ( n69534, n69536, n69121 );
nor U95063 ( n69536, n69463, n6049 );
not U95064 ( n6049, n69469 );
nor U95065 ( n60698, n60700, n60268 );
nor U95066 ( n60700, n60623, n6904 );
not U95067 ( n6904, n60629 );
nand U95068 ( n27476, n27543, n76517 );
nor U95069 ( n27543, n27544, n27545 );
and U95070 ( n27545, n27481, P1_P2_STATE2_REG_3_ );
nor U95071 ( n27544, n27546, n27547 );
nand U95072 ( n34720, n34787, n76461 );
nor U95073 ( n34787, n34788, n34789 );
and U95074 ( n34789, n34726, P1_P3_STATE2_REG_3_ );
nor U95075 ( n34788, n34790, n34791 );
nand U95076 ( n69464, n69531, n76193 );
nor U95077 ( n69531, n69532, n69533 );
and U95078 ( n69533, n69470, P2_P3_STATE2_REG_3_ );
nor U95079 ( n69532, n69534, n69535 );
nand U95080 ( n60625, n60695, n76259 );
nor U95081 ( n60695, n60696, n60697 );
and U95082 ( n60697, n60630, P2_P2_STATE2_REG_3_ );
nor U95083 ( n60696, n60698, n60699 );
nor U95084 ( n60099, n60065, n60110 );
nor U95085 ( n26959, n26925, n26970 );
nor U95086 ( n34204, n34170, n34215 );
nor U95087 ( n68958, n68924, n68969 );
and U95088 ( n67184, n68635, n68636 );
nand U95089 ( n68636, n5817, n68637 );
nand U95090 ( n68635, n5803, n5804 );
nand U95091 ( n68637, n5804, n68638 );
and U95092 ( n25286, n26634, n26635 );
nand U95093 ( n26635, n4048, n26636 );
nand U95094 ( n26634, n4037, n4038 );
nand U95095 ( n26636, n4038, n26637 );
and U95096 ( n58422, n59776, n59777 );
nand U95097 ( n59777, n6680, n59778 );
nand U95098 ( n59776, n6669, n6670 );
nand U95099 ( n59778, n6670, n59779 );
and U95100 ( n46232, n47614, n47615 );
nand U95101 ( n47615, n7604, n47616 );
nand U95102 ( n47614, n7590, n7592 );
nand U95103 ( n47616, n7592, n47617 );
and U95104 ( n12595, n14308, n14309 );
nand U95105 ( n14309, n4950, n14310 );
nand U95106 ( n14308, n4937, n4938 );
nand U95107 ( n14310, n4938, n14312 );
and U95108 ( n32528, n33879, n33880 );
nand U95109 ( n33880, n3218, n33881 );
nand U95110 ( n33879, n3204, n3205 );
nand U95111 ( n33881, n3205, n33882 );
nand U95112 ( n47995, n7414, n47996 );
nand U95113 ( n34249, n3038, n34250 );
nand U95114 ( n27004, n3882, n27005 );
nand U95115 ( n69003, n5639, n69004 );
nand U95116 ( n60147, n6514, n60148 );
nand U95117 ( n26994, n3882, n26995 );
nand U95118 ( n60137, n6514, n60138 );
nand U95119 ( n47985, n7414, n47986 );
nand U95120 ( n34239, n3038, n34240 );
nand U95121 ( n68993, n5639, n68994 );
and U95122 ( n21627, n21629, n76628 );
nand U95123 ( n14765, n4770, n14767 );
not U95124 ( n76610, n76612 );
nand U95125 ( n27309, n27372, n76517 );
nor U95126 ( n27372, n27373, n27374 );
and U95127 ( n27374, n27314, P1_P2_STATE2_REG_3_ );
nor U95128 ( n27373, n27375, n27376 );
nand U95129 ( n60452, n60520, n76259 );
nor U95130 ( n60520, n60521, n60522 );
and U95131 ( n60522, n60457, P2_P2_STATE2_REG_3_ );
nor U95132 ( n60521, n60523, n60524 );
nand U95133 ( n34554, n34617, n76461 );
nor U95134 ( n34617, n34618, n34619 );
and U95135 ( n34619, n34559, P1_P3_STATE2_REG_3_ );
nor U95136 ( n34618, n34620, n34621 );
nand U95137 ( n69302, n69363, n76193 );
nor U95138 ( n69363, n69364, n69365 );
and U95139 ( n69365, n69307, P2_P3_STATE2_REG_3_ );
nor U95140 ( n69364, n69366, n69367 );
nor U95141 ( n27375, n27377, n27124 );
nor U95142 ( n27377, n4277, n27310 );
not U95143 ( n4277, n27311 );
nor U95144 ( n34620, n34622, n34369 );
nor U95145 ( n34622, n3439, n34555 );
not U95146 ( n3439, n34556 );
nor U95147 ( n69366, n69368, n69121 );
nor U95148 ( n69368, n6054, n69303 );
not U95149 ( n6054, n69304 );
nor U95150 ( n60523, n60525, n60268 );
nor U95151 ( n60525, n6909, n60453 );
not U95152 ( n6909, n60454 );
nand U95153 ( n14784, n4770, n14785 );
nand U95154 ( n31725, n3077, n31818 );
nand U95155 ( n31818, n31819, n31820 );
nand U95156 ( n31819, n3137, n31823 );
or U95157 ( n31820, n31821, n31822 );
nor U95158 ( n54151, n7602, n7343 );
nor U95159 ( n21168, n4948, n4711 );
nand U95160 ( n48003, n7414, n48007 );
nand U95161 ( n34257, n3038, n34261 );
nand U95162 ( n27014, n3882, n27018 );
nand U95163 ( n69011, n5639, n69015 );
nand U95164 ( n60155, n6514, n60159 );
nand U95165 ( n14794, n4770, n14799 );
and U95166 ( n27228, n27296, n27127 );
and U95167 ( n34473, n34541, n34371 );
and U95168 ( n60373, n60439, n60271 );
and U95169 ( n69223, n69289, n69123 );
nor U95170 ( n27293, n27295, n27124 );
nor U95171 ( n27295, n4278, n27228 );
not U95172 ( n4278, n27229 );
nor U95173 ( n34538, n34540, n34369 );
nor U95174 ( n34540, n3440, n34473 );
not U95175 ( n3440, n34474 );
nor U95176 ( n69286, n69288, n69121 );
nor U95177 ( n69288, n6055, n69223 );
not U95178 ( n6055, n69224 );
nor U95179 ( n60436, n60438, n60268 );
nor U95180 ( n60438, n6910, n60373 );
not U95181 ( n6910, n60374 );
nor U95182 ( n35653, n3215, n2978 );
nor U95183 ( n28474, n4045, n3822 );
nor U95184 ( n70379, n5814, n5579 );
nor U95185 ( n61779, n6678, n6454 );
buf U95186 ( n76518, n26979 );
buf U95187 ( n76260, n60119 );
nor U95188 ( n34365, n34368, n34369 );
nor U95189 ( n34368, n34281, n3443 );
not U95190 ( n3443, n34288 );
nor U95191 ( n69117, n69120, n69121 );
nor U95192 ( n69120, n69033, n6058 );
not U95193 ( n6058, n69040 );
and U95194 ( n34281, n34370, n34371 );
and U95195 ( n69033, n69122, n69123 );
nor U95196 ( n27041, n27042, n27043 );
nor U95197 ( n60182, n60183, n60184 );
nand U95198 ( n34636, n34699, n76461 );
nor U95199 ( n34699, n34700, n34701 );
and U95200 ( n34701, n34638, P1_P3_STATE2_REG_3_ );
nor U95201 ( n34700, n34702, n34703 );
nand U95202 ( n27391, n27454, n76517 );
nor U95203 ( n27454, n27455, n27456 );
and U95204 ( n27456, n27393, P1_P2_STATE2_REG_3_ );
nor U95205 ( n27455, n27457, n27458 );
nand U95206 ( n69382, n69443, n76193 );
nor U95207 ( n69443, n69444, n69445 );
and U95208 ( n69445, n69384, P2_P3_STATE2_REG_3_ );
nor U95209 ( n69444, n69446, n69447 );
nand U95210 ( n60539, n60603, n76259 );
nor U95211 ( n60603, n60604, n60605 );
and U95212 ( n60605, n60541, P2_P2_STATE2_REG_3_ );
nor U95213 ( n60604, n60606, n60607 );
and U95214 ( n34637, n34370, n34707 );
and U95215 ( n27392, n27126, n27462 );
and U95216 ( n69383, n69122, n69451 );
and U95217 ( n60540, n60270, n60611 );
and U95218 ( n27036, n27126, n27127 );
and U95219 ( n60177, n60270, n60271 );
nor U95220 ( n27120, n27123, n27124 );
nor U95221 ( n27123, n27036, n4280 );
not U95222 ( n4280, n27044 );
nor U95223 ( n34702, n34706, n34369 );
nor U95224 ( n34706, n34637, n3438 );
not U95225 ( n3438, n34642 );
nor U95226 ( n27457, n27461, n27124 );
nor U95227 ( n27461, n27392, n4275 );
not U95228 ( n4275, n27397 );
nor U95229 ( n69446, n69450, n69121 );
nor U95230 ( n69450, n69383, n6053 );
not U95231 ( n6053, n69388 );
nor U95232 ( n60606, n60610, n60268 );
nor U95233 ( n60610, n60540, n6908 );
not U95234 ( n6908, n60545 );
nor U95235 ( n60264, n60267, n60268 );
nor U95236 ( n60267, n60177, n6913 );
not U95237 ( n6913, n60185 );
nor U95238 ( n15679, n14734, n14733 );
nor U95239 ( n15697, n15699, n14947 );
nor U95240 ( n15699, n5184, n15679 );
nor U95241 ( n27395, n27043, n27396 );
nor U95242 ( n60543, n60184, n60544 );
nor U95243 ( n28043, n27043, n28046 );
nor U95244 ( n27718, n27043, n27721 );
nor U95245 ( n61202, n60184, n61205 );
nor U95246 ( n60869, n60184, n60872 );
nand U95247 ( n47171, n47266, n47311 );
nand U95248 ( n69140, n69201, n76193 );
nor U95249 ( n69201, n69202, n69203 );
and U95250 ( n69203, n69145, P2_P3_STATE2_REG_3_ );
nor U95251 ( n69202, n69204, n69205 );
nor U95252 ( n34454, n34456, n34369 );
nor U95253 ( n34456, n3442, n34389 );
not U95254 ( n3442, n34390 );
nor U95255 ( n69204, n69206, n69121 );
nor U95256 ( n69206, n6057, n69141 );
not U95257 ( n6057, n69142 );
nand U95258 ( n34388, n34451, n76461 );
nor U95259 ( n34451, n34452, n34453 );
and U95260 ( n34453, n34393, P1_P3_STATE2_REG_3_ );
nor U95261 ( n34452, n34454, n34455 );
nor U95262 ( n27209, n27211, n27124 );
nor U95263 ( n27211, n4279, n27146 );
not U95264 ( n4279, n27147 );
nor U95265 ( n60354, n60356, n60268 );
nor U95266 ( n60356, n6912, n60288 );
not U95267 ( n6912, n60289 );
nand U95268 ( n27145, n27206, n76517 );
nor U95269 ( n27206, n27207, n27208 );
and U95270 ( n27208, n27150, P1_P2_STATE2_REG_3_ );
nor U95271 ( n27207, n27209, n27210 );
nand U95272 ( n60287, n60351, n76259 );
nor U95273 ( n60351, n60352, n60353 );
and U95274 ( n60353, n60292, P2_P2_STATE2_REG_3_ );
nor U95275 ( n60352, n60354, n60355 );
nor U95276 ( n27132, n27042, n27133 );
nor U95277 ( n27109, n27042, n27110 );
nor U95278 ( n27098, n27042, n27099 );
nor U95279 ( n60242, n60183, n60243 );
nor U95280 ( n60253, n60183, n60254 );
nor U95281 ( n60276, n60183, n60277 );
not U95282 ( n4950, n14285 );
not U95283 ( n5817, n68617 );
not U95284 ( n4048, n26616 );
not U95285 ( n6680, n59758 );
not U95286 ( n7604, n47596 );
not U95287 ( n3218, n33861 );
nor U95288 ( n27466, n27133, n27396 );
nor U95289 ( n27437, n27099, n27396 );
nor U95290 ( n27447, n27110, n27396 );
nor U95291 ( n60588, n60243, n60544 );
nor U95292 ( n60596, n60254, n60544 );
nor U95293 ( n60615, n60277, n60544 );
buf U95294 ( n76462, n34224 );
buf U95295 ( n76194, n68978 );
nor U95296 ( n28113, n27133, n28046 );
nor U95297 ( n27790, n27133, n27721 );
nor U95298 ( n28097, n27110, n28046 );
nor U95299 ( n27774, n27110, n27721 );
nor U95300 ( n28089, n27099, n28046 );
nor U95301 ( n27766, n27099, n27721 );
nor U95302 ( n61244, n60243, n61205 );
nor U95303 ( n60914, n60243, n60872 );
nor U95304 ( n61252, n60254, n61205 );
nor U95305 ( n60922, n60254, n60872 );
nor U95306 ( n61268, n60277, n61205 );
nor U95307 ( n60938, n60277, n60872 );
not U95308 ( n5207, n21114 );
nor U95309 ( n27054, n27042, n27055 );
nor U95310 ( n27076, n27042, n27077 );
nor U95311 ( n27087, n27042, n27088 );
nor U95312 ( n27065, n27042, n27066 );
nor U95313 ( n60217, n60183, n60218 );
nor U95314 ( n60195, n60183, n60196 );
nor U95315 ( n60206, n60183, n60207 );
nor U95316 ( n60228, n60183, n60229 );
nand U95317 ( n67452, n67552, n67553 );
nand U95318 ( n67552, n67413, n67554 );
nand U95319 ( n67553, n64573, n67554 );
nand U95320 ( n32687, n32787, n32788 );
nand U95321 ( n32787, n32648, n32789 );
nand U95322 ( n32788, n30414, n32789 );
nand U95323 ( n46388, n46489, n46490 );
nand U95324 ( n46489, n46349, n46491 );
nand U95325 ( n46490, n43731, n46491 );
nand U95326 ( n25447, n25547, n25548 );
nand U95327 ( n25547, n25408, n25549 );
nand U95328 ( n25548, n23083, n25549 );
nand U95329 ( n58584, n58684, n58685 );
nand U95330 ( n58684, n58545, n58686 );
nand U95331 ( n58685, n56204, n58686 );
not U95332 ( n5202, n18715 );
nor U95333 ( n27405, n27055, n27396 );
nor U95334 ( n27421, n27077, n27396 );
nor U95335 ( n27429, n27088, n27396 );
nor U95336 ( n27413, n27066, n27396 );
nor U95337 ( n60572, n60218, n60544 );
nor U95338 ( n60561, n60207, n60544 );
nor U95339 ( n60580, n60229, n60544 );
nor U95340 ( n60553, n60196, n60544 );
nor U95341 ( n28053, n27055, n28046 );
nor U95342 ( n27728, n27055, n27721 );
nor U95343 ( n28073, n27077, n28046 );
nor U95344 ( n27744, n27077, n27721 );
nor U95345 ( n28081, n27088, n28046 );
nor U95346 ( n27758, n27088, n27721 );
nor U95347 ( n28065, n27066, n28046 );
nor U95348 ( n27736, n27066, n27721 );
nor U95349 ( n61228, n60218, n61205 );
nor U95350 ( n60898, n60218, n60872 );
nor U95351 ( n61212, n60196, n61205 );
nor U95352 ( n60882, n60196, n60872 );
nor U95353 ( n61220, n60207, n61205 );
nor U95354 ( n60890, n60207, n60872 );
nor U95355 ( n61236, n60229, n61205 );
nor U95356 ( n60906, n60229, n60872 );
and U95357 ( n12770, n12759, n12777 );
not U95358 ( n76143, n31624 );
not U95359 ( n76142, n31624 );
not U95360 ( n76144, n31624 );
not U95361 ( n8089, n43471 );
not U95362 ( n8090, n43490 );
not U95363 ( n8092, n43509 );
not U95364 ( n8093, n43528 );
not U95365 ( n8094, n43547 );
not U95366 ( n8095, n43579 );
not U95367 ( n3674, n30169 );
not U95368 ( n3675, n30188 );
not U95369 ( n3677, n30211 );
not U95370 ( n3678, n30230 );
not U95371 ( n3679, n30249 );
not U95372 ( n3680, n30268 );
not U95373 ( n3682, n30287 );
not U95374 ( n3683, n30310 );
not U95375 ( n6308, n64182 );
not U95376 ( n6309, n64254 );
not U95377 ( n6310, n64273 );
not U95378 ( n6312, n64292 );
not U95379 ( n6313, n64311 );
not U95380 ( n6314, n64330 );
not U95381 ( n6315, n64410 );
not U95382 ( n6317, n64429 );
not U95383 ( n3684, n30329 );
not U95384 ( n3685, n30347 );
not U95385 ( n3687, n30364 );
not U95386 ( n4568, n22844 );
not U95387 ( n4569, n22863 );
not U95388 ( n4570, n22884 );
not U95389 ( n4572, n22903 );
not U95390 ( n4573, n22922 );
not U95391 ( n4574, n22941 );
not U95392 ( n4575, n22960 );
not U95393 ( n4577, n22981 );
not U95394 ( n4578, n23000 );
not U95395 ( n4579, n23018 );
not U95396 ( n4580, n23035 );
not U95397 ( n6318, n64448 );
not U95398 ( n6319, n64466 );
not U95399 ( n6320, n64483 );
not U95400 ( n7200, n55961 );
not U95401 ( n7202, n55980 );
not U95402 ( n7203, n55999 );
not U95403 ( n7204, n56018 );
not U95404 ( n7205, n56037 );
not U95405 ( n7207, n56059 );
not U95406 ( n7208, n56078 );
not U95407 ( n7209, n56097 );
not U95408 ( n7210, n56116 );
not U95409 ( n7212, n56134 );
not U95410 ( n7213, n56154 );
not U95411 ( n8097, n43598 );
not U95412 ( n8098, n43617 );
not U95413 ( n8099, n43636 );
not U95414 ( n8100, n43654 );
not U95415 ( n8102, n43685 );
nand U95416 ( n46851, n46954, n46980 );
not U95417 ( n7869, n46491 );
not U95418 ( n7870, n46627 );
not U95419 ( n7872, n46725 );
and U95420 ( n46348, n46366, n7869 );
not U95421 ( n5434, n9514 );
not U95422 ( n5435, n9538 );
not U95423 ( n5437, n9562 );
not U95424 ( n5438, n9585 );
not U95425 ( n5439, n9608 );
not U95426 ( n5442, n9659 );
not U95427 ( n5443, n9683 );
not U95428 ( n5444, n9707 );
not U95429 ( n5445, n9729 );
not U95430 ( n5447, n9750 );
not U95431 ( n5440, n9632 );
nand U95432 ( n13392, n13507, n13539 );
not U95433 ( n5215, n12944 );
not U95434 ( n5218, n13237 );
not U95435 ( n5217, n13098 );
nand U95436 ( n13779, n13888, n13944 );
not U95437 ( n5224, n13880 );
not U95438 ( n5223, n13643 );
and U95439 ( n12817, n12942, n12943 );
nand U95440 ( n12942, n9812, n12944 );
nand U95441 ( n12943, n12777, n12944 );
not U95442 ( n7878, n47260 );
not U95443 ( n910, n42310 );
not U95444 ( n7877, n47068 );
nand U95445 ( n46352, n46366, n7869 );
nor U95446 ( n34950, n34214, n34213 );
nor U95447 ( n69690, n68968, n68967 );
nor U95448 ( n34947, n34949, n34369 );
nor U95449 ( n34949, n3437, n34950 );
nor U95450 ( n69687, n69689, n69121 );
nor U95451 ( n69689, n6052, n69690 );
nor U95452 ( n27702, n27704, n27124 );
nor U95453 ( n27704, n4274, n27705 );
nor U95454 ( n60853, n60855, n60268 );
nor U95455 ( n60855, n6907, n60856 );
nor U95456 ( n27705, n26969, n26968 );
nor U95457 ( n60856, n60109, n60108 );
nand U95458 ( n33451, n33542, n33587 );
nand U95459 ( n68202, n68298, n68343 );
nand U95460 ( n26201, n26297, n26342 );
nand U95461 ( n59340, n59436, n59481 );
nor U95462 ( n44531, n7793, n44507 );
nor U95463 ( n10742, n5138, n10712 );
nor U95464 ( n31152, n3390, n31128 );
nor U95465 ( n65406, n6005, n65382 );
nand U95466 ( n30746, n30802, n30803 );
nor U95467 ( n30803, n30804, n30805 );
nor U95468 ( n30802, n30826, n30827 );
nand U95469 ( n30805, n30806, n30807 );
nand U95470 ( n10232, n10298, n10299 );
nor U95471 ( n10299, n10300, n10302 );
nor U95472 ( n10298, n10328, n10329 );
nand U95473 ( n10302, n10303, n10304 );
nand U95474 ( n64952, n65004, n65005 );
nor U95475 ( n65005, n65006, n65007 );
nor U95476 ( n65004, n65028, n65029 );
nand U95477 ( n65007, n65008, n65009 );
nand U95478 ( n44109, n44162, n44163 );
nor U95479 ( n44163, n44164, n44165 );
nor U95480 ( n44162, n44186, n44187 );
nand U95481 ( n44165, n44166, n44167 );
xnor U95482 ( n30122, n30428, n30429 );
nor U95483 ( n30429, n30430, n30431 );
nand U95484 ( n30428, n30476, n30477 );
nand U95485 ( n30431, n30432, n30433 );
xnor U95486 ( n9455, n9828, n9829 );
nor U95487 ( n9829, n9830, n9832 );
nand U95488 ( n9828, n9888, n9889 );
nand U95489 ( n9832, n9833, n9834 );
xnor U95490 ( n64135, n64587, n64588 );
nor U95491 ( n64588, n64589, n64590 );
nand U95492 ( n64587, n64635, n64636 );
nand U95493 ( n64590, n64591, n64592 );
xnor U95494 ( n43391, n43744, n43745 );
nor U95495 ( n43745, n43746, n43747 );
nand U95496 ( n43744, n43792, n43793 );
nand U95497 ( n43747, n43748, n43749 );
nor U95498 ( n23860, n4228, n23836 );
nor U95499 ( n56984, n6860, n56960 );
nand U95500 ( n23436, n23495, n23496 );
nor U95501 ( n23496, n23497, n23498 );
nor U95502 ( n23495, n23519, n23520 );
nand U95503 ( n23498, n23499, n23500 );
nand U95504 ( n56558, n56617, n56618 );
nor U95505 ( n56618, n56619, n56620 );
nor U95506 ( n56617, n56641, n56642 );
nand U95507 ( n56620, n56621, n56622 );
xnor U95508 ( n22797, n23097, n23098 );
nor U95509 ( n23098, n23099, n23100 );
nand U95510 ( n23097, n23145, n23146 );
nand U95511 ( n23100, n23101, n23102 );
xnor U95512 ( n55911, n56218, n56219 );
nor U95513 ( n56219, n56220, n56221 );
nand U95514 ( n56218, n56266, n56267 );
nand U95515 ( n56221, n56222, n56223 );
nand U95516 ( n44193, n44531, n7812 );
nand U95517 ( n10337, n10742, n5157 );
nand U95518 ( n30833, n31152, n3409 );
nand U95519 ( n65035, n65406, n6024 );
nand U95520 ( n23526, n23860, n4247 );
nand U95521 ( n56648, n56984, n6879 );
nand U95522 ( n44196, n44531, n7807 );
nand U95523 ( n10340, n10742, n5152 );
nand U95524 ( n30836, n31152, n3404 );
nand U95525 ( n65038, n65406, n6019 );
nand U95526 ( n23529, n23860, n4242 );
nand U95527 ( n56651, n56984, n6874 );
xor U95528 ( n15062, n15278, n5202 );
not U95529 ( n912, n42301 );
not U95530 ( n489, n62885 );
not U95531 ( n218, n29163 );
not U95532 ( n455, n54941 );
not U95533 ( n184, n21850 );
not U95534 ( n514, n42376 );
not U95535 ( n243, n8287 );
nand U95536 ( n44202, n44538, n44507 );
nor U95537 ( n44538, n7793, n44509 );
nand U95538 ( n10348, n10750, n10712 );
nor U95539 ( n10750, n5138, n10714 );
nand U95540 ( n30842, n31159, n31128 );
nor U95541 ( n31159, n3390, n31130 );
nand U95542 ( n65044, n65413, n65382 );
nor U95543 ( n65413, n6005, n65384 );
nand U95544 ( n42352, n42310, n42308 );
nand U95545 ( n23535, n23867, n23836 );
nor U95546 ( n23867, n4228, n23838 );
nand U95547 ( n56657, n56991, n56960 );
nor U95548 ( n56991, n6860, n56962 );
nand U95549 ( n44207, n44543, n44507 );
nor U95550 ( n44543, n7793, n44517 );
nand U95551 ( n10354, n10757, n10712 );
nor U95552 ( n10757, n5138, n10724 );
nand U95553 ( n30847, n31164, n31128 );
nor U95554 ( n31164, n3390, n31138 );
nand U95555 ( n65049, n65418, n65382 );
nor U95556 ( n65418, n6005, n65392 );
nand U95557 ( n23540, n23872, n23836 );
nor U95558 ( n23872, n4228, n23846 );
nand U95559 ( n56662, n56996, n56960 );
nor U95560 ( n56996, n6860, n56970 );
not U95561 ( n5205, n14692 );
nand U95562 ( n33142, n33234, n33256 );
nand U95563 ( n67898, n67989, n68015 );
nand U95564 ( n25895, n25986, n26012 );
nand U95565 ( n59033, n59124, n59150 );
not U95566 ( n4302, n25549 );
not U95567 ( n6934, n58686 );
not U95568 ( n3464, n32789 );
not U95569 ( n6079, n67554 );
not U95570 ( n4304, n25769 );
not U95571 ( n6937, n58907 );
not U95572 ( n6082, n67772 );
not U95573 ( n3467, n33016 );
not U95574 ( n4303, n25669 );
not U95575 ( n6935, n58809 );
not U95576 ( n3465, n32913 );
not U95577 ( n6080, n67674 );
and U95578 ( n25407, n25425, n4302 );
and U95579 ( n58544, n58562, n6934 );
and U95580 ( n32647, n32665, n3464 );
and U95581 ( n67412, n67430, n6079 );
nor U95582 ( n49251, n51671, n7838 );
not U95583 ( n4643, n22075 );
not U95584 ( n7275, n55185 );
not U95585 ( n6383, n63157 );
not U95586 ( n3749, n29394 );
not U95587 ( n4288, n28412 );
not U95588 ( n6920, n61721 );
not U95589 ( n3450, n35593 );
not U95590 ( n6065, n70321 );
nand U95591 ( n32651, n32665, n3464 );
nand U95592 ( n25411, n25425, n4302 );
nand U95593 ( n67416, n67430, n6079 );
nand U95594 ( n58548, n58562, n6934 );
not U95595 ( n2979, n31619 );
not U95596 ( n6089, n68291 );
not U95597 ( n3474, n33535 );
not U95598 ( n4312, n26290 );
not U95599 ( n6944, n59429 );
not U95600 ( n6088, n68099 );
not U95601 ( n3473, n33342 );
not U95602 ( n4310, n26096 );
not U95603 ( n6943, n59237 );
not U95604 ( n8164, n42616 );
not U95605 ( n5510, n8558 );
xor U95606 ( n27213, n27379, n4288 );
xor U95607 ( n60358, n60527, n6920 );
nand U95608 ( n21945, n21946, n21947 );
nand U95609 ( n55057, n55058, n55059 );
xor U95610 ( n34458, n34624, n3450 );
xor U95611 ( n69208, n69370, n6065 );
nand U95612 ( n63029, n63030, n63031 );
nand U95613 ( n29262, n29263, n29264 );
nand U95614 ( n44180, n44522, n7810 );
nand U95615 ( n30820, n31143, n3408 );
nand U95616 ( n65022, n65397, n6023 );
nand U95617 ( n23513, n23851, n4245 );
nand U95618 ( n56635, n56975, n6878 );
nand U95619 ( n44181, n44522, n7812 );
nand U95620 ( n30821, n31143, n3409 );
nand U95621 ( n65023, n65397, n6024 );
nand U95622 ( n23514, n23851, n4247 );
nand U95623 ( n56636, n56975, n6879 );
nand U95624 ( n44184, n44522, n7807 );
nand U95625 ( n30824, n31143, n3404 );
nand U95626 ( n65026, n65397, n6019 );
nand U95627 ( n23517, n23851, n4242 );
nand U95628 ( n56639, n56975, n6874 );
nand U95629 ( n44185, n44522, n7808 );
nand U95630 ( n30825, n31143, n3405 );
nand U95631 ( n65027, n65397, n6020 );
nor U95632 ( n16225, n18715, n5183 );
nand U95633 ( n23518, n23851, n4243 );
nand U95634 ( n56640, n56975, n6875 );
nand U95635 ( n10320, n10730, n5155 );
nand U95636 ( n10322, n10730, n5157 );
nand U95637 ( n10325, n10730, n5152 );
nand U95638 ( n10327, n10730, n5153 );
not U95639 ( n6924, n60075 );
not U95640 ( n4292, n26935 );
not U95641 ( n4293, n28413 );
not U95642 ( n6925, n61722 );
not U95643 ( n3454, n34180 );
not U95644 ( n6069, n68934 );
not U95645 ( n3455, n35594 );
not U95646 ( n6070, n70322 );
not U95647 ( n6545, n54900 );
not U95648 ( n3913, n21824 );
not U95649 ( n3069, n29139 );
not U95650 ( n5670, n62806 );
not U95651 ( n7455, n42318 );
not U95652 ( n4812, n8257 );
nand U95653 ( n14730, n5179, n14732 );
nand U95654 ( n14732, n14733, n14734 );
nand U95655 ( n14723, n14724, n14725 );
nand U95656 ( n14725, n14727, n14728 );
nand U95657 ( n14724, n4768, n14730 );
nor U95658 ( n14727, n4769, n4772 );
nand U95659 ( n30464, n30783, n3410 );
nand U95660 ( n9873, n10274, n5158 );
nand U95661 ( n64623, n64985, n6025 );
nand U95662 ( n43780, n44143, n7813 );
not U95663 ( n3395, n30771 );
not U95664 ( n5143, n10259 );
not U95665 ( n6010, n64973 );
not U95666 ( n7798, n44131 );
nand U95667 ( n30745, n30763, n30764 );
nor U95668 ( n30763, n30786, n30787 );
nor U95669 ( n30764, n30765, n30766 );
nand U95670 ( n30786, n30795, n30796 );
nand U95671 ( n10230, n10249, n10250 );
nor U95672 ( n10249, n10278, n10279 );
nor U95673 ( n10250, n10252, n10253 );
nand U95674 ( n10278, n10289, n10290 );
nand U95675 ( n64951, n64965, n64966 );
nor U95676 ( n64965, n64988, n64989 );
nor U95677 ( n64966, n64967, n64968 );
nand U95678 ( n64988, n64997, n64998 );
nand U95679 ( n44108, n44123, n44124 );
nor U95680 ( n44123, n44146, n44147 );
nor U95681 ( n44124, n44125, n44126 );
nand U95682 ( n44146, n44155, n44156 );
nor U95683 ( n42861, n42863, n42864 );
nor U95684 ( n8829, n8832, n8833 );
nand U95685 ( n30461, n30783, n3414 );
nand U95686 ( n9869, n10274, n5162 );
nand U95687 ( n64620, n64985, n6029 );
nand U95688 ( n43777, n44143, n7817 );
nand U95689 ( n23133, n23476, n4248 );
nand U95690 ( n56254, n56598, n6880 );
not U95691 ( n4233, n23464 );
not U95692 ( n6865, n56586 );
nand U95693 ( n23435, n23456, n23457 );
nor U95694 ( n23456, n23479, n23480 );
nor U95695 ( n23457, n23458, n23459 );
nand U95696 ( n23479, n23488, n23489 );
nand U95697 ( n56557, n56578, n56579 );
nor U95698 ( n56578, n56601, n56602 );
nor U95699 ( n56579, n56580, n56581 );
nand U95700 ( n56601, n56610, n56611 );
nand U95701 ( n30460, n30783, n3413 );
nand U95702 ( n9868, n10274, n5160 );
nand U95703 ( n64619, n64985, n6028 );
nand U95704 ( n43776, n44143, n7815 );
nand U95705 ( n23130, n23476, n4252 );
nand U95706 ( n56251, n56598, n6884 );
nand U95707 ( n23129, n23476, n4250 );
nand U95708 ( n56250, n56598, n6883 );
nand U95709 ( n12680, n8294, n14640 );
nand U95710 ( n46293, n42382, n47873 );
and U95711 ( n30671, n30715, n30716 );
nor U95712 ( n30715, n30731, n30732 );
nor U95713 ( n30716, n30717, n30718 );
nand U95714 ( n30731, n30739, n30740 );
and U95715 ( n10135, n10193, n10194 );
nor U95716 ( n10193, n10213, n10214 );
nor U95717 ( n10194, n10195, n10197 );
nand U95718 ( n10213, n10223, n10224 );
and U95719 ( n64877, n64921, n64922 );
nor U95720 ( n64921, n64937, n64938 );
nor U95721 ( n64922, n64923, n64924 );
nand U95722 ( n64937, n64945, n64946 );
and U95723 ( n44032, n44078, n44079 );
nor U95724 ( n44078, n44094, n44095 );
nor U95725 ( n44079, n44080, n44081 );
nand U95726 ( n44094, n44102, n44103 );
and U95727 ( n23360, n23405, n23406 );
nor U95728 ( n23405, n23421, n23422 );
nor U95729 ( n23406, n23407, n23408 );
nand U95730 ( n23421, n23429, n23430 );
and U95731 ( n56484, n56527, n56528 );
nor U95732 ( n56527, n56543, n56544 );
nor U95733 ( n56528, n56529, n56530 );
nand U95734 ( n56543, n56551, n56552 );
nand U95735 ( n35519, n35346, n34624 );
nand U95736 ( n70247, n70078, n69370 );
nor U95737 ( n28111, n28412, n4273 );
nor U95738 ( n70078, n70321, n6050 );
nor U95739 ( n35346, n35593, n3435 );
nor U95740 ( n61266, n61721, n6905 );
not U95741 ( n228, n8314 );
not U95742 ( n4977, n12658 );
not U95743 ( n3243, n32571 );
not U95744 ( n7630, n46275 );
not U95745 ( n4068, n25329 );
not U95746 ( n5843, n67336 );
not U95747 ( n6700, n58468 );
nor U95748 ( n63513, n63515, n63516 );
nor U95749 ( n29614, n29616, n29617 );
nor U95750 ( n22293, n22295, n22296 );
nor U95751 ( n55405, n55407, n55408 );
not U95752 ( n202, n29189 );
not U95753 ( n168, n21872 );
not U95754 ( n473, n62907 );
not U95755 ( n440, n54963 );
not U95756 ( n499, n42398 );
nand U95757 ( n30452, n30792, n3410 );
nand U95758 ( n9858, n10285, n5158 );
nand U95759 ( n64611, n64994, n6025 );
nand U95760 ( n43768, n44152, n7813 );
nand U95761 ( n30449, n30792, n3414 );
nand U95762 ( n9854, n10285, n5162 );
nand U95763 ( n64608, n64994, n6029 );
nand U95764 ( n43765, n44152, n7817 );
nand U95765 ( n23121, n23485, n4248 );
nand U95766 ( n56242, n56607, n6880 );
nand U95767 ( n30448, n30792, n3413 );
nand U95768 ( n9853, n10285, n5160 );
nand U95769 ( n64607, n64994, n6028 );
nand U95770 ( n43764, n44152, n7815 );
nand U95771 ( n23118, n23485, n4252 );
nand U95772 ( n56239, n56607, n6884 );
nand U95773 ( n34390, n34459, n34381 );
nand U95774 ( n69142, n69209, n69133 );
nand U95775 ( n34556, n34381, n34624 );
nand U95776 ( n69304, n69133, n69370 );
nand U95777 ( n23117, n23485, n4250 );
nand U95778 ( n56238, n56607, n6883 );
nand U95779 ( n23122, n23475, n4233 );
nand U95780 ( n56243, n56597, n6865 );
nand U95781 ( n30453, n30782, n3395 );
nand U95782 ( n9859, n10273, n5143 );
nand U95783 ( n64612, n64984, n6010 );
nand U95784 ( n43769, n44142, n7798 );
nand U95785 ( n76130, n3077, n31818 );
nand U95786 ( n76129, n3077, n31818 );
and U95787 ( n27964, n27788, n27379 );
and U95788 ( n27800, n27788, n27214 );
and U95789 ( n61113, n60936, n60527 );
and U95790 ( n60948, n60936, n60359 );
and U95791 ( n35199, n35029, n34624 );
and U95792 ( n35041, n35029, n34459 );
and U95793 ( n69935, n69767, n69370 );
and U95794 ( n69779, n69767, n69209 );
xor U95795 ( n42880, n42864, n42863 );
xor U95796 ( n8853, n8833, n8832 );
and U95797 ( n28122, n28111, n27214 );
and U95798 ( n61277, n61266, n60359 );
and U95799 ( n35357, n35346, n34459 );
and U95800 ( n70089, n70078, n69209 );
not U95801 ( n7953, n42862 );
not U95802 ( n5298, n8830 );
nand U95803 ( n34641, n34378, n3444 );
nand U95804 ( n27396, n27134, n4282 );
nand U95805 ( n69387, n69130, n6059 );
nand U95806 ( n60544, n60278, n6914 );
not U95807 ( n5669, n68893 );
not U95808 ( n3068, n34139 );
not U95809 ( n6544, n60034 );
not U95810 ( n3912, n26894 );
nand U95811 ( n27042, n27134, n27122 );
nand U95812 ( n34286, n34378, n34367 );
nand U95813 ( n69038, n69130, n69119 );
nand U95814 ( n60183, n60278, n60266 );
nand U95815 ( n30657, n30672, n30673 );
nor U95816 ( n30672, n30688, n30689 );
nor U95817 ( n30673, n30674, n30675 );
nand U95818 ( n30688, n30696, n30697 );
nand U95819 ( n10110, n10137, n10138 );
nor U95820 ( n10137, n10157, n10158 );
nor U95821 ( n10138, n10139, n10140 );
nand U95822 ( n10157, n10167, n10168 );
nand U95823 ( n64863, n64878, n64879 );
nor U95824 ( n64878, n64894, n64895 );
nor U95825 ( n64879, n64880, n64881 );
nand U95826 ( n64894, n64902, n64903 );
nand U95827 ( n44016, n44033, n44034 );
nor U95828 ( n44033, n44049, n44050 );
nor U95829 ( n44034, n44035, n44036 );
nand U95830 ( n44049, n44057, n44058 );
nand U95831 ( n23343, n23361, n23362 );
nor U95832 ( n23361, n23377, n23378 );
nor U95833 ( n23362, n23363, n23364 );
nand U95834 ( n23377, n23385, n23386 );
nand U95835 ( n56467, n56485, n56486 );
nor U95836 ( n56485, n56501, n56502 );
nor U95837 ( n56486, n56487, n56488 );
nand U95838 ( n56501, n56509, n56510 );
not U95839 ( n6183, n66678 );
not U95840 ( n3568, n32075 );
not U95841 ( n4405, n24843 );
not U95842 ( n7038, n57977 );
not U95843 ( n4404, n24764 );
not U95844 ( n3567, n31996 );
not U95845 ( n6182, n66599 );
not U95846 ( n7037, n57898 );
not U95847 ( n4403, n24676 );
not U95848 ( n7035, n57810 );
not U95849 ( n3565, n31888 );
not U95850 ( n6180, n66511 );
not U95851 ( n6184, n66798 );
not U95852 ( n6187, n66934 );
not U95853 ( n3569, n32152 );
not U95854 ( n4407, n24920 );
not U95855 ( n4409, n25058 );
not U95856 ( n7039, n58057 );
not U95857 ( n7042, n58193 );
not U95858 ( n3572, n32295 );
nor U95859 ( n42386, n498, n42387 );
nor U95860 ( n42387, n7343, n42388 );
nor U95861 ( n42388, n7620, n7617 );
nor U95862 ( n8299, n227, n8300 );
nor U95863 ( n8300, n4711, n8302 );
nor U95864 ( n8302, n4967, n4963 );
nor U95865 ( n21860, n167, n21861 );
nor U95866 ( n21861, n3822, n21862 );
nor U95867 ( n21862, n4062, n4058 );
nor U95868 ( n29173, n200, n29174 );
nor U95869 ( n29174, n2978, n29175 );
nor U95870 ( n29175, n3234, n3230 );
nor U95871 ( n62895, n472, n62896 );
nor U95872 ( n62896, n5579, n62897 );
nor U95873 ( n62897, n5833, n5829 );
nor U95874 ( n54951, n439, n54952 );
nor U95875 ( n54952, n6454, n54953 );
nor U95876 ( n54953, n6694, n6690 );
nand U95877 ( n30465, n30771, n30782 );
nand U95878 ( n9874, n10259, n10273 );
nand U95879 ( n64624, n64973, n64984 );
nand U95880 ( n43781, n44131, n44142 );
nand U95881 ( n23134, n23464, n23475 );
nand U95882 ( n56255, n56586, n56597 );
and U95883 ( n30582, n30626, n30627 );
nor U95884 ( n30626, n30642, n30643 );
nor U95885 ( n30627, n30628, n30629 );
nand U95886 ( n30642, n30650, n30651 );
and U95887 ( n64741, n64832, n64833 );
nor U95888 ( n64832, n64848, n64849 );
nor U95889 ( n64833, n64834, n64835 );
nand U95890 ( n64848, n64856, n64857 );
and U95891 ( n43941, n43985, n43986 );
nor U95892 ( n43985, n44001, n44002 );
nor U95893 ( n43986, n43987, n43988 );
nand U95894 ( n44001, n44009, n44010 );
and U95895 ( n10025, n10072, n10073 );
nor U95896 ( n10072, n10092, n10093 );
nor U95897 ( n10073, n10074, n10075 );
nand U95898 ( n10092, n10102, n10103 );
and U95899 ( n23261, n23312, n23313 );
nor U95900 ( n23312, n23328, n23329 );
nor U95901 ( n23313, n23314, n23315 );
nand U95902 ( n23328, n23336, n23337 );
and U95903 ( n56385, n56436, n56437 );
nor U95904 ( n56436, n56452, n56453 );
nor U95905 ( n56437, n56438, n56439 );
nand U95906 ( n56452, n56460, n56461 );
and U95907 ( n27474, n27214, n27467 );
and U95908 ( n60623, n60359, n60616 );
and U95909 ( n34719, n34459, n34712 );
and U95910 ( n69463, n69209, n69456 );
not U95911 ( n5317, n12024 );
not U95912 ( n5314, n11838 );
not U95913 ( n5315, n11938 );
not U95914 ( n5318, n12125 );
not U95915 ( n5320, n12307 );
nand U95916 ( n60107, n60108, n60109 );
nand U95917 ( n26967, n26968, n26969 );
nand U95918 ( n34212, n34213, n34214 );
nand U95919 ( n68966, n68967, n68968 );
not U95920 ( n7972, n45770 );
not U95921 ( n7969, n45586 );
not U95922 ( n7970, n45675 );
not U95923 ( n7973, n45847 );
not U95924 ( n7975, n45983 );
buf U95925 ( n76238, n76236 );
buf U95926 ( n76237, n76236 );
buf U95927 ( n76239, n76236 );
buf U95928 ( n76507, n76505 );
buf U95929 ( n76506, n76505 );
buf U95930 ( n76306, n76305 );
buf U95931 ( n76307, n76305 );
buf U95932 ( n76508, n76505 );
buf U95933 ( n76308, n76305 );
buf U95934 ( n76565, n76564 );
buf U95935 ( n76566, n76564 );
buf U95936 ( n76567, n76564 );
nand U95937 ( n28297, n27217, n28398 );
nand U95938 ( n61519, n60362, n61679 );
nand U95939 ( n35523, n34462, n35581 );
nand U95940 ( n70251, n69212, n70309 );
nand U95941 ( n28046, n28108, n27217 );
nand U95942 ( n27721, n27785, n27217 );
nand U95943 ( n27315, n27376, n27217 );
nand U95944 ( n27233, n27294, n27217 );
nand U95945 ( n27151, n27210, n27217 );
nand U95946 ( n34560, n34621, n34462 );
nand U95947 ( n34478, n34539, n34462 );
nand U95948 ( n34394, n34455, n34462 );
nand U95949 ( n35283, n35343, n34462 );
nand U95950 ( n34966, n35026, n34462 );
nand U95951 ( n70017, n70075, n69212 );
nand U95952 ( n69706, n69764, n69212 );
nand U95953 ( n69308, n69367, n69212 );
nand U95954 ( n69228, n69287, n69212 );
nand U95955 ( n69146, n69205, n69212 );
nand U95956 ( n60458, n60524, n60362 );
nand U95957 ( n60378, n60437, n60362 );
nand U95958 ( n60293, n60355, n60362 );
nand U95959 ( n61205, n61263, n60362 );
nand U95960 ( n60872, n60933, n60362 );
nand U95961 ( n28124, n27217, n28191 );
nand U95962 ( n27966, n27217, n28029 );
nand U95963 ( n27884, n27217, n27947 );
nand U95964 ( n27802, n27217, n27869 );
nand U95965 ( n27563, n27217, n27626 );
nand U95966 ( n27477, n27217, n27547 );
nand U95967 ( n35359, n34462, n35424 );
nand U95968 ( n35201, n34462, n35266 );
nand U95969 ( n35123, n34462, n35186 );
nand U95970 ( n35043, n34462, n35108 );
nand U95971 ( n34806, n34462, n34871 );
nand U95972 ( n34721, n34462, n34791 );
nand U95973 ( n70091, n69212, n70154 );
nand U95974 ( n69937, n69212, n70000 );
nand U95975 ( n69859, n69212, n69922 );
nand U95976 ( n69781, n69212, n69844 );
nand U95977 ( n69550, n69212, n69613 );
nand U95978 ( n69465, n69212, n69535 );
nand U95979 ( n61279, n60362, n61355 );
nand U95980 ( n61115, n60362, n61188 );
nand U95981 ( n61031, n60362, n61100 );
nand U95982 ( n60950, n60362, n61016 );
nand U95983 ( n60713, n60362, n60779 );
nand U95984 ( n60626, n60362, n60699 );
nand U95985 ( n28205, n27217, n28272 );
nand U95986 ( n70168, n69212, n70231 );
nand U95987 ( n35438, n34462, n35503 );
nand U95988 ( n61369, n60362, n61494 );
nand U95989 ( n30567, n30583, n30584 );
nor U95990 ( n30583, n30599, n30600 );
nor U95991 ( n30584, n30585, n30586 );
nand U95992 ( n30599, n30607, n30608 );
nand U95993 ( n10012, n10026, n10027 );
nor U95994 ( n10026, n10042, n10043 );
nor U95995 ( n10027, n10028, n10029 );
nand U95996 ( n10042, n10050, n10051 );
nand U95997 ( n64726, n64742, n64743 );
nor U95998 ( n64742, n64758, n64759 );
nor U95999 ( n64743, n64744, n64745 );
nand U96000 ( n64758, n64766, n64767 );
nand U96001 ( n43928, n43942, n43943 );
nor U96002 ( n43942, n43958, n43959 );
nor U96003 ( n43943, n43944, n43945 );
nand U96004 ( n43958, n43966, n43967 );
nand U96005 ( n23247, n23262, n23263 );
nor U96006 ( n23262, n23278, n23279 );
nor U96007 ( n23263, n23264, n23265 );
nand U96008 ( n23278, n23286, n23287 );
nand U96009 ( n56368, n56386, n56387 );
nor U96010 ( n56386, n56402, n56403 );
nor U96011 ( n56387, n56388, n56389 );
nand U96012 ( n56402, n56410, n56411 );
and U96013 ( n27639, n27217, n27703 );
and U96014 ( n34884, n34462, n34948 );
and U96015 ( n69626, n69212, n69688 );
and U96016 ( n60792, n60362, n60854 );
and U96017 ( n30492, n30536, n30537 );
nor U96018 ( n30536, n30552, n30553 );
nor U96019 ( n30537, n30538, n30539 );
nand U96020 ( n30552, n30560, n30561 );
and U96021 ( n9913, n9975, n9977 );
nor U96022 ( n9975, n9995, n9997 );
nor U96023 ( n9977, n9978, n9979 );
nand U96024 ( n9995, n10005, n10006 );
and U96025 ( n64651, n64695, n64696 );
nor U96026 ( n64695, n64711, n64712 );
nor U96027 ( n64696, n64697, n64698 );
nand U96028 ( n64711, n64719, n64720 );
and U96029 ( n43812, n43897, n43898 );
nor U96030 ( n43897, n43913, n43914 );
nor U96031 ( n43898, n43899, n43900 );
nand U96032 ( n43913, n43921, n43922 );
and U96033 ( n23168, n23216, n23217 );
nor U96034 ( n23216, n23232, n23233 );
nor U96035 ( n23217, n23218, n23219 );
nand U96036 ( n23232, n23240, n23241 );
and U96037 ( n56289, n56337, n56338 );
nor U96038 ( n56337, n56353, n56354 );
nor U96039 ( n56338, n56339, n56340 );
nand U96040 ( n56353, n56361, n56362 );
nor U96041 ( n16119, n14934, n16034 );
nor U96042 ( n16020, n14934, n15927 );
nor U96043 ( n15913, n14934, n15822 );
nor U96044 ( n15598, n14934, n15513 );
nor U96045 ( n15500, n14934, n15407 );
nor U96046 ( n48709, n48122, n48625 );
nor U96047 ( n48615, n48122, n48531 );
nor U96048 ( n49075, n48122, n48991 );
nor U96049 ( n48980, n48122, n48892 );
nor U96050 ( n49344, n48122, n49276 );
nor U96051 ( n49437, n48122, n49354 );
nor U96052 ( n16433, n14934, n16342 );
nand U96053 ( n30254, n31119, n31120 );
nor U96054 ( n31120, n31121, n31122 );
nor U96055 ( n31119, n31146, n31147 );
nand U96056 ( n31122, n31123, n31124 );
nand U96057 ( n43565, n44498, n44499 );
nor U96058 ( n44499, n44500, n44501 );
nor U96059 ( n44498, n44525, n44526 );
nand U96060 ( n44501, n44502, n44503 );
nand U96061 ( n64316, n65373, n65374 );
nor U96062 ( n65374, n65375, n65376 );
nor U96063 ( n65373, n65400, n65401 );
nand U96064 ( n65376, n65377, n65378 );
or U96065 ( n34258, n34234, n3394 );
or U96066 ( n27015, n26989, n4232 );
or U96067 ( n69012, n68988, n6009 );
or U96068 ( n60156, n60132, n6864 );
nand U96069 ( n30245, n31073, n31074 );
nor U96070 ( n31074, n31075, n31076 );
nor U96071 ( n31073, n31089, n31090 );
nand U96072 ( n31076, n31077, n31078 );
nand U96073 ( n30193, n30861, n30862 );
nor U96074 ( n30862, n30863, n30864 );
nor U96075 ( n30861, n30877, n30878 );
nand U96076 ( n30864, n30865, n30866 );
nand U96077 ( n30207, n30903, n30904 );
nor U96078 ( n30904, n30905, n30906 );
nor U96079 ( n30903, n30919, n30920 );
nand U96080 ( n30906, n30907, n30908 );
nand U96081 ( n30216, n30946, n30947 );
nor U96082 ( n30947, n30948, n30949 );
nor U96083 ( n30946, n30962, n30963 );
nand U96084 ( n30949, n30950, n30951 );
nand U96085 ( n9580, n10533, n10534 );
nor U96086 ( n10534, n10535, n10537 );
nor U96087 ( n10533, n10553, n10554 );
nand U96088 ( n10537, n10538, n10539 );
nand U96089 ( n9590, n10588, n10589 );
nor U96090 ( n10589, n10590, n10592 );
nor U96091 ( n10588, n10608, n10609 );
nand U96092 ( n10592, n10593, n10594 );
nand U96093 ( n9557, n10427, n10428 );
nor U96094 ( n10428, n10429, n10430 );
nor U96095 ( n10427, n10447, n10448 );
nand U96096 ( n10430, n10432, n10433 );
nand U96097 ( n9544, n10372, n10373 );
nor U96098 ( n10373, n10374, n10375 );
nor U96099 ( n10372, n10392, n10393 );
nand U96100 ( n10375, n10377, n10378 );
nand U96101 ( n43524, n44350, n44351 );
nor U96102 ( n44351, n44352, n44353 );
nor U96103 ( n44350, n44366, n44367 );
nand U96104 ( n44353, n44354, n44355 );
nand U96105 ( n43533, n44408, n44409 );
nor U96106 ( n44409, n44410, n44411 );
nor U96107 ( n44408, n44424, n44425 );
nand U96108 ( n44411, n44412, n44413 );
nand U96109 ( n43495, n44221, n44222 );
nor U96110 ( n44222, n44223, n44224 );
nor U96111 ( n44221, n44237, n44238 );
nand U96112 ( n44224, n44225, n44226 );
nand U96113 ( n43505, n44265, n44266 );
nor U96114 ( n44266, n44267, n44268 );
nor U96115 ( n44265, n44281, n44282 );
nand U96116 ( n44268, n44269, n44270 );
nand U96117 ( n43543, n44450, n44451 );
nor U96118 ( n44451, n44452, n44453 );
nor U96119 ( n44450, n44466, n44467 );
nand U96120 ( n44453, n44454, n44455 );
nand U96121 ( n9603, n10640, n10642 );
nor U96122 ( n10642, n10643, n10644 );
nor U96123 ( n10640, n10660, n10662 );
nand U96124 ( n10644, n10645, n10647 );
nand U96125 ( n64259, n65063, n65064 );
nor U96126 ( n65064, n65065, n65066 );
nor U96127 ( n65063, n65079, n65080 );
nand U96128 ( n65066, n65067, n65068 );
nand U96129 ( n64269, n65105, n65106 );
nor U96130 ( n65106, n65107, n65108 );
nor U96131 ( n65105, n65121, n65122 );
nand U96132 ( n65108, n65109, n65110 );
nand U96133 ( n64278, n65148, n65149 );
nor U96134 ( n65149, n65150, n65151 );
nor U96135 ( n65148, n65164, n65165 );
nand U96136 ( n65151, n65152, n65153 );
nand U96137 ( n64288, n65190, n65191 );
nor U96138 ( n65191, n65192, n65193 );
nor U96139 ( n65190, n65206, n65207 );
nand U96140 ( n65193, n65194, n65195 );
nand U96141 ( n64297, n65233, n65234 );
nor U96142 ( n65234, n65235, n65236 );
nor U96143 ( n65233, n65249, n65250 );
nand U96144 ( n65236, n65237, n65238 );
nand U96145 ( n30226, n30988, n30989 );
nor U96146 ( n30989, n30990, n30991 );
nor U96147 ( n30988, n31004, n31005 );
nand U96148 ( n30991, n30992, n30993 );
nand U96149 ( n30235, n31031, n31032 );
nor U96150 ( n31032, n31033, n31034 );
nor U96151 ( n31031, n31047, n31048 );
nand U96152 ( n31034, n31035, n31036 );
nand U96153 ( n64307, n65275, n65276 );
nor U96154 ( n65276, n65277, n65278 );
nor U96155 ( n65275, n65291, n65292 );
nand U96156 ( n65278, n65279, n65280 );
nand U96157 ( n9614, n10700, n10702 );
nor U96158 ( n10702, n10703, n10704 );
nor U96159 ( n10700, n10734, n10735 );
nand U96160 ( n10704, n10705, n10707 );
nand U96161 ( n9568, n10483, n10484 );
nor U96162 ( n10484, n10485, n10487 );
nor U96163 ( n10483, n10503, n10504 );
nand U96164 ( n10487, n10488, n10489 );
nand U96165 ( n43514, n44310, n44311 );
nor U96166 ( n44311, n44312, n44313 );
nor U96167 ( n44310, n44326, n44327 );
nand U96168 ( n44313, n44314, n44315 );
nand U96169 ( n22889, n23645, n23646 );
nor U96170 ( n23646, n23647, n23648 );
nor U96171 ( n23645, n23661, n23662 );
nand U96172 ( n23648, n23649, n23650 );
nand U96173 ( n22899, n23689, n23690 );
nor U96174 ( n23690, n23691, n23692 );
nor U96175 ( n23689, n23705, n23706 );
nand U96176 ( n23692, n23693, n23694 );
nand U96177 ( n22908, n23734, n23735 );
nor U96178 ( n23735, n23736, n23737 );
nor U96179 ( n23734, n23750, n23751 );
nand U96180 ( n23737, n23738, n23739 );
nand U96181 ( n22880, n23600, n23601 );
nor U96182 ( n23601, n23602, n23603 );
nor U96183 ( n23600, n23616, n23617 );
nand U96184 ( n23603, n23604, n23605 );
nand U96185 ( n22870, n23556, n23557 );
nor U96186 ( n23557, n23558, n23559 );
nor U96187 ( n23556, n23572, n23573 );
nand U96188 ( n23559, n23560, n23561 );
nand U96189 ( n55995, n56722, n56723 );
nor U96190 ( n56723, n56724, n56725 );
nor U96191 ( n56722, n56738, n56739 );
nand U96192 ( n56725, n56726, n56727 );
nand U96193 ( n56004, n56767, n56768 );
nor U96194 ( n56768, n56769, n56770 );
nor U96195 ( n56767, n56783, n56784 );
nand U96196 ( n56770, n56771, n56772 );
nand U96197 ( n55985, n56678, n56679 );
nor U96198 ( n56679, n56680, n56681 );
nor U96199 ( n56678, n56694, n56695 );
nand U96200 ( n56681, n56682, n56683 );
nand U96201 ( n56014, n56811, n56812 );
nor U96202 ( n56812, n56813, n56814 );
nor U96203 ( n56811, n56827, n56828 );
nand U96204 ( n56814, n56815, n56816 );
nand U96205 ( n56023, n56856, n56857 );
nor U96206 ( n56857, n56858, n56859 );
nor U96207 ( n56856, n56872, n56873 );
nand U96208 ( n56859, n56860, n56861 );
nand U96209 ( n22918, n23778, n23779 );
nor U96210 ( n23779, n23780, n23781 );
nor U96211 ( n23778, n23794, n23795 );
nand U96212 ( n23781, n23782, n23783 );
nand U96213 ( n56033, n56903, n56904 );
nor U96214 ( n56904, n56905, n56906 );
nor U96215 ( n56903, n56919, n56920 );
nand U96216 ( n56906, n56907, n56908 );
not U96217 ( n205, n30074 );
not U96218 ( n477, n64091 );
not U96219 ( n2892, n38313 );
and U96220 ( n49451, n76325, n7453 );
and U96221 ( n16450, n76591, n4809 );
not U96222 ( n1775, n48449 );
nand U96223 ( n30477, n30493, n30494 );
nor U96224 ( n30493, n30509, n30510 );
nor U96225 ( n30494, n30495, n30496 );
nand U96226 ( n30509, n30517, n30518 );
nand U96227 ( n9889, n9914, n9915 );
nor U96228 ( n9914, n9934, n9935 );
nor U96229 ( n9915, n9917, n9918 );
nand U96230 ( n9934, n9944, n9945 );
nand U96231 ( n64636, n64652, n64653 );
nor U96232 ( n64652, n64668, n64669 );
nor U96233 ( n64653, n64654, n64655 );
nand U96234 ( n64668, n64676, n64677 );
nand U96235 ( n43793, n43813, n43814 );
nor U96236 ( n43813, n43829, n43830 );
nor U96237 ( n43814, n43815, n43816 );
nand U96238 ( n43829, n43837, n43838 );
nand U96239 ( n23146, n23169, n23170 );
nor U96240 ( n23169, n23185, n23186 );
nor U96241 ( n23170, n23171, n23172 );
nand U96242 ( n23185, n23193, n23194 );
nand U96243 ( n56267, n56290, n56291 );
nor U96244 ( n56290, n56306, n56307 );
nor U96245 ( n56291, n56292, n56293 );
nand U96246 ( n56306, n56314, n56315 );
not U96247 ( n7862, n53885 );
nand U96248 ( n22927, n23827, n23828 );
nor U96249 ( n23828, n23829, n23830 );
nor U96250 ( n23827, n23854, n23855 );
nand U96251 ( n23830, n23831, n23832 );
nand U96252 ( n56042, n56951, n56952 );
nor U96253 ( n56952, n56953, n56954 );
nor U96254 ( n56951, n56978, n56979 );
nand U96255 ( n56954, n56955, n56956 );
nand U96256 ( n51667, n51665, n53884 );
nand U96257 ( n53884, n49247, n7862 );
and U96258 ( n49448, n76325, n76175 );
and U96259 ( n16447, n76591, n76185 );
nand U96260 ( n15733, n5198, n4756 );
nand U96261 ( n48828, n7853, n7400 );
nand U96262 ( n15752, n5198, n4755 );
nand U96263 ( n48836, n7853, n7399 );
nand U96264 ( n15723, n5198, n4757 );
nand U96265 ( n48820, n7853, n7402 );
nand U96266 ( n15762, n5198, n4754 );
nand U96267 ( n48844, n7853, n7398 );
nand U96268 ( n15772, n5198, n4753 );
nand U96269 ( n48852, n7853, n7397 );
not U96270 ( n76557, n76559 );
nand U96271 ( n15708, n5198, n4758 );
nand U96272 ( n48808, n7853, n7403 );
nand U96273 ( n15782, n5198, n4752 );
nand U96274 ( n48860, n7853, n7395 );
nand U96275 ( n49163, n49086, n49168 );
nand U96276 ( n49168, n48878, n7862 );
not U96277 ( n76464, n76466 );
nand U96278 ( n48406, n48350, n48411 );
nand U96279 ( n48411, n48131, n7862 );
nand U96280 ( n30430, n30454, n30455 );
nor U96281 ( n30454, n30466, n30467 );
nor U96282 ( n30455, n30456, n30457 );
nand U96283 ( n30466, n30472, n30473 );
nand U96284 ( n9830, n9860, n9862 );
nor U96285 ( n9860, n9875, n9877 );
nor U96286 ( n9862, n9863, n9864 );
nand U96287 ( n9875, n9883, n9884 );
nand U96288 ( n64589, n64613, n64614 );
nor U96289 ( n64613, n64625, n64626 );
nor U96290 ( n64614, n64615, n64616 );
nand U96291 ( n64625, n64631, n64632 );
nand U96292 ( n43746, n43770, n43771 );
nor U96293 ( n43770, n43782, n43783 );
nor U96294 ( n43771, n43772, n43773 );
nand U96295 ( n43782, n43788, n43789 );
nand U96296 ( n23099, n23123, n23124 );
nor U96297 ( n23123, n23135, n23136 );
nor U96298 ( n23124, n23125, n23126 );
nand U96299 ( n23135, n23141, n23142 );
nand U96300 ( n56220, n56244, n56245 );
nor U96301 ( n56244, n56256, n56257 );
nor U96302 ( n56245, n56246, n56247 );
nand U96303 ( n56256, n56262, n56263 );
nand U96304 ( n16012, n15927, n16018 );
nand U96305 ( n16018, n15804, n15162 );
nand U96306 ( n16110, n16034, n16117 );
nand U96307 ( n16117, n15804, n5209 );
nor U96308 ( n9023, n9025, n9027 );
nor U96309 ( n43030, n43032, n43033 );
not U96310 ( n5192, n15390 );
nand U96311 ( n15589, n15513, n15595 );
nand U96312 ( n15595, n15162, n5192 );
nand U96313 ( n49068, n48991, n49073 );
nand U96314 ( n49073, n48878, n48315 );
not U96315 ( n7847, n48518 );
nand U96316 ( n48702, n48625, n48707 );
nand U96317 ( n48707, n48315, n7847 );
not U96318 ( n76558, n76559 );
not U96319 ( n5293, n9024 );
not U96320 ( n7948, n43031 );
nand U96321 ( n18711, n18709, n20928 );
nand U96322 ( n20928, n16220, n5209 );
nor U96323 ( n15312, n14854, n15292 );
nor U96324 ( n48461, n48051, n48429 );
and U96325 ( n15803, n5208, n15804 );
not U96326 ( n76465, n76466 );
nand U96327 ( n10797, n11165, n5160 );
nand U96328 ( n44570, n44879, n7815 );
nand U96329 ( n31190, n31494, n3413 );
nand U96330 ( n65444, n65744, n6028 );
nor U96331 ( n63729, n63731, n63732 );
nor U96332 ( n29769, n29771, n29772 );
nor U96333 ( n22448, n22450, n22451 );
nor U96334 ( n55563, n55565, n55566 );
nand U96335 ( n30264, n31182, n31183 );
nor U96336 ( n31182, n31206, n31207 );
nor U96337 ( n31183, n31184, n31185 );
nand U96338 ( n31206, n31218, n31219 );
nand U96339 ( n30273, n31239, n31240 );
nor U96340 ( n31239, n31255, n31256 );
nor U96341 ( n31240, n31241, n31242 );
nand U96342 ( n31255, n31263, n31264 );
nand U96343 ( n30283, n31283, n31284 );
nor U96344 ( n31283, n31299, n31300 );
nor U96345 ( n31284, n31285, n31286 );
nand U96346 ( n31299, n31307, n31308 );
nand U96347 ( n30292, n31324, n31325 );
nor U96348 ( n31324, n31340, n31341 );
nor U96349 ( n31325, n31326, n31327 );
nand U96350 ( n31340, n31348, n31349 );
nand U96351 ( n30306, n31364, n31365 );
nor U96352 ( n31364, n31380, n31381 );
nor U96353 ( n31365, n31366, n31367 );
nand U96354 ( n31380, n31388, n31389 );
nand U96355 ( n9638, n10855, n10857 );
nor U96356 ( n10855, n10875, n10877 );
nor U96357 ( n10857, n10858, n10859 );
nand U96358 ( n10875, n10885, n10887 );
nand U96359 ( n9654, n10905, n10907 );
nor U96360 ( n10905, n10925, n10927 );
nor U96361 ( n10907, n10908, n10909 );
nand U96362 ( n10925, n10935, n10937 );
nand U96363 ( n9665, n10957, n10958 );
nor U96364 ( n10957, n10977, n10978 );
nor U96365 ( n10958, n10959, n10960 );
nand U96366 ( n10977, n10987, n10988 );
nand U96367 ( n9678, n11005, n11007 );
nor U96368 ( n11005, n11025, n11027 );
nor U96369 ( n11007, n11008, n11009 );
nand U96370 ( n11025, n11035, n11037 );
nand U96371 ( n9689, n11055, n11057 );
nor U96372 ( n11055, n11075, n11077 );
nor U96373 ( n11057, n11058, n11059 );
nand U96374 ( n11075, n11085, n11087 );
nand U96375 ( n9702, n11107, n11108 );
nor U96376 ( n11107, n11127, n11128 );
nor U96377 ( n11108, n11109, n11110 );
nand U96378 ( n11127, n11137, n11138 );
nand U96379 ( n9713, n11155, n11157 );
nor U96380 ( n11155, n11185, n11187 );
nor U96381 ( n11157, n11158, n11159 );
nand U96382 ( n11185, n11202, n11203 );
nand U96383 ( n64396, n65493, n65494 );
nor U96384 ( n65493, n65509, n65510 );
nor U96385 ( n65494, n65495, n65496 );
nand U96386 ( n65509, n65517, n65518 );
nand U96387 ( n64406, n65533, n65534 );
nor U96388 ( n65533, n65549, n65550 );
nor U96389 ( n65534, n65535, n65536 );
nand U96390 ( n65549, n65557, n65558 );
nand U96391 ( n64415, n65574, n65575 );
nor U96392 ( n65574, n65590, n65591 );
nor U96393 ( n65575, n65576, n65577 );
nand U96394 ( n65590, n65598, n65599 );
nand U96395 ( n64425, n65614, n65615 );
nor U96396 ( n65614, n65630, n65631 );
nor U96397 ( n65615, n65616, n65617 );
nand U96398 ( n65630, n65638, n65639 );
nand U96399 ( n43594, n44657, n44658 );
nor U96400 ( n44657, n44673, n44674 );
nor U96401 ( n44658, n44659, n44660 );
nand U96402 ( n44673, n44681, n44682 );
nand U96403 ( n43603, n44698, n44699 );
nor U96404 ( n44698, n44714, n44715 );
nor U96405 ( n44699, n44700, n44701 );
nand U96406 ( n44714, n44722, n44723 );
nand U96407 ( n43613, n44737, n44738 );
nor U96408 ( n44737, n44753, n44754 );
nor U96409 ( n44738, n44739, n44740 );
nand U96410 ( n44753, n44761, n44762 );
nand U96411 ( n43622, n44777, n44778 );
nor U96412 ( n44777, n44793, n44794 );
nor U96413 ( n44778, n44779, n44780 );
nand U96414 ( n44793, n44801, n44802 );
nand U96415 ( n43641, n44871, n44872 );
nor U96416 ( n44871, n44895, n44896 );
nor U96417 ( n44872, n44873, n44874 );
nand U96418 ( n44895, n44908, n44909 );
nand U96419 ( n43632, n44818, n44819 );
nor U96420 ( n44818, n44834, n44835 );
nor U96421 ( n44819, n44820, n44821 );
nand U96422 ( n44834, n44842, n44843 );
nand U96423 ( n43584, n44617, n44618 );
nor U96424 ( n44617, n44633, n44634 );
nor U96425 ( n44618, n44619, n44620 );
nand U96426 ( n44633, n44641, n44642 );
nand U96427 ( n9627, n10787, n10788 );
nor U96428 ( n10787, n10817, n10818 );
nor U96429 ( n10788, n10789, n10790 );
nand U96430 ( n10817, n10832, n10833 );
nand U96431 ( n64326, n65436, n65437 );
nor U96432 ( n65436, n65460, n65461 );
nor U96433 ( n65437, n65438, n65439 );
nand U96434 ( n65460, n65472, n65473 );
nand U96435 ( n43575, n44562, n44563 );
nor U96436 ( n44562, n44586, n44587 );
nor U96437 ( n44563, n44564, n44565 );
nand U96438 ( n44586, n44598, n44599 );
nand U96439 ( n30315, n31405, n31406 );
nor U96440 ( n31405, n31421, n31422 );
nor U96441 ( n31406, n31407, n31408 );
nand U96442 ( n31421, n31429, n31430 );
nand U96443 ( n30325, n31445, n31446 );
nor U96444 ( n31445, n31461, n31462 );
nor U96445 ( n31446, n31447, n31448 );
nand U96446 ( n31461, n31469, n31470 );
nand U96447 ( n30334, n31486, n31487 );
nor U96448 ( n31486, n31510, n31511 );
nor U96449 ( n31487, n31488, n31489 );
nand U96450 ( n31510, n31523, n31524 );
nand U96451 ( n64434, n65655, n65656 );
nor U96452 ( n65655, n65671, n65672 );
nor U96453 ( n65656, n65657, n65658 );
nand U96454 ( n65671, n65679, n65680 );
nand U96455 ( n64444, n65695, n65696 );
nor U96456 ( n65695, n65711, n65712 );
nor U96457 ( n65696, n65697, n65698 );
nand U96458 ( n65711, n65719, n65720 );
nand U96459 ( n64453, n65736, n65737 );
nor U96460 ( n65736, n65760, n65761 );
nor U96461 ( n65737, n65738, n65739 );
nand U96462 ( n65760, n65773, n65774 );
nor U96463 ( n15323, n14868, n15292 );
nor U96464 ( n48470, n48062, n48429 );
nand U96465 ( n10802, n11165, n5158 );
nand U96466 ( n44574, n44879, n7813 );
nand U96467 ( n31194, n31494, n3410 );
nand U96468 ( n65448, n65744, n6025 );
nor U96469 ( n15300, n14840, n15292 );
nor U96470 ( n48436, n48040, n48429 );
nor U96471 ( n15334, n14882, n15292 );
nor U96472 ( n48479, n48087, n48429 );
nor U96473 ( n9048, n5280, n9025 );
nor U96474 ( n43050, n7935, n43032 );
nor U96475 ( n9075, n5280, n9077 );
nor U96476 ( n9077, n9078, n9079 );
nor U96477 ( n9078, n9080, n9082 );
nor U96478 ( n43072, n7935, n43073 );
nor U96479 ( n43073, n43074, n43075 );
nor U96480 ( n43074, n43076, n43077 );
nor U96481 ( n15352, n14895, n15292 );
nor U96482 ( n48488, n48098, n48429 );
nand U96483 ( n10798, n11165, n5162 );
nand U96484 ( n44571, n44879, n7817 );
nand U96485 ( n31191, n31494, n3414 );
nand U96486 ( n65445, n65744, n6029 );
not U96487 ( n7454, n47873 );
nor U96488 ( n48140, n7450, n7863 );
not U96489 ( n7450, n48227 );
nor U96490 ( n15283, n14824, n15292 );
nor U96491 ( n48422, n48027, n48429 );
not U96492 ( n503, n43346 );
and U96493 ( n48877, n48130, n48878 );
nand U96494 ( n48032, n48140, n48131 );
nand U96495 ( n10803, n11165, n5150 );
nand U96496 ( n44575, n44879, n7805 );
nand U96497 ( n31195, n31494, n3403 );
nand U96498 ( n65449, n65744, n6018 );
nor U96499 ( n15363, n14909, n15292 );
nor U96500 ( n48497, n48109, n48429 );
nand U96501 ( n48346, n48406, n48227 );
not U96502 ( n172, n22753 );
not U96503 ( n444, n55867 );
not U96504 ( n2889, n38345 );
nand U96505 ( n15297, n14955, n5192 );
not U96506 ( n4810, n14640 );
nand U96507 ( n14830, n14955, n14944 );
not U96508 ( n1773, n48679 );
not U96509 ( n232, n9399 );
nand U96510 ( n57019, n57322, n6883 );
nand U96511 ( n23895, n24200, n4250 );
nand U96512 ( n22937, n23887, n23888 );
nor U96513 ( n23887, n23911, n23912 );
nor U96514 ( n23888, n23889, n23890 );
nand U96515 ( n23911, n23923, n23924 );
nand U96516 ( n56055, n57011, n57012 );
nor U96517 ( n57011, n57035, n57036 );
nor U96518 ( n57012, n57013, n57014 );
nand U96519 ( n57035, n57047, n57048 );
nand U96520 ( n57023, n57322, n6880 );
nand U96521 ( n23899, n24200, n4248 );
nand U96522 ( n15264, n15185, n15270 );
nand U96523 ( n15270, n14944, n5209 );
nand U96524 ( n48151, n48226, n48227 );
nand U96525 ( n16424, n16342, n16430 );
nand U96526 ( n16430, n16220, n15162 );
not U96527 ( n6160, n63730 );
not U96528 ( n3545, n29770 );
not U96529 ( n4383, n22449 );
not U96530 ( n7015, n55564 );
nand U96531 ( n57020, n57322, n6884 );
nand U96532 ( n23896, n24200, n4252 );
nand U96533 ( n22956, n23989, n23990 );
nor U96534 ( n23989, n24005, n24006 );
nor U96535 ( n23990, n23991, n23992 );
nand U96536 ( n24005, n24013, n24014 );
nand U96537 ( n22967, n24030, n24031 );
nor U96538 ( n24030, n24046, n24047 );
nor U96539 ( n24031, n24032, n24033 );
nand U96540 ( n24046, n24054, n24055 );
nand U96541 ( n22977, n24070, n24071 );
nor U96542 ( n24070, n24086, n24087 );
nor U96543 ( n24071, n24072, n24073 );
nand U96544 ( n24086, n24094, n24095 );
nand U96545 ( n56064, n57071, n57072 );
nor U96546 ( n57071, n57087, n57088 );
nor U96547 ( n57072, n57073, n57074 );
nand U96548 ( n57087, n57095, n57096 );
nand U96549 ( n56074, n57111, n57112 );
nor U96550 ( n57111, n57127, n57128 );
nor U96551 ( n57112, n57113, n57114 );
nand U96552 ( n57127, n57135, n57136 );
nand U96553 ( n56083, n57152, n57153 );
nor U96554 ( n57152, n57168, n57169 );
nor U96555 ( n57153, n57154, n57155 );
nand U96556 ( n57168, n57176, n57177 );
nand U96557 ( n56093, n57192, n57193 );
nor U96558 ( n57192, n57208, n57209 );
nor U96559 ( n57193, n57194, n57195 );
nand U96560 ( n57208, n57216, n57217 );
nand U96561 ( n22946, n23949, n23950 );
nor U96562 ( n23949, n23965, n23966 );
nor U96563 ( n23950, n23951, n23952 );
nand U96564 ( n23965, n23973, n23974 );
nand U96565 ( n56102, n57233, n57234 );
nor U96566 ( n57233, n57249, n57250 );
nor U96567 ( n57234, n57235, n57236 );
nand U96568 ( n57249, n57257, n57258 );
nand U96569 ( n56112, n57273, n57274 );
nor U96570 ( n57273, n57289, n57290 );
nor U96571 ( n57274, n57275, n57276 );
nand U96572 ( n57289, n57297, n57298 );
nand U96573 ( n56121, n57314, n57315 );
nor U96574 ( n57314, n57338, n57339 );
nor U96575 ( n57315, n57316, n57317 );
nand U96576 ( n57338, n57351, n57352 );
nand U96577 ( n22986, n24111, n24112 );
nor U96578 ( n24111, n24127, n24128 );
nor U96579 ( n24112, n24113, n24114 );
nand U96580 ( n24127, n24135, n24136 );
nand U96581 ( n22996, n24151, n24152 );
nor U96582 ( n24151, n24167, n24168 );
nor U96583 ( n24152, n24153, n24154 );
nand U96584 ( n24167, n24175, n24176 );
nand U96585 ( n23005, n24192, n24193 );
nor U96586 ( n24192, n24216, n24217 );
nor U96587 ( n24193, n24194, n24195 );
nand U96588 ( n24216, n24229, n24230 );
nand U96589 ( n23900, n24200, n4240 );
nand U96590 ( n57024, n57322, n6873 );
nand U96591 ( n49430, n49354, n49435 );
nand U96592 ( n49435, n49247, n48315 );
nor U96593 ( n48517, n7863, n48518 );
nand U96594 ( n30083, n2978, n205 );
nand U96595 ( n27947, n27888, n27949 );
nand U96596 ( n27949, n27793, n27301 );
nand U96597 ( n61100, n61035, n61102 );
nand U96598 ( n61102, n60941, n60444 );
nand U96599 ( n28029, n27970, n28031 );
nand U96600 ( n28031, n27793, n4290 );
nand U96601 ( n61188, n61119, n61190 );
nand U96602 ( n61190, n60941, n6923 );
nand U96603 ( n35186, n35127, n35188 );
nand U96604 ( n35188, n35034, n34546 );
nand U96605 ( n69922, n69863, n69924 );
nand U96606 ( n69924, n69772, n69294 );
nand U96607 ( n35266, n35205, n35268 );
nand U96608 ( n35268, n35034, n3453 );
nand U96609 ( n70000, n69941, n70002 );
nand U96610 ( n70002, n69772, n6068 );
nand U96611 ( n64100, n5579, n477 );
not U96612 ( n4282, n27460 );
not U96613 ( n3444, n34705 );
not U96614 ( n6059, n69449 );
not U96615 ( n6914, n60609 );
buf U96616 ( n76040, n76921 );
nand U96617 ( n27626, n27567, n27628 );
nand U96618 ( n27628, n27301, n4282 );
nand U96619 ( n34871, n34810, n34873 );
nand U96620 ( n34873, n34546, n3444 );
nand U96621 ( n69613, n69554, n69615 );
nand U96622 ( n69615, n69294, n6059 );
nand U96623 ( n60779, n60717, n60781 );
nand U96624 ( n60781, n60444, n6914 );
not U96625 ( n4768, n14688 );
not U96626 ( n5209, n20929 );
nand U96627 ( n60090, n54947, n60105 );
nand U96628 ( n26950, n21856, n26965 );
nand U96629 ( n34195, n29169, n34210 );
nand U96630 ( n68949, n62891, n68964 );
nand U96631 ( n14969, n15044, n15045 );
nand U96632 ( n15073, n15154, n15045 );
nand U96633 ( n15180, n15264, n15045 );
and U96634 ( n16219, n5208, n16220 );
and U96635 ( n14943, n5208, n14944 );
nand U96636 ( n15470, n15045, n15492 );
nand U96637 ( n15577, n15045, n15589 );
nand U96638 ( n48249, n48309, n48227 );
nand U96639 ( n49152, n48227, n49163 );
and U96640 ( n49246, n48130, n49247 );
nor U96641 ( n14722, n14679, n14735 );
and U96642 ( n48129, n48130, n48131 );
nand U96643 ( n48769, n48227, n48779 );
and U96644 ( n27785, n27793, n4294 );
and U96645 ( n60933, n60941, n6927 );
nand U96646 ( n48598, n48227, n48608 );
and U96647 ( n35026, n35034, n3457 );
and U96648 ( n69764, n69772, n6072 );
nor U96649 ( n47940, n47904, n47941 );
nand U96650 ( n49648, n48227, n51667 );
nand U96651 ( n48692, n48227, n48702 );
nand U96652 ( n15712, n15810, n15804 );
nand U96653 ( n16130, n15810, n16220 );
nand U96654 ( n49180, n48883, n49247 );
nand U96655 ( n48811, n48883, n48878 );
nor U96656 ( n48883, n49252, n7863 );
nor U96657 ( n49252, n7453, n48133 );
nand U96658 ( n22762, n3822, n172 );
nand U96659 ( n16098, n15045, n16110 );
nand U96660 ( n15990, n15045, n16012 );
nand U96661 ( n15892, n15045, n15904 );
nand U96662 ( n48963, n48227, n48973 );
nand U96663 ( n49327, n48227, n49337 );
nor U96664 ( n63772, n63773, n63774 );
nor U96665 ( n63773, n63775, n63776 );
nor U96666 ( n29812, n29813, n29814 );
nor U96667 ( n29813, n29815, n29816 );
nor U96668 ( n22493, n22494, n22495 );
nor U96669 ( n22494, n22496, n22497 );
nor U96670 ( n55606, n55607, n55608 );
nor U96671 ( n55607, n55609, n55610 );
nand U96672 ( n49058, n48227, n49068 );
nand U96673 ( n55876, n6454, n444 );
nand U96674 ( n15678, n15045, n15692 );
buf U96675 ( n76326, n47970 );
buf U96676 ( n76592, n14747 );
nand U96677 ( n34621, n34559, n34627 );
nand U96678 ( n34627, n34367, n3453 );
nand U96679 ( n69367, n69307, n69373 );
nand U96680 ( n69373, n69119, n6068 );
nand U96681 ( n27376, n27314, n27382 );
nand U96682 ( n27382, n27122, n4290 );
nand U96683 ( n60524, n60457, n60530 );
nand U96684 ( n60530, n60266, n6923 );
nand U96685 ( n35581, n35516, n35588 );
nand U96686 ( n35588, n35350, n3453 );
nand U96687 ( n28398, n28288, n28407 );
nand U96688 ( n28407, n28115, n4290 );
nand U96689 ( n70309, n70244, n70316 );
nand U96690 ( n70316, n70082, n6068 );
nand U96691 ( n61679, n61510, n61716 );
nand U96692 ( n61716, n61270, n6923 );
nor U96693 ( n9140, n5282, n9142 );
nor U96694 ( n9142, n9143, n9144 );
nor U96695 ( n9143, n9145, n9147 );
nor U96696 ( n43124, n7937, n43125 );
nor U96697 ( n43125, n43126, n43127 );
nor U96698 ( n43126, n43128, n43129 );
nand U96699 ( n28272, n28209, n28274 );
nand U96700 ( n28274, n28115, n27301 );
nand U96701 ( n61494, n61373, n61496 );
nand U96702 ( n61496, n61270, n60444 );
nand U96703 ( n70231, n70172, n70233 );
nand U96704 ( n70233, n70082, n69294 );
nand U96705 ( n35503, n35442, n35505 );
nand U96706 ( n35505, n35350, n34546 );
buf U96707 ( n76050, n76045 );
buf U96708 ( n76053, n76046 );
buf U96709 ( n76047, n76045 );
buf U96710 ( n76052, n76046 );
buf U96711 ( n76049, n76045 );
buf U96712 ( n76051, n76046 );
buf U96713 ( n76048, n76045 );
buf U96714 ( n76033, n76560 );
not U96715 ( n1800, n48911 );
not U96716 ( n2918, n38377 );
buf U96717 ( n76031, n76560 );
buf U96718 ( n76032, n76560 );
buf U96719 ( n76054, n76046 );
buf U96720 ( n76120, n76115 );
buf U96721 ( n76123, n76116 );
buf U96722 ( n76117, n76115 );
buf U96723 ( n76122, n76116 );
buf U96724 ( n76119, n76115 );
buf U96725 ( n76121, n76116 );
buf U96726 ( n76118, n76115 );
buf U96727 ( n76232, n75011 );
buf U96728 ( n76124, n76116 );
buf U96729 ( n76499, n75027 );
nand U96730 ( n18709, n16217, n5204 );
buf U96731 ( n76298, n75029 );
nand U96732 ( n51665, n49244, n7865 );
buf U96733 ( n76056, n70861 );
buf U96734 ( n76020, n76467 );
buf U96735 ( n76055, n70861 );
buf U96736 ( n76018, n76467 );
buf U96737 ( n76019, n76467 );
buf U96738 ( n76126, n36141 );
buf U96739 ( n76642, n75047 );
buf U96740 ( n76125, n36141 );
not U96741 ( n6078, n68253 );
not U96742 ( n7868, n47222 );
not U96743 ( n4300, n26252 );
not U96744 ( n6933, n59391 );
and U96745 ( n28108, n28115, n4294 );
and U96746 ( n61263, n61270, n6927 );
and U96747 ( n35343, n35350, n3457 );
and U96748 ( n70075, n70082, n6072 );
buf U96749 ( n76370, n75048 );
buf U96750 ( n76552, n75049 );
not U96751 ( n5214, n13834 );
and U96752 ( n27121, n4294, n27122 );
and U96753 ( n34366, n3457, n34367 );
and U96754 ( n69118, n6072, n69119 );
and U96755 ( n60265, n6927, n60266 );
nand U96756 ( n9412, n4711, n232 );
nand U96757 ( n16412, n15045, n16424 );
nand U96758 ( n43356, n7343, n503 );
not U96759 ( n3463, n33498 );
nand U96760 ( n49420, n48227, n49430 );
nand U96761 ( n16309, n15045, n16321 );
not U96762 ( n7849, n47941 );
nand U96763 ( n16677, n15045, n18711 );
not U96764 ( n3038, n29169 );
not U96765 ( n3882, n21856 );
not U96766 ( n5639, n62891 );
not U96767 ( n6514, n54947 );
buf U96768 ( n76042, n76926 );
not U96769 ( n3453, n35589 );
not U96770 ( n6068, n70317 );
not U96771 ( n4290, n28408 );
not U96772 ( n6923, n61717 );
not U96773 ( n5194, n14735 );
nand U96774 ( n16237, n16217, n5210 );
not U96775 ( n5197, n16212 );
not U96776 ( n7852, n49240 );
nor U96777 ( n63824, n63825, n63826 );
nor U96778 ( n63825, n63827, n63828 );
nor U96779 ( n29868, n29869, n29870 );
nor U96780 ( n29869, n29871, n29872 );
nor U96781 ( n22545, n22546, n22547 );
nor U96782 ( n22546, n22548, n22549 );
nor U96783 ( n55658, n55659, n55660 );
nor U96784 ( n55659, n55661, n55662 );
not U96785 ( n4284, n26970 );
not U96786 ( n3447, n34215 );
not U96787 ( n6062, n68969 );
not U96788 ( n6917, n60110 );
nor U96789 ( n9178, n5283, n9145 );
nor U96790 ( n43154, n7938, n43128 );
not U96791 ( n1798, n49136 );
not U96792 ( n2915, n38408 );
nand U96793 ( n35363, n35347, n3458 );
nand U96794 ( n70095, n70079, n6073 );
nand U96795 ( n35516, n35347, n3460 );
nand U96796 ( n28288, n28112, n4298 );
nand U96797 ( n70244, n70079, n6075 );
nand U96798 ( n61510, n61267, n6930 );
nor U96799 ( n63885, n63887, n63888 );
nor U96800 ( n29929, n29931, n29932 );
nor U96801 ( n22606, n22608, n22609 );
nor U96802 ( n55719, n55721, n55722 );
nor U96803 ( n43186, n43188, n43189 );
nor U96804 ( n9218, n9220, n9222 );
nor U96805 ( n43205, n7939, n43188 );
nor U96806 ( n9242, n5284, n9220 );
not U96807 ( n2913, n38440 );
not U96808 ( n1795, n49373 );
nor U96809 ( n9282, n5284, n9283 );
nor U96810 ( n9283, n9284, n9285 );
nor U96811 ( n9284, n9287, n9288 );
nor U96812 ( n43251, n7939, n43252 );
nor U96813 ( n43252, n43253, n43254 );
nor U96814 ( n43253, n43255, n43256 );
or U96815 ( n48004, n47980, n7797 );
or U96816 ( n14795, n14759, n5142 );
nand U96817 ( n47930, n42382, n47945 );
nand U96818 ( n14710, n8294, n14729 );
not U96819 ( n1793, n54614 );
not U96820 ( n2910, n38476 );
nor U96821 ( n63937, n63938, n63939 );
nor U96822 ( n63938, n63940, n63941 );
nor U96823 ( n29981, n29982, n29983 );
nor U96824 ( n29982, n29984, n29985 );
nor U96825 ( n22658, n22659, n22660 );
nor U96826 ( n22659, n22661, n22662 );
nor U96827 ( n55771, n55772, n55773 );
nor U96828 ( n55772, n55774, n55775 );
nand U96829 ( n62918, n62987, n62988 );
nor U96830 ( n62988, n62989, n62990 );
nor U96831 ( n62987, n63003, n63004 );
nand U96832 ( n62989, n62997, n62998 );
nand U96833 ( n29200, n29220, n29221 );
nor U96834 ( n29221, n29222, n29223 );
nor U96835 ( n29220, n29236, n29237 );
nand U96836 ( n29222, n29230, n29231 );
nand U96837 ( n42409, n42452, n42453 );
nor U96838 ( n42453, n42454, n42455 );
nor U96839 ( n42452, n42468, n42469 );
nand U96840 ( n42454, n42462, n42463 );
nand U96841 ( n21883, n21903, n21904 );
nor U96842 ( n21904, n21905, n21906 );
nor U96843 ( n21903, n21919, n21920 );
nand U96844 ( n21905, n21913, n21914 );
nand U96845 ( n54974, n55015, n55016 );
nor U96846 ( n55016, n55017, n55018 );
nor U96847 ( n55015, n55031, n55032 );
nand U96848 ( n55017, n55025, n55026 );
nand U96849 ( n8328, n8353, n8354 );
nor U96850 ( n8354, n8355, n8357 );
nor U96851 ( n8353, n8373, n8374 );
nand U96852 ( n8355, n8365, n8367 );
nor U96853 ( n9320, n5285, n9287 );
nor U96854 ( n43282, n7940, n43255 );
not U96855 ( n7414, n42382 );
not U96856 ( n4770, n8294 );
not U96857 ( n1802, n54645 );
not U96858 ( n2919, n38508 );
xor U96859 ( n50009, n49742, n50081 );
xnor U96860 ( n50081, n49743, n49744 );
not U96861 ( n8230, n49940 );
xor U96862 ( n50025, n50079, n50018 );
xnor U96863 ( n50079, n50019, n50017 );
xnor U96864 ( n49661, n49695, n50041 );
xor U96865 ( n50041, n49694, n1278 );
nor U96866 ( n49868, n1738, n50250 );
xor U96867 ( n50168, n50169, n50170 );
xor U96868 ( n50120, n50121, n50122 );
xor U96869 ( n50144, n50145, n50146 );
nor U96870 ( n50304, n50537, n50534 );
nor U96871 ( n50275, n50276, n50273 );
nor U96872 ( n50276, n50277, n49891 );
nor U96873 ( n50277, n1755, n49887 );
nand U96874 ( n49670, n49671, n76476 );
nand U96875 ( n49671, n49672, n49673 );
xor U96876 ( n49672, n49674, n49675 );
nand U96877 ( n49674, n49676, n49677 );
nand U96878 ( n49677, n49661, n49678 );
nand U96879 ( n49678, n1210, n49679 );
nor U96880 ( n15161, n48772, n48773 );
nor U96881 ( n48772, n7832, n48774 );
nand U96882 ( n48774, n48775, n48776 );
nor U96883 ( n15001, n49155, n49156 );
nor U96884 ( n49155, n49158, n49157 );
nand U96885 ( n49157, n49159, n49160 );
nor U96886 ( n15201, n48695, n48696 );
nor U96887 ( n48695, n7835, n48697 );
not U96888 ( n7835, n48629 );
nor U96889 ( n15361, n48302, n48303 );
nor U96890 ( n48302, n48248, n48304 );
nand U96891 ( n48304, n48305, n48306 );
nor U96892 ( n15241, n48601, n48602 );
nor U96893 ( n48601, n7837, n48603 );
not U96894 ( n7837, n48535 );
nor U96895 ( n15281, n48504, n48505 );
nor U96896 ( n48504, n48427, n48506 );
nand U96897 ( n48506, n48507, n48508 );
nor U96898 ( n15441, n48114, n48115 );
nor U96899 ( n48114, n48025, n48117 );
nand U96900 ( n48117, n48118, n48119 );
nor U96901 ( n15401, n48219, n48220 );
nor U96902 ( n48219, n48150, n48221 );
nand U96903 ( n48221, n48222, n48223 );
nor U96904 ( n15041, n49061, n49062 );
nor U96905 ( n49061, n7825, n49063 );
not U96906 ( n7825, n48995 );
nor U96907 ( n14961, n49233, n49234 );
nor U96908 ( n49233, n7828, n49235 );
not U96909 ( n7828, n49184 );
nor U96910 ( n15121, n48864, n48865 );
nor U96911 ( n48864, n7829, n48866 );
not U96912 ( n7829, n48815 );
nor U96913 ( n15081, n48966, n48967 );
nor U96914 ( n48966, n7830, n48968 );
not U96915 ( n7830, n48896 );
nor U96916 ( n15321, n48399, n48400 );
nor U96917 ( n48399, n48345, n48401 );
nand U96918 ( n48401, n48402, n48403 );
nor U96919 ( n14921, n49330, n49331 );
nor U96920 ( n49330, n7827, n49332 );
not U96921 ( n7827, n49280 );
nor U96922 ( n14881, n49423, n49424 );
nor U96923 ( n49423, n7824, n49425 );
not U96924 ( n7824, n49358 );
nor U96925 ( n14841, n49663, n49664 );
nor U96926 ( n49663, n7823, n49665 );
not U96927 ( n7823, n49462 );
or U96928 ( n49963, n50218, n50217 );
and U96929 ( n75778, n76653, n54061 );
not U96930 ( n76930, n76927 );
xor U96931 ( n50216, n50217, n50218 );
or U96932 ( n49983, n50122, n50121 );
nand U96933 ( n49985, n50121, n50122 );
nand U96934 ( n49980, n50145, n50146 );
nand U96935 ( n49812, n50169, n50170 );
nand U96936 ( n49965, n50217, n50218 );
or U96937 ( n49810, n50170, n50169 );
or U96938 ( n49978, n50146, n50145 );
nor U96939 ( n49669, n49681, n49673 );
xor U96940 ( n49681, n49683, n49675 );
nand U96941 ( n49683, n49676, n50039 );
nand U96942 ( n50039, n50040, n49661 );
nand U96943 ( n50293, n50531, n50532 );
nand U96944 ( n50532, n50533, n50303 );
nand U96945 ( n50531, n50536, n50301 );
xor U96946 ( n50533, n50534, n50535 );
xor U96947 ( n49690, n49696, n49697 );
nand U96948 ( n49696, n49707, n49708 );
xor U96949 ( n49697, n49698, n49699 );
nand U96950 ( n49708, n49709, n49710 );
nand U96951 ( n50301, n50534, n50537 );
nand U96952 ( n48501, n49451, n43796 );
nand U96953 ( n15286, n48495, n48496 );
nor U96954 ( n48495, n48502, n48503 );
nor U96955 ( n48496, n48497, n48498 );
nor U96956 ( n48502, n48113, n48433 );
nand U96957 ( n15326, n48391, n48392 );
nor U96958 ( n48391, n48397, n48398 );
nor U96959 ( n48392, n48393, n48394 );
nor U96960 ( n48397, n48109, n48350 );
nand U96961 ( n15406, n48211, n48212 );
nor U96962 ( n48211, n48217, n48218 );
nor U96963 ( n48212, n48213, n48214 );
nor U96964 ( n48217, n48109, n48155 );
nand U96965 ( n15366, n48294, n48295 );
nor U96966 ( n48294, n48300, n48301 );
nor U96967 ( n48295, n48296, n48297 );
nor U96968 ( n48300, n48109, n48253 );
nand U96969 ( n15446, n48103, n48104 );
nor U96970 ( n48103, n48110, n48111 );
nor U96971 ( n48104, n48105, n48106 );
nor U96972 ( n48110, n48032, n48113 );
nor U96973 ( n49886, n49887, n1749 );
nor U96974 ( n50790, n50789, n50788 );
nand U96975 ( n50292, n1758, n50528 );
nand U96976 ( n50528, n50529, n50530 );
nand U96977 ( n50525, n50785, n50786 );
nand U96978 ( n50786, n50787, n50530 );
nand U96979 ( n50785, n50529, n50791 );
nor U96980 ( n50787, n50529, n50790 );
nand U96981 ( n50791, n1758, n50792 );
nand U96982 ( n50792, n50793, n50789 );
xor U96983 ( n17064, n2608, n17131 );
xor U96984 ( n17131, n16779, n17056 );
xnor U96985 ( n17071, n17130, n17064 );
xnor U96986 ( n17130, n17065, n17063 );
xnor U96987 ( n16693, n16739, n17087 );
xor U96988 ( n17087, n16738, n2393 );
and U96989 ( n75779, n76654, n17374 );
nor U96990 ( n16913, n2855, n17304 );
xor U96991 ( n17246, n17247, n17248 );
xor U96992 ( n17222, n17223, n17224 );
xor U96993 ( n17174, n17175, n17176 );
xor U96994 ( n17198, n17199, n17200 );
nor U96995 ( n17358, n17578, n17576 );
or U96996 ( n17008, n17272, n17271 );
or U96997 ( n16958, n17341, n17340 );
nand U96998 ( n8551, n15360, n15362 );
nor U96999 ( n15360, n15369, n15370 );
nor U97000 ( n15362, n15363, n15364 );
nor U97001 ( n15369, n14914, n15297 );
nand U97002 ( n8591, n15245, n15247 );
nor U97003 ( n15245, n15253, n15254 );
nor U97004 ( n15247, n15248, n15249 );
nor U97005 ( n15253, n14909, n15185 );
nand U97006 ( n8631, n15135, n15137 );
nor U97007 ( n15135, n15143, n15144 );
nor U97008 ( n15137, n15138, n15139 );
nor U97009 ( n15143, n14909, n15078 );
nand U97010 ( n8671, n15025, n15027 );
nor U97011 ( n15025, n15033, n15034 );
nor U97012 ( n15027, n15028, n15029 );
nor U97013 ( n15033, n14909, n14974 );
nand U97014 ( n50530, n50788, n50789 );
nand U97015 ( n8711, n14902, n14903 );
nor U97016 ( n14902, n14910, n14912 );
nor U97017 ( n14903, n14904, n14905 );
nor U97018 ( n14910, n14830, n14914 );
nand U97019 ( n16713, n16714, n76613 );
nand U97020 ( n16714, n16715, n16717 );
xor U97021 ( n16715, n16718, n16719 );
nand U97022 ( n16718, n16720, n16721 );
nand U97023 ( n16721, n16693, n16722 );
nand U97024 ( n16722, n2353, n16723 );
nor U97025 ( n8586, n15255, n15257 );
nor U97026 ( n15255, n15179, n15258 );
nand U97027 ( n15258, n15259, n15260 );
nor U97028 ( n8626, n15145, n15147 );
nor U97029 ( n15145, n15072, n15148 );
nand U97030 ( n15148, n15149, n15150 );
nor U97031 ( n8666, n15035, n15037 );
nor U97032 ( n15035, n14968, n15038 );
nand U97033 ( n15038, n15039, n15040 );
nor U97034 ( n8706, n14924, n14925 );
nor U97035 ( n14924, n14822, n14928 );
nand U97036 ( n14928, n14929, n14930 );
nor U97037 ( n8266, n16102, n16103 );
nor U97038 ( n16102, n5175, n16104 );
not U97039 ( n5175, n16039 );
nor U97040 ( n8306, n16003, n16004 );
nor U97041 ( n16003, n5170, n16005 );
not U97042 ( n5170, n15932 );
nor U97043 ( n8346, n15895, n15897 );
nor U97044 ( n15895, n5177, n15898 );
not U97045 ( n5177, n15827 );
nor U97046 ( n8386, n15787, n15788 );
nor U97047 ( n15787, n5174, n15789 );
not U97048 ( n5174, n15717 );
nor U97049 ( n8226, n16203, n16204 );
nor U97050 ( n16203, n5173, n16205 );
not U97051 ( n5173, n16135 );
nor U97052 ( n8546, n15372, n15373 );
nor U97053 ( n15372, n15289, n15374 );
nand U97054 ( n15374, n15375, n15377 );
nor U97055 ( n8466, n15580, n15582 );
nor U97056 ( n15580, n5180, n15583 );
not U97057 ( n5180, n15518 );
nor U97058 ( n8506, n15483, n15484 );
nor U97059 ( n15483, n5182, n15485 );
not U97060 ( n5182, n15412 );
nor U97061 ( n8186, n16313, n16314 );
nor U97062 ( n16313, n5172, n16315 );
not U97063 ( n5172, n16242 );
nor U97064 ( n8146, n16415, n16417 );
nor U97065 ( n16415, n5169, n16418 );
not U97066 ( n5169, n16347 );
nor U97067 ( n8106, n16704, n16705 );
nor U97068 ( n16704, n18701, n16707 );
nand U97069 ( n16707, n18702, n18703 );
xor U97070 ( n17270, n17271, n17272 );
or U97071 ( n17029, n17176, n17175 );
nand U97072 ( n15166, n48763, n48764 );
nor U97073 ( n48763, n48770, n48771 );
nor U97074 ( n48764, n48765, n48766 );
nor U97075 ( n48770, n47941, n48109 );
xor U97076 ( n17339, n17340, n17341 );
nand U97077 ( n16857, n17223, n17224 );
nand U97078 ( n17031, n17175, n17176 );
nand U97079 ( n17026, n17199, n17200 );
nand U97080 ( n17022, n17247, n17248 );
nand U97081 ( n17010, n17271, n17272 );
nor U97082 ( n16712, n16725, n16717 );
xor U97083 ( n16725, n16727, n16719 );
nand U97084 ( n16727, n16720, n17085 );
nand U97085 ( n17085, n17086, n16693 );
nand U97086 ( n14926, n49321, n49322 );
nor U97087 ( n49322, n49323, n49324 );
nor U97088 ( n49321, n49328, n49329 );
nor U97089 ( n49323, n48109, n49276 );
nand U97090 ( n14886, n49414, n49415 );
nor U97091 ( n49415, n49416, n49417 );
nor U97092 ( n49414, n49421, n49422 );
nor U97093 ( n49416, n48109, n49354 );
nand U97094 ( n15006, n49146, n49147 );
nor U97095 ( n49147, n49148, n49149 );
nor U97096 ( n49146, n49153, n49154 );
nor U97097 ( n49148, n48109, n49086 );
nand U97098 ( n15046, n49052, n49053 );
nor U97099 ( n49053, n49054, n49055 );
nor U97100 ( n49052, n49059, n49060 );
nor U97101 ( n49054, n48109, n48991 );
nand U97102 ( n15086, n48957, n48958 );
nor U97103 ( n48958, n48959, n48960 );
nor U97104 ( n48957, n48964, n48965 );
nor U97105 ( n48959, n48109, n48892 );
nand U97106 ( n15206, n48686, n48687 );
nor U97107 ( n48687, n48688, n48689 );
nor U97108 ( n48686, n48693, n48694 );
nor U97109 ( n48688, n48109, n48625 );
nand U97110 ( n15246, n48592, n48593 );
nor U97111 ( n48593, n48594, n48595 );
nor U97112 ( n48592, n48599, n48600 );
nor U97113 ( n48594, n48109, n48531 );
nand U97114 ( n14966, n49225, n49226 );
nor U97115 ( n49226, n49227, n49228 );
nor U97116 ( n49225, n49231, n49232 );
nand U97117 ( n49228, n49229, n49230 );
nand U97118 ( n15126, n48856, n48857 );
nor U97119 ( n48857, n48858, n48859 );
nor U97120 ( n48856, n48862, n48863 );
nand U97121 ( n48859, n48860, n48861 );
or U97122 ( n16855, n17224, n17223 );
or U97123 ( n17024, n17200, n17199 );
or U97124 ( n17020, n17248, n17247 );
nand U97125 ( n16961, n17341, n17340 );
nor U97126 ( n50803, n51053, n51050 );
nand U97127 ( n50526, n50800, n50801 );
nand U97128 ( n50801, n50802, n1750 );
not U97129 ( n1750, n50803 );
nand U97130 ( n17347, n17572, n17573 );
nand U97131 ( n17573, n17574, n17357 );
nand U97132 ( n17572, n17577, n17355 );
xor U97133 ( n17574, n17575, n17576 );
nor U97134 ( n15683, n15679, n15685 );
nand U97135 ( n15685, n15687, n15688 );
nand U97136 ( n17355, n17576, n17578 );
nor U97137 ( n50307, n73402, n49923 );
not U97138 ( n8232, n54061 );
nand U97139 ( n8431, n15670, n15672 );
nor U97140 ( n15670, n15680, n15682 );
nor U97141 ( n15672, n15673, n15674 );
nor U97142 ( n15680, n14735, n14909 );
nand U97143 ( n8151, n16404, n16405 );
nor U97144 ( n16405, n16407, n16408 );
nor U97145 ( n16404, n16413, n16414 );
nor U97146 ( n16407, n14909, n16342 );
nand U97147 ( n8191, n16302, n16303 );
nor U97148 ( n16303, n16304, n16305 );
nor U97149 ( n16302, n16310, n16312 );
nor U97150 ( n16304, n14909, n16237 );
nand U97151 ( n8271, n16090, n16092 );
nor U97152 ( n16092, n16093, n16094 );
nor U97153 ( n16090, n16099, n16100 );
nor U97154 ( n16093, n14909, n16034 );
nand U97155 ( n8311, n15983, n15984 );
nor U97156 ( n15984, n15985, n15987 );
nor U97157 ( n15983, n15992, n15993 );
nor U97158 ( n15985, n14909, n15927 );
nand U97159 ( n8351, n15884, n15885 );
nor U97160 ( n15885, n15887, n15888 );
nor U97161 ( n15884, n15893, n15894 );
nor U97162 ( n15887, n14909, n15822 );
nand U97163 ( n8471, n15569, n15570 );
nor U97164 ( n15570, n15572, n15573 );
nor U97165 ( n15569, n15578, n15579 );
nor U97166 ( n15572, n14909, n15513 );
nand U97167 ( n8511, n15463, n15464 );
nor U97168 ( n15464, n15465, n15467 );
nor U97169 ( n15463, n15472, n15473 );
nor U97170 ( n15465, n14909, n15407 );
nand U97171 ( n8391, n15777, n15778 );
nor U97172 ( n15778, n15779, n15780 );
nor U97173 ( n15777, n15784, n15785 );
nand U97174 ( n15780, n15782, n15783 );
nand U97175 ( n8231, n16193, n16194 );
nor U97176 ( n16194, n16195, n16197 );
nor U97177 ( n16193, n16200, n16202 );
nand U97178 ( n16197, n16198, n16199 );
xor U97179 ( n16734, n16740, n16741 );
nand U97180 ( n16740, n16751, n16752 );
xor U97181 ( n16741, n16742, n16743 );
nand U97182 ( n16752, n16753, n16754 );
and U97183 ( n43795, n43796, n43797 );
nand U97184 ( n16316, n43732, n43733 );
nor U97185 ( n43733, n43734, n43735 );
nor U97186 ( n43732, n43794, n43795 );
nor U97187 ( n43734, n43391, n76362 );
nand U97188 ( n17335, n17563, n17562 );
or U97189 ( n17333, n17562, n17563 );
nand U97190 ( n50800, n51050, n51053 );
nor U97191 ( n17845, n17844, n17843 );
nand U97192 ( n17346, n2873, n17584 );
nand U97193 ( n17584, n17585, n17586 );
nand U97194 ( n17569, n17840, n17841 );
nand U97195 ( n17841, n17842, n17586 );
nand U97196 ( n17840, n17585, n17846 );
nor U97197 ( n17842, n17585, n17845 );
nand U97198 ( n17846, n2873, n17847 );
nand U97199 ( n17847, n17848, n17844 );
xor U97200 ( n20774, n20785, n20734 );
nand U97201 ( n20785, n20735, n20732 );
xnor U97202 ( n20704, n20771, n20721 );
xnor U97203 ( n20771, n20719, n20720 );
xor U97204 ( n19845, n19965, n20098 );
xor U97205 ( n20098, n19964, n19966 );
xnor U97206 ( n20108, n20423, n20424 );
nor U97207 ( n20424, n73418, n20425 );
nand U97208 ( n20425, n20426, n2614 );
not U97209 ( n2614, n20427 );
nor U97210 ( n17964, n18189, n18188 );
nor U97211 ( n20628, n20693, n2688 );
nor U97212 ( n18927, n17028, n2524 );
nand U97213 ( n18905, n18910, n18911 );
or U97214 ( n18910, n18915, n18914 );
nand U97215 ( n18911, n18912, n18913 );
nand U97216 ( n18912, n18914, n18915 );
nor U97217 ( n17696, n17910, n18152 );
and U97218 ( n18152, n18153, n17911 );
nand U97219 ( n18153, n17917, n17915 );
nand U97220 ( n18925, n19393, n19394 );
nand U97221 ( n19393, n19398, n19397 );
nand U97222 ( n19394, n19395, n19396 );
or U97223 ( n19395, n19397, n19398 );
nand U97224 ( n18182, n18199, n8218 );
nor U97225 ( n18199, n2485, n73022 );
nand U97226 ( n17690, n17692, n17693 );
or U97227 ( n17692, n17697, n17696 );
nand U97228 ( n17693, n17694, n17695 );
nand U97229 ( n17694, n17696, n17697 );
nor U97230 ( n18191, n18192, n17962 );
nor U97231 ( n18192, n18193, n17964 );
and U97232 ( n18193, n18189, n18188 );
nand U97233 ( n20732, n20787, n20788 );
nand U97234 ( n16724, n17398, n17399 );
nand U97235 ( n17398, n16655, n16659 );
nand U97236 ( n17399, n16658, n17400 );
or U97237 ( n17400, n16659, n16655 );
nand U97238 ( n20101, n20102, n20103 );
or U97239 ( n20102, n20088, n20085 );
nand U97240 ( n20103, n20087, n20104 );
nand U97241 ( n20104, n20085, n20088 );
nor U97242 ( n17628, n17634, n17635 );
nor U97243 ( n17634, n2392, n17636 );
nand U97244 ( n17636, n17076, n17077 );
nand U97245 ( n20793, n76589, n20794 );
nand U97246 ( n20794, n76655, n75911 );
nor U97247 ( n17910, n17917, n17915 );
nor U97248 ( n49951, n50250, n1729 );
nand U97249 ( n17680, n17907, n8212 );
nor U97250 ( n17907, n2397, n73422 );
or U97251 ( n20735, n20788, n20787 );
nor U97252 ( n20752, n20779, n20774 );
nand U97253 ( n17586, n17843, n17844 );
xor U97254 ( n20887, n20898, n20783 );
nand U97255 ( n20898, n20784, n20781 );
nor U97256 ( n20518, n20525, n2667 );
nand U97257 ( n20781, n20899, n20900 );
nand U97258 ( n20705, n20765, n20766 );
nand U97259 ( n20766, n20767, n20768 );
nand U97260 ( n20905, n76589, n20906 );
nand U97261 ( n20906, n76654, n73404 );
nor U97262 ( n53278, n73017, n53279 );
nand U97263 ( n53279, n53280, n1490 );
not U97264 ( n1490, n53281 );
nor U97265 ( n53070, n53072, n53064 );
nor U97266 ( n50922, n51145, n51144 );
nor U97267 ( n53379, n53381, n53382 );
and U97268 ( n53381, n53383, n1518 );
xor U97269 ( n53613, n53674, n53675 );
nand U97270 ( n53674, n53676, n53677 );
nor U97271 ( n50863, n1282, n73425 );
nor U97272 ( n53382, n53383, n1518 );
nor U97273 ( n53496, n53499, n1567 );
nand U97274 ( n52797, n52925, n52926 );
or U97275 ( n52925, n52787, n52790 );
nand U97276 ( n52926, n52927, n52789 );
nand U97277 ( n52927, n52790, n52787 );
nor U97278 ( n51883, n49982, n1404 );
nand U97279 ( n51881, n52508, n52509 );
nand U97280 ( n52508, n52513, n52512 );
nand U97281 ( n52509, n52510, n52511 );
or U97282 ( n52510, n52512, n52513 );
nand U97283 ( n51138, n51155, n8235 );
nor U97284 ( n51155, n1369, n73424 );
nor U97285 ( n51147, n51148, n50920 );
nor U97286 ( n51148, n51149, n50922 );
nand U97287 ( n51861, n51866, n51867 );
or U97288 ( n51866, n51871, n51870 );
nand U97289 ( n51867, n51868, n51869 );
nand U97290 ( n51868, n51870, n51871 );
nor U97291 ( n50040, n50342, n50343 );
nor U97292 ( n50342, n49633, n50345 );
nor U97293 ( n50345, n50346, n1212 );
nand U97294 ( n53732, n76323, n53733 );
nand U97295 ( n53733, n76652, n73400 );
or U97296 ( n53676, n53725, n53726 );
nor U97297 ( n51117, n1368, n51122 );
nand U97298 ( n50906, n51113, n8239 );
nor U97299 ( n51113, n1325, n73426 );
xor U97300 ( n52650, n52787, n52788 );
xor U97301 ( n52788, n52789, n52790 );
xor U97302 ( n52181, n52330, n52331 );
xor U97303 ( n52331, n52332, n52333 );
xor U97304 ( n51827, n52187, n52188 );
xor U97305 ( n52188, n52189, n52190 );
nand U97306 ( n49501, n50613, n50614 );
nand U97307 ( n50613, n49466, n49469 );
nand U97308 ( n50614, n49468, n50615 );
or U97309 ( n50615, n49469, n49466 );
xnor U97310 ( n20884, n20769, n20768 );
nor U97311 ( n20524, n20525, n2640 );
or U97312 ( n20784, n20900, n20899 );
nor U97313 ( n17086, n17387, n17388 );
nor U97314 ( n17387, n16658, n17390 );
nor U97315 ( n17390, n17391, n2354 );
xor U97316 ( n20097, n20217, n20218 );
xor U97317 ( n20218, n20219, n20220 );
nand U97318 ( n19841, n19969, n19970 );
or U97319 ( n19969, n19831, n19834 );
nand U97320 ( n19970, n19971, n19833 );
nand U97321 ( n19971, n19834, n19831 );
nor U97322 ( n53687, n53689, n53681 );
xor U97323 ( n53681, n53734, n53735 );
nand U97324 ( n53734, n53736, n53737 );
nor U97325 ( n53438, n53441, n1564 );
nor U97326 ( n53552, n53559, n1587 );
nand U97327 ( n53737, n53768, n53767 );
nand U97328 ( n53773, n76323, n53774 );
nand U97329 ( n53774, n76652, n72999 );
nor U97330 ( n20521, n20523, n20524 );
and U97331 ( n20523, n20525, n2640 );
nand U97332 ( n49680, n50354, n50355 );
nand U97333 ( n50355, n49633, n50356 );
nand U97334 ( n17570, n17836, n17837 );
nand U97335 ( n17837, n17838, n2867 );
not U97336 ( n2867, n17839 );
nor U97337 ( n17839, n18099, n18097 );
xor U97338 ( n49709, n49720, n49721 );
xor U97339 ( n49721, n49722, n49723 );
xor U97340 ( n49720, n50026, n50027 );
xor U97341 ( n49723, n49724, n49725 );
xor U97342 ( n50026, n50032, n50033 );
nor U97343 ( n50033, n73424, n50034 );
nand U97344 ( n50032, n50035, n50036 );
nand U97345 ( n50036, n50037, n50038 );
nand U97346 ( n17949, n18156, n8213 );
nor U97347 ( n18156, n2443, n73423 );
or U97348 ( n53736, n53767, n53768 );
xor U97349 ( n51899, n52382, n52032 );
xor U97350 ( n52382, n52034, n52035 );
nor U97351 ( n52395, n50320, n1538 );
nand U97352 ( n53790, n53853, n53854 );
nand U97353 ( n53853, n53857, n53859 );
nand U97354 ( n53854, n53855, n53856 );
nand U97355 ( n53859, n1654, n53860 );
nor U97356 ( n53858, n53862, n53865 );
nand U97357 ( n53571, n53638, n53639 );
nand U97358 ( n53639, n53640, n1584 );
nor U97359 ( n53638, n53642, n53643 );
not U97360 ( n1584, n53641 );
nand U97361 ( n53753, n53784, n53785 );
nand U97362 ( n53785, n53786, n1633 );
nor U97363 ( n53784, n53788, n53789 );
not U97364 ( n1633, n53787 );
nor U97365 ( n53788, n53792, n53793 );
nor U97366 ( n53792, n72999, n49898 );
xor U97367 ( n53793, n53787, n53790 );
nor U97368 ( n53642, n53646, n53647 );
nor U97369 ( n53646, n73410, n50496 );
xor U97370 ( n53647, n53641, n53644 );
nand U97371 ( n52911, n53504, n53503 );
nand U97372 ( n51531, n51885, n51886 );
or U97373 ( n51885, n51890, n51889 );
nand U97374 ( n51886, n51887, n51888 );
nand U97375 ( n51887, n51889, n51890 );
nor U97376 ( n53855, n53857, n53858 );
nor U97377 ( n18160, n2484, n18165 );
and U97378 ( n17957, n17902, n75780 );
xnor U97379 ( n75780, n17900, n17901 );
nand U97380 ( n17695, n17954, n17955 );
nand U97381 ( n17955, n17897, n17900 );
nor U97382 ( n17954, n17956, n17957 );
nor U97383 ( n17956, n17902, n17959 );
xor U97384 ( n53054, n52920, n52922 );
nor U97385 ( n53543, n53545, n53537 );
nor U97386 ( n50651, n50866, n51109 );
nand U97387 ( n51110, n50873, n50871 );
nand U97388 ( n50645, n50647, n50648 );
or U97389 ( n50647, n50652, n50651 );
nand U97390 ( n50648, n50649, n50650 );
nand U97391 ( n50649, n50651, n50652 );
nand U97392 ( n53609, n53667, n53666 );
nor U97393 ( n50585, n50589, n50590 );
nor U97394 ( n50589, n1277, n50591 );
nand U97395 ( n50591, n50030, n50031 );
xor U97396 ( n53537, n53606, n53607 );
nand U97397 ( n53606, n53608, n53609 );
nand U97398 ( n53672, n76323, n53673 );
nand U97399 ( n53673, n76652, n73003 );
nand U97400 ( n53393, n1513, n53407 );
not U97401 ( n1513, n53396 );
nor U97402 ( n49925, n49922, n1764 );
not U97403 ( n1767, n50311 );
nor U97404 ( n50866, n50873, n50871 );
xnor U97405 ( n19718, n20085, n20086 );
xnor U97406 ( n20086, n20087, n20088 );
nand U97407 ( n53677, n53726, n53725 );
xnor U97408 ( n20641, n20722, n20686 );
xnor U97409 ( n20722, n20685, n20684 );
nand U97410 ( n18194, n18189, n2442 );
nor U97411 ( n50303, n49923, n73010 );
and U97412 ( n49676, n50352, n50353 );
nand U97413 ( n50352, n49682, n76835 );
nand U97414 ( n50353, n1214, n49680 );
nor U97415 ( n51524, n51514, n51527 );
or U97416 ( n51527, n1459, n51512 );
xor U97417 ( n20082, n20213, n20214 );
xor U97418 ( n20214, n20215, n20216 );
nor U97419 ( n20081, n20084, n2588 );
nor U97420 ( n53558, n53559, n1565 );
nor U97421 ( n53376, n53383, n1544 );
nor U97422 ( n53555, n53557, n53558 );
and U97423 ( n53557, n53559, n1565 );
nand U97424 ( n19245, n19701, n19702 );
or U97425 ( n19701, n19696, n19699 );
nand U97426 ( n19702, n19703, n19698 );
nand U97427 ( n19703, n19699, n19696 );
xor U97428 ( n53038, n53169, n53170 );
xor U97429 ( n53170, n53171, n53172 );
nor U97430 ( n53037, n53040, n1465 );
or U97431 ( n52909, n53503, n53504 );
nand U97432 ( n51150, n51145, n1324 );
nand U97433 ( n53498, n53499, n53494 );
or U97434 ( n53608, n53666, n53667 );
nand U97435 ( n20725, n20736, n20737 );
nand U97436 ( n20736, n20740, n20676 );
nand U97437 ( n20737, n2774, n20738 );
nand U97438 ( n20740, n20673, n20675 );
nand U97439 ( n20745, n76589, n20746 );
nand U97440 ( n20746, n76655, n73406 );
not U97441 ( n2774, n20676 );
xor U97442 ( n20875, n20919, n20896 );
nand U97443 ( n20919, n20897, n20894 );
nor U97444 ( n20881, n20883, n20875 );
nand U97445 ( n20894, n20920, n20921 );
nand U97446 ( n20926, n76589, n20927 );
nand U97447 ( n20927, n76654, n73009 );
nand U97448 ( n19714, n19974, n19975 );
nand U97449 ( n19974, n19830, n19827 );
nand U97450 ( n19975, n19829, n19976 );
or U97451 ( n19976, n19827, n19830 );
nand U97452 ( n52360, n52657, n52658 );
or U97453 ( n52657, n52652, n52655 );
nand U97454 ( n52658, n52659, n52654 );
nand U97455 ( n52659, n52655, n52652 );
xor U97456 ( n17561, n17562, n17563 );
xor U97457 ( n52344, n52652, n52653 );
xor U97458 ( n52653, n52654, n52655 );
or U97459 ( n51653, n51875, n51876 );
nand U97460 ( n20642, n20716, n20717 );
or U97461 ( n20716, n20721, n20720 );
nand U97462 ( n20717, n20718, n20719 );
nand U97463 ( n20718, n20720, n20721 );
nand U97464 ( n50635, n50874, n50875 );
or U97465 ( n50874, n50626, n50629 );
nand U97466 ( n50875, n50628, n50876 );
nand U97467 ( n50876, n50629, n50626 );
nor U97468 ( n50885, n50625, n50888 );
nor U97469 ( n50888, n50882, n50889 );
nand U97470 ( n50889, n50879, n50624 );
and U97471 ( n50629, n50877, n50878 );
nand U97472 ( n50878, n1250, n50623 );
nand U97473 ( n50877, n50885, n50886 );
not U97474 ( n1250, n50624 );
nand U97475 ( n20510, n20811, n20812 );
or U97476 ( n20811, n20499, n20496 );
nand U97477 ( n20812, n20498, n20813 );
nand U97478 ( n20813, n20496, n20499 );
nor U97479 ( n20407, n20408, n2617 );
nor U97480 ( n20821, n20822, n2670 );
nand U97481 ( n20825, n20841, n20859 );
nand U97482 ( n20859, n20839, n20840 );
nor U97483 ( n20403, n20404, n20405 );
nor U97484 ( n20404, n20406, n20407 );
and U97485 ( n20406, n20408, n2617 );
nor U97486 ( n20818, n20819, n2690 );
nor U97487 ( n20819, n20820, n20821 );
and U97488 ( n20820, n20822, n2670 );
nand U97489 ( n20866, n76589, n20867 );
nand U97490 ( n20867, n76655, n73012 );
or U97491 ( n20840, n20860, n20861 );
xor U97492 ( n51874, n51875, n51876 );
nand U97493 ( n52185, n52204, n52205 );
or U97494 ( n52204, n52174, n52171 );
nand U97495 ( n52205, n52173, n52206 );
nand U97496 ( n52206, n52171, n52174 );
nand U97497 ( n51831, n52055, n52056 );
or U97498 ( n52055, n51819, n51818 );
nand U97499 ( n52056, n51820, n52057 );
nand U97500 ( n52057, n51818, n51819 );
xnor U97501 ( n17625, n17698, n17421 );
xor U97502 ( n17698, n17420, n17419 );
nor U97503 ( n17420, n17897, n17898 );
and U97504 ( n17898, n17899, n17900 );
nand U97505 ( n17899, n17901, n17902 );
nand U97506 ( n52340, n52517, n52518 );
or U97507 ( n52517, n52330, n52333 );
nand U97508 ( n52518, n52519, n52332 );
nand U97509 ( n52519, n52333, n52330 );
and U97510 ( n50915, n50857, n75781 );
xnor U97511 ( n75781, n50855, n50856 );
nand U97512 ( n50650, n50912, n50913 );
nand U97513 ( n50913, n50852, n50855 );
nor U97514 ( n50912, n50914, n50915 );
nor U97515 ( n50914, n50857, n50917 );
or U97516 ( n20897, n20921, n20920 );
nand U97517 ( n52913, n53399, n8238 );
nor U97518 ( n53399, n1534, n73413 );
nand U97519 ( n52493, n52913, n52914 );
nand U97520 ( n52914, n52915, n52916 );
nand U97521 ( n52915, n1534, n50320 );
nand U97522 ( n51655, n51876, n51875 );
nand U97523 ( n20112, n20329, n20330 );
or U97524 ( n20329, n20213, n20216 );
nand U97525 ( n20330, n20331, n20215 );
nand U97526 ( n20331, n20216, n20213 );
xor U97527 ( n19246, n19847, n19397 );
xor U97528 ( n19847, n19396, n19398 );
nand U97529 ( n20803, n20854, n20855 );
or U97530 ( n20854, n20843, n20844 );
nand U97531 ( n20855, n20856, n20845 );
nand U97532 ( n20856, n20844, n20843 );
xor U97533 ( n53502, n53503, n53504 );
xnor U97534 ( n50910, n50651, n50911 );
xor U97535 ( n50911, n50650, n50652 );
nand U97536 ( n50808, n51047, n51048 );
nand U97537 ( n51048, n51049, n50802 );
nand U97538 ( n51047, n51052, n50800 );
xor U97539 ( n51049, n51050, n51051 );
nor U97540 ( n51052, n50802, n50803 );
nand U97541 ( n52636, n1372, n52663 );
not U97542 ( n1372, n52639 );
xnor U97543 ( n51880, n52369, n51890 );
xnor U97544 ( n52369, n51888, n51889 );
xnor U97545 ( n20506, n20842, n20843 );
xnor U97546 ( n20842, n20844, n20845 );
nand U97547 ( n20694, n20693, n20627 );
and U97548 ( n9892, n9893, n9894 );
nand U97549 ( n9581, n9813, n9814 );
nor U97550 ( n9814, n9815, n9817 );
nor U97551 ( n9813, n9890, n9892 );
nor U97552 ( n9815, n9455, n76632 );
nand U97553 ( n50623, n50879, n50880 );
nand U97554 ( n50880, n50881, n50882 );
nand U97555 ( n50881, n50883, n50884 );
nand U97556 ( n52506, n52917, n52918 );
or U97557 ( n52917, n52922, n52921 );
nand U97558 ( n52918, n52919, n52920 );
nand U97559 ( n52919, n52921, n52922 );
xor U97560 ( n19694, n19831, n19832 );
xor U97561 ( n19832, n19833, n19834 );
nor U97562 ( n50632, n50331, n1249 );
xnor U97563 ( n20352, n20496, n20497 );
xnor U97564 ( n20497, n20498, n20499 );
nand U97565 ( n53068, n53183, n53184 );
or U97566 ( n53183, n53169, n53172 );
nand U97567 ( n53184, n53185, n53171 );
nand U97568 ( n53185, n53172, n53169 );
xor U97569 ( n18924, n18934, n19254 );
xor U97570 ( n19254, n18932, n18933 );
nand U97571 ( n19259, n19961, n19962 );
or U97572 ( n19961, n19966, n19965 );
nand U97573 ( n19962, n19963, n19964 );
nand U97574 ( n19963, n19965, n19966 );
nor U97575 ( n53630, n53633, n1601 );
nand U97576 ( n17836, n18097, n18099 );
nand U97577 ( n53741, n53775, n53776 );
nand U97578 ( n53775, n53781, n53780 );
nand U97579 ( n53776, n1644, n53777 );
nand U97580 ( n53781, n53782, n53783 );
nand U97581 ( n53849, n76323, n53850 );
nand U97582 ( n53850, n76652, n73397 );
not U97583 ( n1644, n53780 );
xor U97584 ( n52361, n52803, n52512 );
xor U97585 ( n52803, n52511, n52513 );
nand U97586 ( n50315, n1764, n49922 );
nand U97587 ( n52908, n53653, n53654 );
nand U97588 ( n53654, n53644, n53641 );
nor U97589 ( n53653, n53640, n1583 );
not U97590 ( n1583, n53645 );
or U97591 ( n52486, n52835, n52836 );
nand U97592 ( n20234, n2637, n20533 );
not U97593 ( n2637, n20534 );
nand U97594 ( n20841, n20861, n20860 );
nand U97595 ( n20751, n20781, n20782 );
nand U97596 ( n20782, n20783, n20784 );
xor U97597 ( n52834, n52835, n52836 );
xnor U97598 ( n17650, n17696, n17953 );
xor U97599 ( n17953, n17695, n17697 );
nand U97600 ( n53581, n1585, n53569 );
not U97601 ( n1585, n53567 );
and U97602 ( n53574, n53579, n53580 );
nand U97603 ( n53579, n53567, n1570 );
nand U97604 ( n53580, n53581, n53570 );
not U97605 ( n1570, n53569 );
nor U97606 ( n53261, n53262, n1493 );
nor U97607 ( n53257, n53258, n53259 );
nor U97608 ( n53258, n53260, n53261 );
and U97609 ( n53260, n53262, n1493 );
nand U97610 ( n20115, n20116, n20112 );
nand U97611 ( n20727, n20732, n20733 );
nand U97612 ( n20733, n20734, n20735 );
and U97613 ( n52394, n52827, n8238 );
nor U97614 ( n52827, n1557, n73412 );
xor U97615 ( n51123, n51172, n51173 );
xnor U97616 ( n51173, n51174, n51175 );
xor U97617 ( n51119, n51121, n1368 );
nand U97618 ( n52488, n52836, n52835 );
nand U97619 ( n20432, n20426, n20437 );
nand U97620 ( n20437, n20438, n20423 );
nor U97621 ( n20438, n20427, n73418 );
nor U97622 ( n51845, n51848, n1287 );
nand U97623 ( n52194, n52199, n52200 );
or U97624 ( n52199, n52187, n52190 );
nand U97625 ( n52200, n52189, n52201 );
nand U97626 ( n52201, n52190, n52187 );
xnor U97627 ( n50582, n50653, n50375 );
xor U97628 ( n50653, n50374, n50373 );
nor U97629 ( n50374, n50852, n50853 );
and U97630 ( n50853, n50854, n50855 );
nand U97631 ( n50854, n50856, n50857 );
nand U97632 ( n53856, n53865, n53862 );
nor U97633 ( n20470, n20476, n20477 );
xor U97634 ( n20477, n20838, n20839 );
nand U97635 ( n20838, n20840, n20841 );
nand U97636 ( n53465, n53483, n53521 );
nand U97637 ( n53521, n53481, n53482 );
nor U97638 ( n53202, n53209, n1522 );
nand U97639 ( n53604, n76323, n53605 );
nand U97640 ( n53605, n76652, n73410 );
nand U97641 ( n53528, n76323, n53529 );
nand U97642 ( n53529, n76652, n73008 );
nand U97643 ( n53541, n53533, n53596 );
nand U97644 ( n53596, n53531, n53532 );
or U97645 ( n53482, n53522, n53523 );
or U97646 ( n53532, n53597, n53598 );
nand U97647 ( n52321, n52521, n52522 );
nand U97648 ( n52521, n52317, n52315 );
nand U97649 ( n52522, n52316, n52523 );
or U97650 ( n52523, n52315, n52317 );
nor U97651 ( n52773, n52780, n1437 );
xor U97652 ( n20823, n20868, n20869 );
nand U97653 ( n20868, n20870, n20871 );
nand U97654 ( n20871, n20911, n20910 );
nand U97655 ( n20917, n76589, n20918 );
nand U97656 ( n20918, n76654, n75913 );
nand U97657 ( n19547, n19561, n19562 );
or U97658 ( n19561, n19538, n19539 );
nand U97659 ( n19562, n19563, n19540 );
nand U97660 ( n19563, n19539, n19538 );
nor U97661 ( n53333, n53334, n1523 );
nor U97662 ( n53208, n53209, n1495 );
nor U97663 ( n52779, n52780, n1409 );
nor U97664 ( n52957, n52964, n1470 );
nand U97665 ( n53337, n53353, n53470 );
nand U97666 ( n53470, n53351, n53352 );
nor U97667 ( n53330, n53331, n1548 );
nor U97668 ( n53331, n53332, n53333 );
and U97669 ( n53332, n53334, n1523 );
nor U97670 ( n53204, n53205, n53206 );
nor U97671 ( n53205, n53207, n53208 );
and U97672 ( n53207, n53209, n1495 );
nor U97673 ( n52775, n52776, n52777 );
nor U97674 ( n52776, n52778, n52779 );
and U97675 ( n52778, n52780, n1409 );
nand U97676 ( n53478, n76323, n53479 );
nand U97677 ( n53479, n76652, n73412 );
or U97678 ( n53352, n53471, n53472 );
nand U97679 ( n52380, n52809, n52808 );
nand U97680 ( n50905, n1283, n51124 );
nand U97681 ( n51124, n51125, n50893 );
not U97682 ( n1283, n50892 );
nand U97683 ( n51125, n50899, n50897 );
nor U97684 ( n51135, n51139, n51140 );
nor U97685 ( n51139, n73424, n50089 );
xor U97686 ( n51140, n51141, n51137 );
nor U97687 ( n50892, n50899, n50897 );
nand U97688 ( n53384, n53383, n53385 );
nand U97689 ( n53289, n53280, n53296 );
nand U97690 ( n53296, n53297, n53277 );
nor U97691 ( n53297, n53281, n73017 );
xnor U97692 ( n16657, n16658, n16659 );
nand U97693 ( n8556, n15349, n15350 );
nor U97694 ( n15349, n15358, n15359 );
nor U97695 ( n15350, n15352, n15353 );
nor U97696 ( n15358, n14900, n15297 );
nand U97697 ( n49724, n49726, n49727 );
nand U97698 ( n49726, n49735, n49736 );
nand U97699 ( n49727, n49728, n49729 );
xnor U97700 ( n49736, n49730, n49731 );
nand U97701 ( n8596, n15235, n15237 );
nor U97702 ( n15235, n15243, n15244 );
nor U97703 ( n15237, n15238, n15239 );
nor U97704 ( n15243, n14895, n15185 );
nand U97705 ( n8636, n15125, n15127 );
nor U97706 ( n15125, n15133, n15134 );
nor U97707 ( n15127, n15128, n15129 );
nor U97708 ( n15133, n14895, n15078 );
nand U97709 ( n8676, n15015, n15017 );
nor U97710 ( n15015, n15023, n15024 );
nor U97711 ( n15017, n15018, n15019 );
nor U97712 ( n15023, n14895, n14974 );
nand U97713 ( n20356, n20465, n20466 );
or U97714 ( n20465, n20394, n20391 );
nand U97715 ( n20466, n20393, n20467 );
nand U97716 ( n20467, n20391, n20394 );
nor U97717 ( n20475, n20476, n2645 );
nand U97718 ( n20479, n20495, n20828 );
nand U97719 ( n20828, n20493, n20494 );
nor U97720 ( n20472, n20473, n2672 );
nor U97721 ( n20473, n20474, n20475 );
and U97722 ( n20474, n20476, n2645 );
nand U97723 ( n20836, n76589, n20837 );
nand U97724 ( n20837, n76655, n73414 );
or U97725 ( n20494, n20829, n20830 );
xor U97726 ( n53335, n53480, n53481 );
nand U97727 ( n53480, n53482, n53483 );
nor U97728 ( n53328, n53334, n53335 );
nand U97729 ( n53483, n53523, n53522 );
xor U97730 ( n53566, n53567, n53568 );
xor U97731 ( n53568, n53569, n53570 );
nand U97732 ( n50619, n51676, n51677 );
nand U97733 ( n51676, n49653, n49654 );
nand U97734 ( n51677, n49655, n51678 );
or U97735 ( n51678, n49654, n49653 );
nor U97736 ( n51840, n1287, n51847 );
nand U97737 ( n51847, n51848, n51843 );
nand U97738 ( n53071, n53072, n53068 );
nand U97739 ( n8716, n14888, n14889 );
nor U97740 ( n14888, n14897, n14898 );
nor U97741 ( n14889, n14890, n14892 );
nor U97742 ( n14897, n14830, n14900 );
nor U97743 ( n16996, n17304, n2847 );
xor U97744 ( n49499, n50626, n50627 );
xor U97745 ( n50627, n50628, n50629 );
nand U97746 ( n53685, n53677, n53724 );
nand U97747 ( n53724, n53675, n53676 );
nand U97748 ( n20780, n20779, n20751 );
nand U97749 ( n20879, n20871, n20909 );
nand U97750 ( n20909, n20869, n20870 );
or U97751 ( n20870, n20910, n20911 );
xor U97752 ( n18166, n18216, n18217 );
xnor U97753 ( n18217, n18218, n18219 );
xor U97754 ( n18162, n18164, n2484 );
xor U97755 ( n53466, n53530, n53531 );
nand U97756 ( n53530, n53532, n53533 );
nand U97757 ( n53533, n53598, n53597 );
xor U97758 ( n19574, n19827, n19828 );
xor U97759 ( n19828, n19829, n19830 );
nand U97760 ( n19680, n2488, n19707 );
not U97761 ( n2488, n19683 );
nand U97762 ( n20526, n20525, n20527 );
xnor U97763 ( n52069, n52314, n52315 );
xnor U97764 ( n52314, n52316, n52317 );
xor U97765 ( n52807, n52808, n52809 );
nand U97766 ( n20797, n20894, n20895 );
nand U97767 ( n20895, n20896, n20897 );
nand U97768 ( n20893, n20892, n20797 );
nor U97769 ( n20401, n20408, n2642 );
or U97770 ( n52378, n52808, n52809 );
nand U97771 ( n17679, n17918, n17919 );
or U97772 ( n17918, n17670, n17673 );
nand U97773 ( n17919, n17672, n17920 );
nand U97774 ( n17920, n17673, n17670 );
nor U97775 ( n50310, n1764, n50311 );
nand U97776 ( n53560, n53559, n53561 );
xnor U97777 ( n18943, n19076, n19273 );
xnor U97778 ( n19273, n19079, n19078 );
nand U97779 ( n18575, n18929, n18930 );
or U97780 ( n18929, n18934, n18933 );
nand U97781 ( n18930, n18931, n18932 );
nand U97782 ( n18931, n18933, n18934 );
nand U97783 ( n19277, n19955, n19956 );
or U97784 ( n19955, n19960, n19959 );
nand U97785 ( n19956, n19957, n19958 );
nand U97786 ( n19957, n19959, n19960 );
xor U97787 ( n20564, n20575, n20651 );
xor U97788 ( n20651, n20573, n20574 );
xnor U97789 ( n19278, n19392, n19862 );
xor U97790 ( n19862, n19390, n19391 );
nor U97791 ( n19291, n17014, n2659 );
nor U97792 ( n20655, n20657, n20658 );
nor U97793 ( n20657, n16943, n75911 );
xor U97794 ( n20658, n20585, n20584 );
nand U97795 ( n20584, n20659, n20660 );
nand U97796 ( n20660, n20661, n20604 );
nand U97797 ( n20659, n20603, n20665 );
nor U97798 ( n20661, n20603, n20664 );
nor U97799 ( n20664, n20663, n20662 );
nand U97800 ( n20253, n20550, n20551 );
nand U97801 ( n20551, n20264, n2705 );
nor U97802 ( n20550, n20553, n20554 );
not U97803 ( n2705, n20263 );
nand U97804 ( n20574, n20652, n20653 );
nand U97805 ( n20653, n20586, n2757 );
nor U97806 ( n20652, n20655, n20656 );
not U97807 ( n2757, n20585 );
nor U97808 ( n20553, n20555, n20556 );
nor U97809 ( n20555, n16966, n75913 );
xor U97810 ( n20556, n20263, n20262 );
nand U97811 ( n19949, n20239, n20238 );
nand U97812 ( n20665, n2775, n20666 );
nand U97813 ( n20666, n20667, n20663 );
nand U97814 ( n53617, n53609, n53665 );
nand U97815 ( n53665, n53607, n53608 );
nand U97816 ( n53620, n53621, n53617 );
xnor U97817 ( n51811, n52171, n52172 );
xnor U97818 ( n52172, n52173, n52174 );
nor U97819 ( n19817, n19824, n2558 );
nand U97820 ( n53632, n53633, n53628 );
xor U97821 ( n19551, n19696, n19697 );
xor U97822 ( n19697, n19698, n19699 );
nand U97823 ( n53745, n53737, n53766 );
nand U97824 ( n53766, n53735, n53736 );
xor U97825 ( n51893, n51894, n51895 );
nand U97826 ( n51544, n52030, n52031 );
nand U97827 ( n52030, n52035, n52034 );
nand U97828 ( n52031, n52032, n52033 );
or U97829 ( n52033, n52034, n52035 );
xnor U97830 ( n49632, n49633, n49634 );
nand U97831 ( n15291, n48486, n48487 );
nor U97832 ( n48486, n48493, n48494 );
nor U97833 ( n48487, n48488, n48489 );
nor U97834 ( n48493, n48102, n48433 );
nand U97835 ( n15331, n48383, n48384 );
nor U97836 ( n48383, n48389, n48390 );
nor U97837 ( n48384, n48385, n48386 );
nor U97838 ( n48389, n48098, n48350 );
nand U97839 ( n15371, n48286, n48287 );
nor U97840 ( n48286, n48292, n48293 );
nor U97841 ( n48287, n48288, n48289 );
nor U97842 ( n48292, n48098, n48253 );
nand U97843 ( n15411, n48188, n48189 );
nor U97844 ( n48188, n48194, n48195 );
nor U97845 ( n48189, n48190, n48191 );
nor U97846 ( n48194, n48098, n48155 );
or U97847 ( n18697, n18919, n18920 );
xor U97848 ( n18871, n19231, n19232 );
xor U97849 ( n19232, n19233, n19234 );
xnor U97850 ( n19225, n19537, n19538 );
xnor U97851 ( n19537, n19539, n19540 );
nand U97852 ( n16512, n17657, n17658 );
nand U97853 ( n17657, n16468, n16472 );
nand U97854 ( n17658, n16470, n17659 );
or U97855 ( n17659, n16472, n16468 );
or U97856 ( n51649, n51894, n51895 );
nand U97857 ( n15451, n48092, n48093 );
nor U97858 ( n48092, n48099, n48100 );
nor U97859 ( n48093, n48094, n48095 );
nor U97860 ( n48099, n48032, n48102 );
nand U97861 ( n17321, n17587, n17588 );
nand U97862 ( n17587, n17592, n17591 );
nand U97863 ( n17588, n17589, n17590 );
or U97864 ( n17589, n17591, n17592 );
nand U97865 ( n53688, n53689, n53685 );
nor U97866 ( n50894, n50893, n50898 );
nand U97867 ( n50898, n1329, n50897 );
nand U97868 ( n53353, n53472, n53471 );
nand U97869 ( n53787, n53782, n53844 );
nand U97870 ( n53844, n53783, n53780 );
xor U97871 ( n18918, n18919, n18920 );
nor U97872 ( n18568, n18558, n18571 );
or U97873 ( n18571, n2582, n18556 );
nand U97874 ( n51651, n51895, n51894 );
nand U97875 ( n17948, n17937, n18167 );
nand U97876 ( n18167, n18168, n17936 );
nand U97877 ( n18168, n18175, n17941 );
nand U97878 ( n17937, n2448, n2399 );
not U97879 ( n2399, n17941 );
nor U97880 ( n53699, n50508, n1600 );
nand U97881 ( n18699, n18920, n18919 );
nor U97882 ( n53219, n53225, n53226 );
xor U97883 ( n53226, n53350, n53351 );
nand U97884 ( n53350, n53352, n53353 );
nand U97885 ( n20495, n20830, n20829 );
nand U97886 ( n19229, n19411, n19412 );
or U97887 ( n19411, n19218, n19215 );
nand U97888 ( n19412, n19217, n19413 );
nand U97889 ( n19413, n19215, n19218 );
nand U97890 ( n18875, n19099, n19100 );
nand U97891 ( n19099, n18864, n18862 );
nand U97892 ( n19100, n18863, n19101 );
or U97893 ( n19101, n18862, n18864 );
or U97894 ( n19947, n20238, n20239 );
nor U97895 ( n53255, n53262, n1519 );
nand U97896 ( n20083, n20084, n20079 );
nor U97897 ( n16987, n17369, n17365 );
nand U97898 ( n52354, n52350, n52349 );
nor U97899 ( n53102, n53109, n1497 );
nor U97900 ( n52963, n52964, n1440 );
nor U97901 ( n53224, n53225, n1498 );
nor U97902 ( n52974, n52981, n1473 );
nor U97903 ( n53221, n53222, n1524 );
nor U97904 ( n53222, n53223, n53224 );
and U97905 ( n53223, n53225, n1498 );
nand U97906 ( n53346, n76323, n53347 );
nand U97907 ( n53347, n76652, n73413 );
or U97908 ( n53243, n53341, n53342 );
xnor U97909 ( n49731, n49737, n49738 );
nand U97910 ( n49737, n49745, n49746 );
nor U97911 ( n49738, n49739, n49740 );
nand U97912 ( n49745, n49751, n49752 );
xor U97913 ( n49729, n49730, n49731 );
nor U97914 ( n49740, n49741, n49742 );
nor U97915 ( n49741, n49743, n49744 );
nand U97916 ( n19401, n19557, n19556 );
nor U97917 ( n20816, n20822, n20823 );
nand U97918 ( n53440, n53441, n53436 );
or U97919 ( n49689, n49695, n49694 );
xor U97920 ( n20372, n20492, n20493 );
nand U97921 ( n20492, n20494, n20495 );
nor U97922 ( n20365, n20371, n20372 );
nand U97923 ( n20824, n20822, n20825 );
nor U97924 ( n52543, n52550, n1410 );
nor U97925 ( n49735, n50008, n49734 );
nor U97926 ( n50008, n49733, n50011 );
nand U97927 ( n19859, n20324, n20325 );
or U97928 ( n20324, n20217, n20220 );
nand U97929 ( n20325, n20326, n20219 );
nand U97930 ( n20326, n20220, n20217 );
xor U97931 ( n49466, n50622, n50623 );
xor U97932 ( n50622, n50624, n50625 );
xor U97933 ( n20630, n20549, n20631 );
xor U97934 ( n20631, n20548, n20547 );
nand U97935 ( n19951, n20225, n8217 );
nor U97936 ( n20225, n2657, n73015 );
nand U97937 ( n19390, n19951, n19952 );
nand U97938 ( n19952, n19953, n19954 );
nand U97939 ( n19953, n2657, n17014 );
xor U97940 ( n16753, n16764, n16765 );
xor U97941 ( n16765, n16766, n16767 );
xor U97942 ( n16764, n17072, n17073 );
xor U97943 ( n16767, n16768, n16769 );
xor U97944 ( n17072, n17078, n17079 );
nor U97945 ( n17079, n73022, n17080 );
nand U97946 ( n17078, n17081, n17082 );
nand U97947 ( n17082, n17083, n17084 );
xor U97948 ( n20237, n20238, n20239 );
xor U97949 ( n19085, n19241, n18915 );
xnor U97950 ( n19241, n18914, n18913 );
nand U97951 ( n53039, n53040, n53035 );
xor U97952 ( n49760, n49761, n49762 );
nor U97953 ( n49762, n49763, n49764 );
nand U97954 ( n49761, n49997, n49998 );
nor U97955 ( n49763, n49770, n49766 );
nand U97956 ( n49746, n1482, n49747 );
nand U97957 ( n49747, n49748, n49749 );
not U97958 ( n1482, n49751 );
nand U97959 ( n49749, n1507, n49750 );
xor U97960 ( n51906, n51907, n51908 );
or U97961 ( n51645, n51907, n51908 );
nand U97962 ( n20546, n2703, n20548 );
not U97963 ( n2703, n20549 );
and U97964 ( n20252, n20544, n20545 );
nand U97965 ( n20544, n20549, n2685 );
nand U97966 ( n20545, n20546, n20547 );
not U97967 ( n2685, n20548 );
xor U97968 ( n50896, n50893, n50897 );
nand U97969 ( n50893, n51126, n51127 );
or U97970 ( n51126, n51131, n51130 );
nand U97971 ( n51127, n51128, n51129 );
nand U97972 ( n51128, n51130, n51131 );
or U97973 ( n52353, n52349, n52350 );
nand U97974 ( n51647, n51908, n51907 );
or U97975 ( n51505, n51538, n51539 );
nand U97976 ( n51336, n51509, n51510 );
nand U97977 ( n51510, n51511, n51512 );
nand U97978 ( n51511, n51513, n51514 );
nand U97979 ( n20409, n20408, n20410 );
xor U97980 ( n51537, n51538, n51539 );
or U97981 ( n19399, n19556, n19557 );
nand U97982 ( n50015, n50016, n50017 );
nand U97983 ( n50016, n50018, n50019 );
nand U97984 ( n17833, n18093, n18094 );
nand U97985 ( n18094, n18095, n17838 );
nand U97986 ( n18093, n18098, n17836 );
xor U97987 ( n18095, n18096, n18097 );
nor U97988 ( n18098, n17838, n17839 );
nand U97989 ( n8436, n15660, n15662 );
nor U97990 ( n15660, n15668, n15669 );
nor U97991 ( n15662, n15663, n15664 );
nor U97992 ( n15668, n14735, n14895 );
nand U97993 ( n17857, n18084, n18083 );
nand U97994 ( n50535, n50541, n76648 );
nor U97995 ( n50541, n50542, n73405 );
xor U97996 ( n52041, n52356, n51871 );
xnor U97997 ( n52356, n51870, n51869 );
nor U97998 ( n53108, n53109, n1472 );
nor U97999 ( n53104, n53105, n53106 );
nor U98000 ( n53105, n53107, n53108 );
and U98001 ( n53107, n53109, n1472 );
or U98002 ( n19269, n19852, n19853 );
nor U98003 ( n18889, n18892, n2403 );
nand U98004 ( n19237, n19406, n19407 );
or U98005 ( n19406, n19231, n19234 );
nand U98006 ( n19407, n19233, n19408 );
nand U98007 ( n19408, n19234, n19231 );
nand U98008 ( n53544, n53545, n53541 );
nand U98009 ( n53244, n53342, n53341 );
nand U98010 ( n8156, n16394, n16395 );
nor U98011 ( n16395, n16397, n16398 );
nor U98012 ( n16394, n16402, n16403 );
nor U98013 ( n16397, n14895, n16342 );
nand U98014 ( n8196, n16292, n16293 );
nor U98015 ( n16293, n16294, n16295 );
nor U98016 ( n16292, n16299, n16300 );
nor U98017 ( n16294, n14895, n16237 );
nand U98018 ( n8276, n16080, n16082 );
nor U98019 ( n16082, n16083, n16084 );
nor U98020 ( n16080, n16088, n16089 );
nor U98021 ( n16083, n14895, n16034 );
nand U98022 ( n8316, n15973, n15974 );
nor U98023 ( n15974, n15975, n15977 );
nor U98024 ( n15973, n15980, n15982 );
nor U98025 ( n15975, n14895, n15927 );
nand U98026 ( n8356, n15874, n15875 );
nor U98027 ( n15875, n15877, n15878 );
nor U98028 ( n15874, n15882, n15883 );
nor U98029 ( n15877, n14895, n15822 );
nand U98030 ( n8476, n15559, n15560 );
nor U98031 ( n15560, n15562, n15563 );
nor U98032 ( n15559, n15567, n15568 );
nor U98033 ( n15562, n14895, n15513 );
nand U98034 ( n8516, n15453, n15454 );
nor U98035 ( n15454, n15455, n15457 );
nor U98036 ( n15453, n15460, n15462 );
nor U98037 ( n15455, n14895, n15407 );
nand U98038 ( n8236, n16183, n16184 );
nor U98039 ( n16184, n16185, n16187 );
nor U98040 ( n16183, n16190, n16192 );
nand U98041 ( n16187, n16188, n16189 );
nand U98042 ( n8396, n15767, n15768 );
nor U98043 ( n15768, n15769, n15770 );
nor U98044 ( n15767, n15774, n15775 );
nand U98045 ( n15770, n15772, n15773 );
or U98046 ( n16733, n16739, n16738 );
xor U98047 ( n19851, n19852, n19853 );
nand U98048 ( n19886, n20260, n20261 );
nand U98049 ( n20261, n20262, n20263 );
nor U98050 ( n20260, n20264, n2704 );
not U98051 ( n2704, n20265 );
or U98052 ( n19383, n19873, n19874 );
nand U98053 ( n19528, n19565, n19566 );
or U98054 ( n19565, n19524, n19521 );
nand U98055 ( n19566, n19523, n19567 );
nand U98056 ( n19567, n19521, n19524 );
xor U98057 ( n19872, n19873, n19874 );
nor U98058 ( n17929, n17669, n17932 );
nor U98059 ( n17932, n17926, n17933 );
nand U98060 ( n17933, n17923, n17668 );
and U98061 ( n17673, n17921, n17922 );
nand U98062 ( n17922, n2365, n17667 );
nand U98063 ( n17921, n17929, n17930 );
not U98064 ( n2365, n17668 );
nand U98065 ( n51507, n51539, n51538 );
nand U98066 ( n20313, n20570, n20571 );
or U98067 ( n20570, n20575, n20574 );
nand U98068 ( n20571, n20572, n20573 );
nand U98069 ( n20572, n20574, n20575 );
xor U98070 ( n50883, n51855, n51130 );
xnor U98071 ( n51855, n51129, n51131 );
xnor U98072 ( n19113, n19521, n19522 );
xnor U98073 ( n19522, n19523, n19524 );
nand U98074 ( n19578, n19722, n19723 );
or U98075 ( n19722, n19672, n19675 );
nand U98076 ( n19723, n19674, n19724 );
nand U98077 ( n19724, n19675, n19672 );
nand U98078 ( n19271, n19853, n19852 );
nand U98079 ( n49687, n49694, n49695 );
nand U98080 ( n16731, n16738, n16739 );
nor U98081 ( n52705, n52712, n1442 );
and U98082 ( n19290, n19865, n8217 );
nor U98083 ( n19865, n2678, n73414 );
nand U98084 ( n19385, n19874, n19873 );
nor U98085 ( n20370, n20371, n2624 );
nand U98086 ( n20374, n20390, n20482 );
nand U98087 ( n20482, n20388, n20389 );
nand U98088 ( n20488, n76589, n20489 );
nand U98089 ( n20489, n76655, n73015 );
or U98090 ( n20389, n20483, n20484 );
nor U98091 ( n52858, n50508, n1629 );
xor U98092 ( n51932, n51933, n51934 );
nand U98093 ( n53799, n53842, n53843 );
nand U98094 ( n53843, n53790, n53787 );
nor U98095 ( n53842, n53786, n1632 );
not U98096 ( n1632, n53791 );
nor U98097 ( n52416, n52417, n52414 );
xor U98098 ( n52417, n52413, n1628 );
or U98099 ( n51558, n51934, n51933 );
nor U98100 ( n19818, n2558, n19825 );
nand U98101 ( n19825, n19824, n19826 );
nor U98102 ( n51300, n51476, n51473 );
nand U98103 ( n51042, n51297, n51298 );
nand U98104 ( n51298, n51299, n1730 );
not U98105 ( n1730, n51300 );
nand U98106 ( n16984, n17365, n17369 );
nor U98107 ( n17939, n2448, n17940 );
xor U98108 ( n17940, n17936, n17941 );
nand U98109 ( n20565, n20681, n20682 );
or U98110 ( n20681, n20686, n20685 );
nand U98111 ( n20682, n20683, n20684 );
nand U98112 ( n20683, n20685, n20686 );
nand U98113 ( n15171, n48755, n48756 );
nor U98114 ( n48755, n48761, n48762 );
nor U98115 ( n48756, n48757, n48758 );
nor U98116 ( n48761, n47941, n48098 );
nor U98117 ( n52463, n52886, n52883 );
nand U98118 ( n52442, n52880, n52881 );
nand U98119 ( n52881, n52882, n52462 );
nand U98120 ( n52880, n52885, n52460 );
xor U98121 ( n52882, n52883, n52884 );
nor U98122 ( n52885, n52462, n52463 );
nand U98123 ( n14931, n49313, n49314 );
nor U98124 ( n49314, n49315, n49316 );
nor U98125 ( n49313, n49319, n49320 );
nor U98126 ( n49315, n48098, n49276 );
nand U98127 ( n15011, n49122, n49123 );
nor U98128 ( n49123, n49124, n49125 );
nor U98129 ( n49122, n49128, n49129 );
nor U98130 ( n49124, n48098, n49086 );
nand U98131 ( n15051, n49044, n49045 );
nor U98132 ( n49045, n49046, n49047 );
nor U98133 ( n49044, n49050, n49051 );
nor U98134 ( n49046, n48098, n48991 );
nand U98135 ( n15091, n48949, n48950 );
nor U98136 ( n48950, n48951, n48952 );
nor U98137 ( n48949, n48955, n48956 );
nor U98138 ( n48951, n48098, n48892 );
nand U98139 ( n15211, n48662, n48663 );
nor U98140 ( n48663, n48664, n48665 );
nor U98141 ( n48662, n48668, n48669 );
nor U98142 ( n48664, n48098, n48625 );
nand U98143 ( n15251, n48584, n48585 );
nor U98144 ( n48585, n48586, n48587 );
nor U98145 ( n48584, n48590, n48591 );
nor U98146 ( n48586, n48098, n48531 );
nand U98147 ( n14891, n49406, n49407 );
nor U98148 ( n49407, n49408, n49409 );
nor U98149 ( n49406, n49412, n49413 );
nor U98150 ( n49408, n48098, n49354 );
nand U98151 ( n14971, n49217, n49218 );
nor U98152 ( n49218, n49219, n49220 );
nor U98153 ( n49217, n49223, n49224 );
nand U98154 ( n49220, n49221, n49222 );
nand U98155 ( n15131, n48848, n48849 );
nor U98156 ( n48849, n48850, n48851 );
nor U98157 ( n48848, n48854, n48855 );
nand U98158 ( n48851, n48852, n48853 );
nor U98159 ( n52959, n52960, n52961 );
nor U98160 ( n52960, n52962, n52963 );
and U98161 ( n52962, n52964, n1440 );
nor U98162 ( n53840, n53878, n53875 );
and U98163 ( n52857, n53805, n8227 );
nor U98164 ( n53805, n1645, n72999 );
nand U98165 ( n52873, n53837, n53838 );
nand U98166 ( n53838, n53839, n1665 );
not U98167 ( n1665, n53840 );
nand U98168 ( n51560, n51933, n51934 );
nor U98169 ( n17938, n17936, n17942 );
nand U98170 ( n17942, n2448, n17941 );
or U98171 ( n17855, n18083, n18084 );
nand U98172 ( n17667, n17923, n17924 );
nand U98173 ( n17924, n17925, n17926 );
nand U98174 ( n17925, n17927, n17928 );
nand U98175 ( n18957, n19387, n19388 );
or U98176 ( n19387, n19392, n19391 );
nand U98177 ( n19388, n19389, n19390 );
nand U98178 ( n19389, n19391, n19392 );
nand U98179 ( n20882, n20883, n20879 );
nor U98180 ( n53828, n53827, n53826 );
nand U98181 ( n52874, n53823, n53824 );
nand U98182 ( n53824, n53825, n52879 );
nand U98183 ( n53823, n52878, n53829 );
nor U98184 ( n53825, n52878, n53828 );
nand U98185 ( n53829, n1684, n53830 );
nand U98186 ( n53830, n53831, n53827 );
nand U98187 ( n53263, n53262, n53264 );
nand U98188 ( n20604, n20662, n20663 );
nand U98189 ( n17111, n17416, n17417 );
or U98190 ( n17416, n17421, n17420 );
nand U98191 ( n17417, n17418, n17419 );
nand U98192 ( n17418, n17420, n17421 );
nor U98193 ( n17361, n16988, n73399 );
nor U98194 ( n50309, n50312, n50313 );
nor U98195 ( n52549, n52550, n1375 );
nor U98196 ( n52545, n52546, n52547 );
nor U98197 ( n52546, n52548, n52549 );
and U98198 ( n52548, n52550, n1375 );
nand U98199 ( n53336, n53334, n53337 );
nand U98200 ( n15296, n48477, n48478 );
nor U98201 ( n48477, n48484, n48485 );
nor U98202 ( n48478, n48479, n48480 );
nor U98203 ( n48484, n48091, n48433 );
nand U98204 ( n15336, n48375, n48376 );
nor U98205 ( n48375, n48381, n48382 );
nor U98206 ( n48376, n48377, n48378 );
nor U98207 ( n48381, n48087, n48350 );
nand U98208 ( n15376, n48278, n48279 );
nor U98209 ( n48278, n48284, n48285 );
nor U98210 ( n48279, n48280, n48281 );
nor U98211 ( n48284, n48087, n48253 );
nand U98212 ( n15416, n48180, n48181 );
nor U98213 ( n48180, n48186, n48187 );
nor U98214 ( n48181, n48182, n48183 );
nor U98215 ( n48186, n48087, n48155 );
nor U98216 ( n53124, n53125, n1474 );
nor U98217 ( n52980, n52981, n1443 );
nor U98218 ( n53121, n53122, n1499 );
nor U98219 ( n53122, n53123, n53124 );
and U98220 ( n53123, n53125, n1474 );
nand U98221 ( n53239, n76323, n53240 );
nand U98222 ( n53240, n76652, n73017 );
nand U98223 ( n53128, n53231, n53232 );
nand U98224 ( n53231, n53144, n53141 );
nand U98225 ( n53232, n53143, n53233 );
or U98226 ( n53233, n53141, n53144 );
nor U98227 ( n50799, n49930, n73014 );
xnor U98228 ( n20150, n20391, n20392 );
xnor U98229 ( n20392, n20393, n20394 );
xnor U98230 ( n53713, n52903, n53714 );
xor U98231 ( n53714, n52902, n52904 );
nand U98232 ( n15456, n48081, n48082 );
nor U98233 ( n48081, n48088, n48089 );
nor U98234 ( n48082, n48083, n48084 );
nor U98235 ( n48088, n48032, n48091 );
nand U98236 ( n20478, n20476, n20479 );
xor U98237 ( n50920, n51176, n51107 );
xor U98238 ( n51176, n51108, n51105 );
nor U98239 ( n50921, n51145, n1364 );
nand U98240 ( n51108, n51342, n51343 );
or U98241 ( n51342, n51172, n51175 );
nand U98242 ( n51343, n51344, n51174 );
nand U98243 ( n51344, n51175, n51172 );
nand U98244 ( n52073, n52209, n52210 );
or U98245 ( n52209, n52169, n52168 );
nand U98246 ( n52210, n52170, n52211 );
nand U98247 ( n52211, n52168, n52169 );
nor U98248 ( n53119, n53125, n53126 );
xor U98249 ( n51703, n52167, n52168 );
xor U98250 ( n52167, n52169, n52170 );
nand U98251 ( n51815, n52060, n52061 );
or U98252 ( n52060, n51803, n51802 );
nand U98253 ( n52061, n51804, n52062 );
nand U98254 ( n52062, n51802, n51803 );
nand U98255 ( n51707, n52077, n52078 );
nand U98256 ( n52077, n51798, n51799 );
nand U98257 ( n52078, n51800, n52079 );
or U98258 ( n52079, n51799, n51798 );
nor U98259 ( n52577, n52584, n1415 );
nor U98260 ( n52087, n52094, n1339 );
nor U98261 ( n52976, n52977, n52978 );
nor U98262 ( n52977, n52979, n52980 );
and U98263 ( n52979, n52981, n1443 );
xnor U98264 ( n18855, n19215, n19216 );
xnor U98265 ( n19216, n19217, n19218 );
xor U98266 ( n16509, n17670, n17671 );
xor U98267 ( n17671, n17672, n17673 );
nor U98268 ( n53877, n53839, n53840 );
nand U98269 ( n53820, n53872, n53873 );
nand U98270 ( n53873, n53874, n53839 );
nand U98271 ( n53872, n53877, n53837 );
xor U98272 ( n53874, n53875, n53876 );
xor U98273 ( n18937, n18938, n18939 );
nor U98274 ( n17963, n18189, n2480 );
nand U98275 ( n18151, n18386, n18387 );
or U98276 ( n18386, n18216, n18219 );
nand U98277 ( n18387, n18388, n18218 );
nand U98278 ( n18388, n18219, n18216 );
nand U98279 ( n18588, n19074, n19075 );
or U98280 ( n19074, n19079, n19078 );
nand U98281 ( n19075, n19076, n19077 );
nand U98282 ( n19077, n19078, n19079 );
nand U98283 ( n20390, n20484, n20483 );
nand U98284 ( n50065, n50370, n50371 );
or U98285 ( n50370, n50375, n50374 );
nand U98286 ( n50371, n50372, n50373 );
nand U98287 ( n50372, n50374, n50375 );
or U98288 ( n18693, n18938, n18939 );
nand U98289 ( n53210, n53209, n53211 );
nand U98290 ( n52781, n52780, n52782 );
nor U98291 ( n20001, n20008, n2593 );
xor U98292 ( n16468, n17666, n17667 );
xor U98293 ( n17666, n17668, n17669 );
nor U98294 ( n52711, n52712, n1414 );
nor U98295 ( n52722, n52729, n1444 );
nor U98296 ( n52707, n52708, n52709 );
nor U98297 ( n52708, n52710, n52711 );
and U98298 ( n52710, n52712, n1414 );
nand U98299 ( n51985, n52460, n52461 );
nand U98300 ( n52461, n52462, n1689 );
not U98301 ( n1689, n52463 );
nand U98302 ( n52441, n1684, n52877 );
nand U98303 ( n52877, n52878, n52879 );
xor U98304 ( n19857, n19960, n20222 );
xor U98305 ( n20222, n19958, n19959 );
nor U98306 ( n19823, n19824, n2529 );
nor U98307 ( n19820, n19822, n19823 );
and U98308 ( n19822, n19824, n2529 );
nand U98309 ( n8561, n15332, n15333 );
nor U98310 ( n15332, n15340, n15342 );
nor U98311 ( n15333, n15334, n15335 );
nor U98312 ( n15340, n14887, n15297 );
nand U98313 ( n8601, n15225, n15227 );
nor U98314 ( n15225, n15233, n15234 );
nor U98315 ( n15227, n15228, n15229 );
nor U98316 ( n15233, n14882, n15185 );
nand U98317 ( n8641, n15115, n15117 );
nor U98318 ( n15115, n15123, n15124 );
nor U98319 ( n15117, n15118, n15119 );
nor U98320 ( n15123, n14882, n15078 );
nand U98321 ( n8681, n15005, n15007 );
nor U98322 ( n15005, n15013, n15014 );
nor U98323 ( n15007, n15008, n15009 );
nor U98324 ( n15013, n14882, n14974 );
nand U98325 ( n18695, n18939, n18938 );
nand U98326 ( n18891, n18892, n18887 );
nand U98327 ( n8721, n14874, n14875 );
nor U98328 ( n14874, n14883, n14884 );
nor U98329 ( n14875, n14877, n14878 );
nor U98330 ( n14883, n14830, n14887 );
nand U98331 ( n20585, n20673, n20674 );
nand U98332 ( n20674, n20675, n20676 );
xor U98333 ( n20022, n20189, n20190 );
xor U98334 ( n20190, n20191, n20192 );
nor U98335 ( n20007, n20008, n2562 );
nor U98336 ( n20367, n20368, n2647 );
nor U98337 ( n20368, n20369, n20370 );
and U98338 ( n20369, n20371, n2624 );
nand U98339 ( n51554, n52022, n52023 );
nand U98340 ( n52023, n52024, n52025 );
nor U98341 ( n16772, n16776, n16777 );
nor U98342 ( n16776, n2574, n16778 );
not U98343 ( n2574, n16779 );
xor U98344 ( n52348, n52349, n52350 );
xnor U98345 ( n17555, n17591, n17828 );
xnor U98346 ( n17828, n17590, n17592 );
not U98347 ( n1764, n50312 );
not U98348 ( n76929, n76927 );
buf U98349 ( n76319, n49931 );
nor U98350 ( n53009, n53010, n1445 );
nor U98351 ( n52728, n52729, n1417 );
nor U98352 ( n52093, n52094, n1297 );
nor U98353 ( n52265, n52272, n1382 );
nand U98354 ( n53012, n53131, n53132 );
nand U98355 ( n53131, n53000, n52997 );
nand U98356 ( n53132, n52999, n53133 );
or U98357 ( n53133, n52997, n53000 );
nor U98358 ( n53005, n53006, n53007 );
nor U98359 ( n53006, n53008, n53009 );
and U98360 ( n53008, n53010, n1445 );
nor U98361 ( n52724, n52725, n52726 );
nor U98362 ( n52725, n52727, n52728 );
and U98363 ( n52727, n52729, n1417 );
nand U98364 ( n53139, n76323, n53140 );
nand U98365 ( n53140, n76651, n73419 );
nand U98366 ( n53227, n53225, n53228 );
nand U98367 ( n52418, n52413, n52414 );
nand U98368 ( n53819, n1654, n53864 );
nand U98369 ( n53864, n53857, n53856 );
nand U98370 ( n52879, n53826, n53827 );
xor U98371 ( n51380, n51548, n51501 );
xor U98372 ( n51548, n51503, n51504 );
xor U98373 ( n18950, n18951, n18952 );
nand U98374 ( n51297, n51473, n51476 );
or U98375 ( n18689, n18951, n18952 );
xor U98376 ( n49549, n51817, n51818 );
xor U98377 ( n51817, n51819, n51820 );
nand U98378 ( n52460, n52883, n52886 );
nor U98379 ( n52583, n52584, n1380 );
nand U98380 ( n50664, n51103, n51104 );
nand U98381 ( n51103, n51107, n51108 );
nand U98382 ( n51104, n51105, n51106 );
or U98383 ( n51106, n51107, n51108 );
nand U98384 ( n52477, n52899, n52900 );
or U98385 ( n52899, n52903, n52904 );
nand U98386 ( n52900, n52901, n52902 );
nand U98387 ( n52901, n52903, n52904 );
nand U98388 ( n18691, n18952, n18951 );
or U98389 ( n18549, n18582, n18583 );
nand U98390 ( n53837, n53875, n53878 );
xor U98391 ( n18581, n18582, n18583 );
nand U98392 ( n15176, n48747, n48748 );
nor U98393 ( n48747, n48753, n48754 );
nor U98394 ( n48748, n48749, n48750 );
nor U98395 ( n48753, n47941, n48087 );
xor U98396 ( n19425, n19672, n19673 );
xor U98397 ( n19673, n19674, n19675 );
nand U98398 ( n14936, n49305, n49306 );
nor U98399 ( n49306, n49307, n49308 );
nor U98400 ( n49305, n49311, n49312 );
nor U98401 ( n49307, n48087, n49276 );
nand U98402 ( n15016, n49114, n49115 );
nor U98403 ( n49115, n49116, n49117 );
nor U98404 ( n49114, n49120, n49121 );
nor U98405 ( n49116, n48087, n49086 );
nand U98406 ( n15056, n49036, n49037 );
nor U98407 ( n49037, n49038, n49039 );
nor U98408 ( n49036, n49042, n49043 );
nor U98409 ( n49038, n48087, n48991 );
nand U98410 ( n15096, n48941, n48942 );
nor U98411 ( n48942, n48943, n48944 );
nor U98412 ( n48941, n48947, n48948 );
nor U98413 ( n48943, n48087, n48892 );
nand U98414 ( n15216, n48654, n48655 );
nor U98415 ( n48655, n48656, n48657 );
nor U98416 ( n48654, n48660, n48661 );
nor U98417 ( n48656, n48087, n48625 );
nand U98418 ( n15256, n48576, n48577 );
nor U98419 ( n48577, n48578, n48579 );
nor U98420 ( n48576, n48582, n48583 );
nor U98421 ( n48578, n48087, n48531 );
nand U98422 ( n14896, n49398, n49399 );
nor U98423 ( n49399, n49400, n49401 );
nor U98424 ( n49398, n49404, n49405 );
nor U98425 ( n49400, n48087, n49354 );
nand U98426 ( n14976, n49209, n49210 );
nor U98427 ( n49210, n49211, n49212 );
nor U98428 ( n49209, n49215, n49216 );
nand U98429 ( n49212, n49213, n49214 );
nand U98430 ( n15136, n48840, n48841 );
nor U98431 ( n48841, n48842, n48843 );
nor U98432 ( n48840, n48846, n48847 );
nand U98433 ( n48843, n48844, n48845 );
xor U98434 ( n17927, n18899, n18173 );
xnor U98435 ( n18899, n18172, n18174 );
nor U98436 ( n49764, n49765, n1577 );
not U98437 ( n1577, n49766 );
nor U98438 ( n49765, n49767, n49768 );
nor U98439 ( n49767, n1555, n49769 );
nand U98440 ( n15301, n48468, n48469 );
nor U98441 ( n48468, n48475, n48476 );
nor U98442 ( n48469, n48470, n48471 );
nor U98443 ( n48475, n48066, n48433 );
nand U98444 ( n15341, n48367, n48368 );
nor U98445 ( n48367, n48373, n48374 );
nor U98446 ( n48368, n48369, n48370 );
nor U98447 ( n48373, n48062, n48350 );
nand U98448 ( n15381, n48270, n48271 );
nor U98449 ( n48270, n48276, n48277 );
nor U98450 ( n48271, n48272, n48273 );
nor U98451 ( n48276, n48062, n48253 );
nand U98452 ( n15421, n48172, n48173 );
nor U98453 ( n48172, n48178, n48179 );
nor U98454 ( n48173, n48174, n48175 );
nor U98455 ( n48178, n48062, n48155 );
xor U98456 ( n19555, n19556, n19557 );
nand U98457 ( n17936, n18169, n18170 );
or U98458 ( n18169, n18174, n18173 );
nand U98459 ( n18170, n18171, n18172 );
nand U98460 ( n18171, n18173, n18174 );
nand U98461 ( n20154, n20360, n20361 );
nand U98462 ( n20360, n20192, n20189 );
nand U98463 ( n20361, n20191, n20362 );
or U98464 ( n20362, n20189, n20192 );
nand U98465 ( n15461, n48056, n48057 );
nor U98466 ( n48056, n48063, n48064 );
nor U98467 ( n48057, n48058, n48059 );
nor U98468 ( n48063, n48032, n48066 );
nand U98469 ( n50793, n50797, n76648 );
nor U98470 ( n50797, n50798, n73010 );
nor U98471 ( n17357, n16988, n73409 );
nand U98472 ( n18551, n18583, n18582 );
nor U98473 ( n19587, n19594, n2530 );
nor U98474 ( n52579, n52580, n52581 );
nor U98475 ( n52580, n52582, n52583 );
and U98476 ( n52582, n52584, n1380 );
nand U98477 ( n20309, n20582, n20583 );
nand U98478 ( n20583, n20584, n20585 );
nor U98479 ( n20582, n20586, n2755 );
not U98480 ( n2755, n20587 );
xor U98481 ( n18963, n18964, n18965 );
xor U98482 ( n20277, n20278, n20279 );
xor U98483 ( n18976, n18977, n18978 );
nor U98484 ( n20291, n20595, n20593 );
nand U98485 ( n19382, n19907, n19908 );
nand U98486 ( n19908, n19909, n19910 );
nor U98487 ( n19907, n19911, n19912 );
nor U98488 ( n19327, n19328, n19325 );
xor U98489 ( n19328, n19324, n2750 );
nand U98490 ( n19923, n20288, n20289 );
nand U98491 ( n20289, n20290, n2788 );
not U98492 ( n2788, n20291 );
xor U98493 ( n20578, n20579, n20580 );
nand U98494 ( n20285, n20589, n20590 );
nand U98495 ( n20590, n20591, n20290 );
nand U98496 ( n20589, n20594, n20288 );
xor U98497 ( n20591, n20592, n20593 );
nor U98498 ( n20594, n20290, n20291 );
or U98499 ( n18679, n18964, n18965 );
xnor U98500 ( n16775, n16782, n16783 );
nand U98501 ( n16782, n16790, n16791 );
nor U98502 ( n16783, n16784, n16785 );
nand U98503 ( n16790, n16796, n16797 );
xor U98504 ( n16773, n16774, n16775 );
nand U98505 ( n51279, n51470, n51471 );
nand U98506 ( n51471, n51472, n51299 );
nand U98507 ( n51470, n51475, n51297 );
xor U98508 ( n51472, n51473, n51474 );
nor U98509 ( n51475, n51299, n51300 );
nand U98510 ( n19945, n20279, n20278 );
nand U98511 ( n20308, n20580, n20579 );
nor U98512 ( n20297, n20296, n20295 );
nand U98513 ( n20298, n2802, n20299 );
nand U98514 ( n20299, n20300, n20296 );
nand U98515 ( n19924, n20292, n20293 );
nand U98516 ( n20293, n20294, n19942 );
nand U98517 ( n20292, n19941, n20298 );
nor U98518 ( n20294, n19941, n20297 );
or U98519 ( n20306, n20579, n20580 );
xor U98520 ( n19205, n19517, n19518 );
xor U98521 ( n19517, n19519, n19520 );
nand U98522 ( n19117, n19416, n19417 );
or U98523 ( n19416, n19213, n19212 );
nand U98524 ( n19417, n19214, n19418 );
nand U98525 ( n19418, n19212, n19213 );
nor U98526 ( n19593, n19594, n2492 );
nor U98527 ( n20003, n20004, n20005 );
nor U98528 ( n20004, n20006, n20007 );
and U98529 ( n20006, n20008, n2562 );
nor U98530 ( n19589, n19590, n19591 );
nor U98531 ( n19590, n19592, n19593 );
and U98532 ( n19592, n19594, n2492 );
nor U98533 ( n52271, n52272, n1343 );
nor U98534 ( n52751, n52752, n1420 );
nor U98535 ( n52612, n52613, n1384 );
nor U98536 ( n52608, n52609, n52610 );
nor U98537 ( n52609, n52611, n52612 );
and U98538 ( n52611, n52613, n1384 );
nor U98539 ( n52747, n52748, n52749 );
nor U98540 ( n52748, n52750, n52751 );
and U98541 ( n52750, n52752, n1420 );
nor U98542 ( n52267, n52268, n52269 );
nor U98543 ( n52268, n52270, n52271 );
and U98544 ( n52270, n52272, n1343 );
nand U98545 ( n53980, n76323, n53981 );
nand U98546 ( n53981, n76653, n73019 );
nand U98547 ( n52754, n52991, n52992 );
nand U98548 ( n52991, n52996, n52995 );
nand U98549 ( n52992, n52993, n52994 );
or U98550 ( n52994, n52995, n52996 );
or U98551 ( n18602, n18978, n18977 );
nand U98552 ( n53110, n53109, n53111 );
nand U98553 ( n18681, n18965, n18964 );
nand U98554 ( n18604, n18977, n18978 );
or U98555 ( n19943, n20278, n20279 );
xnor U98556 ( n16781, n16774, n16775 );
nand U98557 ( n19429, n19582, n19583 );
or U98558 ( n19582, n19519, n19518 );
nand U98559 ( n19583, n19520, n19584 );
nand U98560 ( n19584, n19518, n19519 );
xor U98561 ( n53007, n53141, n53142 );
xor U98562 ( n53142, n53143, n53144 );
nor U98563 ( n53003, n53010, n1475 );
nand U98564 ( n18380, n18553, n18554 );
nand U98565 ( n18554, n18555, n18556 );
nand U98566 ( n18555, n18557, n18558 );
nor U98567 ( n19378, n19933, n19931 );
nand U98568 ( n19357, n19927, n19928 );
nand U98569 ( n19928, n19929, n19377 );
nand U98570 ( n19927, n19932, n19375 );
xor U98571 ( n19929, n19930, n19931 );
nor U98572 ( n19932, n19377, n19378 );
or U98573 ( n19343, n19917, n19918 );
nand U98574 ( n17061, n17062, n17063 );
nand U98575 ( n17062, n17064, n17065 );
nor U98576 ( n20168, n20169, n2600 );
nand U98577 ( n20172, n20377, n20378 );
nand U98578 ( n20377, n20187, n20186 );
nand U98579 ( n20378, n20188, n20379 );
or U98580 ( n20379, n20186, n20187 );
nor U98581 ( n20165, n20166, n2625 );
nor U98582 ( n20166, n20167, n20168 );
and U98583 ( n20167, n20169, n2600 );
nand U98584 ( n20385, n76589, n20386 );
nand U98585 ( n20386, n76655, n73418 );
nand U98586 ( n20026, n20158, n20159 );
or U98587 ( n20158, n20060, n20057 );
nand U98588 ( n20159, n20059, n20160 );
nand U98589 ( n20160, n20057, n20060 );
xor U98590 ( n16805, n16806, n16807 );
nor U98591 ( n16807, n16808, n16809 );
nand U98592 ( n16806, n17043, n17044 );
nor U98593 ( n16808, n16815, n16811 );
nand U98594 ( n16791, n2605, n16792 );
nand U98595 ( n16792, n16793, n16794 );
not U98596 ( n2605, n16796 );
nand U98597 ( n16794, n2629, n16795 );
and U98598 ( n9953, n9954, n9894 );
nand U98599 ( n9576, n9898, n9899 );
nor U98600 ( n9899, n9900, n9902 );
nor U98601 ( n9898, n9952, n9953 );
nor U98602 ( n9900, n9464, n76632 );
nand U98603 ( n8441, n15650, n15652 );
nor U98604 ( n15650, n15658, n15659 );
nor U98605 ( n15652, n15653, n15654 );
nor U98606 ( n15658, n14735, n14882 );
xor U98607 ( n19916, n19917, n19918 );
xor U98608 ( n53777, n53778, n53779 );
nand U98609 ( n53779, n53851, n8229 );
nor U98610 ( n53851, n73397, n72999 );
nor U98611 ( n18344, n18512, n18510 );
nand U98612 ( n18089, n18341, n18342 );
nand U98613 ( n18342, n18343, n2849 );
not U98614 ( n2849, n18344 );
nand U98615 ( n8201, n16282, n16283 );
nor U98616 ( n16283, n16284, n16285 );
nor U98617 ( n16282, n16289, n16290 );
nor U98618 ( n16284, n14882, n16237 );
nand U98619 ( n8281, n16070, n16072 );
nor U98620 ( n16072, n16073, n16074 );
nor U98621 ( n16070, n16078, n16079 );
nor U98622 ( n16073, n14882, n16034 );
nand U98623 ( n8321, n15963, n15964 );
nor U98624 ( n15964, n15965, n15967 );
nor U98625 ( n15963, n15970, n15972 );
nor U98626 ( n15965, n14882, n15927 );
nand U98627 ( n8361, n15858, n15859 );
nor U98628 ( n15859, n15860, n15862 );
nor U98629 ( n15858, n15865, n15867 );
nor U98630 ( n15860, n14882, n15822 );
nand U98631 ( n8481, n15549, n15550 );
nor U98632 ( n15550, n15552, n15553 );
nor U98633 ( n15549, n15557, n15558 );
nor U98634 ( n15552, n14882, n15513 );
nand U98635 ( n8521, n15443, n15444 );
nor U98636 ( n15444, n15445, n15447 );
nor U98637 ( n15443, n15450, n15452 );
nor U98638 ( n15445, n14882, n15407 );
nand U98639 ( n8161, n16378, n16379 );
nor U98640 ( n16379, n16380, n16382 );
nor U98641 ( n16378, n16385, n16387 );
nor U98642 ( n16380, n14882, n16342 );
nand U98643 ( n8241, n16173, n16174 );
nor U98644 ( n16174, n16175, n16177 );
nor U98645 ( n16173, n16180, n16182 );
nand U98646 ( n16177, n16178, n16179 );
nand U98647 ( n8401, n15757, n15758 );
nor U98648 ( n15758, n15759, n15760 );
nor U98649 ( n15757, n15764, n15765 );
nand U98650 ( n15760, n15762, n15763 );
nor U98651 ( n17897, n17902, n17901 );
nor U98652 ( n17055, n16777, n16779 );
xor U98653 ( n18082, n18083, n18084 );
nand U98654 ( n51208, n51499, n51500 );
nand U98655 ( n51499, n51504, n51503 );
nand U98656 ( n51500, n51501, n51502 );
or U98657 ( n51502, n51503, n51504 );
or U98658 ( n51329, n51362, n51363 );
or U98659 ( n51325, n51375, n51376 );
nand U98660 ( n19345, n19918, n19917 );
xor U98661 ( n51361, n51362, n51363 );
or U98662 ( n53782, n53779, n53778 );
xor U98663 ( n51374, n51375, n51376 );
nand U98664 ( n52551, n52550, n52552 );
nor U98665 ( n20163, n20169, n20170 );
xor U98666 ( n20170, n20387, n20388 );
nand U98667 ( n20387, n20389, n20390 );
nand U98668 ( n19072, n2679, n19292 );
not U98669 ( n2679, n19284 );
nand U98670 ( n51331, n51363, n51362 );
nand U98671 ( n52965, n52964, n52966 );
nand U98672 ( n53127, n53125, n53128 );
xor U98673 ( n18747, n19211, n19212 );
xor U98674 ( n19211, n19213, n19214 );
nand U98675 ( n18859, n19104, n19105 );
or U98676 ( n19104, n18847, n18846 );
nand U98677 ( n19105, n18848, n19106 );
nand U98678 ( n19106, n18846, n18847 );
xnor U98679 ( n51924, n52397, n52024 );
nand U98680 ( n52397, n52025, n52022 );
nand U98681 ( n51327, n51376, n51375 );
nand U98682 ( n53783, n53779, n53778 );
nor U98683 ( n50852, n50857, n50856 );
and U98684 ( n43844, n43845, n43797 );
nand U98685 ( n16311, n43800, n43801 );
nor U98686 ( n43801, n43802, n43803 );
nor U98687 ( n43800, n43843, n43844 );
nor U98688 ( n43802, n43398, n76362 );
nand U98689 ( n20284, n2775, n20602 );
nand U98690 ( n20602, n20603, n20604 );
nand U98691 ( n8566, n15320, n15322 );
nor U98692 ( n15320, n15329, n15330 );
nor U98693 ( n15322, n15323, n15324 );
nor U98694 ( n15329, n14873, n15297 );
nand U98695 ( n8606, n15215, n15217 );
nor U98696 ( n15215, n15223, n15224 );
nor U98697 ( n15217, n15218, n15219 );
nor U98698 ( n15223, n14868, n15185 );
nand U98699 ( n8646, n15105, n15107 );
nor U98700 ( n15105, n15113, n15114 );
nor U98701 ( n15107, n15108, n15109 );
nor U98702 ( n15113, n14868, n15078 );
nand U98703 ( n8686, n14995, n14997 );
nor U98704 ( n14995, n15003, n15004 );
nor U98705 ( n14997, n14998, n14999 );
nor U98706 ( n15003, n14868, n14974 );
nand U98707 ( n51051, n51057, n76648 );
nor U98708 ( n51057, n51058, n73014 );
nand U98709 ( n8726, n14860, n14862 );
nor U98710 ( n14860, n14869, n14870 );
nor U98711 ( n14862, n14863, n14864 );
nor U98712 ( n14869, n14830, n14873 );
xor U98713 ( n51387, n51388, n51389 );
nor U98714 ( n19749, n19756, n2563 );
xor U98715 ( n19349, n19350, n19351 );
nand U98716 ( n19034, n19375, n19376 );
nand U98717 ( n19376, n19377, n2809 );
not U98718 ( n2809, n19378 );
nor U98719 ( n51783, n51790, n1298 );
or U98720 ( n51321, n51388, n51389 );
nand U98721 ( n20288, n20593, n20595 );
nand U98722 ( n19023, n19351, n19350 );
or U98723 ( n19021, n19350, n19351 );
nand U98724 ( n19356, n2802, n19940 );
nand U98725 ( n19940, n19941, n19942 );
nor U98726 ( n19755, n19756, n2534 );
nor U98727 ( n19751, n19752, n19753 );
nor U98728 ( n19752, n19754, n19755 );
and U98729 ( n19754, n19756, n2534 );
nand U98730 ( n52713, n52712, n52714 );
nand U98731 ( n50886, n50887, n50883 );
nor U98732 ( n50887, n50006, n8239 );
nor U98733 ( n52089, n52090, n52091 );
nor U98734 ( n52090, n52092, n52093 );
and U98735 ( n52092, n52094, n1297 );
nand U98736 ( n51323, n51389, n51388 );
nand U98737 ( n19900, n20268, n20269 );
nand U98738 ( n20269, n19911, n2752 );
nor U98739 ( n20268, n20271, n20272 );
nor U98740 ( n20271, n20273, n20274 );
nand U98741 ( n52982, n52981, n52983 );
nand U98742 ( n15181, n48739, n48740 );
nor U98743 ( n48739, n48745, n48746 );
nor U98744 ( n48740, n48741, n48742 );
nor U98745 ( n48745, n47941, n48062 );
nand U98746 ( n20373, n20371, n20374 );
nor U98747 ( n51469, n51615, n51612 );
nand U98748 ( n51278, n51466, n51467 );
nand U98749 ( n51467, n51468, n1720 );
not U98750 ( n1720, n51469 );
nand U98751 ( n14901, n49390, n49391 );
nor U98752 ( n49391, n49392, n49393 );
nor U98753 ( n49390, n49396, n49397 );
nor U98754 ( n49392, n48062, n49354 );
nand U98755 ( n14941, n49297, n49298 );
nor U98756 ( n49298, n49299, n49300 );
nor U98757 ( n49297, n49303, n49304 );
nor U98758 ( n49299, n48062, n49276 );
nand U98759 ( n15021, n49106, n49107 );
nor U98760 ( n49107, n49108, n49109 );
nor U98761 ( n49106, n49112, n49113 );
nor U98762 ( n49108, n48062, n49086 );
nand U98763 ( n15061, n49012, n49013 );
nor U98764 ( n49013, n49014, n49015 );
nor U98765 ( n49012, n49018, n49019 );
nor U98766 ( n49014, n48062, n48991 );
nand U98767 ( n15101, n48929, n48930 );
nor U98768 ( n48930, n48931, n48932 );
nor U98769 ( n48929, n48935, n48936 );
nor U98770 ( n48931, n48062, n48892 );
nand U98771 ( n15221, n48646, n48647 );
nor U98772 ( n48647, n48648, n48649 );
nor U98773 ( n48646, n48652, n48653 );
nor U98774 ( n48648, n48062, n48625 );
nand U98775 ( n15261, n48552, n48553 );
nor U98776 ( n48553, n48554, n48555 );
nor U98777 ( n48552, n48558, n48559 );
nor U98778 ( n48554, n48062, n48531 );
nand U98779 ( n15141, n48832, n48833 );
nor U98780 ( n48833, n48834, n48835 );
nor U98781 ( n48832, n48838, n48839 );
nand U98782 ( n48835, n48836, n48837 );
nand U98783 ( n14981, n49201, n49202 );
nor U98784 ( n49202, n49203, n49204 );
nor U98785 ( n49201, n49207, n49208 );
nand U98786 ( n49204, n49205, n49206 );
xnor U98787 ( n19770, n20057, n20058 );
xnor U98788 ( n20058, n20059, n20060 );
nor U98789 ( n51789, n51790, n1259 );
xor U98790 ( n18424, n18592, n18545 );
xor U98791 ( n18592, n18547, n18548 );
nand U98792 ( n19375, n19931, n19933 );
nand U98793 ( n53011, n53010, n53012 );
nand U98794 ( n19309, n19888, n19889 );
nand U98795 ( n19888, n19893, n2715 );
nand U98796 ( n19889, n19890, n19891 );
nand U98797 ( n19890, n2734, n19892 );
nor U98798 ( n19621, n19628, n2535 );
nor U98799 ( n52606, n52613, n1418 );
nor U98800 ( n52115, n1344, n52118 );
nand U98801 ( n19329, n19324, n19325 );
nand U98802 ( n18078, n18317, n18316 );
nand U98803 ( n19209, n19433, n19434 );
nand U98804 ( n19433, n19197, n19196 );
nand U98805 ( n19434, n19198, n19435 );
or U98806 ( n19435, n19196, n19197 );
nand U98807 ( n18751, n19121, n19122 );
nand U98808 ( n19121, n18842, n18843 );
nand U98809 ( n19122, n18844, n19123 );
or U98810 ( n19123, n18843, n18842 );
nor U98811 ( n19131, n19138, n2457 );
nand U98812 ( n49551, n51688, n51689 );
nand U98813 ( n51688, n49520, n49521 );
nand U98814 ( n51689, n49522, n51690 );
or U98815 ( n51690, n49521, n49520 );
nand U98816 ( n18598, n19066, n19067 );
nand U98817 ( n19067, n19068, n19069 );
nor U98818 ( n53727, n49930, n73400 );
nor U98819 ( n50954, n49989, n1458 );
and U98820 ( n51101, n51179, n51180 );
nand U98821 ( n51180, n50953, n1458 );
nor U98822 ( n51179, n51182, n51183 );
nor U98823 ( n51182, n51184, n51185 );
or U98824 ( n50848, n50927, n50928 );
nand U98825 ( n53731, n76649, n72999 );
nand U98826 ( n53772, n76650, n73397 );
nand U98827 ( n19942, n20295, n20296 );
xor U98828 ( n50926, n50927, n50928 );
nand U98829 ( n19774, n20030, n20031 );
or U98830 ( n20030, n19800, n19802 );
nand U98831 ( n20031, n19801, n20032 );
nand U98832 ( n20032, n19802, n19800 );
nor U98833 ( n20053, n20054, n2570 );
nand U98834 ( n20056, n20175, n20176 );
nand U98835 ( n20175, n20043, n20042 );
nand U98836 ( n20176, n20044, n20177 );
or U98837 ( n20177, n20042, n20043 );
nor U98838 ( n20049, n20050, n20051 );
nor U98839 ( n20050, n20052, n20053 );
and U98840 ( n20052, n20054, n2570 );
nand U98841 ( n20183, n76589, n20184 );
nand U98842 ( n20184, n76655, n73018 );
xor U98843 ( n52749, n52997, n52998 );
xor U98844 ( n52998, n52999, n53000 );
nor U98845 ( n52745, n52752, n1447 );
nand U98846 ( n50850, n50928, n50927 );
nor U98847 ( n19137, n19138, n2413 );
nor U98848 ( n19472, n19479, n2498 );
nand U98849 ( n52730, n52729, n52731 );
nor U98850 ( n19627, n19628, n2497 );
nand U98851 ( n18341, n18510, n18512 );
nor U98852 ( n19623, n19624, n19625 );
nor U98853 ( n19624, n19626, n19627 );
and U98854 ( n19626, n19628, n2497 );
nand U98855 ( n19658, n19778, n19779 );
or U98856 ( n19778, n19645, n19647 );
nand U98857 ( n19779, n19646, n19780 );
nand U98858 ( n19780, n19647, n19645 );
nor U98859 ( n19478, n19479, n2462 );
nor U98860 ( n19795, n19796, n2540 );
nand U98861 ( n19798, n20035, n20036 );
nand U98862 ( n20035, n20040, n20039 );
nand U98863 ( n20036, n20037, n20038 );
or U98864 ( n20038, n20039, n20040 );
nor U98865 ( n19474, n19475, n19476 );
nor U98866 ( n19475, n19477, n19478 );
and U98867 ( n19477, n19479, n2462 );
nor U98868 ( n19791, n19792, n19793 );
nor U98869 ( n19792, n19794, n19795 );
and U98870 ( n19794, n19796, n2540 );
nand U98871 ( n21084, n76589, n21085 );
nand U98872 ( n21085, n76654, n73420 );
nand U98873 ( n53671, n76649, n73400 );
xnor U98874 ( n16572, n18861, n18862 );
xnor U98875 ( n18861, n18863, n18864 );
nor U98876 ( n53866, n49930, n73002 );
or U98877 ( n18076, n18316, n18317 );
nor U98878 ( n50936, n50937, n50938 );
nand U98879 ( n50938, n50939, n50940 );
nor U98880 ( n52742, n53962, n1388 );
nor U98881 ( n52292, n52293, n1347 );
nor U98882 ( n53964, n53965, n52739 );
nor U98883 ( n53965, n53966, n52742 );
and U98884 ( n53966, n53962, n1388 );
nand U98885 ( n54062, n76323, n54063 );
nand U98886 ( n54063, n76653, n73421 );
nand U98887 ( n52740, n53968, n53969 );
nand U98888 ( n53968, n53973, n53972 );
nand U98889 ( n53969, n53970, n53971 );
or U98890 ( n53971, n53972, n53973 );
nor U98891 ( n53599, n49930, n73410 );
nand U98892 ( n52585, n52584, n52586 );
nand U98893 ( n8446, n15640, n15642 );
nor U98894 ( n15640, n15648, n15649 );
nor U98895 ( n15642, n15643, n15644 );
nor U98896 ( n15648, n14735, n14868 );
or U98897 ( n19066, n17525, n19295 );
xor U98898 ( n51400, n51497, n51557 );
xor U98899 ( n51557, n51496, n51498 );
xnor U98900 ( n18969, n19068, n75782 );
nand U98901 ( n75782, n19066, n19069 );
nand U98902 ( n8166, n16368, n16369 );
nor U98903 ( n16369, n16370, n16372 );
nor U98904 ( n16368, n16375, n16377 );
nor U98905 ( n16370, n14868, n16342 );
nand U98906 ( n8206, n16272, n16273 );
nor U98907 ( n16273, n16274, n16275 );
nor U98908 ( n16272, n16279, n16280 );
nor U98909 ( n16274, n14868, n16237 );
nand U98910 ( n8286, n16060, n16062 );
nor U98911 ( n16062, n16063, n16064 );
nor U98912 ( n16060, n16068, n16069 );
nor U98913 ( n16063, n14868, n16034 );
nand U98914 ( n8326, n15953, n15954 );
nor U98915 ( n15954, n15955, n15957 );
nor U98916 ( n15953, n15960, n15962 );
nor U98917 ( n15955, n14868, n15927 );
nand U98918 ( n8366, n15848, n15849 );
nor U98919 ( n15849, n15850, n15852 );
nor U98920 ( n15848, n15855, n15857 );
nor U98921 ( n15850, n14868, n15822 );
nand U98922 ( n8486, n15539, n15540 );
nor U98923 ( n15540, n15542, n15543 );
nor U98924 ( n15539, n15547, n15548 );
nor U98925 ( n15542, n14868, n15513 );
nand U98926 ( n8526, n15433, n15434 );
nor U98927 ( n15434, n15435, n15437 );
nor U98928 ( n15433, n15440, n15442 );
nor U98929 ( n15435, n14868, n15407 );
nand U98930 ( n8246, n16163, n16164 );
nor U98931 ( n16164, n16165, n16167 );
nor U98932 ( n16163, n16170, n16172 );
nand U98933 ( n16167, n16168, n16169 );
nand U98934 ( n8406, n15747, n15748 );
nor U98935 ( n15748, n15749, n15750 );
nor U98936 ( n15747, n15754, n15755 );
nand U98937 ( n15750, n15752, n15753 );
and U98938 ( n43884, n43893, n43797 );
nand U98939 ( n16306, n43882, n43883 );
nor U98940 ( n43882, n43894, n43895 );
nor U98941 ( n43883, n43884, n43885 );
nor U98942 ( n43894, n43408, n76362 );
nand U98943 ( n52753, n52752, n52754 );
nand U98944 ( n52273, n52272, n52274 );
nand U98945 ( n19595, n19594, n19596 );
nand U98946 ( n51463, n51609, n51610 );
nand U98947 ( n51610, n51611, n51468 );
nand U98948 ( n51609, n51614, n51466 );
xor U98949 ( n51611, n51612, n51613 );
nor U98950 ( n51614, n51468, n51469 );
not U98951 ( n8222, n17374 );
nand U98952 ( n18323, n18506, n18507 );
nand U98953 ( n18507, n18508, n18343 );
nand U98954 ( n18506, n18511, n18341 );
xor U98955 ( n18508, n18509, n18510 );
nor U98956 ( n18511, n18343, n18344 );
nand U98957 ( n49977, n50196, n50197 );
or U98958 ( n50196, n50200, n50201 );
nand U98959 ( n50197, n50198, n50199 );
nand U98960 ( n50198, n50200, n50201 );
nor U98961 ( n52286, n52293, n1385 );
nand U98962 ( n20009, n20008, n20010 );
nand U98963 ( n20171, n20169, n20172 );
xor U98964 ( n18315, n18316, n18317 );
not U98965 ( n2758, n20747 );
xor U98966 ( n52739, n52995, n53974 );
xor U98967 ( n53974, n52993, n52996 );
nor U98968 ( n52741, n53962, n1419 );
nor U98969 ( n16809, n16810, n2698 );
not U98970 ( n2698, n16811 );
nor U98971 ( n16810, n16812, n16813 );
nor U98972 ( n16812, n2675, n16814 );
xnor U98973 ( n20051, n20185, n20186 );
xnor U98974 ( n20185, n20187, n20188 );
nor U98975 ( n20047, n20054, n2602 );
nand U98976 ( n51466, n51612, n51615 );
nand U98977 ( n52614, n52613, n52615 );
xor U98978 ( n18431, n18432, n18433 );
nand U98979 ( n18366, n18442, n18443 );
nand U98980 ( n18442, n18447, n18446 );
nand U98981 ( n18443, n18444, n18445 );
or U98982 ( n18445, n18446, n18447 );
or U98983 ( n18373, n18406, n18407 );
or U98984 ( n18243, n18419, n18420 );
nand U98985 ( n18256, n18543, n18544 );
nand U98986 ( n18543, n18548, n18547 );
nand U98987 ( n18544, n18545, n18546 );
or U98988 ( n18546, n18547, n18548 );
xor U98989 ( n18405, n18406, n18407 );
or U98990 ( n18369, n18432, n18433 );
xor U98991 ( n18418, n18419, n18420 );
nand U98992 ( n18375, n18407, n18406 );
nand U98993 ( n18245, n18420, n18419 );
nand U98994 ( n18371, n18433, n18432 );
nand U98995 ( n50471, n50743, n50742 );
nand U98996 ( n53603, n76649, n73003 );
and U98997 ( n9959, n9970, n9894 );
nand U98998 ( n9571, n9957, n9958 );
nor U98999 ( n9957, n9972, n9973 );
nor U99000 ( n9958, n9959, n9960 );
nor U99001 ( n9972, n9477, n76632 );
nor U99002 ( n53473, n49930, n73412 );
nor U99003 ( n52288, n52289, n52290 );
nor U99004 ( n52289, n52291, n52292 );
and U99005 ( n52291, n52293, n1347 );
nand U99006 ( n15306, n48459, n48460 );
nor U99007 ( n48459, n48466, n48467 );
nor U99008 ( n48460, n48461, n48462 );
nor U99009 ( n48466, n48055, n48433 );
nand U99010 ( n15346, n48359, n48360 );
nor U99011 ( n48359, n48365, n48366 );
nor U99012 ( n48360, n48361, n48362 );
nor U99013 ( n48365, n48051, n48350 );
nand U99014 ( n15386, n48262, n48263 );
nor U99015 ( n48262, n48268, n48269 );
nor U99016 ( n48263, n48264, n48265 );
nor U99017 ( n48268, n48051, n48253 );
nand U99018 ( n15426, n48164, n48165 );
nor U99019 ( n48164, n48170, n48171 );
nor U99020 ( n48165, n48166, n48167 );
nor U99021 ( n48170, n48051, n48155 );
nor U99022 ( n17854, n73013, n18105 );
nand U99023 ( n53861, n53870, n76648 );
nor U99024 ( n53870, n53871, n73002 );
nand U99025 ( n15466, n48045, n48046 );
nor U99026 ( n48045, n48052, n48053 );
nor U99027 ( n48046, n48047, n48048 );
nor U99028 ( n48052, n48032, n48055 );
or U99029 ( n50469, n50742, n50743 );
xor U99030 ( n50656, n50657, n50658 );
nand U99031 ( n20675, n20747, n2759 );
not U99032 ( n2759, n20739 );
nor U99033 ( n20786, n73404, n18105 );
or U99034 ( n50574, n50657, n50658 );
nand U99035 ( n51218, n51493, n51494 );
or U99036 ( n51493, n51497, n51498 );
nand U99037 ( n51494, n51495, n51496 );
nand U99038 ( n51495, n51497, n51498 );
nand U99039 ( n19757, n19756, n19758 );
and U99040 ( n51061, n51296, n8229 );
nor U99041 ( n51296, n73415, n73016 );
nor U99042 ( n51062, n51291, n1742 );
not U99043 ( n1752, n51288 );
nand U99044 ( n53527, n76649, n73410 );
nand U99045 ( n53848, n76650, n73002 );
nand U99046 ( n18311, n18497, n18496 );
or U99047 ( n50286, n76322, n73014 );
buf U99048 ( n76322, n76320 );
nor U99049 ( n17978, n17979, n17980 );
nand U99050 ( n17980, n17981, n17982 );
nand U99051 ( n50847, n50949, n50950 );
nand U99052 ( n50950, n50951, n50952 );
nor U99053 ( n50949, n50953, n50954 );
nand U99054 ( n53477, n76649, n73008 );
nand U99055 ( n18769, n19126, n19127 );
or U99056 ( n19126, n18839, n18838 );
nand U99057 ( n19127, n18840, n19128 );
nand U99058 ( n19128, n18838, n18839 );
nor U99059 ( n18833, n18834, n2374 );
nand U99060 ( n16574, n18732, n18733 );
nand U99061 ( n18732, n16535, n16537 );
nand U99062 ( n18733, n16538, n18734 );
or U99063 ( n18734, n16537, n16535 );
nand U99064 ( n50576, n50658, n50657 );
nor U99065 ( n51992, n73411, n52001 );
nor U99066 ( n19786, n21067, n2504 );
nand U99067 ( n21104, n76589, n21105 );
nand U99068 ( n21105, n76654, n73020 );
nand U99069 ( n19784, n21073, n21074 );
nand U99070 ( n21073, n21078, n21077 );
nand U99071 ( n21074, n21075, n21076 );
or U99072 ( n21076, n21077, n21078 );
xnor U99073 ( n19654, n19799, n19800 );
xnor U99074 ( n19799, n19801, n19802 );
and U99075 ( n53242, n53343, n8229 );
nor U99076 ( n53343, n73413, n73017 );
nor U99077 ( n19159, n2463, n19162 );
nor U99078 ( n52447, n73401, n52001 );
nor U99079 ( n18522, n18655, n18653 );
nand U99080 ( n18322, n18519, n18520 );
nand U99081 ( n18520, n18521, n2840 );
not U99082 ( n2840, n18522 );
xnor U99083 ( n50467, n50200, n50468 );
xor U99084 ( n50468, n50199, n50201 );
nor U99085 ( n53987, n54039, n1348 );
nand U99086 ( n54053, n76323, n54054 );
nand U99087 ( n54054, n76653, n73021 );
nand U99088 ( n53985, n54045, n54046 );
nand U99089 ( n54045, n54036, n54033 );
nand U99090 ( n54046, n54035, n54047 );
or U99091 ( n54047, n54033, n54036 );
nor U99092 ( n50935, n1429, n50941 );
nand U99093 ( n50941, n50001, n50089 );
nor U99094 ( n19133, n19134, n19135 );
nor U99095 ( n19134, n19136, n19137 );
and U99096 ( n19136, n19138, n2413 );
nor U99097 ( n52301, n53947, n1305 );
nor U99098 ( n54041, n54042, n53984 );
nor U99099 ( n54042, n54043, n53987 );
and U99100 ( n54043, n54039, n1348 );
nand U99101 ( n52095, n52094, n52096 );
or U99102 ( n18309, n18496, n18497 );
nand U99103 ( n19501, n19638, n19639 );
or U99104 ( n19638, n19643, n19642 );
nand U99105 ( n19639, n19640, n19641 );
nand U99106 ( n19641, n19642, n19643 );
nor U99107 ( n21069, n21070, n19783 );
nor U99108 ( n21070, n21071, n19786 );
and U99109 ( n21071, n21067, n2504 );
and U99110 ( n43973, n43974, n43797 );
nand U99111 ( n16301, n43929, n43930 );
nor U99112 ( n43930, n43931, n43932 );
nor U99113 ( n43929, n43972, n43973 );
nor U99114 ( n43931, n43416, n76362 );
nand U99115 ( n20055, n20054, n20056 );
nor U99116 ( n18827, n18834, n2414 );
xor U99117 ( n50741, n50742, n50743 );
xor U99118 ( n18444, n18541, n18601 );
xor U99119 ( n18601, n18540, n18542 );
nand U99120 ( n19629, n19628, n19630 );
nand U99121 ( n19797, n19796, n19798 );
xnor U99122 ( n19793, n20041, n20042 );
xnor U99123 ( n20041, n20043, n20044 );
nor U99124 ( n19789, n19796, n2572 );
nand U99125 ( n19480, n19479, n19481 );
nand U99126 ( n17023, n17250, n17251 );
or U99127 ( n17250, n17254, n17255 );
nand U99128 ( n17251, n17252, n17253 );
nand U99129 ( n17252, n17254, n17255 );
xor U99130 ( n53984, n53972, n54055 );
xor U99131 ( n54055, n53970, n53973 );
nor U99132 ( n53986, n54039, n1387 );
xor U99133 ( n18495, n18496, n18497 );
nor U99134 ( n50298, n49898, n73010 );
and U99135 ( n49493, n51694, n51695 );
or U99136 ( n51694, n49457, n49456 );
nand U99137 ( n51695, n49458, n51696 );
nand U99138 ( n51696, n49456, n49457 );
xor U99139 ( n17701, n17702, n17703 );
xnor U99140 ( n18765, n19195, n19196 );
xnor U99141 ( n19195, n19197, n19198 );
or U99142 ( n17617, n17702, n17703 );
xnor U99143 ( n19783, n21079, n20039 );
xnor U99144 ( n21079, n20037, n20040 );
nor U99145 ( n19785, n21067, n2539 );
xnor U99146 ( n49490, n51801, n51802 );
xor U99147 ( n51801, n51803, n51804 );
nand U99148 ( n53967, n53962, n52740 );
nor U99149 ( n20831, n73414, n18105 );
xnor U99150 ( n18437, n18444, n18594 );
xnor U99151 ( n18594, n18447, n18446 );
nor U99152 ( n17365, n73004, n76575 );
buf U99153 ( n76575, n76574 );
nand U99154 ( n17619, n17703, n17702 );
nand U99155 ( n53349, n76649, n73412 );
nand U99156 ( n50951, n51186, n51187 );
nand U99157 ( n51187, n1485, n51188 );
nand U99158 ( n51186, n51191, n51096 );
xor U99159 ( n51188, n51189, n51190 );
or U99160 ( n51093, n51189, n51190 );
or U99161 ( n50969, n51202, n51203 );
nor U99162 ( n17996, n17035, n2580 );
xor U99163 ( n17968, n17969, n17970 );
and U99164 ( n18144, n18223, n18224 );
nand U99165 ( n18224, n17995, n2580 );
nor U99166 ( n18223, n18226, n18227 );
nor U99167 ( n18226, n18228, n18229 );
nand U99168 ( n15186, n48731, n48732 );
nor U99169 ( n48731, n48737, n48738 );
nor U99170 ( n48732, n48733, n48734 );
nor U99171 ( n48737, n47941, n48051 );
or U99172 ( n17893, n17969, n17970 );
nand U99173 ( n14906, n49382, n49383 );
nor U99174 ( n49383, n49384, n49385 );
nor U99175 ( n49382, n49388, n49389 );
nor U99176 ( n49384, n48051, n49354 );
nand U99177 ( n14946, n49289, n49290 );
nor U99178 ( n49290, n49291, n49292 );
nor U99179 ( n49289, n49295, n49296 );
nor U99180 ( n49291, n48051, n49276 );
nand U99181 ( n15026, n49098, n49099 );
nor U99182 ( n49099, n49100, n49101 );
nor U99183 ( n49098, n49104, n49105 );
nor U99184 ( n49100, n48051, n49086 );
nand U99185 ( n15066, n49004, n49005 );
nor U99186 ( n49005, n49006, n49007 );
nor U99187 ( n49004, n49010, n49011 );
nor U99188 ( n49006, n48051, n48991 );
nand U99189 ( n15106, n48921, n48922 );
nor U99190 ( n48922, n48923, n48924 );
nor U99191 ( n48921, n48927, n48928 );
nor U99192 ( n48923, n48051, n48892 );
nand U99193 ( n15226, n48638, n48639 );
nor U99194 ( n48639, n48640, n48641 );
nor U99195 ( n48638, n48644, n48645 );
nor U99196 ( n48640, n48051, n48625 );
nand U99197 ( n15266, n48544, n48545 );
nor U99198 ( n48545, n48546, n48547 );
nor U99199 ( n48544, n48550, n48551 );
nor U99200 ( n48546, n48051, n48531 );
nand U99201 ( n14986, n49193, n49194 );
nor U99202 ( n49194, n49195, n49196 );
nor U99203 ( n49193, n49199, n49200 );
nand U99204 ( n49196, n49197, n49198 );
nand U99205 ( n15146, n48824, n48825 );
nor U99206 ( n48825, n48826, n48827 );
nor U99207 ( n48824, n48830, n48831 );
nand U99208 ( n48827, n48828, n48829 );
xor U99209 ( n49782, n49788, n49789 );
or U99210 ( n49788, n49982, n73400 );
xor U99211 ( n49789, n49790, n49791 );
nand U99212 ( n49791, n49792, n49793 );
or U99213 ( n51305, n51409, n51410 );
and U99214 ( n53143, n53234, n8229 );
nor U99215 ( n53234, n73017, n73419 );
nor U99216 ( n17364, n17365, n17366 );
xor U99217 ( n51201, n51202, n51203 );
nand U99218 ( n18503, n18649, n18650 );
nand U99219 ( n18650, n18651, n18521 );
nand U99220 ( n18649, n18654, n18519 );
xor U99221 ( n18651, n18652, n18653 );
nor U99222 ( n18654, n18521, n18522 );
xnor U99223 ( n19497, n19644, n19645 );
xnor U99224 ( n19644, n19646, n19647 );
xor U99225 ( n51408, n51409, n51410 );
nor U99226 ( n51774, n51765, n52119 );
and U99227 ( n52119, n52120, n51766 );
nand U99228 ( n52120, n1303, n51771 );
nand U99229 ( n51059, n1742, n51291 );
nor U99230 ( n20912, n75913, n18105 );
nand U99231 ( n50971, n51203, n51202 );
nand U99232 ( n8571, n15309, n15310 );
nor U99233 ( n15309, n15318, n15319 );
nor U99234 ( n15310, n15312, n15313 );
nor U99235 ( n15318, n14859, n15297 );
nand U99236 ( n8611, n15197, n15198 );
nor U99237 ( n15197, n15204, n15205 );
nor U99238 ( n15198, n15199, n15200 );
nor U99239 ( n15204, n14854, n15185 );
nand U99240 ( n8651, n15095, n15097 );
nor U99241 ( n15095, n15103, n15104 );
nor U99242 ( n15097, n15098, n15099 );
nor U99243 ( n15103, n14854, n15078 );
nand U99244 ( n8691, n14985, n14987 );
nor U99245 ( n14985, n14993, n14994 );
nor U99246 ( n14987, n14988, n14989 );
nor U99247 ( n14993, n14854, n14974 );
nand U99248 ( n51307, n51410, n51409 );
nand U99249 ( n17895, n17970, n17969 );
and U99250 ( n10057, n10058, n9894 );
nand U99251 ( n9566, n10013, n10014 );
nor U99252 ( n10014, n10015, n10016 );
nor U99253 ( n10013, n10056, n10057 );
nor U99254 ( n10015, n9487, n76632 );
nand U99255 ( n8731, n14847, n14848 );
nor U99256 ( n14847, n14855, n14857 );
nor U99257 ( n14848, n14849, n14850 );
nor U99258 ( n14855, n14830, n14859 );
nand U99259 ( n17516, n17784, n17783 );
nand U99260 ( n51095, n51190, n51189 );
nor U99261 ( n51765, n51771, n1303 );
or U99262 ( n50391, n50670, n50671 );
nor U99263 ( n52300, n53947, n1345 );
nand U99264 ( n18525, n18640, n18639 );
xor U99265 ( n50669, n50670, n50671 );
or U99266 ( n17514, n17783, n17784 );
not U99267 ( n1709, n52001 );
nand U99268 ( n51601, n52006, n52007 );
nand U99269 ( n52007, n52008, n1709 );
nor U99270 ( n52008, n52009, n73401 );
nand U99271 ( n18519, n18653, n18655 );
xnor U99272 ( n18367, n18448, n18264 );
xor U99273 ( n18448, n18266, n18267 );
nand U99274 ( n18266, n18537, n18538 );
or U99275 ( n18537, n18541, n18542 );
nand U99276 ( n18538, n18539, n18540 );
nand U99277 ( n18539, n18541, n18542 );
nand U99278 ( n50393, n50671, n50670 );
nand U99279 ( n15311, n48434, n48435 );
nor U99280 ( n48434, n48441, n48442 );
nor U99281 ( n48435, n48436, n48437 );
nor U99282 ( n48441, n48044, n48433 );
nor U99283 ( n51608, n52000, n1708 );
not U99284 ( n1724, n51996 );
nand U99285 ( n15351, n48351, n48352 );
nor U99286 ( n48351, n48357, n48358 );
nor U99287 ( n48352, n48353, n48354 );
nor U99288 ( n48357, n48040, n48350 );
nand U99289 ( n15391, n48254, n48255 );
nor U99290 ( n48254, n48260, n48261 );
nor U99291 ( n48255, n48256, n48257 );
nor U99292 ( n48260, n48040, n48253 );
nand U99293 ( n15431, n48156, n48157 );
nor U99294 ( n48156, n48162, n48163 );
nor U99295 ( n48157, n48158, n48159 );
nor U99296 ( n48162, n48040, n48155 );
nand U99297 ( n53860, n53861, n53862 );
nor U99298 ( n52009, n52455, n1700 );
not U99299 ( n1710, n52451 );
nand U99300 ( n50826, n51006, n51005 );
xnor U99301 ( n17505, n17254, n17513 );
xor U99302 ( n17513, n17253, n17255 );
nand U99303 ( n17242, n17505, n17504 );
or U99304 ( n50332, n50381, n50382 );
nand U99305 ( n15471, n48034, n48035 );
nor U99306 ( n48034, n48041, n48042 );
nor U99307 ( n48035, n48036, n48037 );
nor U99308 ( n48041, n48032, n48044 );
or U99309 ( n18523, n18639, n18640 );
nor U99310 ( n18109, n18335, n18331 );
nand U99311 ( n17832, n18106, n18107 );
nand U99312 ( n18107, n18108, n2858 );
not U99313 ( n2858, n18109 );
xor U99314 ( n50380, n50381, n50382 );
nand U99315 ( n50334, n50382, n50381 );
or U99316 ( n50824, n51005, n51006 );
nand U99317 ( n52294, n52293, n52295 );
or U99318 ( n17240, n17504, n17505 );
nor U99319 ( n52892, n49930, n73005 );
xor U99320 ( n18638, n18639, n18640 );
nand U99321 ( n50164, n50447, n50446 );
nand U99322 ( n19506, n21034, n21035 );
or U99323 ( n21034, n21023, n21025 );
nand U99324 ( n21035, n21024, n21036 );
nand U99325 ( n21036, n21025, n21023 );
nor U99326 ( n21060, n21061, n2465 );
nand U99327 ( n21063, n21089, n21090 );
nand U99328 ( n21089, n21050, n21049 );
nand U99329 ( n21090, n21051, n21091 );
or U99330 ( n21091, n21049, n21050 );
nor U99331 ( n21056, n21057, n21058 );
nor U99332 ( n21057, n21059, n21060 );
and U99333 ( n21059, n21061, n2465 );
nand U99334 ( n21097, n76589, n21098 );
nand U99335 ( n21098, n76654, n75919 );
xor U99336 ( n17782, n17783, n17784 );
and U99337 ( n52999, n53134, n8229 );
nor U99338 ( n53134, n73419, n73019 );
nor U99339 ( n50294, n49898, n73014 );
nand U99340 ( n53238, n76649, n73413 );
nand U99341 ( n52117, n52118, n52113 );
nor U99342 ( n17576, n73409, n76575 );
nor U99343 ( n51482, n49930, n73416 );
nand U99344 ( n54044, n54039, n53985 );
nand U99345 ( n19139, n19138, n19140 );
nor U99346 ( n53949, n53950, n52298 );
nor U99347 ( n53950, n53951, n52301 );
and U99348 ( n53951, n53947, n1305 );
nand U99349 ( n21072, n21067, n19784 );
xnor U99350 ( n16498, n18845, n18846 );
xor U99351 ( n18845, n18847, n18848 );
or U99352 ( n50162, n50446, n50447 );
xor U99353 ( n50958, n50959, n50960 );
or U99354 ( n50693, n50959, n50960 );
nand U99355 ( n8451, n15630, n15632 );
nor U99356 ( n15630, n15638, n15639 );
nor U99357 ( n15632, n15633, n15634 );
nor U99358 ( n15638, n14735, n14854 );
or U99359 ( n18353, n18453, n18454 );
nor U99360 ( n54001, n54002, n1307 );
nand U99361 ( n54004, n54020, n54024 );
nand U99362 ( n54024, n54018, n54019 );
nand U99363 ( n54031, n76323, n54032 );
nand U99364 ( n54032, n76653, n73424 );
or U99365 ( n54019, n54025, n54026 );
nand U99366 ( n8171, n16358, n16359 );
nor U99367 ( n16359, n16360, n16362 );
nor U99368 ( n16358, n16365, n16367 );
nor U99369 ( n16360, n14854, n16342 );
nand U99370 ( n8211, n16253, n16254 );
nor U99371 ( n16254, n16255, n16257 );
nor U99372 ( n16253, n16260, n16262 );
nor U99373 ( n16255, n14854, n16237 );
nand U99374 ( n8291, n16050, n16052 );
nor U99375 ( n16052, n16053, n16054 );
nor U99376 ( n16050, n16058, n16059 );
nor U99377 ( n16053, n14854, n16034 );
nand U99378 ( n8331, n15943, n15944 );
nor U99379 ( n15944, n15945, n15947 );
nor U99380 ( n15943, n15950, n15952 );
nor U99381 ( n15945, n14854, n15927 );
nand U99382 ( n8371, n15838, n15839 );
nor U99383 ( n15839, n15840, n15842 );
nor U99384 ( n15838, n15845, n15847 );
nor U99385 ( n15840, n14854, n15822 );
nand U99386 ( n8491, n15529, n15530 );
nor U99387 ( n15530, n15532, n15533 );
nor U99388 ( n15529, n15537, n15538 );
nor U99389 ( n15532, n14854, n15513 );
nand U99390 ( n8531, n15423, n15424 );
nor U99391 ( n15424, n15425, n15427 );
nor U99392 ( n15423, n15430, n15432 );
nor U99393 ( n15425, n14854, n15407 );
nand U99394 ( n8251, n16153, n16154 );
nor U99395 ( n16154, n16155, n16157 );
nor U99396 ( n16153, n16160, n16162 );
nand U99397 ( n16157, n16158, n16159 );
nand U99398 ( n8411, n15728, n15729 );
nor U99399 ( n15729, n15730, n15732 );
nor U99400 ( n15728, n15735, n15737 );
nand U99401 ( n15732, n15733, n15734 );
nand U99402 ( n51605, n1708, n52000 );
nand U99403 ( n50695, n50960, n50959 );
nand U99404 ( n18090, n18326, n18327 );
nand U99405 ( n18327, n18108, n18328 );
nand U99406 ( n18326, n18334, n18106 );
nand U99407 ( n18328, n18329, n18330 );
nor U99408 ( n18334, n18108, n18109 );
xor U99409 ( n18452, n18453, n18454 );
nand U99410 ( n17892, n17991, n17992 );
nand U99411 ( n17992, n17993, n17994 );
nor U99412 ( n17991, n17995, n17996 );
or U99413 ( n50518, n76322, n73415 );
nand U99414 ( n52006, n1700, n52455 );
nand U99415 ( n18355, n18454, n18453 );
buf U99416 ( n76318, n49931 );
nor U99417 ( n20601, n73408, n18105 );
xor U99418 ( n50976, n51212, n51089 );
xor U99419 ( n51212, n51091, n51092 );
xnor U99420 ( n21058, n21099, n21077 );
xnor U99421 ( n21099, n21078, n21075 );
nor U99422 ( n21054, n21061, n2503 );
nor U99423 ( n17977, n2550, n17983 );
nand U99424 ( n17983, n17047, n17052 );
nand U99425 ( n53138, n76649, n73017 );
xor U99426 ( n53999, n54033, n54034 );
xor U99427 ( n54034, n54035, n54036 );
nor U99428 ( n53995, n54002, n1349 );
nand U99429 ( n15191, n48723, n48724 );
nor U99430 ( n48723, n48729, n48730 );
nor U99431 ( n48724, n48725, n48726 );
nor U99432 ( n48729, n47941, n48040 );
and U99433 ( n52993, n53975, n8229 );
nor U99434 ( n53975, n73019, n73421 );
not U99435 ( n2882, n17366 );
or U99436 ( n18136, n18233, n18234 );
or U99437 ( n18011, n18250, n18251 );
nand U99438 ( n14951, n49281, n49282 );
nor U99439 ( n49282, n49283, n49284 );
nor U99440 ( n49281, n49287, n49288 );
nor U99441 ( n49283, n48040, n49276 );
nand U99442 ( n15031, n49090, n49091 );
nor U99443 ( n49091, n49092, n49093 );
nor U99444 ( n49090, n49096, n49097 );
nor U99445 ( n49092, n48040, n49086 );
nand U99446 ( n15071, n48996, n48997 );
nor U99447 ( n48997, n48998, n48999 );
nor U99448 ( n48996, n49002, n49003 );
nor U99449 ( n48998, n48040, n48991 );
nand U99450 ( n15111, n48897, n48898 );
nor U99451 ( n48898, n48899, n48900 );
nor U99452 ( n48897, n48903, n48904 );
nor U99453 ( n48899, n48040, n48892 );
nand U99454 ( n15231, n48630, n48631 );
nor U99455 ( n48631, n48632, n48633 );
nor U99456 ( n48630, n48636, n48637 );
nor U99457 ( n48632, n48040, n48625 );
nand U99458 ( n15271, n48536, n48537 );
nor U99459 ( n48537, n48538, n48539 );
nor U99460 ( n48536, n48542, n48543 );
nor U99461 ( n48538, n48040, n48531 );
nand U99462 ( n14911, n49359, n49360 );
nor U99463 ( n49360, n49361, n49362 );
nor U99464 ( n49359, n49365, n49366 );
nor U99465 ( n49361, n48040, n49354 );
nand U99466 ( n14991, n49185, n49186 );
nor U99467 ( n49186, n49187, n49188 );
nor U99468 ( n49185, n49191, n49192 );
nand U99469 ( n49188, n49189, n49190 );
nand U99470 ( n15151, n48816, n48817 );
nor U99471 ( n48817, n48818, n48819 );
nor U99472 ( n48816, n48822, n48823 );
nand U99473 ( n48819, n48820, n48821 );
nand U99474 ( n51079, n51226, n51225 );
nand U99475 ( n53876, n53882, n76648 );
nor U99476 ( n53882, n53883, n73403 );
nand U99477 ( n18106, n18331, n18335 );
xor U99478 ( n18249, n18250, n18251 );
xor U99479 ( n18232, n18233, n18234 );
nand U99480 ( n51285, n51288, n51289 );
nand U99481 ( n51474, n51480, n76648 );
nor U99482 ( n51480, n51481, n73016 );
xor U99483 ( n17503, n17504, n17505 );
xnor U99484 ( n19505, n21064, n19643 );
xnor U99485 ( n21064, n19640, n19642 );
or U99486 ( n51077, n51225, n51226 );
nand U99487 ( n18013, n18251, n18250 );
nand U99488 ( n54020, n54026, n54025 );
xor U99489 ( n50842, n50701, n50973 );
xnor U99490 ( n50973, n50704, n50703 );
nand U99491 ( n18138, n18234, n18233 );
nor U99492 ( n18818, n18809, n19163 );
and U99493 ( n19163, n19164, n18810 );
nand U99494 ( n19164, n2419, n18815 );
and U99495 ( n44018, n44019, n43797 );
nand U99496 ( n52884, n52890, n76649 );
nor U99497 ( n52890, n52891, n73401 );
nor U99498 ( n51995, n1708, n51996 );
and U99499 ( n16502, n18738, n18739 );
or U99500 ( n18738, n16458, n16457 );
nand U99501 ( n18739, n16459, n18740 );
nand U99502 ( n18740, n16457, n16458 );
nor U99503 ( n18809, n18815, n2419 );
nor U99504 ( n52450, n1700, n52451 );
nand U99505 ( n53831, n53835, n76648 );
nor U99506 ( n53835, n53836, n73005 );
xor U99507 ( n50445, n50446, n50447 );
or U99508 ( n17436, n17715, n17716 );
xor U99509 ( n45513, n51797, n51798 );
xor U99510 ( n51797, n51799, n51800 );
xor U99511 ( n17714, n17715, n17716 );
xor U99512 ( n16827, n16833, n16834 );
or U99513 ( n16833, n17028, n73404 );
xor U99514 ( n16834, n16835, n16836 );
nand U99515 ( n16836, n16837, n16838 );
nand U99516 ( n17438, n17716, n17715 );
xor U99517 ( n51004, n51005, n51006 );
nand U99518 ( n17595, n17771, n17770 );
nand U99519 ( n45515, n51712, n51713 );
nand U99520 ( n51712, n45503, n45502 );
nand U99521 ( n51713, n45504, n51714 );
or U99522 ( n51714, n45502, n45503 );
nor U99523 ( n51785, n51786, n51787 );
nor U99524 ( n51786, n51788, n51789 );
and U99525 ( n51788, n51790, n1259 );
nand U99526 ( n53979, n76650, n73419 );
nand U99527 ( n17867, n18048, n18047 );
nor U99528 ( n19057, n19370, n19366 );
or U99529 ( n17593, n17770, n17771 );
nor U99530 ( n20787, n73404, n76576 );
buf U99531 ( n76576, n76574 );
nand U99532 ( n21062, n21061, n21063 );
nand U99533 ( n17218, n17492, n17491 );
or U99534 ( n17865, n18047, n18048 );
not U99535 ( n8227, n50508 );
not U99536 ( n1747, n49887 );
not U99537 ( n1742, n51289 );
xnor U99538 ( n49467, n49468, n49469 );
nand U99539 ( n15316, n48420, n48421 );
nor U99540 ( n48420, n48430, n48431 );
nor U99541 ( n48421, n48422, n48423 );
nor U99542 ( n48430, n48033, n48433 );
nand U99543 ( n15356, n48338, n48339 );
nor U99544 ( n48338, n48347, n48348 );
nor U99545 ( n48339, n48340, n48341 );
nor U99546 ( n48347, n48027, n48350 );
nand U99547 ( n15396, n48241, n48242 );
nor U99548 ( n48241, n48250, n48251 );
nor U99549 ( n48242, n48243, n48244 );
nor U99550 ( n48250, n48027, n48253 );
nand U99551 ( n15436, n48143, n48144 );
nor U99552 ( n48143, n48152, n48153 );
nor U99553 ( n48144, n48145, n48146 );
nor U99554 ( n48152, n48027, n48155 );
nor U99555 ( n21002, n21003, n2424 );
nand U99556 ( n21005, n21021, n21039 );
nand U99557 ( n21039, n21019, n21020 );
nand U99558 ( n21046, n76589, n21047 );
nand U99559 ( n21047, n76654, n73022 );
or U99560 ( n21020, n21040, n21041 );
nand U99561 ( n17127, n17427, n17426 );
nand U99562 ( n19161, n19162, n19157 );
nand U99563 ( n15476, n48018, n48019 );
nor U99564 ( n48018, n48028, n48029 );
nor U99565 ( n48019, n48020, n48021 );
nor U99566 ( n48028, n48032, n48033 );
nor U99567 ( n18664, n19048, n19044 );
xor U99568 ( n19027, n19028, n19029 );
nand U99569 ( n53952, n53947, n52299 );
xor U99570 ( n18000, n18001, n18002 );
or U99571 ( n17885, n18001, n18002 );
nand U99572 ( n18667, n19029, n19028 );
or U99573 ( n18665, n19028, n19029 );
and U99574 ( n53970, n54056, n8229 );
nor U99575 ( n54056, n73421, n73021 );
nand U99576 ( n18645, n19054, n19055 );
nand U99577 ( n19055, n19056, n2826 );
nor U99578 ( n19056, n19057, n73407 );
xor U99579 ( n49799, n49805, n49806 );
xor U99580 ( n49805, n49814, n49815 );
xor U99581 ( n49806, n49807, n49808 );
nor U99582 ( n49815, n73397, n49816 );
or U99583 ( n17216, n17491, n17492 );
nor U99584 ( n53940, n53941, n1263 );
nor U99585 ( n53997, n53998, n53999 );
nor U99586 ( n53998, n54000, n54001 );
and U99587 ( n54000, n54002, n1307 );
and U99588 ( n50104, n50422, n50423 );
nand U99589 ( n50422, n50427, n50426 );
nand U99590 ( n50423, n50424, n50425 );
or U99591 ( n50425, n50426, n50427 );
or U99592 ( n50321, n50399, n50400 );
nand U99593 ( n17887, n18002, n18001 );
xor U99594 ( n51224, n51225, n51226 );
nand U99595 ( n51286, n1742, n51287 );
nand U99596 ( n50140, n50434, n50433 );
xor U99597 ( n17769, n17770, n17771 );
xor U99598 ( n50398, n50399, n50400 );
nor U99599 ( n20739, n75911, n76576 );
or U99600 ( n17125, n17426, n17427 );
nand U99601 ( n50556, n50717, n50716 );
nand U99602 ( n18122, n18274, n18273 );
nor U99603 ( n20899, n73009, n76577 );
buf U99604 ( n76577, n76574 );
nand U99605 ( n19054, n19366, n19370 );
nor U99606 ( n19362, n73407, n19049 );
nand U99607 ( n50323, n50400, n50399 );
nand U99608 ( n8576, n15298, n15299 );
nor U99609 ( n15298, n15307, n15308 );
nor U99610 ( n15299, n15300, n15302 );
nor U99611 ( n15307, n14845, n15297 );
nor U99612 ( n53934, n53941, n1304 );
nand U99613 ( n8616, n15187, n15188 );
nor U99614 ( n15187, n15194, n15195 );
nor U99615 ( n15188, n15189, n15190 );
nor U99616 ( n15194, n14840, n15185 );
nand U99617 ( n8656, n15085, n15087 );
nor U99618 ( n15085, n15093, n15094 );
nor U99619 ( n15087, n15088, n15089 );
nor U99620 ( n15093, n14840, n15078 );
nand U99621 ( n8696, n14975, n14977 );
nor U99622 ( n14975, n14983, n14984 );
nor U99623 ( n14977, n14978, n14979 );
nor U99624 ( n14983, n14840, n14974 );
xor U99625 ( n17425, n17426, n17427 );
or U99626 ( n17844, n73013, n76577 );
or U99627 ( n50554, n50716, n50717 );
nand U99628 ( n8736, n14833, n14834 );
nor U99629 ( n14833, n14842, n14843 );
nor U99630 ( n14834, n14835, n14837 );
nor U99631 ( n14842, n14830, n14845 );
xor U99632 ( n18132, n18260, n18126 );
xor U99633 ( n18260, n18128, n18129 );
or U99634 ( n18120, n18273, n18274 );
xnor U99635 ( n21000, n21048, n21049 );
xnor U99636 ( n21048, n21050, n21051 );
nor U99637 ( n20996, n21003, n2467 );
or U99638 ( n50138, n50433, n50434 );
nand U99639 ( n21021, n21041, n21040 );
and U99640 ( n10113, n10114, n9894 );
nor U99641 ( n51994, n51997, n51998 );
nand U99642 ( n20792, n8222, n73406 );
not U99643 ( n8233, n49898 );
nor U99644 ( n52449, n52452, n52453 );
nand U99645 ( n50710, n51087, n51088 );
nand U99646 ( n51087, n51092, n51091 );
nand U99647 ( n51088, n51089, n51090 );
or U99648 ( n51090, n51091, n51092 );
nand U99649 ( n18661, n19044, n19048 );
nor U99650 ( n18097, n75916, n76575 );
nand U99651 ( n54060, n76650, n73019 );
nor U99652 ( n19040, n73398, n19049 );
not U99653 ( n1569, n53545 );
xor U99654 ( n53925, n54017, n54018 );
nand U99655 ( n54017, n54019, n54020 );
nor U99656 ( n53918, n53924, n53925 );
nor U99657 ( n50514, n76321, n73016 );
buf U99658 ( n76321, n76320 );
and U99659 ( n44064, n44065, n43797 );
nand U99660 ( n16291, n44021, n44022 );
nor U99661 ( n44022, n44023, n44024 );
nor U99662 ( n44021, n44063, n44064 );
nor U99663 ( n44023, n43467, n76362 );
nor U99664 ( n20920, n75913, n76576 );
xnor U99665 ( n17883, n18015, n17742 );
xor U99666 ( n18015, n17744, n17745 );
not U99667 ( n1603, n53689 );
xor U99668 ( n50715, n50716, n50717 );
nor U99669 ( n20861, n73414, n76577 );
xor U99670 ( n17490, n17491, n17492 );
not U99671 ( n1589, n53621 );
nand U99672 ( n15196, n48712, n48713 );
nor U99673 ( n48712, n48720, n48721 );
nor U99674 ( n48713, n48714, n48715 );
nor U99675 ( n48720, n47941, n48027 );
nand U99676 ( n20904, n8222, n75911 );
nand U99677 ( n50567, n50699, n50700 );
nand U99678 ( n50699, n50704, n50703 );
nand U99679 ( n50700, n50701, n50702 );
or U99680 ( n50702, n50703, n50704 );
nand U99681 ( n14916, n49347, n49348 );
nor U99682 ( n49348, n49349, n49350 );
nor U99683 ( n49347, n49355, n49356 );
nor U99684 ( n49349, n48027, n49354 );
nand U99685 ( n14956, n49269, n49270 );
nor U99686 ( n49270, n49271, n49272 );
nor U99687 ( n49269, n49277, n49278 );
nor U99688 ( n49271, n48027, n49276 );
nand U99689 ( n15036, n49079, n49080 );
nor U99690 ( n49080, n49081, n49082 );
nor U99691 ( n49079, n49087, n49088 );
nor U99692 ( n49081, n48027, n49086 );
nand U99693 ( n15076, n48984, n48985 );
nor U99694 ( n48985, n48986, n48987 );
nor U99695 ( n48984, n48992, n48993 );
nor U99696 ( n48986, n48027, n48991 );
nand U99697 ( n15116, n48885, n48886 );
nor U99698 ( n48886, n48887, n48888 );
nor U99699 ( n48885, n48893, n48894 );
nor U99700 ( n48887, n48027, n48892 );
nand U99701 ( n15236, n48618, n48619 );
nor U99702 ( n48619, n48620, n48621 );
nor U99703 ( n48618, n48626, n48627 );
nor U99704 ( n48620, n48027, n48625 );
nand U99705 ( n15276, n48524, n48525 );
nor U99706 ( n48525, n48526, n48527 );
nor U99707 ( n48524, n48532, n48533 );
nor U99708 ( n48526, n48027, n48531 );
nand U99709 ( n14996, n49173, n49174 );
nor U99710 ( n49174, n49175, n49176 );
nor U99711 ( n49173, n49181, n49182 );
nand U99712 ( n49176, n49177, n49178 );
nand U99713 ( n15156, n48804, n48805 );
nor U99714 ( n48805, n48806, n48807 );
nor U99715 ( n48804, n48812, n48813 );
nand U99716 ( n48807, n48808, n48809 );
nand U99717 ( n51462, n51605, n51606 );
nand U99718 ( n51606, n51607, n1709 );
nor U99719 ( n51607, n51608, n73411 );
nand U99720 ( n11713, n18774, n18775 );
nand U99721 ( n18774, n11702, n11699 );
nand U99722 ( n18775, n11700, n18776 );
or U99723 ( n18776, n11699, n11702 );
nor U99724 ( n18829, n18830, n18831 );
nor U99725 ( n18830, n18832, n18833 );
and U99726 ( n18832, n18834, n2374 );
and U99727 ( n11742, n18756, n18757 );
nand U99728 ( n18756, n11725, n11724 );
nand U99729 ( n18757, n11727, n18758 );
or U99730 ( n18758, n11724, n11725 );
xnor U99731 ( n50418, n50697, n50424 );
xor U99732 ( n50697, n50426, n50427 );
nand U99733 ( n51791, n51790, n51792 );
nor U99734 ( n19939, n73011, n18105 );
not U99735 ( n1708, n51997 );
nor U99736 ( n50523, n49898, n73415 );
nand U99737 ( n50128, n50558, n50559 );
nand U99738 ( n50558, n50562, n50563 );
nand U99739 ( n50559, n50560, n50561 );
or U99740 ( n50561, n50562, n50563 );
nor U99741 ( n53923, n53924, n1264 );
nand U99742 ( n53927, n53915, n54007 );
nand U99743 ( n54007, n53913, n53914 );
nand U99744 ( n54015, n76323, n54016 );
nand U99745 ( n54016, n76653, n73426 );
or U99746 ( n53914, n54008, n54009 );
not U99747 ( n1700, n52452 );
nand U99748 ( n49235, n49236, n49237 );
nor U99749 ( n49237, n49238, n49239 );
nor U99750 ( n49236, n49249, n49250 );
nor U99751 ( n49239, n48122, n49240 );
nand U99752 ( n48866, n48867, n48868 );
nor U99753 ( n48868, n48869, n48870 );
nor U99754 ( n48867, n48880, n48881 );
nor U99755 ( n48870, n48122, n48871 );
nor U99756 ( n48305, n48317, n48318 );
nor U99757 ( n48317, n48122, n48253 );
nor U99758 ( n48318, n48136, n48252 );
xor U99759 ( n18046, n18047, n18048 );
nand U99760 ( n51613, n51619, n76648 );
nor U99761 ( n51619, n51620, n73416 );
nand U99762 ( n8456, n15620, n15622 );
nor U99763 ( n15620, n15628, n15629 );
nor U99764 ( n15622, n15623, n15624 );
nor U99765 ( n15628, n14735, n14840 );
nand U99766 ( n8176, n16348, n16349 );
nor U99767 ( n16349, n16350, n16352 );
nor U99768 ( n16348, n16355, n16357 );
nor U99769 ( n16350, n14840, n16342 );
nand U99770 ( n8216, n16243, n16244 );
nor U99771 ( n16244, n16245, n16247 );
nor U99772 ( n16243, n16250, n16252 );
nor U99773 ( n16245, n14840, n16237 );
nand U99774 ( n8296, n16040, n16042 );
nor U99775 ( n16042, n16043, n16044 );
nor U99776 ( n16040, n16048, n16049 );
nor U99777 ( n16043, n14840, n16034 );
nand U99778 ( n8336, n15933, n15934 );
nor U99779 ( n15934, n15935, n15937 );
nor U99780 ( n15933, n15940, n15942 );
nor U99781 ( n15935, n14840, n15927 );
nand U99782 ( n8376, n15828, n15829 );
nor U99783 ( n15829, n15830, n15832 );
nor U99784 ( n15828, n15835, n15837 );
nor U99785 ( n15830, n14840, n15822 );
nand U99786 ( n8496, n15519, n15520 );
nor U99787 ( n15520, n15522, n15523 );
nor U99788 ( n15519, n15527, n15528 );
nor U99789 ( n15522, n14840, n15513 );
nand U99790 ( n8536, n15413, n15414 );
nor U99791 ( n15414, n15415, n15417 );
nor U99792 ( n15413, n15420, n15422 );
nor U99793 ( n15415, n14840, n15407 );
nand U99794 ( n8256, n16143, n16144 );
nor U99795 ( n16144, n16145, n16147 );
nor U99796 ( n16143, n16150, n16152 );
nand U99797 ( n16147, n16148, n16149 );
nand U99798 ( n8416, n15718, n15719 );
nor U99799 ( n15719, n15720, n15722 );
nor U99800 ( n15718, n15725, n15727 );
nand U99801 ( n15722, n15723, n15724 );
xor U99802 ( n18272, n18273, n18274 );
and U99803 ( n54035, n54048, n8229 );
nor U99804 ( n54048, n73021, n73424 );
xnor U99805 ( n50708, n50981, n50836 );
xnor U99806 ( n50981, n50837, n50834 );
nand U99807 ( n17599, n17758, n17757 );
nor U99808 ( n51037, n76321, n73416 );
nand U99809 ( n17871, n18035, n18034 );
nand U99810 ( n18021, n18262, n18263 );
nand U99811 ( n18262, n18267, n18266 );
nand U99812 ( n18263, n18264, n18265 );
or U99813 ( n18265, n18266, n18267 );
nand U99814 ( n50439, n50832, n50833 );
or U99815 ( n50832, n50836, n50837 );
nand U99816 ( n50833, n50834, n50835 );
nand U99817 ( n50835, n50836, n50837 );
or U99818 ( n53549, n76322, n73008 );
and U99819 ( n17158, n17467, n17468 );
nand U99820 ( n17467, n17472, n17471 );
nand U99821 ( n17468, n17469, n17470 );
or U99822 ( n17470, n17471, n17472 );
or U99823 ( n17132, n17444, n17445 );
or U99824 ( n17597, n17757, n17758 );
nand U99825 ( n20925, n8222, n73404 );
nor U99826 ( n18518, n73000, n18105 );
nand U99827 ( n20744, n8222, n73408 );
nor U99828 ( n20911, n73012, n76576 );
xor U99829 ( n17443, n17444, n17445 );
nor U99830 ( n20830, n73015, n76576 );
xnor U99831 ( n11738, n18841, n18842 );
xor U99832 ( n18841, n18843, n18844 );
nand U99833 ( n54003, n54002, n54004 );
or U99834 ( n53693, n76322, n73003 );
nand U99835 ( n17134, n17445, n17444 );
nand U99836 ( n17194, n17479, n17478 );
xor U99837 ( n11710, n18837, n18838 );
xor U99838 ( n18837, n18839, n18840 );
nand U99839 ( n20865, n8222, n75913 );
xnor U99840 ( n50105, n50428, n50114 );
xor U99841 ( n50428, n50116, n50117 );
nand U99842 ( n53915, n54009, n54008 );
xnor U99843 ( n50568, n50562, n50705 );
xnor U99844 ( n50705, n50560, n50563 );
xor U99845 ( n50432, n50433, n50434 );
or U99846 ( n17869, n18034, n18035 );
not U99847 ( n2826, n19049 );
nor U99848 ( n20998, n20999, n21000 );
nor U99849 ( n20999, n21001, n21002 );
and U99850 ( n21001, n21003, n2424 );
nand U99851 ( n20986, n20991, n20992 );
or U99852 ( n20991, n20974, n20973 );
nand U99853 ( n20992, n20975, n20993 );
nand U99854 ( n20993, n20973, n20974 );
xnor U99855 ( n18022, n18268, n18029 );
xnor U99856 ( n18268, n18030, n18027 );
nor U99857 ( n53748, n49898, n73400 );
or U99858 ( n17192, n17478, n17479 );
buf U99859 ( n76583, n76584 );
xor U99860 ( n16844, n16850, n16851 );
xor U99861 ( n16850, n16859, n16860 );
xor U99862 ( n16851, n16852, n16853 );
nor U99863 ( n16860, n73406, n16861 );
xor U99864 ( n17756, n17757, n17758 );
or U99865 ( n18329, n18333, n18331 );
xnor U99866 ( n20982, n21022, n21023 );
xnor U99867 ( n21022, n21024, n21025 );
nand U99868 ( n17751, n18124, n18125 );
nand U99869 ( n18124, n18129, n18128 );
nand U99870 ( n18125, n18126, n18127 );
or U99871 ( n18127, n18128, n18129 );
nor U99872 ( n53357, n76321, n73413 );
nand U99873 ( n54052, n76650, n73421 );
and U99874 ( n20037, n21086, n8220 );
nor U99875 ( n21086, n73020, n73420 );
nand U99876 ( n17764, n18025, n18026 );
or U99877 ( n18025, n18029, n18030 );
nand U99878 ( n18026, n18027, n18028 );
nand U99879 ( n18028, n18029, n18030 );
xnor U99880 ( n16469, n16470, n16472 );
nand U99881 ( n8581, n15280, n15282 );
nor U99882 ( n15280, n15293, n15294 );
nor U99883 ( n15282, n15283, n15284 );
nor U99884 ( n15293, n14832, n15297 );
nand U99885 ( n8621, n15170, n15172 );
nor U99886 ( n15170, n15182, n15183 );
nor U99887 ( n15172, n15173, n15174 );
nor U99888 ( n15182, n14824, n15185 );
nand U99889 ( n8661, n15063, n15064 );
nor U99890 ( n15063, n15074, n15075 );
nor U99891 ( n15064, n15065, n15067 );
nor U99892 ( n15074, n14824, n15078 );
nand U99893 ( n8701, n14959, n14960 );
nor U99894 ( n14959, n14970, n14972 );
nor U99895 ( n14960, n14962, n14963 );
nor U99896 ( n14970, n14824, n14974 );
nand U99897 ( n17610, n17740, n17741 );
nand U99898 ( n17740, n17745, n17744 );
nand U99899 ( n17741, n17742, n17743 );
or U99900 ( n17743, n17744, n17745 );
nor U99901 ( n53464, n49898, n73412 );
nand U99902 ( n8741, n14813, n14814 );
nor U99903 ( n14813, n14825, n14827 );
nor U99904 ( n14814, n14815, n14817 );
nor U99905 ( n14825, n14830, n14832 );
xor U99906 ( n17463, n17738, n17469 );
xor U99907 ( n17738, n17471, n17472 );
nand U99908 ( n17182, n17601, n17602 );
nand U99909 ( n17601, n17605, n17606 );
nand U99910 ( n17602, n17603, n17604 );
or U99911 ( n17604, n17605, n17606 );
nor U99912 ( n20484, n73418, n76576 );
nand U99913 ( n20916, n8222, n73009 );
nor U99914 ( n50262, n76316, n73016 );
buf U99915 ( n76316, n76315 );
nand U99916 ( n49994, n50112, n50113 );
nand U99917 ( n50112, n50117, n50116 );
nand U99918 ( n50113, n50114, n50115 );
or U99919 ( n50115, n50116, n50117 );
nand U99920 ( n18835, n18834, n18836 );
xor U99921 ( n20969, n21018, n21019 );
nand U99922 ( n21018, n21020, n21021 );
nor U99923 ( n20962, n20968, n20969 );
or U99924 ( n20663, n73406, n76577 );
nand U99925 ( n20835, n8222, n73012 );
nor U99926 ( n53248, n76321, n73017 );
nor U99927 ( n50809, n49898, n73016 );
and U99928 ( n44111, n44112, n43797 );
nand U99929 ( n16286, n44067, n44068 );
nor U99930 ( n44068, n44069, n44070 );
nor U99931 ( n44067, n44110, n44111 );
nor U99932 ( n44069, n43476, n76362 );
nor U99933 ( n17352, n73409, n16943 );
nand U99934 ( n18502, n18661, n18662 );
nand U99935 ( n18662, n18663, n2826 );
nor U99936 ( n18663, n18664, n73398 );
xnor U99937 ( n17749, n17877, n18017 );
xnor U99938 ( n18017, n17875, n17878 );
nor U99939 ( n20967, n20968, n2379 );
nand U99940 ( n21016, n76589, n21017 );
nand U99941 ( n21017, n76654, n73423 );
nand U99942 ( n20971, n20959, n21008 );
nand U99943 ( n21008, n20957, n20958 );
or U99944 ( n20958, n21009, n21010 );
nand U99945 ( n17484, n17873, n17874 );
nand U99946 ( n17873, n17877, n17878 );
nand U99947 ( n17874, n17875, n17876 );
or U99948 ( n17876, n17877, n17878 );
nor U99949 ( n53487, n76321, n73412 );
xnor U99950 ( n17159, n17473, n17168 );
xor U99951 ( n17473, n17170, n17171 );
xor U99952 ( n18033, n18034, n18035 );
xnor U99953 ( n17611, n17605, n17746 );
xnor U99954 ( n17746, n17603, n17606 );
and U99955 ( n10175, n10177, n9894 );
nand U99956 ( n9556, n10122, n10123 );
nor U99957 ( n10123, n10124, n10125 );
nor U99958 ( n10122, n10174, n10175 );
nor U99959 ( n10124, n9509, n76632 );
nor U99960 ( n54010, n49930, n73426 );
nand U99961 ( n18330, n18331, n18332 );
xor U99962 ( n49839, n49847, n49848 );
xor U99963 ( n49847, n49967, n49968 );
xor U99964 ( n49848, n49849, n49850 );
nor U99965 ( n49968, n73005, n76091 );
xor U99966 ( n49824, n49830, n49831 );
nand U99967 ( n49830, n49974, n49975 );
xor U99968 ( n49831, n49832, n49833 );
nand U99969 ( n49975, n49976, n49977 );
nor U99970 ( n18331, n73417, n76576 );
nand U99971 ( n8461, n15602, n15603 );
nor U99972 ( n15602, n15610, n15612 );
nor U99973 ( n15603, n15604, n15605 );
nor U99974 ( n15610, n14735, n14824 );
nand U99975 ( n54030, n76650, n73021 );
xor U99976 ( n17477, n17478, n17479 );
nand U99977 ( n8181, n16333, n16334 );
nor U99978 ( n16334, n16335, n16337 );
nor U99979 ( n16333, n16343, n16344 );
nor U99980 ( n16335, n14824, n16342 );
nand U99981 ( n8221, n16228, n16229 );
nor U99982 ( n16229, n16230, n16232 );
nor U99983 ( n16228, n16238, n16239 );
nor U99984 ( n16230, n14824, n16237 );
nand U99985 ( n8301, n16025, n16027 );
nor U99986 ( n16027, n16028, n16029 );
nor U99987 ( n16025, n16035, n16037 );
nor U99988 ( n16028, n14824, n16034 );
nand U99989 ( n8341, n15918, n15919 );
nor U99990 ( n15919, n15920, n15922 );
nor U99991 ( n15918, n15928, n15929 );
nor U99992 ( n15920, n14824, n15927 );
nand U99993 ( n8381, n15813, n15814 );
nor U99994 ( n15814, n15815, n15817 );
nor U99995 ( n15813, n15823, n15824 );
nor U99996 ( n15815, n14824, n15822 );
nand U99997 ( n8501, n15504, n15505 );
nor U99998 ( n15505, n15507, n15508 );
nor U99999 ( n15504, n15514, n15515 );
nor U100000 ( n15507, n14824, n15513 );
nand U100001 ( n8541, n15398, n15399 );
nor U100002 ( n15399, n15400, n15402 );
nor U100003 ( n15398, n15408, n15409 );
nor U100004 ( n15400, n14824, n15407 );
nand U100005 ( n8261, n16122, n16123 );
nor U100006 ( n16123, n16124, n16125 );
nor U100007 ( n16122, n16132, n16133 );
nand U100008 ( n16125, n16127, n16128 );
nand U100009 ( n8421, n15703, n15704 );
nor U100010 ( n15704, n15705, n15707 );
nor U100011 ( n15703, n15713, n15714 );
nand U100012 ( n15707, n15708, n15709 );
nand U100013 ( n21004, n21003, n21005 );
nand U100014 ( n20959, n21010, n21009 );
or U100015 ( n53813, n76322, n73397 );
or U100016 ( n53750, n76322, n73400 );
nand U100017 ( n15789, n15790, n15792 );
nor U100018 ( n15792, n15793, n15794 );
nor U100019 ( n15790, n15807, n15808 );
nor U100020 ( n15794, n14934, n15795 );
nand U100021 ( n16205, n16207, n16208 );
nor U100022 ( n16208, n16209, n16210 );
nor U100023 ( n16207, n16223, n16224 );
nor U100024 ( n16210, n14934, n16212 );
nor U100025 ( n15149, n15164, n15165 );
nor U100026 ( n15164, n14934, n15078 );
nor U100027 ( n15165, n14950, n15077 );
or U100028 ( n53587, n76322, n73410 );
nor U100029 ( n51044, n49898, n73416 );
nor U100030 ( n51980, n76321, n73005 );
nand U100031 ( n20491, n8222, n73414 );
nor U100032 ( n53148, n76321, n73419 );
nor U100033 ( n16936, n75916, n76587 );
buf U100034 ( n76587, n76585 );
or U100035 ( n52867, n76322, n73002 );
or U100036 ( n52435, n76322, n73403 );
nand U100037 ( n17040, n17166, n17167 );
nand U100038 ( n17166, n17171, n17170 );
nand U100039 ( n17167, n17168, n17169 );
or U100040 ( n17169, n17170, n17171 );
or U100041 ( n51272, n76322, n73411 );
not U100042 ( n8225, n16943 );
not U100043 ( n2722, n20779 );
not U100044 ( n2707, n20892 );
nor U100045 ( n53016, n76321, n73019 );
nor U100046 ( n52875, n49898, n73002 );
or U100047 ( n53797, n76322, n72999 );
nor U100048 ( n17348, n73013, n16943 );
nor U100049 ( n20593, n73408, n76576 );
nor U100050 ( n51768, n51769, n51770 );
xor U100051 ( n51770, n51766, n51771 );
nor U100052 ( n19366, n73407, n76576 );
nor U100053 ( n50269, n50508, n73016 );
xor U100054 ( n49652, n49654, n49655 );
nor U100055 ( n19931, n73011, n76576 );
nor U100056 ( n18510, n73000, n76575 );
or U100057 ( n50500, n76317, n73416 );
buf U100058 ( n76317, n76315 );
nor U100059 ( n19365, n19366, n19367 );
nor U100060 ( n20187, n73018, n76576 );
not U100061 ( n2692, n20883 );
nor U100062 ( n19044, n73006, n76576 );
nor U100063 ( n53821, n49898, n73397 );
or U100064 ( n20296, n73007, n76577 );
and U100065 ( n10234, n10235, n9894 );
nand U100066 ( n9551, n10179, n10180 );
nor U100067 ( n10180, n10182, n10183 );
nor U100068 ( n10179, n10233, n10234 );
nor U100069 ( n10182, n9520, n76632 );
xor U100070 ( n16869, n16875, n16876 );
nand U100071 ( n16875, n17020, n17021 );
xor U100072 ( n16876, n16877, n16878 );
nand U100073 ( n17021, n17022, n17023 );
xor U100074 ( n16883, n16884, n16885 );
nor U100075 ( n19043, n19044, n19045 );
and U100076 ( n44209, n44210, n43797 );
buf U100077 ( n76581, n76584 );
nor U100078 ( n20043, n76575, n73420 );
nor U100079 ( n20726, n73404, n16943 );
nand U100080 ( n51772, n51769, n51771 );
xnor U100081 ( n16891, n16885, n16884 );
nand U100082 ( n20384, n8222, n73015 );
nor U100083 ( n52443, n49898, n73403 );
nor U100084 ( n20040, n76575, n73020 );
nor U100085 ( n51603, n49898, n73401 );
nor U100086 ( n51987, n49898, n73005 );
nor U100087 ( n51280, n49898, n73411 );
not U100088 ( n1549, n53499 );
or U100089 ( n51456, n76322, n73001 );
nand U100090 ( n54014, n76650, n73424 );
nor U100091 ( n18812, n18813, n18814 );
xor U100092 ( n18814, n18810, n18815 );
not U100093 ( n1590, n53633 );
nor U100094 ( n52757, n76321, n73421 );
not U100095 ( n2827, n19367 );
nor U100096 ( n50780, n50508, n73416 );
buf U100097 ( n76582, n76584 );
nor U100098 ( n17567, n75916, n16943 );
nand U100099 ( n20182, n8222, n73418 );
nand U100100 ( n21083, n8222, n73018 );
nor U100101 ( n21011, n73423, n18105 );
not U100102 ( n2839, n19045 );
nor U100103 ( n53936, n53937, n53938 );
nor U100104 ( n53937, n53939, n53940 );
and U100105 ( n53939, n53941, n1263 );
nand U100106 ( n18816, n18813, n18815 );
nor U100107 ( n52602, n76321, n73021 );
nor U100108 ( n18653, n73398, n76575 );
nor U100109 ( n21078, n76575, n75919 );
nor U100110 ( n53367, n50508, n73413 );
or U100111 ( n50768, n76317, n73411 );
not U100112 ( n8234, n50496 );
not U100113 ( n1725, n50250 );
or U100114 ( n51595, n76322, n73401 );
or U100115 ( n53565, n76317, n73008 );
and U100116 ( n44252, n44253, n43797 );
nand U100117 ( n16276, n44211, n44212 );
nor U100118 ( n44212, n44213, n44214 );
nor U100119 ( n44211, n44251, n44252 );
nor U100120 ( n44213, n7567, n76361 );
nor U100121 ( n17323, n73417, n76587 );
nor U100122 ( n20710, n75913, n76588 );
buf U100123 ( n76588, n76585 );
nor U100124 ( n20763, n73012, n76588 );
nor U100125 ( n20848, n73414, n76588 );
nor U100126 ( n51464, n49898, n73001 );
or U100127 ( n53707, n76317, n73003 );
and U100128 ( n10357, n10358, n9894 );
nand U100129 ( n21103, n8222, n73420 );
nor U100130 ( n53252, n76316, n73017 );
nor U100131 ( n20509, n73015, n76588 );
or U100132 ( n53373, n76317, n73413 );
or U100133 ( n51020, n76317, n73001 );
nor U100134 ( n52596, n76322, n73424 );
or U100135 ( n52850, n76317, n72999 );
nor U100136 ( n51967, n76316, n73002 );
or U100137 ( n52422, n76317, n73397 );
or U100138 ( n53637, n76317, n73410 );
nor U100139 ( n53757, n50508, n73400 );
and U100140 ( n49739, n49744, n49743 );
nand U100141 ( n53942, n53941, n53943 );
nor U100142 ( n21050, n76575, n73022 );
nor U100143 ( n17316, n73417, n76579 );
buf U100144 ( n76579, n76578 );
nor U100145 ( n53152, n76316, n73419 );
nor U100146 ( n17834, n73417, n16943 );
nor U100147 ( n53920, n53921, n1308 );
nor U100148 ( n53921, n53922, n53923 );
and U100149 ( n53922, n53924, n1264 );
nor U100150 ( n20355, n73418, n76588 );
nor U100151 ( n53020, n76316, n73019 );
or U100152 ( n53444, n76317, n73412 );
and U100153 ( n44296, n44297, n43797 );
nand U100154 ( n16271, n44254, n44255 );
nor U100155 ( n44255, n44256, n44257 );
nor U100156 ( n44254, n44295, n44296 );
nor U100157 ( n44256, n7575, n76361 );
and U100158 ( n10410, n10412, n9894 );
nand U100159 ( n9541, n10359, n10360 );
nor U100160 ( n10360, n10362, n10363 );
nor U100161 ( n10359, n10409, n10410 );
nor U100162 ( n10362, n4916, n76631 );
xor U100163 ( n49866, n49871, n49872 );
xor U100164 ( n49871, n49944, n49945 );
xor U100165 ( n49872, n49873, n49874 );
or U100166 ( n49944, n76311, n73411 );
nor U100167 ( n17825, n73000, n76587 );
nor U100168 ( n50773, n50508, n73411 );
or U100169 ( n50239, n76314, n73411 );
buf U100170 ( n76314, n76312 );
nor U100171 ( n53700, n73003, n50508 );
nor U100172 ( n52895, n76316, n73400 );
xor U100173 ( n16635, n20972, n20973 );
xor U100174 ( n20972, n20974, n20975 );
nand U100175 ( n21096, n8222, n73020 );
nor U100176 ( n53955, n76321, n73426 );
nor U100177 ( n18091, n73000, n16943 );
nor U100178 ( n51028, n50508, n73001 );
or U100179 ( n51255, n76317, n73401 );
nor U100180 ( n52430, n50508, n73397 );
nor U100181 ( n19925, n73408, n16943 );
nor U100182 ( n21041, n73423, n76575 );
nor U100183 ( n52762, n76316, n73421 );
nor U100184 ( n51974, n50508, n73002 );
nand U100185 ( n16638, n20940, n20941 );
or U100186 ( n20940, n16600, n16603 );
nand U100187 ( n20941, n16602, n20942 );
nand U100188 ( n20942, n16603, n16600 );
nor U100189 ( n20964, n20965, n2425 );
nor U100190 ( n20965, n20966, n20967 );
and U100191 ( n20966, n20968, n2379 );
nand U100192 ( n53926, n53924, n53927 );
nor U100193 ( n51590, n50508, n73403 );
nor U100194 ( n17551, n73000, n76579 );
nand U100195 ( n49882, n49883, n49884 );
nand U100196 ( n49883, n1749, n49887 );
or U100197 ( n49884, n49885, n49886 );
xnor U100198 ( n49542, n53912, n53913 );
nand U100199 ( n53912, n53914, n53915 );
and U100200 ( n10465, n10467, n9894 );
nand U100201 ( n9536, n10413, n10414 );
nor U100202 ( n10414, n10415, n10417 );
nor U100203 ( n10413, n10464, n10465 );
nor U100204 ( n10415, n4923, n76631 );
nor U100205 ( n52619, n76316, n73021 );
nor U100206 ( n20315, n73404, n76588 );
or U100207 ( n51439, n76317, n73005 );
nor U100208 ( n49959, n76310, n73001 );
buf U100209 ( n76310, n76309 );
or U100210 ( n20636, n73012, n76580 );
buf U100211 ( n76580, n76578 );
xor U100212 ( n16911, n16916, n16917 );
xor U100213 ( n16916, n16989, n16990 );
xor U100214 ( n16917, n16918, n16919 );
or U100215 ( n16989, n73398, n76570 );
nor U100216 ( n53808, n72999, n50508 );
or U100217 ( n50482, n76314, n73001 );
nand U100218 ( n44301, n44302, n44303 );
nand U100219 ( n44303, n44261, n74965 );
nand U100220 ( n44302, n43797, n44305 );
nand U100221 ( n21045, n8222, n75919 );
buf U100222 ( n76586, n76585 );
nor U100223 ( n20286, n73406, n16943 );
nor U100224 ( n20153, n76586, n73018 );
nor U100225 ( n53930, n76322, n73425 );
nand U100226 ( n53910, n76323, n53911 );
nand U100227 ( n53911, n76652, n73425 );
nand U100228 ( n49544, n53902, n53903 );
nand U100229 ( n53902, n49515, n49512 );
nand U100230 ( n53903, n49514, n53904 );
or U100231 ( n53904, n49512, n49515 );
nor U100232 ( n19358, n73007, n16943 );
xor U100233 ( n49881, n49892, n49893 );
xor U100234 ( n49892, n49916, n49917 );
xor U100235 ( n49893, n49894, n49895 );
xor U100236 ( n49916, n49941, n49942 );
nand U100237 ( n49900, n49901, n49902 );
nand U100238 ( n49902, n49903, n49904 );
nand U100239 ( n49904, n1760, n49905 );
xor U100240 ( n49895, n49896, n49897 );
nor U100241 ( n49897, n73405, n49898 );
nand U100242 ( n49896, n49899, n49900 );
nand U100243 ( n49899, n1754, n49906 );
nor U100244 ( n19036, n73011, n16943 );
nor U100245 ( n51263, n50508, n73401 );
nor U100246 ( n20025, n76586, n73420 );
nand U100247 ( n20970, n20968, n20971 );
nor U100248 ( n50247, n50496, n73411 );
nor U100249 ( n20647, n76586, n73009 );
nor U100250 ( n53388, n76313, n73413 );
buf U100251 ( n76313, n76312 );
nor U100252 ( n17818, n73398, n76587 );
nor U100253 ( n18324, n73398, n16943 );
nor U100254 ( n18647, n73407, n16943 );
nor U100255 ( n53425, n76313, n73412 );
nor U100256 ( n52279, n76316, n73424 );
xnor U100257 ( n16563, n20956, n20957 );
nand U100258 ( n20956, n20958, n20959 );
nor U100259 ( n53651, n76313, n73410 );
or U100260 ( n20515, n73015, n76580 );
or U100261 ( n51951, n76314, n72999 );
nor U100262 ( n19019, n73408, n76587 );
not U100263 ( n1550, n53441 );
nor U100264 ( n51447, n50508, n73005 );
nor U100265 ( n53573, n76313, n73008 );
nor U100266 ( n20397, n76579, n73418 );
or U100267 ( n50755, n76314, n73401 );
nor U100268 ( n18074, n73006, n76587 );
nor U100269 ( n20700, n73414, n76580 );
not U100270 ( n8219, n16966 );
not U100271 ( n2844, n17304 );
nor U100272 ( n19341, n73406, n76587 );
nor U100273 ( n18634, n73007, n76587 );
nor U100274 ( n52474, n76313, n73003 );
not U100275 ( n1625, n52414 );
nor U100276 ( n20560, n73009, n76580 );
nor U100277 ( n53188, n76313, n73017 );
nand U100278 ( n10472, n10473, n10474 );
nand U100279 ( n10474, n10422, n74966 );
nand U100280 ( n10473, n9894, n10477 );
nor U100281 ( n50823, n76313, n73005 );
nor U100282 ( n21010, n76575, n73422 );
nor U100283 ( n19773, n76586, n73020 );
nor U100284 ( n52129, n76316, n73426 );
or U100285 ( n17813, n73398, n76580 );
nor U100286 ( n19657, n76586, n75919 );
or U100287 ( n51582, n76317, n73403 );
nor U100288 ( n53023, n76313, n73019 );
or U100289 ( n52402, n76314, n73400 );
nor U100290 ( n20273, n76586, n75911 );
nor U100291 ( n18504, n73006, n16943 );
xor U100292 ( n16940, n16941, n16942 );
nor U100293 ( n16942, n16943, n73004 );
nand U100294 ( n16941, n16944, n16945 );
nand U100295 ( n16944, n2874, n16951 );
nand U100296 ( n16945, n16946, n16947 );
nand U100297 ( n16947, n16948, n16949 );
nand U100298 ( n16949, n2877, n16950 );
or U100299 ( n20609, n75913, n76580 );
nor U100300 ( n51961, n50496, n73397 );
nor U100301 ( n52485, n76311, n73410 );
buf U100302 ( n76311, n76309 );
or U100303 ( n19904, n75911, n76580 );
nor U100304 ( n50549, n76310, n73005 );
nor U100305 ( n50487, n50496, n73001 );
or U100306 ( n19333, n73406, n76580 );
nand U100307 ( n20954, n76589, n20955 );
nand U100308 ( n20955, n76654, n73422 );
nand U100309 ( n16564, n20946, n20947 );
nand U100310 ( n20946, n16529, n16527 );
nand U100311 ( n20947, n16528, n20948 );
or U100312 ( n20948, n16527, n16529 );
nor U100313 ( n52843, n76310, n73008 );
or U100314 ( n18066, n73006, n76580 );
nor U100315 ( n50222, n76310, n73401 );
nor U100316 ( n20195, n76579, n73018 );
nand U100317 ( n21015, n8222, n73022 );
nor U100318 ( n51631, n76310, n73400 );
nor U100319 ( n53155, n76313, n73419 );
nor U100320 ( n53274, n76311, n73017 );
nor U100321 ( n18307, n73407, n76587 );
or U100322 ( n19011, n73408, n76580 );
nor U100323 ( n20063, n76579, n73420 );
nor U100324 ( n19500, n76586, n73022 );
nor U100325 ( n53092, n50496, n73419 );
nor U100326 ( n19897, n73404, n76580 );
nor U100327 ( n52765, n76313, n73421 );
nor U100328 ( n53415, n73412, n76311 );
nor U100329 ( n53303, n76311, n73413 );
nor U100330 ( n50763, n50496, n73401 );
nor U100331 ( n52947, n76311, n73019 );
or U100332 ( n17293, n73398, n76573 );
buf U100333 ( n76573, n76571 );
nor U100334 ( n52622, n76313, n73021 );
nor U100335 ( n18491, n73011, n76587 );
nand U100336 ( n16261, n44340, n44341 );
nor U100337 ( n44341, n44342, n44343 );
nor U100338 ( n44340, n44380, n44381 );
nor U100339 ( n44342, n7599, n76361 );
and U100340 ( n44381, n44382, n43797 );
nor U100341 ( n51072, n50496, n73005 );
nor U100342 ( n53166, n76311, n73419 );
nor U100343 ( n52410, n50496, n73400 );
not U100344 ( n2665, n20693 );
and U100345 ( n49514, n53905, n8229 );
nor U100346 ( n53905, n73425, n76834 );
or U100347 ( n18299, n73407, n76580 );
nor U100348 ( n20529, n76572, n73015 );
buf U100349 ( n76572, n76571 );
nor U100350 ( n21032, n73423, n76587 );
nor U100351 ( n19805, n76579, n73020 );
or U100352 ( n51238, n76314, n73403 );
nand U100353 ( n53909, n76650, n73426 );
nor U100354 ( n52304, n76313, n73424 );
nor U100355 ( n51938, n76311, n73003 );
nor U100356 ( n17534, n73006, n76572 );
nor U100357 ( n51426, n76314, n73002 );
xor U100358 ( n49519, n49521, n49522 );
nor U100359 ( n19662, n76579, n75919 );
nor U100360 ( n52695, n76311, n73421 );
nor U100361 ( n52123, n76316, n73425 );
nor U100362 ( n17004, n73006, n76569 );
buf U100363 ( n76569, n76568 );
or U100364 ( n18483, n73011, n76580 );
nor U100365 ( n52567, n76311, n73021 );
nor U100366 ( n52133, n76314, n73426 );
nor U100367 ( n20622, n76572, n73414 );
nor U100368 ( n50750, n76310, n73403 );
nor U100369 ( n17301, n73398, n16966 );
not U100370 ( n1302, n52118 );
or U100371 ( n51567, n76314, n73397 );
nand U100372 ( n9526, n10520, n10522 );
nor U100373 ( n10522, n10523, n10524 );
nor U100374 ( n10520, n10570, n10572 );
nor U100375 ( n10523, n4945, n76631 );
and U100376 ( n10572, n10573, n9894 );
nor U100377 ( n20250, n73012, n76573 );
not U100378 ( n2715, n19892 );
or U100379 ( n20334, n76573, n73418 );
xor U100380 ( n49917, n49918, n49919 );
nor U100381 ( n49918, n49926, n49927 );
nor U100382 ( n49919, n49920, n49921 );
nor U100383 ( n49926, n49932, n49933 );
nor U100384 ( n49920, n49923, n49924 );
or U100385 ( n49924, n73402, n49925 );
nor U100386 ( n49927, n1769, n49928 );
nor U100387 ( n49928, n49929, n73402 );
not U100388 ( n1769, n49932 );
xor U100389 ( n49929, n49930, n76318 );
or U100390 ( n18995, n75911, n76573 );
nor U100391 ( n19487, n76579, n73022 );
nor U100392 ( n17796, n73407, n76572 );
not U100393 ( n8237, n50543 );
nor U100394 ( n52255, n76311, n73424 );
not U100395 ( n2748, n19325 );
and U100396 ( n44439, n44440, n43797 );
nand U100397 ( n16256, n44397, n44398 );
nor U100398 ( n44398, n44399, n44400 );
nor U100399 ( n44397, n44438, n44439 );
nor U100400 ( n44399, n7613, n76361 );
or U100401 ( n20257, n75913, n76573 );
nor U100402 ( n51243, n50496, n73403 );
nor U100403 ( n20420, n73418, n76570 );
buf U100404 ( n76570, n76568 );
nor U100405 ( n20199, n76572, n73018 );
nor U100406 ( n49936, n73431, n49939 );
xor U100407 ( n16534, n16537, n16538 );
nor U100408 ( n52144, n76310, n73426 );
nor U100409 ( n19306, n73009, n76573 );
or U100410 ( n18626, n73007, n76580 );
nor U100411 ( n51417, n76310, n72999 );
nor U100412 ( n19174, n73423, n76579 );
nor U100413 ( n20067, n76572, n73420 );
nor U100414 ( n51013, n76310, n73002 );
nor U100415 ( n19005, n73406, n16966 );
or U100416 ( n19313, n73404, n76573 );
nor U100417 ( n20136, n16966, n73018 );
xor U100418 ( n49455, n49457, n49458 );
nor U100419 ( n17864, n73011, n76573 );
nor U100420 ( n20985, n76586, n73422 );
nor U100421 ( n17538, n73006, n16966 );
not U100422 ( n552, n41769 );
not U100423 ( n812, n41449 );
nand U100424 ( n40880, n41379, n41380 );
nand U100425 ( n41379, n41383, n41382 );
nand U100426 ( n41380, n41381, n40826 );
or U100427 ( n41381, n41382, n41383 );
not U100428 ( n815, n11399 );
not U100429 ( n844, n12652 );
not U100430 ( n909, n16703 );
not U100431 ( n883, n15745 );
not U100432 ( n899, n16270 );
not U100433 ( n848, n14375 );
not U100434 ( n860, n15214 );
not U100435 ( n869, n15482 );
not U100436 ( n855, n14923 );
not U100437 ( n889, n16002 );
and U100438 ( n49921, n49922, n1764 );
nor U100439 ( n51233, n76310, n73397 );
nor U100440 ( n20210, n73018, n76570 );
nand U100441 ( n2001, n40698, n40699 );
nor U100442 ( n40698, n40709, n40710 );
nor U100443 ( n40699, n40700, n40701 );
nor U100444 ( n40709, P3_STATE_REG, n74736 );
nor U100445 ( n51433, n50496, n73002 );
nor U100446 ( n20444, n73015, n76569 );
or U100447 ( n51775, n76314, n73425 );
nor U100448 ( n19881, n73012, n76570 );
or U100449 ( n19302, n75913, n76570 );
nor U100450 ( n18675, n73404, n76569 );
not U100451 ( n1754, n49901 );
not U100452 ( n1893, n37764 );
not U100453 ( n2153, n37080 );
nand U100454 ( n40547, n39501, n73035 );
not U100455 ( n1849, n37016 );
nand U100456 ( n40524, n40450, n73496 );
nand U100457 ( n40489, n40346, n73051 );
nor U100458 ( n40342, n40488, n40479 );
nor U100459 ( n40488, n73519, n2154 );
not U100460 ( n2209, n40289 );
not U100461 ( n2203, n39856 );
not U100462 ( n2205, n40035 );
not U100463 ( n2208, n40205 );
not U100464 ( n2202, n39755 );
not U100465 ( n2204, n39955 );
not U100466 ( n2207, n40128 );
nor U100467 ( n17524, n73011, n76569 );
xnor U100468 ( n41383, n40826, n42276 );
nor U100469 ( n42276, n42277, n42278 );
nor U100470 ( n42277, n40665, n73579 );
nand U100471 ( n42278, n42279, n42280 );
nand U100472 ( n42280, n41769, n41264 );
nand U100473 ( n1946, n40936, n40937 );
nor U100474 ( n40936, n40946, n40947 );
nor U100475 ( n40937, n40938, n40939 );
nor U100476 ( n40946, P3_STATE_REG, n74674 );
and U100477 ( n16528, n20949, n8220 );
nor U100478 ( n20949, n76788, n73422 );
nand U100479 ( n3226, n36294, n36295 );
nor U100480 ( n36294, n36306, n36307 );
nor U100481 ( n36295, n36296, n36297 );
nor U100482 ( n36306, P4_STATE_REG, n74708 );
nor U100483 ( n17276, n73407, n76569 );
and U100484 ( n10627, n10628, n9894 );
nand U100485 ( n9521, n10574, n10575 );
nor U100486 ( n10575, n10577, n10578 );
nor U100487 ( n10574, n10625, n10627 );
nor U100488 ( n10577, n4959, n76631 );
and U100489 ( n44481, n44482, n43797 );
not U100490 ( n814, n41972 );
nor U100491 ( n20539, n76569, n73414 );
xor U100492 ( n16962, n16968, n16969 );
nor U100493 ( n16969, n16970, n16971 );
nand U100494 ( n16968, n16984, n16985 );
nor U100495 ( n16970, n16975, n16976 );
nor U100496 ( n17803, n73407, n16966 );
nor U100497 ( n19809, n76572, n73020 );
nor U100498 ( n49972, n50320, n73005 );
nor U100499 ( n50210, n50543, n73005 );
nor U100500 ( n19991, n73420, n76570 );
not U100501 ( n1525, n53407 );
nor U100502 ( n51748, n76310, n73425 );
nor U100503 ( n19321, n73404, n16966 );
nor U100504 ( n19666, n76572, n75919 );
xnor U100505 ( n36487, n37019, n2040 );
nand U100506 ( n37019, n37020, n37021 );
nand U100507 ( n37020, n76828, n37023 );
nand U100508 ( n37021, n37022, n2035 );
nand U100509 ( n37015, n37016, n36481 );
nor U100510 ( n18119, n73011, n16966 );
not U100511 ( n2069, n37300 );
nand U100512 ( n37297, n2069, n37102 );
nor U100513 ( n18286, n73007, n76573 );
xor U100514 ( n40421, n73047, n40530 );
nor U100515 ( n16971, n2884, n16972 );
not U100516 ( n2884, n16975 );
nor U100517 ( n16972, n16973, n73399 );
xor U100518 ( n16973, n76577, n8220 );
xor U100519 ( n36485, n36481, n37759 );
nor U100520 ( n37759, n37760, n37761 );
nor U100521 ( n37760, n36265, n73798 );
nand U100522 ( n37761, n37762, n37763 );
nand U100523 ( n37763, n37764, n2035 );
not U100524 ( n2197, n37609 );
nor U100525 ( n40347, n73051, n40346 );
nor U100526 ( n40345, n40346, n40347 );
and U100527 ( n44485, n44493, n43797 );
nand U100528 ( n16246, n44483, n44484 );
nor U100529 ( n44483, n44496, n44497 );
nor U100530 ( n44484, n44485, n44486 );
nor U100531 ( n44497, n7634, n76361 );
xor U100532 ( n16455, n16458, n16459 );
nand U100533 ( n36486, n37024, n37025 );
nand U100534 ( n37025, n76807, n37023 );
nand U100535 ( n37024, n76828, n37022 );
nor U100536 ( n19511, n76572, n73022 );
nor U100537 ( n18982, n73009, n76570 );
nand U100538 ( n37283, n37284, n37285 );
nand U100539 ( n37284, n37287, n2157 );
nand U100540 ( n37285, n37286, n37022 );
or U100541 ( n37286, n2157, n37287 );
nor U100542 ( n37278, n37280, n37281 );
nor U100543 ( n37281, n2158, n37007 );
nor U100544 ( n37280, n37282, n37283 );
nor U100545 ( n37282, n1909, n36381 );
nand U100546 ( n37122, n37123, n37124 );
nand U100547 ( n37123, n37301, n1850 );
nand U100548 ( n37124, n2060, n37125 );
nor U100549 ( n37301, n37303, n37304 );
nor U100550 ( n18470, n73408, n76573 );
nand U100551 ( n3171, n36538, n36539 );
nor U100552 ( n36538, n36552, n36553 );
nor U100553 ( n36539, n36540, n36541 );
nor U100554 ( n36552, P4_STATE_REG, n74627 );
not U100555 ( n8238, n50320 );
nor U100556 ( n49942, n73415, n76317 );
nor U100557 ( n19739, n73020, n76570 );
xnor U100558 ( n40877, n41384, n593 );
nand U100559 ( n41384, n41385, n41386 );
nand U100560 ( n41385, n76845, n41377 );
nand U100561 ( n41386, n41378, n41264 );
nor U100562 ( n19178, n76572, n73423 );
nor U100563 ( n52769, n50543, n73421 );
nor U100564 ( n19611, n75919, n76570 );
nor U100565 ( n52830, n73412, n50320 );
not U100566 ( n2098, n37022 );
not U100567 ( n1477, n53072 );
nor U100568 ( n19167, n76579, n73422 );
not U100569 ( n2418, n19162 );
nor U100570 ( n49543, n49898, n76835 );
xnor U100571 ( n41163, n41366, n593 );
nand U100572 ( n41366, n41367, n41368 );
nand U100573 ( n41367, n76845, n40784 );
nand U100574 ( n41368, n41369, n41264 );
or U100575 ( n18615, n73406, n76573 );
nand U100576 ( n38136, n38775, n38776 );
nor U100577 ( n38775, n38801, n38802 );
nor U100578 ( n38776, n38777, n38778 );
nor U100579 ( n38801, n2190, n38822 );
and U100580 ( n10679, n10680, n9894 );
nand U100581 ( n37401, n2155, n37764 );
nand U100582 ( n37384, n2157, n37022 );
nand U100583 ( n2811, n38121, n38122 );
nor U100584 ( n38122, n38123, n38124 );
nor U100585 ( n38121, n38131, n38132 );
nor U100586 ( n38123, n37600, n38108 );
nor U100587 ( n51927, n50320, n73008 );
not U100588 ( n1448, n53040 );
xnor U100589 ( n36780, n37004, n2040 );
nand U100590 ( n37004, n37005, n37006 );
nand U100591 ( n37005, n76828, n36381 );
nand U100592 ( n37006, n37007, n2035 );
nor U100593 ( n17791, n73007, n76569 );
not U100594 ( n8215, n17525 );
nor U100595 ( n53403, n50320, n73413 );
not U100596 ( n1909, n37007 );
nor U100597 ( n18290, n73007, n16966 );
nand U100598 ( n39902, n40021, n40022 );
nand U100599 ( n40022, n36462, n36293 );
nor U100600 ( n40021, n40023, n40024 );
nor U100601 ( n40024, n40025, n40026 );
xor U100602 ( n40783, n41389, n40826 );
nand U100603 ( n41389, n41390, n41391 );
nand U100604 ( n41390, n76845, n41036 );
nand U100605 ( n41391, n40789, n41264 );
nor U100606 ( n53292, n50320, n73017 );
nor U100607 ( n51556, n50320, n73410 );
nand U100608 ( n41162, n41370, n41371 );
nand U100609 ( n41371, n76847, n40784 );
nand U100610 ( n41370, n76845, n41369 );
nor U100611 ( n19462, n73022, n76570 );
nand U100612 ( n37276, n2159, n36386 );
nor U100613 ( n53027, n50543, n73019 );
nand U100614 ( n37472, n2158, n37007 );
nand U100615 ( n20953, n8222, n73423 );
xor U100616 ( n36380, n37028, n36481 );
nand U100617 ( n37028, n37029, n37030 );
nand U100618 ( n37029, n76828, n36649 );
nand U100619 ( n37030, n36386, n2035 );
nor U100620 ( n52626, n50543, n73021 );
nand U100621 ( n36779, n37008, n37009 );
nand U100622 ( n37009, n76807, n36381 );
nand U100623 ( n37008, n76828, n37007 );
nand U100624 ( n1991, n40733, n40734 );
nor U100625 ( n40733, n40743, n40744 );
nor U100626 ( n40734, n40735, n40736 );
nor U100627 ( n40743, P3_STATE_REG, n74567 );
nand U100628 ( n40879, n41375, n41376 );
nand U100629 ( n41376, n76847, n41377 );
nand U100630 ( n41375, n76845, n41378 );
not U100631 ( n785, n41378 );
nor U100632 ( n66367, n41574, n66369 );
and U100633 ( n66369, n66370, n66371 );
nand U100634 ( n66370, n635, n40789 );
nand U100635 ( n1586, n45485, n45486 );
nor U100636 ( n45485, n45494, n45406 );
nor U100637 ( n45486, n45487, n45488 );
nor U100638 ( n45494, n76855, n74862 );
and U100639 ( n45493, n61393, n61394 );
nor U100640 ( n61393, n61420, n61421 );
nor U100641 ( n61394, n61395, n61396 );
nor U100642 ( n61420, n775, n61441 );
nand U100643 ( n42011, n624, n41769 );
nor U100644 ( n51489, n50543, n73400 );
and U100645 ( n10684, n10694, n9894 );
nand U100646 ( n9511, n10682, n10683 );
nor U100647 ( n10682, n10698, n10699 );
nor U100648 ( n10683, n10684, n10685 );
nor U100649 ( n10698, n2, n9897 );
nor U100650 ( n19188, n73423, n76570 );
nor U100651 ( n50466, n50320, n73002 );
nand U100652 ( n3216, n36328, n36329 );
nor U100653 ( n36328, n36340, n36341 );
nor U100654 ( n36329, n36330, n36331 );
nor U100655 ( n36340, P4_STATE_REG, n74578 );
nand U100656 ( n41990, n623, n41378 );
not U100657 ( n2635, n20533 );
buf U100658 ( n76091, n49969 );
or U100659 ( n50193, n76091, n73403 );
nor U100660 ( n37412, n36386, n2159 );
nand U100661 ( n40782, n41387, n41388 );
nand U100662 ( n41388, n76847, n41036 );
nand U100663 ( n41387, n76845, n40789 );
nor U100664 ( n18461, n75911, n76569 );
nor U100665 ( n18477, n73408, n16966 );
nor U100666 ( n18055, n73408, n76569 );
nand U100667 ( n1956, n40889, n40890 );
nor U100668 ( n40889, n40909, n40910 );
nor U100669 ( n40890, n40891, n40892 );
nor U100670 ( n40909, P3_STATE_REG, n74492 );
nor U100671 ( n18281, n73406, n76570 );
not U100672 ( n1919, n36655 );
not U100673 ( n786, n41369 );
nor U100674 ( n52309, n50543, n73424 );
nand U100675 ( n36379, n37026, n37027 );
nand U100676 ( n37027, n76807, n36649 );
nand U100677 ( n37026, n76828, n36386 );
not U100678 ( n1928, n36822 );
nand U100679 ( n37268, n2162, n36594 );
nor U100680 ( n52150, n50543, n73426 );
buf U100681 ( n76087, n49969 );
nor U100682 ( n51920, n76087, n73008 );
nand U100683 ( n41989, n628, n41369 );
not U100684 ( n2072, n37097 );
nand U100685 ( n40230, n37023, n37022 );
nand U100686 ( n40665, n70973, n70968 );
nor U100687 ( n70973, n620, n67262 );
not U100688 ( n622, n70976 );
or U100689 ( n18819, n76573, n73422 );
not U100690 ( n1913, n36386 );
nand U100691 ( n3181, n36493, n36494 );
nor U100692 ( n36493, n36513, n36514 );
nor U100693 ( n36494, n36495, n36496 );
nor U100694 ( n36513, P4_STATE_REG, n74485 );
nand U100695 ( n66116, n66193, n66194 );
nand U100696 ( n66194, n40989, n41198 );
nor U100697 ( n66193, n66195, n66196 );
nor U100698 ( n66196, n66197, n66198 );
nand U100699 ( n65945, n66018, n66019 );
nand U100700 ( n66019, n66020, n40697 );
nor U100701 ( n66018, n66021, n66022 );
nor U100702 ( n66022, n654, n66023 );
nor U100703 ( n66021, n66024, n66025 );
nor U100704 ( n66024, n40697, n40864 );
or U100705 ( n66025, n543, n66026 );
nor U100706 ( n17018, n73011, n17014 );
nor U100707 ( n45508, n44560, n45391 );
nor U100708 ( n52388, n76088, n73412 );
buf U100709 ( n76088, n49969 );
nor U100710 ( n44559, n44560, n44561 );
nand U100711 ( n16241, n44549, n44550 );
nor U100712 ( n44550, n44551, n44552 );
nor U100713 ( n44549, n44558, n44559 );
nor U100714 ( n44551, n44556, n44557 );
nor U100715 ( n49618, n50508, n76835 );
not U100716 ( n1925, n36594 );
nor U100717 ( n51314, n50320, n73400 );
nor U100718 ( n50459, n76088, n73002 );
nor U100719 ( n49829, n76096, n73002 );
buf U100720 ( n76096, n49970 );
nor U100721 ( n16979, n73430, n16982 );
not U100722 ( n2874, n16946 );
nor U100723 ( n52495, n76092, n73413 );
buf U100724 ( n76092, n49969 );
nand U100725 ( n1576, n45993, n45994 );
nor U100726 ( n45994, n45995, n45996 );
nor U100727 ( n45993, n45406, n46000 );
nor U100728 ( n45995, n40715, n76336 );
not U100729 ( n620, n70965 );
nor U100730 ( n17264, n73011, n17525 );
nor U100731 ( n67237, n76248, n73579 );
not U100732 ( n783, n67249 );
nand U100733 ( n42184, n67233, n67234 );
nor U100734 ( n67234, n67235, n67236 );
nor U100735 ( n67233, n67237, n67238 );
nor U100736 ( n67235, n76246, n73633 );
nand U100737 ( n61294, n783, n67248 );
nor U100738 ( n49945, n73416, n76314 );
not U100739 ( n787, n40789 );
not U100740 ( n8217, n17014 );
nand U100741 ( n40226, n37007, n36381 );
nor U100742 ( n52238, n50320, n73424 );
xnor U100743 ( n41032, n41392, n593 );
nand U100744 ( n41392, n41393, n41394 );
nand U100745 ( n41393, n76845, n40984 );
nand U100746 ( n41394, n41042, n41264 );
or U100747 ( n52823, n76088, n73017 );
nor U100748 ( n41574, n40789, n635 );
nor U100749 ( n67236, n76241, n73637 );
nand U100750 ( n61595, n67248, n67249 );
nor U100751 ( n50737, n50320, n73397 );
nor U100752 ( n18792, n76569, n73422 );
not U100753 ( n2597, n20116 );
nor U100754 ( n51403, n76090, n73410 );
buf U100755 ( n76090, n49969 );
nor U100756 ( n52501, n76096, n73017 );
nor U100757 ( n37265, n2163, n36822 );
buf U100758 ( n76089, n49969 );
or U100759 ( n53176, n76089, n73419 );
nor U100760 ( n53044, n76086, n73019 );
buf U100761 ( n76086, n49969 );
not U100762 ( n838, n41466 );
not U100763 ( n843, n67316 );
nand U100764 ( n40111, n36386, n36649 );
nand U100765 ( n71104, n72890, n6259 );
nor U100766 ( n72923, n72924, n72925 );
nand U100767 ( n72924, n73407, n73006 );
nand U100768 ( n72925, n73011, n73422 );
not U100769 ( n2362, n71021 );
nor U100770 ( n72900, n72915, n72916 );
nand U100771 ( n72916, n72917, n72918 );
nand U100772 ( n72915, n72922, n72923 );
nor U100773 ( n72918, n72919, n72920 );
buf U100774 ( n76796, n76791 );
buf U100775 ( n76791, n76792 );
nand U100776 ( n71105, n72890, n72801 );
nor U100777 ( n72760, n73027, n71105 );
not U100778 ( n2567, n20084 );
or U100779 ( n16976, n73399, n76577 );
nor U100780 ( n61291, n67249, n67248 );
nor U100781 ( n72909, n72913, n72914 );
nand U100782 ( n72913, n75919, n73020 );
nand U100783 ( n72914, n73423, n73022 );
nor U100784 ( n20431, n17014, n73418 );
nor U100785 ( n45386, n43798, n45391 );
xnor U100786 ( n45501, n45503, n45504 );
nand U100787 ( n71283, n72830, n3632 );
nand U100788 ( n72880, n73005, n73425 );
not U100789 ( n1244, n71012 );
nand U100790 ( n71429, n72776, n72777 );
nor U100791 ( n72776, n72780, n72781 );
nor U100792 ( n72777, n72778, n72779 );
nor U100793 ( n72781, n73446, n73025 );
nand U100794 ( n72855, n72856, n72857 );
nor U100795 ( n72857, n72858, n72859 );
nor U100796 ( n72856, n72870, n72871 );
nand U100797 ( n72858, n72865, n72866 );
xor U100798 ( n71087, n71092, n71093 );
xor U100799 ( n71093, n71094, n71095 );
xor U100800 ( n71092, n71109, n71110 );
nand U100801 ( n71094, n71098, n71099 );
nand U100802 ( n71284, n72830, n72831 );
nor U100803 ( n72778, n73444, n71284 );
nand U100804 ( n71303, n72765, n72766 );
nor U100805 ( n72765, n72769, n72770 );
nor U100806 ( n72766, n72767, n72768 );
nor U100807 ( n72770, n73442, n73025 );
nand U100808 ( n71108, n2362, n73026 );
nor U100809 ( n72762, n73028, n71108 );
not U100810 ( n842, n41493 );
nor U100811 ( n72767, n73031, n71284 );
nand U100812 ( n42287, n840, n41466 );
nand U100813 ( n72862, n73010, n73426 );
nor U100814 ( n51915, n76098, n73413 );
buf U100815 ( n76098, n49970 );
nor U100816 ( n44616, n43798, n44561 );
nand U100817 ( n71022, n6259, n71021 );
not U100818 ( n1209, n71274 );
nand U100819 ( n71017, n72801, n71021 );
not U100820 ( n789, n40989 );
nor U100821 ( n40355, n76414, n73798 );
nand U100822 ( n37288, n40349, n40350 );
nor U100823 ( n40350, n40351, n40352 );
nor U100824 ( n40349, n40355, n40356 );
nor U100825 ( n40351, n76412, n73799 );
not U100826 ( n2195, n40354 );
nand U100827 ( n38756, n2195, n40353 );
nor U100828 ( n43794, n43798, n43799 );
nand U100829 ( n72774, n1227, n71274 );
nor U100830 ( n51219, n76091, n73003 );
nand U100831 ( n3201, n36387, n36388 );
nor U100832 ( n36387, n36399, n36400 );
nor U100833 ( n36388, n36389, n36390 );
nor U100834 ( n36399, P4_STATE_REG, n74459 );
nor U100835 ( n72910, n72911, n72912 );
nand U100836 ( n72911, n73418, n73015 );
nand U100837 ( n72912, n73420, n73018 );
nand U100838 ( n71287, n1244, n73025 );
nor U100839 ( n72780, n73445, n71287 );
nor U100840 ( n72769, n73032, n71287 );
nand U100841 ( n71413, n72745, n72746 );
nor U100842 ( n72745, n72749, n72750 );
nor U100843 ( n72746, n72747, n72748 );
nor U100844 ( n72750, n73440, n73025 );
nand U100845 ( n71244, n72783, n72784 );
nor U100846 ( n72783, n72787, n72788 );
nor U100847 ( n72784, n72785, n72786 );
nor U100848 ( n72788, n73448, n73025 );
nor U100849 ( n19868, n73414, n17014 );
nor U100850 ( n72866, n72867, n72868 );
nand U100851 ( n72867, n73017, n73413 );
nand U100852 ( n72868, n73019, n73419 );
xnor U100853 ( n40980, n41395, n593 );
nand U100854 ( n41395, n41396, n41397 );
nand U100855 ( n41396, n76845, n41198 );
nand U100856 ( n41397, n40989, n41264 );
nor U100857 ( n72747, n73029, n71284 );
nor U100858 ( n72785, n73033, n71284 );
xnor U100859 ( n36645, n36993, n2040 );
nand U100860 ( n36993, n36994, n36995 );
nand U100861 ( n36994, n76828, n36589 );
nand U100862 ( n36995, n36655, n2035 );
xor U100863 ( n40412, n40547, n73479 );
not U100864 ( n2042, n37303 );
nand U100865 ( n36648, n36996, n36997 );
nand U100866 ( n36997, n76807, n36589 );
nand U100867 ( n36996, n76828, n36655 );
nor U100868 ( n40352, n76403, n73800 );
nand U100869 ( n38843, n40353, n40354 );
nor U100870 ( n18972, n17014, n73012 );
nand U100871 ( n1976, n40790, n40791 );
nor U100872 ( n40790, n40802, n40803 );
nor U100873 ( n40791, n40792, n40793 );
nor U100874 ( n40802, P3_STATE_REG, n74462 );
nand U100875 ( n1571, n46214, n46215 );
nor U100876 ( n46215, n46216, n46217 );
nor U100877 ( n46214, n45406, n46222 );
nand U100878 ( n46217, n46218, n46219 );
nand U100879 ( n66750, n41377, n41378 );
not U100880 ( n2094, n40442 );
nor U100881 ( n40461, n40523, n40496 );
nor U100882 ( n40523, n73050, n2095 );
nand U100883 ( n36265, n40453, n40445 );
nor U100884 ( n40453, n40437, n2094 );
nand U100885 ( n72741, n1228, n71274 );
nor U100886 ( n72749, n73030, n71287 );
nor U100887 ( n72787, n73034, n71287 );
nand U100888 ( n41035, n41358, n41359 );
nand U100889 ( n41359, n76847, n40984 );
nand U100890 ( n41358, n76845, n41042 );
xnor U100891 ( n40359, n73058, n40479 );
nand U100892 ( n37023, n40330, n40331 );
nor U100893 ( n40331, n40332, n40333 );
nor U100894 ( n40330, n40334, n40335 );
nor U100895 ( n40332, n76412, n73802 );
nor U100896 ( n40334, n76414, n73804 );
not U100897 ( n788, n41042 );
nor U100898 ( n11732, n10784, n11594 );
nand U100899 ( n72876, n73412, n73008 );
nor U100900 ( n20071, n73420, n17525 );
nor U100901 ( n10783, n10784, n10785 );
nand U100902 ( n9506, n10770, n10772 );
nor U100903 ( n10772, n10773, n10774 );
nor U100904 ( n10770, n10782, n10783 );
nor U100905 ( n10773, n10779, n10780 );
nor U100906 ( n20229, n17014, n73015 );
nand U100907 ( n72712, n71272, n72713 );
nand U100908 ( n72713, n1229, n71274 );
nand U100909 ( n72919, n73404, n75911 );
nor U100910 ( n19813, n73020, n17525 );
nand U100911 ( n42084, n639, n41042 );
nand U100912 ( n1556, n47410, n47411 );
nor U100913 ( n47411, n47412, n47413 );
nor U100914 ( n47410, n45406, n47417 );
nor U100915 ( n47412, n40748, n76336 );
nor U100916 ( n40106, n36817, n36594 );
nand U100917 ( n72920, n75913, n73009 );
nor U100918 ( n51780, n50543, n73425 );
nand U100919 ( n72546, n1225, n71274 );
nand U100920 ( n38124, n38125, n38126 );
nand U100921 ( n38126, n76448, n2905 );
nand U100922 ( n38125, n76444, n1878 );
not U100923 ( n2905, n38128 );
nand U100924 ( n72875, n73410, n73003 );
nor U100925 ( n40333, n76403, n73801 );
nor U100926 ( n51644, n76099, n73412 );
buf U100927 ( n76099, n49970 );
nand U100928 ( n71246, n72549, n72550 );
nor U100929 ( n72549, n72553, n72554 );
nor U100930 ( n72550, n72551, n72552 );
nor U100931 ( n72554, n73456, n73025 );
nor U100932 ( n72551, n73454, n71284 );
nor U100933 ( n41577, n41203, n650 );
or U100934 ( n51320, n76098, n73410 );
nor U100935 ( n38753, n40354, n40353 );
xnor U100936 ( n36585, n37031, n2040 );
nand U100937 ( n37031, n37032, n37033 );
nand U100938 ( n37032, n76828, n36817 );
nand U100939 ( n37033, n36594, n2035 );
nand U100940 ( n71278, n72789, n72790 );
nand U100941 ( n72790, n71024, n73026 );
xnor U100942 ( n41196, n41400, n593 );
nand U100943 ( n41400, n41401, n41402 );
nand U100944 ( n41401, n76846, n40690 );
nand U100945 ( n41402, n41264, n41203 );
nor U100946 ( n16964, n76579, n75916 );
nand U100947 ( n71574, n72721, n72722 );
nor U100948 ( n72721, n72725, n72726 );
nor U100949 ( n72722, n72723, n72724 );
nor U100950 ( n72726, n73452, n73025 );
nor U100951 ( n16565, n16943, n76789 );
nor U100952 ( n18600, n75913, n17014 );
nor U100953 ( n72723, n73450, n71284 );
nor U100954 ( n72553, n73455, n71287 );
nor U100955 ( n72905, n72906, n72907 );
nand U100956 ( n72906, n73409, n73004 );
nand U100957 ( n72907, n75916, n73013 );
nand U100958 ( n41377, n67244, n67245 );
nor U100959 ( n67245, n67246, n67247 );
nor U100960 ( n67244, n67250, n67251 );
nor U100961 ( n67246, n76246, n73827 );
nand U100962 ( n72879, n73401, n73001 );
nor U100963 ( n67250, n76248, n73825 );
or U100964 ( n50729, n76090, n73397 );
nand U100965 ( n76043, n72789, n72790 );
nand U100966 ( n41562, n648, n40989 );
not U100967 ( n845, n41908 );
buf U100968 ( n76097, n49970 );
nor U100969 ( n51396, n76097, n73008 );
nand U100970 ( n72339, n71272, n72340 );
nand U100971 ( n72340, n1234, n71274 );
nand U100972 ( n71312, n72471, n72472 );
nor U100973 ( n72471, n72475, n72476 );
nor U100974 ( n72472, n72473, n72474 );
nor U100975 ( n72476, n73468, n73025 );
not U100976 ( n790, n41203 );
nand U100977 ( n76044, n72789, n72790 );
nor U100978 ( n72473, n73466, n71284 );
nand U100979 ( n72908, n73000, n73417 );
nand U100980 ( n40784, n66999, n67000 );
nor U100981 ( n67000, n67001, n67002 );
nor U100982 ( n66999, n67003, n67004 );
nor U100983 ( n67001, n76246, n73826 );
nor U100984 ( n67003, n76248, n73829 );
nor U100985 ( n72725, n73451, n71287 );
nor U100986 ( n52631, n76086, n73021 );
nand U100987 ( n37304, n2072, n37300 );
nand U100988 ( n72863, n73415, n73014 );
nor U100989 ( n45382, n43846, n45391 );
nand U100990 ( n71308, n72826, n72827 );
nor U100991 ( n72826, n72832, n72833 );
nor U100992 ( n72827, n72828, n72829 );
nor U100993 ( n72833, n73459, n73025 );
nor U100994 ( n72828, n73036, n71284 );
nor U100995 ( n52312, n76087, n73424 );
nor U100996 ( n44656, n43846, n44561 );
nand U100997 ( n16231, n44647, n44648 );
nor U100998 ( n44648, n44649, n44650 );
nor U100999 ( n44647, n44655, n44656 );
nor U101000 ( n44649, n43808, n44652 );
nor U101001 ( n50996, n50320, n72999 );
nor U101002 ( n67247, n76241, n73823 );
nor U101003 ( n52785, n76086, n73421 );
not U101004 ( n1933, n36293 );
buf U101005 ( n76095, n49970 );
nor U101006 ( n50177, n76095, n73397 );
nor U101007 ( n43843, n43846, n43799 );
not U101008 ( n829, n41471 );
nor U101009 ( n72475, n73467, n71287 );
buf U101010 ( n76093, n49970 );
nor U101011 ( n52816, n76093, n73419 );
nor U101012 ( n19670, n75919, n17525 );
nand U101013 ( n37106, n2032, n37097 );
nand U101014 ( n40983, n41353, n41354 );
nand U101015 ( n41354, n76847, n41198 );
nand U101016 ( n41353, n76845, n40989 );
nand U101017 ( n37260, n2164, n36293 );
nor U101018 ( n66197, n41198, n40989 );
nor U101019 ( n67002, n76241, n73833 );
nor U101020 ( n72832, n73038, n71287 );
xnor U101021 ( n36815, n37036, n2040 );
nand U101022 ( n37036, n37037, n37038 );
nand U101023 ( n37037, n76829, n36286 );
nand U101024 ( n37038, n2035, n36822 );
nor U101025 ( n18533, n73404, n17525 );
xnor U101026 ( n40689, n41405, n593 );
nand U101027 ( n41405, n41406, n41407 );
nand U101028 ( n41406, n76846, n40864 );
nand U101029 ( n41407, n41264, n40697 );
nand U101030 ( n36649, n40258, n40259 );
nor U101031 ( n40259, n40260, n40261 );
nor U101032 ( n40258, n40262, n40263 );
nor U101033 ( n40260, n76412, n73997 );
nor U101034 ( n53051, n73019, n76093 );
nand U101035 ( n71371, n72383, n72384 );
nor U101036 ( n72383, n72387, n72388 );
nor U101037 ( n72384, n72385, n72386 );
nor U101038 ( n72388, n73470, n73025 );
nand U101039 ( n72453, n72808, n72809 );
nor U101040 ( n72808, n72812, n72813 );
nor U101041 ( n72809, n72810, n72811 );
nor U101042 ( n72813, n73458, n73025 );
nand U101043 ( n41195, n41398, n41399 );
nand U101044 ( n41399, n76847, n40690 );
nand U101045 ( n41398, n76845, n41203 );
nand U101046 ( n72499, n72686, n72687 );
nor U101047 ( n72686, n72690, n72691 );
nor U101048 ( n72687, n72688, n72689 );
nor U101049 ( n72691, n73464, n73025 );
nor U101050 ( n72688, n73460, n71284 );
nor U101051 ( n72810, n73037, n71284 );
nand U101052 ( n72454, n1223, n71274 );
nor U101053 ( n72385, n73040, n71284 );
nand U101054 ( n66198, n40984, n41042 );
nor U101055 ( n11588, n9895, n11594 );
xnor U101056 ( n11723, n11725, n11727 );
nor U101057 ( n52153, n76089, n73426 );
nor U101058 ( n40029, n36286, n36822 );
nor U101059 ( n66732, n76248, n73911 );
nand U101060 ( n41036, n66728, n66729 );
nor U101061 ( n66729, n66730, n66731 );
nor U101062 ( n66728, n66732, n66733 );
nor U101063 ( n66730, n76246, n73910 );
nor U101064 ( n52372, n49816, n73419 );
nand U101065 ( n72665, n71272, n72666 );
nand U101066 ( n72666, n1230, n71274 );
nor U101067 ( n10854, n9895, n10785 );
nor U101068 ( n50992, n76090, n72999 );
nor U101069 ( n72387, n73041, n71287 );
nor U101070 ( n72812, n73039, n71287 );
nor U101071 ( n17512, n73408, n17014 );
nor U101072 ( n9890, n9895, n9897 );
nor U101073 ( n72690, n73463, n71287 );
nand U101074 ( n36381, n40299, n40300 );
nor U101075 ( n40300, n40301, n40302 );
nor U101076 ( n40299, n40303, n40304 );
nor U101077 ( n40301, n76412, n73897 );
nor U101078 ( n40303, n76414, n73896 );
nor U101079 ( n52533, n76096, n73021 );
nor U101080 ( n52673, n76095, n73421 );
nor U101081 ( n51383, n49816, n73413 );
buf U101082 ( n76094, n49970 );
nand U101083 ( n72241, n71272, n72242 );
nand U101084 ( n72242, n1235, n71274 );
nor U101085 ( n51759, n50496, n76835 );
nand U101086 ( n36587, n36988, n36989 );
nand U101087 ( n36989, n76807, n36817 );
nand U101088 ( n36988, n76828, n36594 );
buf U101089 ( n76166, n17015 );
nand U101090 ( n72627, n1232, n71274 );
not U101091 ( n1937, n36467 );
nor U101092 ( n40302, n76403, n73895 );
nand U101093 ( n41578, n654, n40697 );
nand U101094 ( n37422, n2168, n36360 );
nand U101095 ( n36814, n37034, n37035 );
nand U101096 ( n37035, n76807, n36286 );
nand U101097 ( n37034, n76828, n36822 );
xnor U101098 ( n36285, n37041, n2040 );
nand U101099 ( n37041, n37042, n37043 );
nand U101100 ( n37042, n76829, n36462 );
nand U101101 ( n37043, n2035, n36293 );
xor U101102 ( n71122, n71127, n71128 );
xor U101103 ( n71127, n71323, n71324 );
xor U101104 ( n71128, n71129, n71130 );
nand U101105 ( n71323, n71326, n71327 );
nand U101106 ( n40688, n41403, n41404 );
nand U101107 ( n41404, n76847, n40864 );
nand U101108 ( n41403, n76846, n40697 );
nand U101109 ( n1561, n46931, n46932 );
nor U101110 ( n46932, n46933, n46934 );
nor U101111 ( n46931, n45406, n46939 );
nand U101112 ( n46934, n46935, n46936 );
or U101113 ( n45488, n75783, n75784 );
nor U101114 ( n75783, n573, n45492 );
nor U101115 ( n75784, n76336, n45491 );
not U101116 ( n792, n40697 );
nand U101117 ( n37445, n2167, n36672 );
not U101118 ( n1940, n36672 );
nand U101119 ( n37583, n2165, n36467 );
nor U101120 ( n66023, n66020, n40697 );
nor U101121 ( n19515, n73022, n17525 );
nand U101122 ( n71245, n72751, n72752 );
nor U101123 ( n72751, n72755, n72756 );
nor U101124 ( n72752, n72753, n72754 );
nor U101125 ( n72756, n73475, n73026 );
nor U101126 ( n72753, n73472, n71105 );
nor U101127 ( n52221, n76094, n73424 );
nand U101128 ( n40026, n36286, n36822 );
not U101129 ( n795, n40765 );
nor U101130 ( n40025, n36293, n36462 );
not U101131 ( n794, n41059 );
nor U101132 ( n37257, n36467, n76802 );
nor U101133 ( n50454, n76094, n72999 );
nor U101134 ( n19193, n73423, n17525 );
buf U101135 ( n76169, n17015 );
nand U101136 ( n72573, n71272, n72574 );
nand U101137 ( n72574, n1224, n71274 );
nor U101138 ( n18362, n73404, n17014 );
nor U101139 ( n49804, n49816, n72999 );
not U101140 ( n1237, n71143 );
nor U101141 ( n72755, n73473, n71108 );
nor U101142 ( n72287, n73476, n71284 );
nor U101143 ( n51546, n49816, n73017 );
nor U101144 ( n11583, n9955, n11594 );
buf U101145 ( n76171, n17015 );
nor U101146 ( n10904, n9955, n10785 );
nand U101147 ( n9496, n10893, n10894 );
nor U101148 ( n10894, n10895, n10897 );
nor U101149 ( n10893, n10903, n10904 );
nor U101150 ( n10895, n9908, n10899 );
nand U101151 ( n42058, n679, n41150 );
nand U101152 ( n64814, n672, n40765 );
nand U101153 ( n36817, n40180, n40181 );
nor U101154 ( n40181, n40182, n40183 );
nor U101155 ( n40180, n40184, n40185 );
nor U101156 ( n40183, n76412, n74165 );
nor U101157 ( n9952, n9955, n9897 );
nor U101158 ( n45378, n43896, n45391 );
nor U101159 ( n72289, n73477, n71287 );
nor U101160 ( n44697, n43896, n44561 );
nand U101161 ( n16226, n44687, n44688 );
nor U101162 ( n44688, n44689, n44690 );
nor U101163 ( n44687, n44696, n44697 );
nor U101164 ( n44689, n44694, n44695 );
nor U101165 ( n43895, n43896, n43799 );
nor U101166 ( n52164, n76097, n73426 );
nand U101167 ( n1546, n48067, n48068 );
nor U101168 ( n48068, n48069, n48070 );
nor U101169 ( n48067, n45406, n48076 );
nor U101170 ( n48069, n40914, n76336 );
not U101171 ( n1947, n36360 );
nand U101172 ( n36284, n37039, n37040 );
nand U101173 ( n37040, n76807, n36462 );
nand U101174 ( n37039, n76829, n36293 );
not U101175 ( n793, n40869 );
xnor U101176 ( n40860, n41408, n593 );
nand U101177 ( n41408, n41409, n41410 );
nand U101178 ( n41409, n76846, n41054 );
nand U101179 ( n41410, n40869, n41264 );
nand U101180 ( n72022, n72127, n72128 );
nand U101181 ( n72127, n72131, n71143 );
nand U101182 ( n72128, n72129, n71371 );
nand U101183 ( n72131, n71276, n72132 );
nand U101184 ( n72129, n71272, n72130 );
nand U101185 ( n72130, n1237, n71274 );
nor U101186 ( n66026, n40690, n41203 );
nor U101187 ( n19445, n17014, n73022 );
nor U101188 ( n52507, n49816, n73019 );
not U101189 ( n2655, n19292 );
buf U101190 ( n76167, n17015 );
nor U101191 ( n42281, n41466, n604 );
not U101192 ( n1953, n36767 );
nor U101193 ( n40182, n38527, n76405 );
buf U101194 ( n76165, n17015 );
xor U101195 ( n40464, n40457, n73505 );
nor U101196 ( n41482, n41490, n41491 );
nand U101197 ( n41491, n41492, n41493 );
nand U101198 ( n41492, n41494, n41495 );
nand U101199 ( n41495, n845, n41496 );
nand U101200 ( n41733, n41752, n41753 );
nand U101201 ( n41753, n40784, n76378 );
nand U101202 ( n41752, n76010, n41369 );
nor U101203 ( n41494, n41600, n41601 );
nor U101204 ( n41600, n41466, n41907 );
nor U101205 ( n41601, n41489, n41602 );
nand U101206 ( n41907, n41599, n41908 );
and U101207 ( n41732, n41750, n41751 );
nand U101208 ( n41750, n76010, n40784 );
nand U101209 ( n41751, n41369, n76378 );
nand U101210 ( n1861, n41480, n41481 );
nor U101211 ( n41480, n41964, n41965 );
nor U101212 ( n41481, n41482, n41483 );
nor U101213 ( n41965, n41966, n74537 );
nand U101214 ( n41735, n41756, n41757 );
nand U101215 ( n41757, n41036, n76378 );
nand U101216 ( n41756, n76010, n40789 );
and U101217 ( n41734, n41754, n41755 );
nand U101218 ( n41754, n76010, n41036 );
nand U101219 ( n41755, n40789, n76378 );
nand U101220 ( n42081, n660, n40869 );
nor U101221 ( n51795, n76087, n73425 );
nor U101222 ( n50985, n76092, n73400 );
nor U101223 ( n16874, n73408, n76161 );
buf U101224 ( n76161, n17016 );
nor U101225 ( n16965, n16966, n73417 );
nand U101226 ( n36286, n40138, n40139 );
nor U101227 ( n40139, n40140, n40141 );
nor U101228 ( n40138, n40143, n40144 );
nor U101229 ( n40141, n76412, n74234 );
nor U101230 ( n17778, n73406, n17014 );
nand U101231 ( n36481, n37774, n37775 );
nand U101232 ( n37775, n37300, n37097 );
nand U101233 ( n37774, n37765, n37776 );
nor U101234 ( n37765, n37097, n2088 );
and U101235 ( n41730, n41760, n41761 );
nand U101236 ( n41760, n76010, n41377 );
nand U101237 ( n41761, n41378, n76379 );
nand U101238 ( n41767, n624, n41768 );
nand U101239 ( n41768, n76010, n41769 );
nand U101240 ( n41731, n41762, n41763 );
nand U101241 ( n41763, n41377, n76378 );
nand U101242 ( n41762, n76010, n41378 );
nand U101243 ( n71357, n72177, n72178 );
nor U101244 ( n72177, n72181, n72182 );
nor U101245 ( n72178, n72179, n72180 );
nor U101246 ( n72182, n73484, n73025 );
nand U101247 ( n41743, n41774, n41775 );
nand U101248 ( n41774, n76011, n41198 );
nand U101249 ( n41775, n40989, n76378 );
nand U101250 ( n36589, n40215, n40216 );
nor U101251 ( n40216, n40217, n40218 );
nor U101252 ( n40215, n40219, n40220 );
nor U101253 ( n40218, n76412, n74218 );
nor U101254 ( n40219, n76414, n74220 );
not U101255 ( n6259, n72801 );
nor U101256 ( n72179, n73043, n71284 );
xnor U101257 ( n36458, n37044, n2040 );
nand U101258 ( n37044, n37045, n37046 );
nand U101259 ( n37045, n76829, n36667 );
nand U101260 ( n37046, n36467, n2035 );
nor U101261 ( n37253, n36672, n76801 );
nor U101262 ( n51210, n49816, n73412 );
and U101263 ( n41742, n41776, n41777 );
nand U101264 ( n41777, n41198, n76379 );
nand U101265 ( n41776, n76011, n40989 );
nor U101266 ( n51086, n76095, n73003 );
nor U101267 ( n72181, n73044, n71287 );
nand U101268 ( n40826, n42289, n42290 );
nand U101269 ( n42290, n41493, n41466 );
nand U101270 ( n42289, n42281, n42291 );
nor U101271 ( n16990, n76572, n73000 );
nand U101272 ( n41737, n41744, n41745 );
nand U101273 ( n41744, n76010, n40984 );
nand U101274 ( n41745, n41042, n76378 );
not U101275 ( n797, n41150 );
buf U101276 ( n76162, n17016 );
or U101277 ( n19279, n73418, n76162 );
nand U101278 ( n39899, n36467, n36667 );
nor U101279 ( n52800, n49816, n73421 );
nand U101280 ( n40984, n66424, n66425 );
nor U101281 ( n66425, n66426, n66427 );
nor U101282 ( n66424, n66428, n66429 );
nor U101283 ( n66427, n76246, n74217 );
nor U101284 ( n66428, n76248, n74219 );
nor U101285 ( n40217, n2930, n76405 );
not U101286 ( n2930, n36654 );
nand U101287 ( n72017, n71272, n72018 );
nand U101288 ( n72018, n1238, n71274 );
and U101289 ( n71887, n72015, n72016 );
nand U101290 ( n72015, n72019, n71357 );
nand U101291 ( n72016, n72017, n71143 );
nand U101292 ( n72019, n71276, n72020 );
nor U101293 ( n18959, n73015, n76163 );
buf U101294 ( n76163, n17016 );
and U101295 ( n41736, n41746, n41747 );
nand U101296 ( n41747, n40984, n76378 );
nand U101297 ( n41746, n76010, n41042 );
nand U101298 ( n42079, n667, n41059 );
nand U101299 ( n40863, n41346, n41347 );
nand U101300 ( n41347, n76847, n41054 );
nand U101301 ( n41346, n76845, n40869 );
nand U101302 ( n37420, n2169, n36767 );
nor U101303 ( n37245, n36360, n76801 );
xnor U101304 ( n41050, n41411, n593 );
nand U101305 ( n41411, n41412, n41413 );
nand U101306 ( n41412, n76846, n40760 );
nand U101307 ( n41413, n41059, n41264 );
buf U101308 ( n76168, n17015 );
nor U101309 ( n65343, n41145, n40765 );
not U101310 ( n1959, n36537 );
nor U101311 ( n65824, n40760, n41059 );
nor U101312 ( n50979, n49816, n73008 );
not U101313 ( n7799, n44548 );
nand U101314 ( n43287, n48005, n48006 );
or U101315 ( n48006, n73497, n44142 );
nor U101316 ( n45630, n46440, n76005 );
not U101317 ( n7544, n47204 );
nor U101318 ( n47770, n73538, n47381 );
not U101319 ( n7538, n46875 );
nand U101320 ( n46581, n46613, n46614 );
nor U101321 ( n46613, n46615, n46616 );
nor U101322 ( n46616, n76005, n46617 );
nor U101323 ( n46615, n46618, n73159 );
not U101324 ( n7539, n47021 );
not U101325 ( n7534, n46692 );
nand U101326 ( n46914, n46962, n46963 );
nor U101327 ( n46962, n46964, n46965 );
nor U101328 ( n46965, n76005, n74417 );
nor U101329 ( n46964, n46966, n46967 );
nand U101330 ( n46871, n46879, n76341 );
nand U101331 ( n46879, n7538, n73118 );
nand U101332 ( n46967, n46968, n7539 );
nand U101333 ( n47766, n47767, n47768 );
nor U101334 ( n47767, n47771, n47772 );
nor U101335 ( n47768, n47769, n47770 );
nor U101336 ( n47771, n73549, n47386 );
nand U101337 ( n46304, n76657, n45546 );
nor U101338 ( n46478, n46521, n46522 );
and U101339 ( n46522, n46482, n76342 );
and U101340 ( n46618, n46617, n76006 );
not U101341 ( n1967, n36735 );
nor U101342 ( n47776, n73541, n47391 );
nand U101343 ( n47765, n47773, n47774 );
nor U101344 ( n47773, n47777, n47778 );
nor U101345 ( n47774, n47775, n47776 );
nor U101346 ( n47777, n73550, n47396 );
nor U101347 ( n47769, n73543, n47382 );
not U101348 ( n3632, n72831 );
nor U101349 ( n47775, n73546, n47392 );
nor U101350 ( n11578, n9974, n11594 );
xnor U101351 ( n11698, n11700, n11702 );
nor U101352 ( n66426, n1813, n76243 );
not U101353 ( n1813, n41041 );
nor U101354 ( n47772, n73552, n47385 );
nand U101355 ( n72518, n71574, n71243 );
nor U101356 ( n47778, n73548, n47395 );
nor U101357 ( n72701, n73045, n71105 );
nor U101358 ( n50724, n76099, n73400 );
nor U101359 ( n10955, n9974, n10785 );
nand U101360 ( n9491, n10943, n10944 );
nor U101361 ( n10944, n10945, n10947 );
nor U101362 ( n10943, n10954, n10955 );
nor U101363 ( n10945, n10952, n10953 );
nor U101364 ( n9973, n9974, n9897 );
not U101365 ( n7805, n44894 );
nand U101366 ( n39896, n36355, n36672 );
not U101367 ( n7533, n45627 );
nor U101368 ( n47849, n44132, n54215 );
nor U101369 ( n54215, n73511, n7805 );
nor U101370 ( n47756, n73534, n47359 );
nand U101371 ( n47752, n47753, n47754 );
nor U101372 ( n47753, n47757, n47758 );
nor U101373 ( n47754, n47755, n47756 );
nor U101374 ( n47757, n73545, n47364 );
nor U101375 ( n47755, n73537, n47360 );
nor U101376 ( n47758, n73539, n47363 );
nand U101377 ( n39893, n36360, n36762 );
not U101378 ( n1975, n36955 );
buf U101379 ( n76842, n76837 );
buf U101380 ( n76837, n76838 );
not U101381 ( n6012, n65423 );
nand U101382 ( n63972, n69013, n69014 );
or U101383 ( n69014, n73502, n64984 );
not U101384 ( n5758, n68235 );
nor U101385 ( n68791, n73588, n68413 );
nor U101386 ( n11196, n67355, n67356 );
nor U101387 ( n67356, n67357, n67358 );
nor U101388 ( n67355, n67359, n67360 );
nand U101389 ( n67359, n67386, n67387 );
nand U101390 ( n67961, n67997, n67998 );
nor U101391 ( n67997, n67999, n68000 );
nor U101392 ( n68000, n75989, n74431 );
nor U101393 ( n67999, n68001, n68002 );
nand U101394 ( n68787, n68788, n68789 );
nor U101395 ( n68788, n68792, n68793 );
nor U101396 ( n68789, n68790, n68791 );
nor U101397 ( n68792, n73612, n68418 );
not U101398 ( n4234, n23877 );
not U101399 ( n6867, n57001 );
nand U101400 ( n22693, n27016, n27017 );
or U101401 ( n27017, n73503, n23475 );
nand U101402 ( n55809, n60157, n60158 );
or U101403 ( n60158, n73504, n56597 );
nor U101404 ( n24719, n25499, n76026 );
nor U101405 ( n66554, n67504, n75989 );
nor U101406 ( n57853, n58636, n75997 );
not U101407 ( n4000, n26234 );
not U101408 ( n6633, n59373 );
not U101409 ( n5752, n67922 );
not U101410 ( n3994, n25919 );
not U101411 ( n6627, n59057 );
nand U101412 ( n67628, n67660, n67661 );
nor U101413 ( n67660, n67662, n67663 );
nor U101414 ( n67663, n75989, n67664 );
nor U101415 ( n67662, n67665, n74637 );
not U101416 ( n5753, n68056 );
nand U101417 ( n25623, n25655, n25656 );
nor U101418 ( n25655, n25657, n25658 );
nor U101419 ( n25658, n76026, n25659 );
nor U101420 ( n25657, n25660, n74638 );
nand U101421 ( n58760, n58795, n58796 );
nor U101422 ( n58795, n58797, n58798 );
nor U101423 ( n58798, n75997, n58799 );
nor U101424 ( n58797, n58800, n74639 );
not U101425 ( n3995, n26053 );
not U101426 ( n6628, n59194 );
nor U101427 ( n25361, n24633, n25364 );
nor U101428 ( n67366, n66470, n67369 );
nor U101429 ( n58498, n57765, n58501 );
not U101430 ( n5748, n67739 );
nor U101431 ( n6706, n25350, n25351 );
nor U101432 ( n25351, n25352, n25353 );
nor U101433 ( n25350, n25354, n25355 );
nand U101434 ( n25354, n25381, n25382 );
nor U101435 ( n13441, n58487, n58488 );
nor U101436 ( n58488, n58489, n58490 );
nor U101437 ( n58487, n58491, n58492 );
nand U101438 ( n58491, n58518, n58519 );
nand U101439 ( n25958, n25994, n25995 );
nor U101440 ( n25994, n25996, n25997 );
nor U101441 ( n25997, n76026, n74432 );
nor U101442 ( n25996, n25998, n25999 );
nand U101443 ( n59096, n59132, n59133 );
nor U101444 ( n59132, n59134, n59135 );
nor U101445 ( n59135, n75997, n74433 );
nor U101446 ( n59134, n59136, n59137 );
nand U101447 ( n67360, n67361, n485 );
not U101448 ( n485, n67358 );
nor U101449 ( n67361, n67366, n67367 );
and U101450 ( n67367, n66472, n76708 );
nand U101451 ( n67918, n67926, n76197 );
nand U101452 ( n67926, n5752, n73130 );
nand U101453 ( n25915, n25923, n76521 );
nand U101454 ( n25923, n3994, n73131 );
nand U101455 ( n59053, n59061, n76263 );
nand U101456 ( n59061, n6627, n73132 );
nand U101457 ( n26788, n26789, n26790 );
nor U101458 ( n26789, n26793, n26794 );
nor U101459 ( n26790, n26791, n26792 );
nor U101460 ( n26793, n73630, n26417 );
nand U101461 ( n59928, n59929, n59930 );
nor U101462 ( n59929, n59933, n59934 );
nor U101463 ( n59930, n59931, n59932 );
nor U101464 ( n59933, n73629, n59556 );
nand U101465 ( n25355, n25356, n180 );
not U101466 ( n180, n25353 );
nor U101467 ( n25356, n25361, n25362 );
and U101468 ( n25362, n24635, n76754 );
nand U101469 ( n58492, n58493, n452 );
not U101470 ( n452, n58490 );
nor U101471 ( n58493, n58498, n58499 );
and U101472 ( n58499, n57767, n76687 );
nor U101473 ( n67541, n67582, n67583 );
and U101474 ( n67583, n67545, n76198 );
nor U101475 ( n26792, n73605, n26412 );
nor U101476 ( n59932, n73604, n59551 );
not U101477 ( n3990, n25734 );
not U101478 ( n6623, n58874 );
nand U101479 ( n68002, n68003, n5753 );
nand U101480 ( n25999, n26000, n3995 );
nand U101481 ( n59137, n59138, n6628 );
nor U101482 ( n25536, n25577, n25578 );
and U101483 ( n25578, n25540, n76522 );
nor U101484 ( n58673, n58714, n58715 );
and U101485 ( n58715, n58677, n76264 );
and U101486 ( n67665, n67664, n75990 );
and U101487 ( n25660, n25659, n76027 );
and U101488 ( n58800, n58799, n75998 );
nor U101489 ( n68797, n73592, n68423 );
nand U101490 ( n68786, n68794, n68795 );
nor U101491 ( n68794, n68798, n68799 );
nor U101492 ( n68795, n68796, n68797 );
nor U101493 ( n68798, n73621, n68428 );
nor U101494 ( n26798, n73614, n26422 );
nor U101495 ( n59938, n73613, n59561 );
nand U101496 ( n26787, n26795, n26796 );
nor U101497 ( n26795, n26799, n26800 );
nor U101498 ( n26796, n26797, n26798 );
nor U101499 ( n26799, n73632, n26427 );
nand U101500 ( n59927, n59935, n59936 );
nor U101501 ( n59935, n59939, n59940 );
nor U101502 ( n59936, n59937, n59938 );
nor U101503 ( n59939, n73631, n59566 );
nand U101504 ( n71882, n71272, n71883 );
nand U101505 ( n71883, n1239, n71274 );
and U101506 ( n71741, n71880, n71881 );
nand U101507 ( n71880, n71884, n71327 );
nand U101508 ( n71881, n71882, n71357 );
nand U101509 ( n71884, n71276, n71885 );
nor U101510 ( n68790, n73595, n68414 );
nor U101511 ( n72060, n73489, n71284 );
nor U101512 ( n26791, n73618, n26413 );
nor U101513 ( n59931, n73617, n59552 );
nor U101514 ( n68796, n73602, n68424 );
nor U101515 ( n26797, n73623, n26423 );
nor U101516 ( n59937, n73622, n59562 );
nand U101517 ( n71267, n71608, n71609 );
nor U101518 ( n71608, n71612, n71613 );
nor U101519 ( n71609, n71610, n71611 );
nor U101520 ( n71613, n73480, n73025 );
nor U101521 ( n68793, n73628, n68417 );
nor U101522 ( n26794, n73635, n26416 );
nor U101523 ( n59934, n73634, n59555 );
buf U101524 ( n76159, n17016 );
nor U101525 ( n18688, n73414, n76159 );
nor U101526 ( n68799, n73610, n68427 );
nor U101527 ( n26800, n73627, n26426 );
nor U101528 ( n59940, n73626, n59565 );
nor U101529 ( n51724, n76098, n73425 );
nor U101530 ( n20095, n76158, n73420 );
buf U101531 ( n76158, n17016 );
nor U101532 ( n72703, n73046, n71108 );
not U101533 ( n4240, n24215 );
not U101534 ( n6873, n57337 );
not U101535 ( n6018, n65759 );
nor U101536 ( n18823, n73422, n17525 );
nor U101537 ( n47717, n73576, n47381 );
nand U101538 ( n47713, n47714, n47715 );
nor U101539 ( n47714, n47718, n47719 );
nor U101540 ( n47715, n47716, n47717 );
nor U101541 ( n47718, n73593, n47386 );
nand U101542 ( n71605, n1233, n71274 );
nor U101543 ( n47723, n73580, n47391 );
nand U101544 ( n47712, n47720, n47721 );
nor U101545 ( n47720, n47724, n47725 );
nor U101546 ( n47721, n47722, n47723 );
nor U101547 ( n47724, n73599, n47396 );
nor U101548 ( n47716, n73582, n47382 );
nor U101549 ( n47722, n73586, n47392 );
nor U101550 ( n47719, n73611, n47385 );
nor U101551 ( n47725, n73591, n47395 );
not U101552 ( n3989, n24717 );
not U101553 ( n5747, n66552 );
not U101554 ( n6622, n57851 );
nor U101555 ( n52649, n49816, n73021 );
or U101556 ( n18368, n75913, n76163 );
nor U101557 ( n47760, n47761, n47762 );
nor U101558 ( n47761, n73540, n47370 );
nor U101559 ( n47762, n73536, n47369 );
nor U101560 ( n68869, n64974, n70443 );
nor U101561 ( n70443, n73515, n6018 );
nor U101562 ( n68777, n73564, n68391 );
nand U101563 ( n68773, n68774, n68775 );
nor U101564 ( n68774, n68778, n68779 );
nor U101565 ( n68775, n68776, n68777 );
nor U101566 ( n68778, n73596, n68396 );
nor U101567 ( n26870, n23465, n28538 );
nor U101568 ( n28538, n73516, n4240 );
nor U101569 ( n60010, n56587, n61843 );
nor U101570 ( n61843, n73517, n6873 );
nor U101571 ( n26778, n73569, n26390 );
nor U101572 ( n59918, n73568, n59529 );
nand U101573 ( n26774, n26775, n26776 );
nor U101574 ( n26775, n26779, n26780 );
nor U101575 ( n26776, n26777, n26778 );
nor U101576 ( n26779, n73620, n26395 );
nand U101577 ( n59914, n59915, n59916 );
nor U101578 ( n59915, n59919, n59920 );
nor U101579 ( n59916, n59917, n59918 );
nor U101580 ( n59919, n73619, n59534 );
nor U101581 ( n68776, n73585, n68392 );
nor U101582 ( n26777, n73601, n26391 );
nor U101583 ( n59917, n73600, n59530 );
nand U101584 ( n36461, n36981, n36982 );
nand U101585 ( n36982, n76807, n36667 );
nand U101586 ( n36981, n76828, n36467 );
nand U101587 ( n37569, n2170, n36537 );
nor U101588 ( n47759, n47763, n47764 );
nor U101589 ( n47763, n73547, n47374 );
nor U101590 ( n47764, n73542, n47373 );
nor U101591 ( n68779, n73589, n68395 );
nor U101592 ( n26780, n73607, n26394 );
nor U101593 ( n59920, n73606, n59533 );
nor U101594 ( n72062, n73490, n71287 );
nor U101595 ( n47703, n73558, n47359 );
nand U101596 ( n47699, n47700, n47701 );
nor U101597 ( n47700, n47704, n47705 );
nor U101598 ( n47701, n47702, n47703 );
nor U101599 ( n47704, n73584, n47364 );
xnor U101600 ( n41113, n41426, n593 );
nand U101601 ( n41426, n41427, n41428 );
nand U101602 ( n41427, n76846, n40727 );
nand U101603 ( n41428, n41119, n41264 );
nor U101604 ( n47702, n73575, n47360 );
xor U101605 ( n40926, n41433, n593 );
nand U101606 ( n41433, n41434, n41435 );
nand U101607 ( n41434, n76846, n41114 );
nand U101608 ( n41435, n40935, n41264 );
nor U101609 ( n47705, n73577, n47363 );
nand U101610 ( n41773, n41778, n41779 );
nand U101611 ( n41778, n76011, n40690 );
nand U101612 ( n41779, n41203, n76379 );
nor U101613 ( n26737, n73713, n26412 );
nor U101614 ( n68738, n73710, n68413 );
nor U101615 ( n59879, n73712, n59551 );
nand U101616 ( n26733, n26734, n26735 );
nor U101617 ( n26734, n26738, n26739 );
nor U101618 ( n26735, n26736, n26737 );
nor U101619 ( n26738, n73742, n26417 );
nand U101620 ( n68734, n68735, n68736 );
nor U101621 ( n68735, n68739, n68740 );
nor U101622 ( n68736, n68737, n68738 );
nor U101623 ( n68739, n73740, n68418 );
nand U101624 ( n59875, n59876, n59877 );
nor U101625 ( n59876, n59880, n59881 );
nor U101626 ( n59877, n59878, n59879 );
nor U101627 ( n59880, n73741, n59556 );
nor U101628 ( n26743, n73721, n26422 );
nor U101629 ( n68744, n73719, n68423 );
nor U101630 ( n59885, n73720, n59561 );
nand U101631 ( n26732, n26740, n26741 );
nor U101632 ( n26740, n26744, n26745 );
nor U101633 ( n26741, n26742, n26743 );
nor U101634 ( n26744, n73745, n26427 );
nand U101635 ( n68733, n68741, n68742 );
nor U101636 ( n68741, n68745, n68746 );
nor U101637 ( n68742, n68743, n68744 );
nor U101638 ( n68745, n73743, n68428 );
nand U101639 ( n59874, n59882, n59883 );
nor U101640 ( n59882, n59886, n59887 );
nor U101641 ( n59883, n59884, n59885 );
nor U101642 ( n59886, n73744, n59566 );
nor U101643 ( n26736, n73727, n26413 );
nor U101644 ( n68737, n73725, n68414 );
nor U101645 ( n59878, n73726, n59552 );
nor U101646 ( n26742, n73733, n26423 );
nor U101647 ( n68743, n73731, n68424 );
nor U101648 ( n59884, n73732, n59562 );
nand U101649 ( n38351, n38352, n38353 );
nand U101650 ( n38353, n76816, n36577 );
nand U101651 ( n38352, n76812, n38354 );
nor U101652 ( n26739, n73748, n26416 );
nor U101653 ( n68740, n73746, n68417 );
nor U101654 ( n59881, n73747, n59555 );
nor U101655 ( n26745, n73739, n26426 );
nor U101656 ( n68746, n73737, n68427 );
nor U101657 ( n59887, n73738, n59565 );
nand U101658 ( n47121, n47157, n47158 );
nand U101659 ( n47158, n47159, n76341 );
nand U101660 ( n47159, n7544, n73078 );
nor U101661 ( n18440, n73012, n76162 );
nand U101662 ( n71624, n71243, n71413 );
buf U101663 ( n76170, n17015 );
and U101664 ( n41772, n41780, n41781 );
nand U101665 ( n41781, n76380, n40690 );
nand U101666 ( n41780, n76011, n41203 );
nor U101667 ( n68781, n68782, n68783 );
nor U101668 ( n68782, n73590, n68402 );
nor U101669 ( n68783, n73583, n68401 );
nor U101670 ( n26782, n26783, n26784 );
nor U101671 ( n26783, n73609, n26401 );
nor U101672 ( n26784, n73598, n26400 );
nor U101673 ( n59922, n59923, n59924 );
nor U101674 ( n59923, n73608, n59540 );
nor U101675 ( n59924, n73597, n59539 );
not U101676 ( n798, n40935 );
nor U101677 ( n68780, n68784, n68785 );
nor U101678 ( n68784, n73603, n68406 );
nor U101679 ( n68785, n73594, n68405 );
nor U101680 ( n26781, n26785, n26786 );
nor U101681 ( n26785, n73625, n26405 );
nor U101682 ( n26786, n73616, n26404 );
nor U101683 ( n59921, n59925, n59926 );
nor U101684 ( n59925, n73624, n59544 );
nor U101685 ( n59926, n73615, n59543 );
nor U101686 ( n50153, n49816, n73400 );
nor U101687 ( n47707, n47708, n47709 );
nor U101688 ( n47708, n73578, n47370 );
nor U101689 ( n47709, n73573, n47369 );
nand U101690 ( n39747, n36767, n36532 );
nor U101691 ( n26723, n73671, n26390 );
nor U101692 ( n68724, n73666, n68391 );
nor U101693 ( n59865, n73670, n59529 );
nand U101694 ( n26719, n26720, n26721 );
nor U101695 ( n26720, n26724, n26725 );
nor U101696 ( n26721, n26722, n26723 );
nor U101697 ( n26724, n73730, n26395 );
nand U101698 ( n68720, n68721, n68722 );
nor U101699 ( n68721, n68725, n68726 );
nor U101700 ( n68722, n68723, n68724 );
nor U101701 ( n68725, n73728, n68396 );
nand U101702 ( n59861, n59862, n59863 );
nor U101703 ( n59862, n59866, n59867 );
nor U101704 ( n59863, n59864, n59865 );
nor U101705 ( n59866, n73729, n59534 );
nor U101706 ( n52328, n49816, n73424 );
nor U101707 ( n26722, n73709, n26391 );
nor U101708 ( n68723, n73707, n68392 );
nor U101709 ( n59864, n73708, n59530 );
nor U101710 ( n44142, n44894, n73511 );
nand U101711 ( n41198, n66351, n66352 );
nor U101712 ( n66352, n66353, n66354 );
nor U101713 ( n66351, n66355, n66356 );
nor U101714 ( n66354, n76246, n74259 );
nor U101715 ( n66355, n76248, n74263 );
nor U101716 ( n47706, n47710, n47711 );
nor U101717 ( n47710, n73587, n47374 );
nor U101718 ( n47711, n73581, n47373 );
nor U101719 ( n26725, n73716, n26394 );
nor U101720 ( n68726, n73714, n68395 );
nor U101721 ( n59867, n73715, n59533 );
nand U101722 ( n41685, n41710, n41711 );
nand U101723 ( n41710, n76011, n40760 );
nand U101724 ( n41711, n41059, n76378 );
nand U101725 ( n40690, n66274, n66275 );
nor U101726 ( n66275, n66276, n66277 );
nor U101727 ( n66274, n66279, n66280 );
nor U101728 ( n66277, n76246, n74281 );
nor U101729 ( n66279, n76248, n74282 );
nand U101730 ( n71447, n1240, n71274 );
nand U101731 ( n72146, n71143, n71245 );
nor U101732 ( n45454, n50543, n76835 );
nand U101733 ( n41694, n41706, n41707 );
nand U101734 ( n41706, n76010, n41054 );
nand U101735 ( n41707, n40869, n76378 );
nand U101736 ( n41697, n41708, n41709 );
nand U101737 ( n41709, n76380, n41054 );
nand U101738 ( n41708, n76010, n40869 );
nand U101739 ( n39749, n36730, n36537 );
nand U101740 ( n68152, n68188, n68189 );
nand U101741 ( n68189, n68190, n76197 );
nand U101742 ( n68190, n5758, n73084 );
not U101743 ( n1383, n52663 );
nor U101744 ( n19860, n73018, n76164 );
nand U101745 ( n26151, n26187, n26188 );
nand U101746 ( n26188, n26189, n76521 );
nand U101747 ( n26189, n4000, n73085 );
nand U101748 ( n59290, n59326, n59327 );
nand U101749 ( n59327, n59328, n76263 );
nand U101750 ( n59328, n6633, n73086 );
buf U101751 ( n76164, n17016 );
nand U101752 ( n42045, n684, n40935 );
nand U101753 ( n66467, n66468, n66469 );
nand U101754 ( n66468, n76720, n66472 );
or U101755 ( n66469, n66470, n66471 );
nand U101756 ( n11356, n66447, n66448 );
nor U101757 ( n66448, n66449, n66450 );
nor U101758 ( n66447, n66466, n66467 );
nand U101759 ( n66449, n66458, n66459 );
nand U101760 ( n24630, n24631, n24632 );
nand U101761 ( n24631, n76768, n24635 );
or U101762 ( n24632, n24633, n24634 );
nand U101763 ( n57762, n57763, n57764 );
nand U101764 ( n57763, n76701, n57767 );
or U101765 ( n57764, n57765, n57766 );
nand U101766 ( n6866, n24610, n24611 );
nor U101767 ( n24611, n24612, n24613 );
nor U101768 ( n24610, n24629, n24630 );
nand U101769 ( n24612, n24621, n24622 );
nand U101770 ( n13601, n57742, n57743 );
nor U101771 ( n57743, n57744, n57745 );
nor U101772 ( n57742, n57761, n57762 );
nand U101773 ( n57744, n57753, n57754 );
nor U101774 ( n18039, n75911, n17014 );
nor U101775 ( n37241, n36767, n76801 );
nor U101776 ( n51533, n49982, n73019 );
xor U101777 ( n36528, n37066, n2040 );
nand U101778 ( n37066, n37067, n37068 );
nand U101779 ( n37067, n76829, n36730 );
nand U101780 ( n37068, n36537, n2035 );
nor U101781 ( n19717, n73020, n76158 );
and U101782 ( n41684, n41712, n41713 );
nand U101783 ( n41713, n40760, n76378 );
nand U101784 ( n41712, n76010, n41059 );
nor U101785 ( n26727, n26728, n26729 );
nor U101786 ( n26728, n73718, n26401 );
nor U101787 ( n26729, n73706, n26400 );
nor U101788 ( n68728, n68729, n68730 );
nor U101789 ( n68729, n73711, n68402 );
nor U101790 ( n68730, n73701, n68401 );
nor U101791 ( n59869, n59870, n59871 );
nor U101792 ( n59870, n73717, n59540 );
nor U101793 ( n59871, n73705, n59539 );
nand U101794 ( n45543, n45544, n45545 );
nand U101795 ( n45544, n76672, n45547 );
nand U101796 ( n45545, n45546, n76662 );
nand U101797 ( n15846, n45523, n45524 );
nor U101798 ( n45524, n45525, n45526 );
nor U101799 ( n45523, n45542, n45543 );
nand U101800 ( n45525, n45534, n45535 );
nor U101801 ( n47640, n73638, n47381 );
nand U101802 ( n47636, n47637, n47638 );
nor U101803 ( n47637, n47641, n47642 );
nor U101804 ( n47638, n47639, n47640 );
nor U101805 ( n47641, n73650, n47386 );
nand U101806 ( n41052, n41341, n41342 );
nand U101807 ( n41342, n76847, n40760 );
nand U101808 ( n41341, n76844, n41059 );
nand U101809 ( n44889, n73052, n73512 );
nand U101810 ( n47864, n44889, n44894 );
not U101811 ( n7807, n44515 );
nor U101812 ( n47646, n73647, n47391 );
nand U101813 ( n47635, n47643, n47644 );
nor U101814 ( n47643, n47647, n47648 );
nor U101815 ( n47644, n47645, n47646 );
nor U101816 ( n47647, n73664, n47396 );
nor U101817 ( n64984, n65759, n73515 );
nor U101818 ( n23475, n24215, n73516 );
nor U101819 ( n56597, n57337, n73517 );
nor U101820 ( n47639, n73646, n47382 );
nor U101821 ( n47645, n73662, n47392 );
nand U101822 ( n44517, n7809, n73512 );
nor U101823 ( n26726, n26730, n26731 );
nor U101824 ( n26730, n73736, n26405 );
nor U101825 ( n26731, n73724, n26404 );
nor U101826 ( n68727, n68731, n68732 );
nor U101827 ( n68731, n73734, n68406 );
nor U101828 ( n68732, n73722, n68405 );
nor U101829 ( n59868, n59872, n59873 );
nor U101830 ( n59872, n73735, n59544 );
nor U101831 ( n59873, n73723, n59543 );
xnor U101832 ( n36729, n37059, n2040 );
nand U101833 ( n37059, n37060, n37061 );
nand U101834 ( n37060, n76829, n36322 );
nand U101835 ( n37061, n36735, n2035 );
nor U101836 ( n47642, n73640, n47385 );
nor U101837 ( n47648, n73651, n47395 );
nand U101838 ( n39748, n36735, n36322 );
xnor U101839 ( n40756, n41414, n593 );
nand U101840 ( n41414, n41415, n41416 );
nand U101841 ( n41415, n76846, n41145 );
nand U101842 ( n41416, n40765, n41264 );
xor U101843 ( n36663, n36973, n36481 );
nand U101844 ( n36973, n36974, n36975 );
nand U101845 ( n36974, n76827, n36355 );
nand U101846 ( n36975, n36672, n2035 );
not U101847 ( n1969, n36327 );
xnor U101848 ( n41142, n41423, n593 );
nand U101849 ( n41423, n41424, n41425 );
nand U101850 ( n41424, n76846, n40930 );
nand U101851 ( n41425, n41150, n41264 );
nand U101852 ( n37567, n2172, n36735 );
nand U101853 ( n38319, n38320, n38321 );
nand U101854 ( n38321, n76815, n36802 );
nand U101855 ( n38320, n76812, n38322 );
nand U101856 ( n71266, n71450, n71451 );
nor U101857 ( n71450, n71454, n71455 );
nor U101858 ( n71451, n71452, n71453 );
nor U101859 ( n71455, n73492, n73025 );
nor U101860 ( n71452, n73048, n71284 );
nor U101861 ( n47626, n73636, n47359 );
nand U101862 ( n47622, n47623, n47624 );
nor U101863 ( n47623, n47627, n47628 );
nor U101864 ( n47624, n47625, n47626 );
nor U101865 ( n47627, n73648, n47364 );
nor U101866 ( n47625, n73644, n47360 );
nand U101867 ( n41112, n41429, n41430 );
nand U101868 ( n41430, n76847, n40727 );
nand U101869 ( n41429, n76846, n41119 );
nand U101870 ( n36665, n36976, n36977 );
nand U101871 ( n36977, n76807, n36355 );
nand U101872 ( n36976, n76827, n36672 );
nor U101873 ( n47628, n73639, n47363 );
and U101874 ( n40925, n41431, n41432 );
nand U101875 ( n41432, n76847, n41114 );
nand U101876 ( n41431, n76846, n40935 );
nor U101877 ( n52072, n49816, n73426 );
nor U101878 ( n64514, n41114, n40935 );
not U101879 ( n799, n41119 );
nor U101880 ( n66353, n54672, n76243 );
nor U101881 ( n68661, n73752, n68413 );
nor U101882 ( n26660, n73753, n26412 );
nor U101883 ( n59802, n73754, n59551 );
nand U101884 ( n68657, n68658, n68659 );
nor U101885 ( n68658, n68662, n68663 );
nor U101886 ( n68659, n68660, n68661 );
nor U101887 ( n68662, n73779, n68418 );
nand U101888 ( n26656, n26657, n26658 );
nor U101889 ( n26657, n26661, n26662 );
nor U101890 ( n26658, n26659, n26660 );
nor U101891 ( n26661, n73780, n26417 );
nand U101892 ( n59798, n59799, n59800 );
nor U101893 ( n59799, n59803, n59804 );
nor U101894 ( n59800, n59801, n59802 );
nor U101895 ( n59803, n73781, n59556 );
nand U101896 ( n65754, n73053, n73518 );
nand U101897 ( n26885, n24210, n24215 );
nand U101898 ( n60025, n57332, n57337 );
nand U101899 ( n68884, n65754, n65759 );
not U101900 ( n4242, n23844 );
not U101901 ( n6874, n56968 );
not U101902 ( n6019, n65390 );
nor U101903 ( n68667, n73768, n68423 );
nor U101904 ( n26666, n73771, n26422 );
nor U101905 ( n59808, n73772, n59561 );
nand U101906 ( n68656, n68664, n68665 );
nor U101907 ( n68664, n68668, n68669 );
nor U101908 ( n68665, n68666, n68667 );
nor U101909 ( n68668, n73794, n68428 );
nand U101910 ( n26655, n26663, n26664 );
nor U101911 ( n26663, n26667, n26668 );
nor U101912 ( n26664, n26665, n26666 );
nor U101913 ( n26667, n73795, n26427 );
nand U101914 ( n59797, n59805, n59806 );
nor U101915 ( n59805, n59809, n59810 );
nor U101916 ( n59806, n59807, n59808 );
nor U101917 ( n59809, n73796, n59566 );
nand U101918 ( n24210, n73055, n73520 );
nand U101919 ( n57332, n73054, n73521 );
nor U101920 ( n68660, n73767, n68414 );
nor U101921 ( n26659, n73769, n26413 );
nor U101922 ( n59801, n73770, n59552 );
nor U101923 ( n68666, n73788, n68424 );
nor U101924 ( n26665, n73789, n26423 );
nor U101925 ( n59807, n73790, n59562 );
nand U101926 ( n65392, n6022, n73518 );
nand U101927 ( n23846, n4244, n73520 );
nand U101928 ( n56970, n6877, n73521 );
nor U101929 ( n68663, n73758, n68417 );
nor U101930 ( n26662, n73759, n26416 );
nor U101931 ( n59804, n73760, n59555 );
nor U101932 ( n68669, n73782, n68427 );
nor U101933 ( n26668, n73783, n26426 );
nor U101934 ( n59810, n73784, n59565 );
nand U101935 ( n37501, n2173, n36327 );
nor U101936 ( n19263, n16861, n73018 );
xnor U101937 ( n45563, n46311, n46370 );
xor U101938 ( n46370, n75016, n76342 );
nor U101939 ( n46337, n46339, n76330 );
nor U101940 ( n46339, n46340, n46341 );
nand U101941 ( n46341, n46342, n46343 );
nand U101942 ( n46340, n46344, n46345 );
nor U101943 ( n37496, n36577, n2175 );
nor U101944 ( n17231, n73406, n76159 );
xnor U101945 ( n24651, n25371, n25429 );
xor U101946 ( n25429, n75038, n76522 );
xnor U101947 ( n57787, n58508, n58566 );
xor U101948 ( n58566, n75040, n76264 );
xnor U101949 ( n66488, n67376, n67434 );
xor U101950 ( n67434, n75039, n76198 );
nor U101951 ( n25396, n25398, n76905 );
nor U101952 ( n25398, n25399, n25400 );
nand U101953 ( n25400, n25401, n25402 );
nand U101954 ( n25399, n25403, n25404 );
nor U101955 ( n58533, n58535, n76879 );
nor U101956 ( n58535, n58536, n58537 );
nand U101957 ( n58537, n58538, n58539 );
nand U101958 ( n58536, n58540, n58541 );
nor U101959 ( n67401, n67403, n76870 );
nor U101960 ( n67403, n67404, n67405 );
nand U101961 ( n67405, n67406, n67407 );
nand U101962 ( n67404, n67408, n67409 );
nor U101963 ( n64382, n40727, n41119 );
buf U101964 ( n76789, n76787 );
nand U101965 ( n41689, n41701, n41702 );
nand U101966 ( n41701, n76010, n40864 );
nand U101967 ( n41702, n76380, n40697 );
nor U101968 ( n71454, n73049, n71287 );
nor U101969 ( n47630, n47631, n47632 );
nor U101970 ( n47631, n73656, n47370 );
nor U101971 ( n47632, n73645, n47369 );
nor U101972 ( n68647, n73749, n68391 );
nor U101973 ( n26646, n73750, n26390 );
nor U101974 ( n59788, n73751, n59529 );
nand U101975 ( n68643, n68644, n68645 );
nor U101976 ( n68644, n68648, n68649 );
nor U101977 ( n68645, n68646, n68647 );
nor U101978 ( n68648, n73773, n68396 );
nand U101979 ( n26642, n26643, n26644 );
nor U101980 ( n26643, n26647, n26648 );
nor U101981 ( n26644, n26645, n26646 );
nor U101982 ( n26647, n73774, n26395 );
nand U101983 ( n59784, n59785, n59786 );
nor U101984 ( n59785, n59789, n59790 );
nor U101985 ( n59786, n59787, n59788 );
nor U101986 ( n59789, n73775, n59534 );
nor U101987 ( n68646, n73761, n68392 );
nor U101988 ( n26645, n73763, n26391 );
nor U101989 ( n59787, n73764, n59530 );
nor U101990 ( n72692, n72696, n72697 );
nor U101991 ( n72693, n72694, n72695 );
nor U101992 ( n72697, n73501, n73026 );
nor U101993 ( n47629, n47633, n47634 );
nor U101994 ( n47633, n73663, n47374 );
nor U101995 ( n47634, n73649, n47373 );
nor U101996 ( n68649, n73755, n68395 );
nor U101997 ( n26648, n73756, n26394 );
nor U101998 ( n59790, n73757, n59533 );
nor U101999 ( n46429, n46433, n7493 );
and U102000 ( n46433, n45627, n46434 );
nor U102001 ( n46419, n46421, n76330 );
nor U102002 ( n46421, n46422, n46423 );
nand U102003 ( n46422, n46442, n46443 );
nand U102004 ( n46423, n46424, n46425 );
and U102005 ( n45623, n46454, n46455 );
xor U102006 ( n46455, n74974, n76341 );
nor U102007 ( n46454, n45630, n46456 );
nor U102008 ( n46456, n7533, n74930 );
nor U102009 ( n67493, n67497, n5707 );
and U102010 ( n67497, n66552, n67498 );
nor U102011 ( n25488, n25492, n3949 );
and U102012 ( n25492, n24717, n25493 );
nor U102013 ( n58625, n58629, n6582 );
and U102014 ( n58629, n57851, n58630 );
nor U102015 ( n67483, n67485, n76870 );
nor U102016 ( n67485, n67486, n67487 );
nand U102017 ( n67486, n67506, n67507 );
nand U102018 ( n67487, n67488, n67489 );
nor U102019 ( n25478, n25480, n76905 );
nor U102020 ( n25480, n25481, n25482 );
nand U102021 ( n25481, n25501, n25502 );
nand U102022 ( n25482, n25483, n25484 );
nor U102023 ( n58615, n58617, n76879 );
nor U102024 ( n58617, n58618, n58619 );
nand U102025 ( n58618, n58638, n58639 );
nand U102026 ( n58619, n58620, n58621 );
and U102027 ( n66548, n67517, n67518 );
xor U102028 ( n67518, n74976, n76197 );
nor U102029 ( n67517, n66554, n67519 );
nor U102030 ( n67519, n5747, n74962 );
and U102031 ( n24713, n25512, n25513 );
xor U102032 ( n25513, n74975, n76521 );
nor U102033 ( n25512, n24719, n25514 );
nor U102034 ( n25514, n3989, n74960 );
and U102035 ( n57847, n58649, n58650 );
xor U102036 ( n58650, n74977, n76263 );
nor U102037 ( n58649, n57853, n58651 );
nor U102038 ( n58651, n6622, n74963 );
nor U102039 ( n37233, n36537, n76801 );
buf U102040 ( n76788, n76787 );
not U102041 ( n7812, n44511 );
nor U102042 ( n51370, n49982, n73419 );
nand U102043 ( n36462, n40091, n40092 );
nor U102044 ( n40092, n40093, n40094 );
nor U102045 ( n40091, n40096, n40097 );
nor U102046 ( n40094, n76412, n74314 );
not U102047 ( n800, n40732 );
nand U102048 ( n71295, n71259, n71246 );
nor U102049 ( n72694, n73498, n71105 );
nand U102050 ( n46443, n46444, n74974 );
nand U102051 ( n46444, n46445, n7503 );
not U102052 ( n7503, n46403 );
nor U102053 ( n46445, n46451, n46452 );
nor U102054 ( n18427, n16861, n73015 );
and U102055 ( n41690, n41703, n41704 );
nand U102056 ( n41704, n40864, n76378 );
nand U102057 ( n41703, n76010, n40697 );
nand U102058 ( n67507, n67508, n74976 );
nand U102059 ( n67508, n67509, n5717 );
not U102060 ( n5717, n67467 );
nor U102061 ( n67509, n67515, n67516 );
nand U102062 ( n25502, n25503, n74975 );
nand U102063 ( n25503, n25504, n3959 );
not U102064 ( n3959, n25462 );
nor U102065 ( n25504, n25510, n25511 );
nand U102066 ( n58639, n58640, n74977 );
nand U102067 ( n58640, n58641, n6592 );
not U102068 ( n6592, n58599 );
nor U102069 ( n58641, n58647, n58648 );
nand U102070 ( n44509, n47864, n73512 );
nor U102071 ( n72696, n73499, n71108 );
nor U102072 ( n68651, n68652, n68653 );
nor U102073 ( n68652, n73785, n68402 );
nor U102074 ( n68653, n73762, n68401 );
nor U102075 ( n26650, n26651, n26652 );
nor U102076 ( n26651, n73786, n26401 );
nor U102077 ( n26652, n73765, n26400 );
nor U102078 ( n59792, n59793, n59794 );
nor U102079 ( n59793, n73787, n59540 );
nor U102080 ( n59794, n73766, n59539 );
nand U102081 ( n48455, n48456, n48457 );
nand U102082 ( n48457, n569, n41183 );
nand U102083 ( n48456, n76857, n48458 );
nor U102084 ( n68650, n68654, n68655 );
nor U102085 ( n68654, n73791, n68406 );
nor U102086 ( n68655, n73776, n68405 );
nor U102087 ( n26649, n26653, n26654 );
nor U102088 ( n26653, n73792, n26405 );
nor U102089 ( n26654, n73777, n26404 );
nor U102090 ( n59791, n59795, n59796 );
nor U102091 ( n59795, n73793, n59544 );
nor U102092 ( n59796, n73778, n59543 );
nand U102093 ( n41542, n689, n41119 );
xnor U102094 ( n36759, n37056, n2040 );
nand U102095 ( n37056, n37057, n37058 );
nand U102096 ( n37057, n76829, n36532 );
nand U102097 ( n37058, n36767, n2035 );
and U102098 ( n36527, n37064, n37065 );
nand U102099 ( n37065, n76807, n36730 );
nand U102100 ( n37064, n76829, n36537 );
nand U102101 ( n72596, n72453, n71243 );
nand U102102 ( n36728, n37062, n37063 );
nand U102103 ( n37063, n76807, n36322 );
nand U102104 ( n37062, n76829, n36735 );
not U102105 ( n6024, n65386 );
not U102106 ( n4247, n23840 );
not U102107 ( n6879, n56964 );
nand U102108 ( n71013, n3632, n71012 );
nor U102109 ( n18803, n16966, n76788 );
nand U102110 ( n65384, n68884, n73518 );
nand U102111 ( n23838, n26885, n73520 );
nand U102112 ( n56962, n60025, n73521 );
xnor U102113 ( n36351, n37047, n2040 );
nand U102114 ( n37047, n37048, n37049 );
nand U102115 ( n37048, n76829, n36762 );
nand U102116 ( n37049, n36360, n2035 );
nor U102117 ( n51194, n49982, n73017 );
nand U102118 ( n41144, n41421, n41422 );
nand U102119 ( n41422, n76847, n40930 );
nand U102120 ( n41421, n76846, n41150 );
nor U102121 ( n50711, n49816, n73410 );
nor U102122 ( n19577, n75919, n76160 );
buf U102123 ( n76160, n17016 );
nand U102124 ( n72615, n72499, n71243 );
nand U102125 ( n71009, n72831, n71012 );
nor U102126 ( n45374, n43975, n45391 );
nor U102127 ( n44736, n43975, n44561 );
nor U102128 ( n40093, n38495, n76405 );
nor U102129 ( n47562, n73806, n47381 );
nand U102130 ( n47558, n47559, n47560 );
nor U102131 ( n47559, n47563, n47564 );
nor U102132 ( n47560, n47561, n47562 );
nor U102133 ( n47563, n73815, n47386 );
nor U102134 ( n47568, n73812, n47391 );
nand U102135 ( n47557, n47565, n47566 );
nor U102136 ( n47565, n47569, n47570 );
nor U102137 ( n47566, n47567, n47568 );
nor U102138 ( n47569, n73820, n47396 );
nand U102139 ( n41683, n41802, n41803 );
nand U102140 ( n41803, n41145, n76379 );
nand U102141 ( n41802, n76011, n40765 );
nor U102142 ( n47561, n73811, n47382 );
nor U102143 ( n47567, n73818, n47392 );
nor U102144 ( n50441, n49816, n73003 );
nor U102145 ( n42099, n40972, n707 );
nor U102146 ( n47564, n73808, n47385 );
nor U102147 ( n47570, n73816, n47395 );
nand U102148 ( n42042, n700, n41323 );
nor U102149 ( n43972, n43975, n43799 );
nand U102150 ( n41596, n707, n40972 );
buf U102151 ( n76834, n76833 );
nand U102152 ( n40864, n66181, n66182 );
nor U102153 ( n66182, n66183, n66184 );
nor U102154 ( n66181, n66186, n66187 );
nor U102155 ( n66184, n76246, n74336 );
nor U102156 ( n66186, n76248, n74337 );
nor U102157 ( n47548, n73805, n47359 );
nand U102158 ( n47544, n47545, n47546 );
nor U102159 ( n47545, n47549, n47550 );
nor U102160 ( n47546, n47547, n47548 );
nor U102161 ( n47549, n73813, n47364 );
nor U102162 ( n47547, n73809, n47360 );
nor U102163 ( n47550, n73807, n47363 );
nand U102164 ( n41682, n41791, n41792 );
nand U102165 ( n41791, n76011, n41145 );
nand U102166 ( n41792, n40765, n76379 );
nand U102167 ( n36762, n39966, n39967 );
nor U102168 ( n39967, n39968, n39969 );
nor U102169 ( n39966, n39971, n39972 );
nor U102170 ( n39969, n76411, n74356 );
nor U102171 ( n68583, n73834, n68413 );
nor U102172 ( n26582, n73835, n26412 );
nor U102173 ( n59724, n73836, n59551 );
nand U102174 ( n68579, n68580, n68581 );
nor U102175 ( n68580, n68584, n68585 );
nor U102176 ( n68581, n68582, n68583 );
nor U102177 ( n68584, n73861, n68418 );
nand U102178 ( n26578, n26579, n26580 );
nor U102179 ( n26579, n26583, n26584 );
nor U102180 ( n26580, n26581, n26582 );
nor U102181 ( n26583, n73862, n26417 );
nand U102182 ( n59720, n59721, n59722 );
nor U102183 ( n59721, n59725, n59726 );
nor U102184 ( n59722, n59723, n59724 );
nor U102185 ( n59725, n73863, n59556 );
nor U102186 ( n68589, n73850, n68423 );
nor U102187 ( n26588, n73853, n26422 );
nor U102188 ( n59730, n73854, n59561 );
nand U102189 ( n68578, n68586, n68587 );
nor U102190 ( n68586, n68590, n68591 );
nor U102191 ( n68587, n68588, n68589 );
nor U102192 ( n68590, n73877, n68428 );
nand U102193 ( n26577, n26585, n26586 );
nor U102194 ( n26585, n26589, n26590 );
nor U102195 ( n26586, n26587, n26588 );
nor U102196 ( n26589, n73878, n26427 );
nand U102197 ( n59719, n59727, n59728 );
nor U102198 ( n59727, n59731, n59732 );
nor U102199 ( n59728, n59729, n59730 );
nor U102200 ( n59731, n73879, n59566 );
nor U102201 ( n68582, n73849, n68414 );
nor U102202 ( n26581, n73851, n26413 );
nor U102203 ( n59723, n73852, n59552 );
nor U102204 ( n68588, n73871, n68424 );
nor U102205 ( n26587, n73872, n26423 );
nor U102206 ( n59729, n73873, n59562 );
nor U102207 ( n68585, n73840, n68417 );
nor U102208 ( n26584, n73841, n26416 );
nor U102209 ( n59726, n73842, n59555 );
nor U102210 ( n68591, n73864, n68427 );
nor U102211 ( n26590, n73865, n26426 );
nor U102212 ( n59732, n73866, n59565 );
nand U102213 ( n41785, n41796, n41797 );
nand U102214 ( n41796, n76011, n40930 );
nand U102215 ( n41797, n41150, n76379 );
nand U102216 ( n40759, n41336, n41337 );
nand U102217 ( n41337, n76848, n41145 );
nand U102218 ( n41336, n76844, n40765 );
not U102219 ( n1987, n36618 );
nor U102220 ( n45464, n50320, n76835 );
and U102221 ( n41788, n41800, n41801 );
nand U102222 ( n41800, n76011, n41114 );
nand U102223 ( n41801, n40935, n76379 );
nand U102224 ( n36355, n40000, n40001 );
nor U102225 ( n40001, n40002, n40003 );
nor U102226 ( n40000, n40005, n40006 );
nor U102227 ( n40003, n76411, n74360 );
nor U102228 ( n18590, n16861, n73418 );
nand U102229 ( n36761, n37054, n37055 );
nand U102230 ( n37055, n76807, n36532 );
nand U102231 ( n37054, n76829, n36767 );
nor U102232 ( n19260, n16861, n73420 );
nor U102233 ( n47552, n47553, n47554 );
nor U102234 ( n47553, n73817, n47370 );
nor U102235 ( n47554, n73810, n47369 );
nor U102236 ( n68569, n73830, n68391 );
nor U102237 ( n26568, n73831, n26390 );
nor U102238 ( n59710, n73832, n59529 );
nand U102239 ( n68565, n68566, n68567 );
nor U102240 ( n68566, n68570, n68571 );
nor U102241 ( n68567, n68568, n68569 );
nor U102242 ( n68570, n73855, n68396 );
nand U102243 ( n26564, n26565, n26566 );
nor U102244 ( n26565, n26569, n26570 );
nor U102245 ( n26566, n26567, n26568 );
nor U102246 ( n26569, n73856, n26395 );
nand U102247 ( n59706, n59707, n59708 );
nor U102248 ( n59707, n59711, n59712 );
nor U102249 ( n59708, n59709, n59710 );
nor U102250 ( n59711, n73857, n59534 );
nor U102251 ( n19428, n73022, n76161 );
nor U102252 ( n68568, n73843, n68392 );
nor U102253 ( n26567, n73845, n26391 );
nor U102254 ( n59709, n73846, n59530 );
nand U102255 ( n41789, n41798, n41799 );
nand U102256 ( n41799, n41114, n76379 );
nand U102257 ( n41798, n76011, n40935 );
nor U102258 ( n51706, n49816, n73425 );
nor U102259 ( n47551, n47555, n47556 );
nor U102260 ( n47555, n73819, n47374 );
nor U102261 ( n47556, n73814, n47373 );
nor U102262 ( n68571, n73837, n68395 );
nor U102263 ( n26570, n73838, n26394 );
nor U102264 ( n59712, n73839, n59533 );
nor U102265 ( n47470, n73880, n47381 );
nand U102266 ( n47466, n47467, n47468 );
nor U102267 ( n47467, n47471, n47472 );
nor U102268 ( n47468, n47469, n47470 );
nor U102269 ( n47471, n73889, n47386 );
nor U102270 ( n47476, n73886, n47391 );
nand U102271 ( n47465, n47473, n47474 );
nor U102272 ( n47473, n47477, n47478 );
nor U102273 ( n47474, n47475, n47476 );
nor U102274 ( n47477, n73894, n47396 );
nor U102275 ( n47469, n73885, n47382 );
nor U102276 ( n47475, n73892, n47392 );
nor U102277 ( n47472, n73882, n47385 );
nand U102278 ( n41782, n41794, n41795 );
nand U102279 ( n41795, n40930, n76379 );
nand U102280 ( n41794, n76011, n41150 );
nor U102281 ( n47478, n73890, n47395 );
nand U102282 ( n41535, n695, n40732 );
nor U102283 ( n19844, n16861, n73020 );
nand U102284 ( n36667, n40045, n40046 );
nor U102285 ( n40046, n40047, n40048 );
nor U102286 ( n40045, n40050, n40051 );
nor U102287 ( n40048, n76411, n74371 );
nor U102288 ( n40050, n76414, n74372 );
nor U102289 ( n66183, n54632, n76243 );
nor U102290 ( n52365, n73421, n49982 );
nor U102291 ( n47456, n73867, n47359 );
nand U102292 ( n47452, n47453, n47454 );
nor U102293 ( n47453, n47457, n47458 );
nor U102294 ( n47454, n47455, n47456 );
nor U102295 ( n47457, n73887, n47364 );
nor U102296 ( n37229, n36735, n76801 );
nor U102297 ( n47455, n73883, n47360 );
nor U102298 ( n68573, n68574, n68575 );
nor U102299 ( n68574, n73868, n68402 );
nor U102300 ( n68575, n73844, n68401 );
nor U102301 ( n26572, n26573, n26574 );
nor U102302 ( n26573, n73869, n26401 );
nor U102303 ( n26574, n73847, n26400 );
nor U102304 ( n59714, n59715, n59716 );
nor U102305 ( n59715, n73870, n59540 );
nor U102306 ( n59716, n73848, n59539 );
nor U102307 ( n65807, n76248, n74379 );
nand U102308 ( n40930, n65802, n65803 );
nor U102309 ( n65803, n65804, n65805 );
nor U102310 ( n65802, n65807, n65808 );
nor U102311 ( n65805, n76245, n74378 );
nor U102312 ( n47458, n73881, n47363 );
nor U102313 ( n68572, n68576, n68577 );
nor U102314 ( n68576, n73874, n68406 );
nor U102315 ( n68577, n73858, n68405 );
nor U102316 ( n26571, n26575, n26576 );
nor U102317 ( n26575, n73875, n26405 );
nor U102318 ( n26576, n73859, n26404 );
nor U102319 ( n59713, n59717, n59718 );
nor U102320 ( n59717, n73876, n59544 );
nor U102321 ( n59718, n73860, n59543 );
nand U102322 ( n37776, n2042, n37102 );
nor U102323 ( n16849, n16861, n75911 );
nor U102324 ( n68491, n73901, n68413 );
nor U102325 ( n26490, n73902, n26412 );
nor U102326 ( n59629, n73903, n59551 );
nand U102327 ( n68487, n68488, n68489 );
nor U102328 ( n68488, n68492, n68493 );
nor U102329 ( n68489, n68490, n68491 );
nor U102330 ( n68492, n73930, n68418 );
nand U102331 ( n26486, n26487, n26488 );
nor U102332 ( n26487, n26491, n26492 );
nor U102333 ( n26488, n26489, n26490 );
nor U102334 ( n26491, n73931, n26417 );
nand U102335 ( n59625, n59626, n59627 );
nor U102336 ( n59626, n59630, n59631 );
nor U102337 ( n59627, n59628, n59629 );
nor U102338 ( n59630, n73932, n59556 );
nor U102339 ( n68497, n73919, n68423 );
nor U102340 ( n26496, n73922, n26422 );
nor U102341 ( n59635, n73923, n59561 );
nand U102342 ( n68486, n68494, n68495 );
nor U102343 ( n68494, n68498, n68499 );
nor U102344 ( n68495, n68496, n68497 );
nor U102345 ( n68498, n73945, n68428 );
nand U102346 ( n26485, n26493, n26494 );
nor U102347 ( n26493, n26497, n26498 );
nor U102348 ( n26494, n26495, n26496 );
nor U102349 ( n26497, n73946, n26427 );
nand U102350 ( n59624, n59632, n59633 );
nor U102351 ( n59632, n59636, n59637 );
nor U102352 ( n59633, n59634, n59635 );
nor U102353 ( n59636, n73947, n59566 );
nor U102354 ( n68490, n73918, n68414 );
nor U102355 ( n26489, n73920, n26413 );
nor U102356 ( n59628, n73921, n59552 );
nor U102357 ( n68496, n73939, n68424 );
nor U102358 ( n26495, n73940, n26423 );
nor U102359 ( n59634, n73941, n59562 );
nor U102360 ( n68493, n73907, n68417 );
nor U102361 ( n26492, n73908, n26416 );
nor U102362 ( n59631, n73909, n59555 );
nor U102363 ( n68499, n73933, n68427 );
nor U102364 ( n26498, n73934, n26426 );
nor U102365 ( n59637, n73935, n59565 );
nand U102366 ( n37453, n2175, n36577 );
nor U102367 ( n17499, n75911, n76158 );
nand U102368 ( n48572, n48573, n48574 );
nand U102369 ( n48574, n569, n41011 );
nand U102370 ( n48573, n76857, n48575 );
nor U102371 ( n40002, n38456, n76405 );
nand U102372 ( n41145, n65926, n65927 );
nor U102373 ( n65927, n65928, n65929 );
nor U102374 ( n65926, n65931, n65932 );
nor U102375 ( n65929, n76245, n74381 );
nor U102376 ( n65931, n76248, n74380 );
nand U102377 ( n42291, n845, n41471 );
not U102378 ( n1982, n36577 );
and U102379 ( n39485, n39493, n39494 );
nand U102380 ( n39493, n36618, n36797 );
nand U102381 ( n39494, n39495, n39492 );
nand U102382 ( n45550, n45561, n45562 );
nand U102383 ( n45561, n45537, n74931 );
nand U102384 ( n45562, n76662, n45563 );
nand U102385 ( n15841, n45548, n45549 );
nor U102386 ( n45548, n45570, n45571 );
nor U102387 ( n45549, n45550, n45551 );
nor U102388 ( n45570, n75237, n76669 );
nand U102389 ( n24638, n24649, n24650 );
nand U102390 ( n24649, n24624, n75186 );
nand U102391 ( n24650, n76758, n24651 );
nand U102392 ( n57774, n57785, n57786 );
nand U102393 ( n57785, n57756, n75187 );
nand U102394 ( n57786, n76691, n57787 );
nand U102395 ( n66475, n66486, n66487 );
nand U102396 ( n66486, n66461, n75188 );
nand U102397 ( n66487, n76710, n66488 );
nand U102398 ( n6861, n24636, n24637 );
nor U102399 ( n24636, n24658, n24659 );
nor U102400 ( n24637, n24638, n24639 );
nor U102401 ( n24658, n75064, n76765 );
nand U102402 ( n13596, n57772, n57773 );
nor U102403 ( n57772, n57794, n57795 );
nor U102404 ( n57773, n57774, n57775 );
nor U102405 ( n57794, n75063, n76698 );
nand U102406 ( n11351, n66473, n66474 );
nor U102407 ( n66473, n66495, n66496 );
nor U102408 ( n66474, n66475, n66476 );
nor U102409 ( n66495, n75070, n76717 );
nor U102410 ( n49787, n49982, n73003 );
nor U102411 ( n47460, n47461, n47462 );
nor U102412 ( n47461, n73891, n47370 );
nor U102413 ( n47462, n73884, n47369 );
nor U102414 ( n68477, n73898, n68391 );
nor U102415 ( n26476, n73899, n26390 );
nor U102416 ( n59615, n73900, n59529 );
nand U102417 ( n68473, n68474, n68475 );
nor U102418 ( n68474, n68478, n68479 );
nor U102419 ( n68475, n68476, n68477 );
nor U102420 ( n68478, n73924, n68396 );
nand U102421 ( n26472, n26473, n26474 );
nor U102422 ( n26473, n26477, n26478 );
nor U102423 ( n26474, n26475, n26476 );
nor U102424 ( n26477, n73925, n26395 );
nand U102425 ( n59611, n59612, n59613 );
nor U102426 ( n59612, n59616, n59617 );
nor U102427 ( n59613, n59614, n59615 );
nor U102428 ( n59616, n73926, n59534 );
nor U102429 ( n68476, n73912, n68392 );
nor U102430 ( n26475, n73914, n26391 );
nor U102431 ( n59614, n73915, n59530 );
nor U102432 ( n47459, n47463, n47464 );
nor U102433 ( n47463, n73893, n47374 );
nor U102434 ( n47464, n73888, n47373 );
nor U102435 ( n68479, n73904, n68395 );
nor U102436 ( n26478, n73905, n26394 );
nor U102437 ( n59617, n73906, n59533 );
nand U102438 ( n38288, n38289, n38290 );
nand U102439 ( n38289, n76815, n36403 );
nand U102440 ( n38290, n38291, n76442 );
nand U102441 ( n72426, n71308, n71243 );
nand U102442 ( n39666, n36327, n36961 );
and U102443 ( n72151, n71143, n71243 );
nand U102444 ( n71872, n71327, n71245 );
nor U102445 ( n19208, n73423, n76160 );
nor U102446 ( n65804, n49259, n76242 );
nor U102447 ( n46376, n46378, n76330 );
nor U102448 ( n46378, n46379, n46380 );
nand U102449 ( n46379, n46399, n46400 );
nand U102450 ( n46380, n46381, n46382 );
nand U102451 ( n46381, n76659, n45605 );
nor U102452 ( n52362, n49982, n73021 );
nor U102453 ( n67440, n67442, n76870 );
nor U102454 ( n67442, n67443, n67444 );
nand U102455 ( n67443, n67463, n67464 );
nand U102456 ( n67444, n67445, n67446 );
nor U102457 ( n25435, n25437, n76905 );
nor U102458 ( n25437, n25438, n25439 );
nand U102459 ( n25438, n25458, n25459 );
nand U102460 ( n25439, n25440, n25441 );
nor U102461 ( n58572, n58574, n76879 );
nor U102462 ( n58574, n58575, n58576 );
nand U102463 ( n58575, n58595, n58596 );
nand U102464 ( n58576, n58577, n58578 );
nand U102465 ( n67445, n76705, n66530 );
nand U102466 ( n25440, n76751, n24695 );
nand U102467 ( n58577, n76684, n57829 );
nor U102468 ( n50967, n49982, n73413 );
nand U102469 ( n36354, n36968, n36969 );
nand U102470 ( n36969, n76807, n36762 );
nand U102471 ( n36968, n76827, n36360 );
nor U102472 ( n45370, n44020, n45391 );
nor U102473 ( n44776, n44020, n44561 );
nand U102474 ( n16216, n44767, n44768 );
nor U102475 ( n44768, n44769, n44770 );
nor U102476 ( n44767, n44775, n44776 );
nor U102477 ( n44769, n43808, n44772 );
nand U102478 ( n48325, n48326, n48327 );
nand U102479 ( n48326, n569, n40806 );
nand U102480 ( n48327, n48328, n45754 );
nor U102481 ( n68481, n68482, n68483 );
nor U102482 ( n68482, n73936, n68402 );
nor U102483 ( n68483, n73913, n68401 );
nor U102484 ( n26480, n26481, n26482 );
nor U102485 ( n26481, n73937, n26401 );
nor U102486 ( n26482, n73916, n26400 );
nor U102487 ( n59619, n59620, n59621 );
nor U102488 ( n59620, n73938, n59540 );
nor U102489 ( n59621, n73917, n59539 );
nor U102490 ( n68480, n68484, n68485 );
nor U102491 ( n68484, n73942, n68406 );
nor U102492 ( n68485, n73927, n68405 );
nor U102493 ( n26479, n26483, n26484 );
nor U102494 ( n26483, n73943, n26405 );
nor U102495 ( n26484, n73928, n26404 );
nor U102496 ( n59618, n59622, n59623 );
nor U102497 ( n59622, n73944, n59544 );
nor U102498 ( n59623, n73929, n59543 );
nor U102499 ( n44017, n44020, n43799 );
nor U102500 ( n37221, n36327, n76801 );
and U102501 ( n72263, n71371, n71243 );
nor U102502 ( n11567, n10059, n11594 );
nor U102503 ( n11004, n10059, n10785 );
nand U102504 ( n72360, n71312, n71243 );
nand U102505 ( n46424, n46440, n46441 );
nand U102506 ( n67488, n67504, n67505 );
nand U102507 ( n25483, n25499, n25500 );
nand U102508 ( n58620, n58636, n58637 );
nor U102509 ( n47380, n73966, n47381 );
nand U102510 ( n47376, n47377, n47378 );
nor U102511 ( n47377, n47383, n47384 );
nor U102512 ( n47378, n47379, n47380 );
nor U102513 ( n47383, n73976, n47386 );
nor U102514 ( n10056, n10059, n9897 );
nor U102515 ( n47390, n73973, n47391 );
nand U102516 ( n47375, n47387, n47388 );
nor U102517 ( n47387, n47393, n47394 );
nor U102518 ( n47388, n47389, n47390 );
nor U102519 ( n47393, n73996, n47396 );
nor U102520 ( n47379, n73972, n47382 );
nor U102521 ( n47389, n73993, n47392 );
nor U102522 ( n47384, n73968, n47385 );
nor U102523 ( n47394, n73977, n47395 );
nand U102524 ( n41496, n41497, n41498 );
or U102525 ( n41497, n41599, n41466 );
nand U102526 ( n41498, n41499, n41500 );
nor U102527 ( n41499, n41598, n40664 );
nand U102528 ( n48800, n48801, n48802 );
nand U102529 ( n48802, n569, n41323 );
nand U102530 ( n48801, n76857, n48803 );
nand U102531 ( n41054, n66092, n66093 );
nor U102532 ( n66093, n66094, n66095 );
nor U102533 ( n66092, n66097, n66098 );
nor U102534 ( n66095, n76245, n74382 );
nor U102535 ( n18258, n16861, n73414 );
nor U102536 ( n47358, n73950, n47359 );
nand U102537 ( n47354, n47355, n47356 );
nor U102538 ( n47355, n47361, n47362 );
nor U102539 ( n47356, n47357, n47358 );
nor U102540 ( n47361, n73974, n47364 );
nor U102541 ( n47357, n73970, n47360 );
not U102542 ( n804, n41011 );
nor U102543 ( n47362, n73967, n47363 );
nor U102544 ( n68412, n74049, n68413 );
nor U102545 ( n26411, n74051, n26412 );
nor U102546 ( n59550, n74050, n59551 );
nand U102547 ( n68408, n68409, n68410 );
nor U102548 ( n68409, n68415, n68416 );
nor U102549 ( n68410, n68411, n68412 );
nor U102550 ( n68415, n74090, n68418 );
nand U102551 ( n26407, n26408, n26409 );
nor U102552 ( n26408, n26414, n26415 );
nor U102553 ( n26409, n26410, n26411 );
nor U102554 ( n26414, n74092, n26417 );
nand U102555 ( n59546, n59547, n59548 );
nor U102556 ( n59547, n59553, n59554 );
nor U102557 ( n59548, n59549, n59550 );
nor U102558 ( n59553, n74091, n59556 );
nand U102559 ( n32780, n32860, n32861 );
nor U102560 ( n32860, n32862, n32863 );
nor U102561 ( n32863, n76021, n74671 );
nor U102562 ( n32862, n32864, n32865 );
not U102563 ( n3397, n31169 );
nand U102564 ( n30016, n34259, n34260 );
or U102565 ( n34260, n73524, n30782 );
nor U102566 ( n31951, n32739, n76021 );
nor U102567 ( n32229, n33165, n76022 );
nand U102568 ( n33299, n33371, n33370 );
nor U102569 ( n34035, n73953, n33657 );
nor U102570 ( n32601, n31847, n32604 );
nor U102571 ( n33297, n33299, n33300 );
nand U102572 ( n33300, n33301, n33302 );
nor U102573 ( n4461, n32590, n32591 );
nor U102574 ( n32591, n32592, n32593 );
nor U102575 ( n32590, n32594, n32595 );
nand U102576 ( n32594, n32621, n32622 );
nand U102577 ( n32865, n32866, n32867 );
nand U102578 ( n32866, n76022, n74671 );
nand U102579 ( n34031, n34032, n34033 );
nor U102580 ( n34032, n34036, n34037 );
nor U102581 ( n34033, n34034, n34035 );
nor U102582 ( n34036, n73963, n33662 );
nand U102583 ( n32595, n32596, n214 );
not U102584 ( n214, n32593 );
nor U102585 ( n32596, n32601, n32602 );
and U102586 ( n32602, n31849, n76774 );
nand U102587 ( n33245, n33293, n33294 );
nor U102588 ( n33294, n3159, n33295 );
nor U102589 ( n33293, n33297, n33298 );
not U102590 ( n3159, n33296 );
nor U102591 ( n68422, n74074, n68423 );
nor U102592 ( n26421, n74078, n26422 );
nor U102593 ( n59560, n74077, n59561 );
nand U102594 ( n68407, n68419, n68420 );
nor U102595 ( n68419, n68425, n68426 );
nor U102596 ( n68420, n68421, n68422 );
nor U102597 ( n68425, n74118, n68428 );
nand U102598 ( n26406, n26418, n26419 );
nor U102599 ( n26418, n26424, n26425 );
nor U102600 ( n26419, n26420, n26421 );
nor U102601 ( n26424, n74120, n26427 );
nand U102602 ( n59545, n59557, n59558 );
nor U102603 ( n59557, n59563, n59564 );
nor U102604 ( n59558, n59559, n59560 );
nor U102605 ( n59563, n74119, n59566 );
nand U102606 ( n71754, n71245, n71096 );
nor U102607 ( n68411, n74073, n68414 );
nor U102608 ( n26410, n74076, n26413 );
nor U102609 ( n59549, n74075, n59552 );
nor U102610 ( n34041, n73956, n33667 );
nand U102611 ( n34030, n34038, n34039 );
nor U102612 ( n34038, n34042, n34043 );
nor U102613 ( n34039, n34040, n34041 );
nor U102614 ( n34042, n73965, n33672 );
nor U102615 ( n34034, n73958, n33658 );
nor U102616 ( n68421, n74112, n68424 );
nor U102617 ( n26420, n74114, n26423 );
nor U102618 ( n59559, n74113, n59562 );
nor U102619 ( n34040, n73960, n33668 );
nor U102620 ( n68416, n74056, n68417 );
nor U102621 ( n26415, n74058, n26416 );
nor U102622 ( n59554, n74057, n59555 );
nor U102623 ( n34037, n73969, n33661 );
nor U102624 ( n68426, n74094, n68427 );
nor U102625 ( n26425, n74096, n26426 );
nor U102626 ( n59564, n74095, n59565 );
nor U102627 ( n34043, n73962, n33671 );
nand U102628 ( n38383, n38384, n38385 );
nand U102629 ( n38385, n76816, n36327 );
nand U102630 ( n38384, n76812, n38386 );
nand U102631 ( n41593, n714, n41011 );
and U102632 ( n41862, n41632, n41897 );
nand U102633 ( n41897, n41510, n76380 );
not U102634 ( n3403, n31509 );
nand U102635 ( n41863, n41635, n41898 );
nand U102636 ( n41898, n76383, n41510 );
nand U102637 ( n71466, n71243, n71303 );
nand U102638 ( n39609, n36955, n36572 );
not U102639 ( n3150, n31949 );
nor U102640 ( n66011, n76248, n74386 );
nand U102641 ( n40760, n66006, n66007 );
nor U102642 ( n66007, n66008, n66009 );
nor U102643 ( n66006, n66011, n66012 );
nor U102644 ( n66009, n76245, n74384 );
not U102645 ( n3152, n32227 );
nor U102646 ( n18023, n73009, n76163 );
xnor U102647 ( n40723, n41436, n593 );
nand U102648 ( n41436, n41437, n41438 );
nand U102649 ( n41437, n76846, n41329 );
nand U102650 ( n41438, n40732, n41264 );
nor U102651 ( n47366, n47367, n47368 );
nor U102652 ( n47367, n73990, n47370 );
nor U102653 ( n47368, n73971, n47369 );
nor U102654 ( n68390, n74027, n68391 );
nor U102655 ( n26389, n74029, n26390 );
nor U102656 ( n59528, n74028, n59529 );
nand U102657 ( n68386, n68387, n68388 );
nor U102658 ( n68387, n68393, n68394 );
nor U102659 ( n68388, n68389, n68390 );
nor U102660 ( n68393, n74079, n68396 );
nand U102661 ( n26385, n26386, n26387 );
nor U102662 ( n26386, n26392, n26393 );
nor U102663 ( n26387, n26388, n26389 );
nor U102664 ( n26392, n74081, n26395 );
nand U102665 ( n59524, n59525, n59526 );
nor U102666 ( n59525, n59531, n59532 );
nor U102667 ( n59526, n59527, n59528 );
nor U102668 ( n59531, n74080, n59534 );
nor U102669 ( n34115, n30772, n35717 );
nor U102670 ( n35717, n73526, n3403 );
nor U102671 ( n34021, n73949, n33635 );
nand U102672 ( n34017, n34018, n34019 );
nor U102673 ( n34018, n34022, n34023 );
nor U102674 ( n34019, n34020, n34021 );
nor U102675 ( n34022, n73959, n33640 );
nor U102676 ( n68389, n74065, n68392 );
nor U102677 ( n26388, n74068, n26391 );
nor U102678 ( n59527, n74067, n59530 );
nor U102679 ( n34020, n73952, n33636 );
nor U102680 ( n47365, n47371, n47372 );
nor U102681 ( n47371, n73994, n47374 );
nor U102682 ( n47372, n73975, n47373 );
nor U102683 ( n68394, n74053, n68395 );
nor U102684 ( n26393, n74055, n26394 );
nor U102685 ( n59532, n74054, n59533 );
nor U102686 ( n34023, n73954, n33639 );
or U102687 ( n50843, n49982, n73412 );
nor U102688 ( n33982, n74023, n33657 );
nand U102689 ( n33978, n33979, n33980 );
nor U102690 ( n33979, n33983, n33984 );
nor U102691 ( n33980, n33981, n33982 );
nor U102692 ( n33983, n74044, n33662 );
nor U102693 ( n33988, n74030, n33667 );
nand U102694 ( n33977, n33985, n33986 );
nor U102695 ( n33985, n33989, n33990 );
nor U102696 ( n33986, n33987, n33988 );
nor U102697 ( n33989, n74047, n33672 );
nor U102698 ( n33981, n74033, n33658 );
nor U102699 ( n33984, n74048, n33661 );
nor U102700 ( n33987, n74036, n33668 );
nor U102701 ( n33990, n74042, n33671 );
not U102702 ( n1432, n51514 );
nand U102703 ( n45602, n45603, n45604 );
nand U102704 ( n45603, n7434, n7960 );
nand U102705 ( n45604, n76663, n45605 );
nand U102706 ( n15836, n45576, n45577 );
nor U102707 ( n45577, n45578, n45579 );
nor U102708 ( n45576, n45601, n45602 );
nand U102709 ( n45579, n45580, n45581 );
nand U102710 ( n66527, n66528, n66529 );
nand U102711 ( n66528, n5660, n6173 );
nand U102712 ( n66529, n76710, n66530 );
nand U102713 ( n24692, n24693, n24694 );
nand U102714 ( n24693, n3903, n4395 );
nand U102715 ( n24694, n76758, n24695 );
nand U102716 ( n57826, n57827, n57828 );
nand U102717 ( n57827, n6535, n7028 );
nand U102718 ( n57828, n76691, n57829 );
nand U102719 ( n11346, n66501, n66502 );
nor U102720 ( n66502, n66503, n66504 );
nor U102721 ( n66501, n66526, n66527 );
nand U102722 ( n66504, n66505, n66506 );
nand U102723 ( n6856, n24666, n24667 );
nor U102724 ( n24667, n24668, n24669 );
nor U102725 ( n24666, n24691, n24692 );
nand U102726 ( n24669, n24670, n24671 );
nand U102727 ( n13591, n57800, n57801 );
nor U102728 ( n57801, n57802, n57803 );
nor U102729 ( n57800, n57825, n57826 );
nand U102730 ( n57803, n57804, n57805 );
nor U102731 ( n68398, n68399, n68400 );
nor U102732 ( n68399, n74108, n68402 );
nor U102733 ( n68400, n74066, n68401 );
nor U102734 ( n26397, n26398, n26399 );
nor U102735 ( n26398, n74110, n26401 );
nor U102736 ( n26399, n74070, n26400 );
nor U102737 ( n59536, n59537, n59538 );
nor U102738 ( n59537, n74109, n59540 );
nor U102739 ( n59538, n74069, n59539 );
nor U102740 ( n34025, n34026, n34027 );
nor U102741 ( n34026, n73955, n33646 );
nor U102742 ( n34027, n73951, n33645 );
nand U102743 ( n42028, n42029, n42030 );
nand U102744 ( n42029, n42060, n41510 );
nand U102745 ( n42030, n42031, n749 );
nand U102746 ( n42060, n41507, n76385 );
and U102747 ( n71993, n71357, n71243 );
nor U102748 ( n68397, n68403, n68404 );
nor U102749 ( n68403, n74115, n68406 );
nor U102750 ( n68404, n74083, n68405 );
nor U102751 ( n26396, n26402, n26403 );
nor U102752 ( n26402, n74117, n26405 );
nor U102753 ( n26403, n74087, n26404 );
nor U102754 ( n59535, n59541, n59542 );
nor U102755 ( n59541, n74116, n59544 );
nor U102756 ( n59542, n74086, n59543 );
nor U102757 ( n34024, n34028, n34029 );
nor U102758 ( n34028, n73961, n33650 );
nor U102759 ( n34029, n73957, n33649 );
nor U102760 ( n30782, n31509, n73526 );
nor U102761 ( n47821, n74133, n47381 );
nand U102762 ( n47817, n47818, n47819 );
nor U102763 ( n47818, n47822, n47823 );
nor U102764 ( n47819, n47820, n47821 );
nor U102765 ( n47822, n74147, n47386 );
nor U102766 ( n47827, n74145, n47391 );
nand U102767 ( n47816, n47824, n47825 );
nor U102768 ( n47824, n47828, n47829 );
nor U102769 ( n47825, n47826, n47827 );
nor U102770 ( n47828, n74160, n47396 );
nor U102771 ( n47820, n74144, n47382 );
nor U102772 ( n47826, n74158, n47392 );
nor U102773 ( n47823, n74132, n47385 );
nor U102774 ( n33968, n74012, n33635 );
nand U102775 ( n33964, n33965, n33966 );
nor U102776 ( n33965, n33969, n33970 );
nor U102777 ( n33966, n33967, n33968 );
nor U102778 ( n33969, n74034, n33640 );
nor U102779 ( n47829, n74148, n47395 );
nor U102780 ( n33967, n74022, n33636 );
nor U102781 ( n33970, n74024, n33639 );
not U102782 ( n802, n41323 );
nand U102783 ( n64230, n40732, n41329 );
nor U102784 ( n66008, n49568, n76243 );
xnor U102785 ( n36318, n37069, n2040 );
nand U102786 ( n37069, n37070, n37071 );
nand U102787 ( n37070, n76829, n36961 );
nand U102788 ( n37071, n36327, n2035 );
nor U102789 ( n47807, n74106, n47359 );
nand U102790 ( n47803, n47804, n47805 );
nor U102791 ( n47804, n47808, n47809 );
nor U102792 ( n47805, n47806, n47807 );
nor U102793 ( n47808, n74141, n47364 );
nand U102794 ( n31844, n31845, n31846 );
nand U102795 ( n31845, n76786, n31849 );
or U102796 ( n31846, n31847, n31848 );
nand U102797 ( n4621, n31824, n31825 );
nor U102798 ( n31825, n31826, n31827 );
nor U102799 ( n31824, n31843, n31844 );
nand U102800 ( n31826, n31835, n31836 );
nor U102801 ( n47806, n74135, n47360 );
nand U102802 ( n48917, n48918, n48919 );
nand U102803 ( n48919, n569, n40732 );
nand U102804 ( n48918, n76857, n48920 );
nor U102805 ( n47809, n74130, n47363 );
nand U102806 ( n71305, n71243, n71429 );
nand U102807 ( n71253, n1208, n71254 );
not U102808 ( n1208, n71260 );
nand U102809 ( n71254, n71255, n71256 );
nand U102810 ( n71255, n71258, n71259 );
nor U102811 ( n68841, n74174, n68413 );
nor U102812 ( n26842, n74175, n26412 );
nor U102813 ( n59982, n74176, n59551 );
nand U102814 ( n68837, n68838, n68839 );
nor U102815 ( n68838, n68842, n68843 );
nor U102816 ( n68839, n68840, n68841 );
nor U102817 ( n68842, n74199, n68418 );
nand U102818 ( n26838, n26839, n26840 );
nor U102819 ( n26839, n26843, n26844 );
nor U102820 ( n26840, n26841, n26842 );
nor U102821 ( n26843, n74200, n26417 );
nand U102822 ( n59978, n59979, n59980 );
nor U102823 ( n59979, n59983, n59984 );
nor U102824 ( n59980, n59981, n59982 );
nor U102825 ( n59983, n74201, n59556 );
nor U102826 ( n68847, n74192, n68423 );
nor U102827 ( n26848, n74193, n26422 );
nor U102828 ( n59988, n74194, n59561 );
nand U102829 ( n68836, n68844, n68845 );
nor U102830 ( n68844, n68848, n68849 );
nor U102831 ( n68845, n68846, n68847 );
nor U102832 ( n68848, n74214, n68428 );
nand U102833 ( n26837, n26845, n26846 );
nor U102834 ( n26845, n26849, n26850 );
nor U102835 ( n26846, n26847, n26848 );
nor U102836 ( n26849, n74215, n26427 );
nand U102837 ( n59977, n59985, n59986 );
nor U102838 ( n59985, n59989, n59990 );
nor U102839 ( n59986, n59987, n59988 );
nor U102840 ( n59989, n74216, n59566 );
nor U102841 ( n68840, n74189, n68414 );
nor U102842 ( n26841, n74190, n26413 );
nor U102843 ( n59981, n74191, n59552 );
nand U102844 ( n36532, n39923, n39924 );
nor U102845 ( n39924, n39925, n39926 );
nor U102846 ( n39923, n39928, n39929 );
nor U102847 ( n39926, n76411, n74393 );
nor U102848 ( n68846, n74208, n68424 );
nor U102849 ( n26847, n74209, n26423 );
nor U102850 ( n59987, n74210, n59562 );
nor U102851 ( n45622, n45623, n45624 );
nor U102852 ( n45624, n76341, n45626 );
nand U102853 ( n45626, n7917, n45627 );
nand U102854 ( n15831, n45607, n45608 );
nor U102855 ( n45607, n45633, n45634 );
nor U102856 ( n45608, n45609, n45610 );
nor U102857 ( n45633, n75302, n76669 );
nor U102858 ( n37217, n36955, n76802 );
nor U102859 ( n68843, n74177, n68417 );
nor U102860 ( n26844, n74178, n26416 );
nor U102861 ( n59984, n74179, n59555 );
nor U102862 ( n33972, n33973, n33974 );
nor U102863 ( n33973, n74025, n33646 );
nor U102864 ( n33974, n74021, n33645 );
nor U102865 ( n24712, n24713, n24714 );
nor U102866 ( n24714, n76521, n24716 );
nand U102867 ( n24716, n4352, n24717 );
nor U102868 ( n66547, n66548, n66549 );
nor U102869 ( n66549, n76197, n66551 );
nand U102870 ( n66551, n6129, n66552 );
nor U102871 ( n57846, n57847, n57848 );
nor U102872 ( n57848, n76263, n57850 );
nand U102873 ( n57850, n6984, n57851 );
nand U102874 ( n6851, n24697, n24698 );
nor U102875 ( n24697, n24722, n24723 );
nor U102876 ( n24698, n24699, n24700 );
nor U102877 ( n24722, n75301, n76765 );
nand U102878 ( n11341, n66532, n66533 );
nor U102879 ( n66532, n66557, n66558 );
nor U102880 ( n66533, n66534, n66535 );
nor U102881 ( n66557, n75361, n76717 );
nand U102882 ( n13586, n57831, n57832 );
nor U102883 ( n57831, n57856, n57857 );
nor U102884 ( n57832, n57833, n57834 );
nor U102885 ( n57856, n75300, n76698 );
nor U102886 ( n68849, n74202, n68427 );
nor U102887 ( n26850, n74203, n26426 );
nor U102888 ( n59990, n74204, n59565 );
nor U102889 ( n17765, n73404, n76161 );
nor U102890 ( n33971, n33975, n33976 );
nor U102891 ( n33975, n74040, n33650 );
nor U102892 ( n33976, n74032, n33649 );
xnor U102893 ( n41272, n41439, n593 );
nand U102894 ( n41439, n41440, n41441 );
nand U102895 ( n41440, n76846, n40967 );
nand U102896 ( n41441, n41323, n41264 );
nor U102897 ( n19693, n16861, n75919 );
not U102898 ( n1994, n36802 );
nor U102899 ( n47811, n47812, n47813 );
nor U102900 ( n47812, n74151, n47370 );
nor U102901 ( n47813, n74138, n47369 );
nor U102902 ( n68827, n74167, n68391 );
nor U102903 ( n26828, n74168, n26390 );
nor U102904 ( n59968, n74169, n59529 );
nand U102905 ( n68823, n68824, n68825 );
nor U102906 ( n68824, n68828, n68829 );
nor U102907 ( n68825, n68826, n68827 );
nor U102908 ( n68828, n74186, n68396 );
nand U102909 ( n26824, n26825, n26826 );
nor U102910 ( n26825, n26829, n26830 );
nor U102911 ( n26826, n26827, n26828 );
nor U102912 ( n26829, n74187, n26395 );
nand U102913 ( n59964, n59965, n59966 );
nor U102914 ( n59965, n59969, n59970 );
nor U102915 ( n59966, n59967, n59968 );
nor U102916 ( n59969, n74188, n59534 );
nand U102917 ( n37553, n2178, n36802 );
nand U102918 ( n38326, n38327, n38328 );
nand U102919 ( n38327, n76815, n36618 );
nand U102920 ( n38328, n1868, n76442 );
not U102921 ( n1868, n38329 );
nor U102922 ( n68826, n74180, n68392 );
nor U102923 ( n26827, n74182, n26391 );
nor U102924 ( n59967, n74183, n59530 );
nor U102925 ( n18135, n16861, n73012 );
nor U102926 ( n47810, n47814, n47815 );
nor U102927 ( n47814, n74159, n47374 );
nor U102928 ( n47815, n74146, n47373 );
nor U102929 ( n68829, n74171, n68395 );
nor U102930 ( n26830, n74172, n26394 );
nor U102931 ( n59970, n74173, n59533 );
nor U102932 ( n11562, n10115, n11594 );
nor U102933 ( n46966, n46969, n76341 );
nor U102934 ( n46969, n74417, n72948 );
nor U102935 ( n33905, n74102, n33657 );
nand U102936 ( n33901, n33902, n33903 );
nor U102937 ( n33902, n33906, n33907 );
nor U102938 ( n33903, n33904, n33905 );
nor U102939 ( n33906, n74129, n33662 );
nor U102940 ( n52184, n49982, n73426 );
nor U102941 ( n33907, n74107, n33661 );
nor U102942 ( n18768, n73422, n76164 );
xnor U102943 ( n40962, n41261, n593 );
nand U102944 ( n41261, n41262, n41263 );
nand U102945 ( n41262, n76844, n41006 );
nand U102946 ( n41263, n40972, n41264 );
nor U102947 ( n33911, n74125, n33667 );
nand U102948 ( n33900, n33908, n33909 );
nor U102949 ( n33908, n33912, n33913 );
nor U102950 ( n33909, n33910, n33911 );
nor U102951 ( n33912, n74142, n33672 );
nand U102952 ( n31504, n73059, n73532 );
nand U102953 ( n34130, n31504, n31509 );
not U102954 ( n3404, n31136 );
nor U102955 ( n33904, n74124, n33658 );
nor U102956 ( n33910, n74136, n33668 );
nor U102957 ( n11054, n10115, n10785 );
nand U102958 ( n9481, n11043, n11044 );
nor U102959 ( n11044, n11045, n11047 );
nor U102960 ( n11043, n11053, n11054 );
nor U102961 ( n11045, n9908, n11049 );
nand U102962 ( n31138, n3407, n73532 );
nor U102963 ( n33913, n74131, n33671 );
not U102964 ( n805, n41183 );
nor U102965 ( n10112, n10115, n9897 );
nor U102966 ( n39925, n38424, n76404 );
xnor U102967 ( n31865, n32611, n32669 );
xor U102968 ( n32669, n75042, n76470 );
nor U102969 ( n32636, n32638, n76896 );
nor U102970 ( n32638, n32639, n32640 );
nand U102971 ( n32640, n32641, n32642 );
nand U102972 ( n32639, n32643, n32644 );
not U102973 ( n2502, n19707 );
nor U102974 ( n68831, n68832, n68833 );
nor U102975 ( n68832, n74205, n68402 );
nor U102976 ( n68833, n74181, n68401 );
nor U102977 ( n26832, n26833, n26834 );
nor U102978 ( n26833, n74206, n26401 );
nor U102979 ( n26834, n74184, n26400 );
nor U102980 ( n59972, n59973, n59974 );
nor U102981 ( n59973, n74207, n59540 );
nor U102982 ( n59974, n74185, n59539 );
nor U102983 ( n39765, n39821, n36767 );
nand U102984 ( n39999, n40090, n40089 );
nor U102985 ( n40090, n36822, n36594 );
nor U102986 ( n39866, n39922, n36672 );
nor U102987 ( n39965, n39999, n36293 );
and U102988 ( n40178, n40257, n1893 );
nor U102989 ( n40257, n37007, n37022 );
and U102990 ( n39572, n39695, n39694 );
nor U102991 ( n39695, n36327, n36735 );
and U102992 ( n39334, n39444, n39443 );
nor U102993 ( n39444, n36802, n36618 );
and U102994 ( n39443, n39573, n39572 );
nor U102995 ( n39573, n36577, n36955 );
and U102996 ( n40089, n40179, n40178 );
nor U102997 ( n40179, n36655, n36386 );
and U102998 ( n39209, n39335, n39334 );
nor U102999 ( n39335, n2102, n36403 );
nor U103000 ( n51357, n49989, n73421 );
nor U103001 ( n68830, n68834, n68835 );
nor U103002 ( n68834, n74211, n68406 );
nor U103003 ( n68835, n74195, n68405 );
nor U103004 ( n26831, n26835, n26836 );
nor U103005 ( n26835, n74212, n26405 );
nor U103006 ( n26836, n74196, n26404 );
nor U103007 ( n59971, n59975, n59976 );
nor U103008 ( n59975, n74213, n59544 );
nor U103009 ( n59976, n74197, n59543 );
not U103010 ( n803, n40972 );
not U103011 ( n807, n40806 );
nor U103012 ( n33891, n74063, n33635 );
nand U103013 ( n33887, n33888, n33889 );
nor U103014 ( n33888, n33892, n33893 );
nor U103015 ( n33889, n33890, n33891 );
nor U103016 ( n33892, n74126, n33640 );
nand U103017 ( n71302, n72802, n72803 );
nor U103018 ( n72802, n72806, n72807 );
nor U103019 ( n72803, n72804, n72805 );
nor U103020 ( n72807, n73523, n73026 );
nor U103021 ( n68001, n68004, n76197 );
nor U103022 ( n68004, n74431, n72950 );
nor U103023 ( n25998, n26001, n76521 );
nor U103024 ( n26001, n74432, n72951 );
nor U103025 ( n59136, n59139, n76263 );
nor U103026 ( n59139, n74433, n72952 );
nor U103027 ( n33890, n74121, n33636 );
nor U103028 ( n72804, n73056, n71105 );
nand U103029 ( n71273, n1242, n71274 );
nor U103030 ( n33893, n74104, n33639 );
nor U103031 ( n19535, n16861, n73022 );
nor U103032 ( n37209, n36577, n76802 );
nor U103033 ( n46467, n46469, n76330 );
nor U103034 ( n46469, n46470, n46471 );
nand U103035 ( n46471, n46472, n46473 );
nand U103036 ( n46470, n46474, n46475 );
nand U103037 ( n46475, n76659, n45653 );
nor U103038 ( n32728, n32732, n3105 );
and U103039 ( n32732, n31949, n32733 );
nor U103040 ( n32718, n32720, n76896 );
nor U103041 ( n32720, n32721, n32722 );
nand U103042 ( n32721, n32741, n32742 );
nand U103043 ( n32722, n32723, n32724 );
and U103044 ( n31945, n32752, n32753 );
xor U103045 ( n32753, n74973, n76471 );
nor U103046 ( n32752, n31951, n32754 );
nor U103047 ( n32754, n3150, n74961 );
nor U103048 ( n25525, n25527, n76905 );
nor U103049 ( n25527, n25528, n25529 );
nand U103050 ( n25529, n25530, n25531 );
nand U103051 ( n25528, n25532, n25533 );
nor U103052 ( n67530, n67532, n76870 );
nor U103053 ( n67532, n67533, n67534 );
nand U103054 ( n67534, n67535, n67536 );
nand U103055 ( n67533, n67537, n67538 );
nor U103056 ( n58662, n58664, n76879 );
nor U103057 ( n58664, n58665, n58666 );
nand U103058 ( n58666, n58667, n58668 );
nand U103059 ( n58665, n58669, n58670 );
nand U103060 ( n25533, n76753, n24742 );
nand U103061 ( n67538, n76707, n66577 );
nand U103062 ( n58670, n76686, n57876 );
nand U103063 ( n41594, n720, n41183 );
nor U103064 ( n52343, n49982, n73424 );
nand U103065 ( n32742, n32743, n74973 );
nand U103066 ( n32743, n32744, n3115 );
not U103067 ( n3115, n32702 );
nor U103068 ( n32744, n32750, n32751 );
nor U103069 ( n39872, n76415, n74399 );
nand U103070 ( n36730, n39867, n39868 );
nor U103071 ( n39868, n39869, n39870 );
nor U103072 ( n39867, n39872, n39873 );
nor U103073 ( n39870, n76411, n74398 );
nand U103074 ( n63312, n41006, n40972 );
nand U103075 ( n40726, n41327, n41328 );
nand U103076 ( n41328, n76848, n41329 );
nand U103077 ( n41327, n76844, n40732 );
nand U103078 ( n63309, n709, n41011 );
nand U103079 ( n41664, n41670, n41671 );
nand U103080 ( n41670, n76010, n40727 );
nand U103081 ( n41671, n41119, n76378 );
xnor U103082 ( n36885, n37072, n2040 );
nand U103083 ( n37072, n37073, n37074 );
nand U103084 ( n37073, n76829, n36572 );
nand U103085 ( n37074, n36955, n2035 );
not U103086 ( n3409, n31132 );
nor U103087 ( n46963, n47022, n47023 );
and U103088 ( n47023, n47024, n76342 );
nand U103089 ( n47024, n73099, n72948 );
nand U103090 ( n64022, n41323, n40967 );
nor U103091 ( n33895, n33896, n33897 );
nor U103092 ( n33896, n74134, n33646 );
nor U103093 ( n33897, n74122, n33645 );
nand U103094 ( n71271, n71279, n71280 );
nor U103095 ( n71279, n71285, n71286 );
nor U103096 ( n71280, n71281, n71282 );
nor U103097 ( n71286, n73509, n73025 );
nor U103098 ( n71281, n73507, n71284 );
nor U103099 ( n51860, n49989, n73021 );
nor U103100 ( n45621, n45628, n45629 );
and U103101 ( n45628, n74974, n45630 );
nor U103102 ( n33894, n33898, n33899 );
nor U103103 ( n33898, n74137, n33650 );
nor U103104 ( n33899, n74127, n33649 );
nor U103105 ( n24711, n24718, n24634 );
and U103106 ( n24718, n74975, n24719 );
nor U103107 ( n66546, n66553, n66471 );
and U103108 ( n66553, n74976, n66554 );
nor U103109 ( n57845, n57852, n57766 );
and U103110 ( n57852, n74977, n57853 );
nor U103111 ( n72806, n73057, n71108 );
nor U103112 ( n49840, n76097, n73403 );
nand U103113 ( n31130, n34130, n73532 );
xnor U103114 ( n36567, n36875, n2040 );
nand U103115 ( n36875, n36876, n36877 );
nand U103116 ( n36876, n76826, n36613 );
nand U103117 ( n36877, n36577, n2035 );
nand U103118 ( n38117, n38744, n38737 );
nand U103119 ( n38744, n2149, n38747 );
nand U103120 ( n38747, n38746, n37600 );
nor U103121 ( n17207, n16861, n73404 );
nand U103122 ( n41271, n41321, n41322 );
nand U103123 ( n41322, n76848, n40967 );
nand U103124 ( n41321, n76844, n41323 );
nor U103125 ( n18577, n17028, n73420 );
xor U103126 ( n41005, n41275, n40826 );
nand U103127 ( n41275, n41276, n41277 );
nand U103128 ( n41276, n76844, n41178 );
nand U103129 ( n41277, n41011, n41264 );
nand U103130 ( n41114, n65319, n65320 );
nor U103131 ( n65320, n65321, n65322 );
nor U103132 ( n65319, n65324, n65325 );
nor U103133 ( n65322, n76245, n74396 );
nor U103134 ( n65324, n76249, n74397 );
not U103135 ( n2102, n36915 );
nand U103136 ( n71894, n71327, n71243 );
nor U103137 ( n67998, n68057, n68058 );
and U103138 ( n68058, n68059, n76198 );
nand U103139 ( n68059, n73104, n72950 );
nor U103140 ( n25995, n26054, n26055 );
and U103141 ( n26055, n26056, n76522 );
nand U103142 ( n26056, n73105, n72951 );
nor U103143 ( n59133, n59195, n59196 );
and U103144 ( n59196, n59197, n76264 );
nand U103145 ( n59197, n73106, n72952 );
and U103146 ( n71760, n71243, n71096 );
nor U103147 ( n71285, n73508, n71287 );
nor U103148 ( n11675, n17525, n76789 );
nor U103149 ( n50129, n49982, n73410 );
nand U103150 ( n40961, n41265, n41266 );
nand U103151 ( n41266, n76848, n41006 );
nand U103152 ( n41265, n76844, n40972 );
nor U103153 ( n38150, n38746, n38832 );
nor U103154 ( n38832, n36425, n1892 );
nor U103155 ( n50569, n49982, n73008 );
nand U103156 ( n62781, n41284, n40806 );
nand U103157 ( n39322, n36702, n36403 );
xnor U103158 ( n38135, n37600, n38746 );
nand U103159 ( n36321, n36959, n36960 );
nand U103160 ( n36960, n76807, n36961 );
nand U103161 ( n36959, n76827, n36327 );
nand U103162 ( n36322, n39822, n39823 );
nor U103163 ( n39823, n39824, n39825 );
nor U103164 ( n39822, n39827, n39828 );
nor U103165 ( n39825, n76411, n74402 );
not U103166 ( n2113, n39260 );
nor U103167 ( n33827, n74222, n33657 );
nand U103168 ( n33823, n33824, n33825 );
nor U103169 ( n33824, n33828, n33829 );
nor U103170 ( n33825, n33826, n33827 );
nor U103171 ( n33828, n74233, n33662 );
not U103172 ( n2054, n36403 );
nor U103173 ( n33829, n74224, n33661 );
nand U103174 ( n2821, n38104, n38105 );
nor U103175 ( n38104, n38111, n38112 );
nor U103176 ( n38105, n38106, n38107 );
nor U103177 ( n38112, n76811, n74773 );
nor U103178 ( n19116, n16861, n73423 );
nand U103179 ( n40517, n73479, n73042 );
and U103180 ( n40511, n40513, n40514 );
nor U103181 ( n40514, n40515, n40516 );
nor U103182 ( n40513, n40517, n40518 );
nand U103183 ( n40516, n73494, n73047 );
nor U103184 ( n18414, n17028, n73018 );
nor U103185 ( n33826, n74228, n33658 );
nor U103186 ( n33833, n74229, n33667 );
nand U103187 ( n33822, n33830, n33831 );
nor U103188 ( n33830, n33834, n33835 );
nor U103189 ( n33831, n33832, n33833 );
nor U103190 ( n33834, n74242, n33672 );
nor U103191 ( n33832, n74238, n33668 );
nand U103192 ( n48673, n48674, n48675 );
nand U103193 ( n48674, n569, n40972 );
nand U103194 ( n48675, n48676, n45754 );
nor U103195 ( n64790, n76249, n74406 );
nand U103196 ( n40727, n64785, n64786 );
nor U103197 ( n64786, n64787, n64788 );
nor U103198 ( n64785, n64790, n64791 );
nor U103199 ( n64788, n76245, n74401 );
nor U103200 ( n46558, n46560, n76330 );
nor U103201 ( n46560, n46561, n46562 );
nand U103202 ( n46561, n46582, n46583 );
nand U103203 ( n46562, n46563, n46564 );
nand U103204 ( n45718, n46573, n46574 );
nand U103205 ( n46574, n46521, n46482 );
nor U103206 ( n46573, n46575, n46576 );
nor U103207 ( n46576, n46482, n46529 );
nor U103208 ( n33835, n74235, n33671 );
nand U103209 ( n38414, n38415, n38416 );
nand U103210 ( n38416, n76816, n36537 );
nand U103211 ( n38415, n76812, n38417 );
nor U103212 ( n67605, n67607, n76870 );
nor U103213 ( n67607, n67608, n67609 );
nand U103214 ( n67608, n67629, n67630 );
nand U103215 ( n67609, n67610, n67611 );
nor U103216 ( n25600, n25602, n76905 );
nor U103217 ( n25602, n25603, n25604 );
nand U103218 ( n25603, n25624, n25625 );
nand U103219 ( n25604, n25605, n25606 );
nor U103220 ( n58737, n58739, n76879 );
nor U103221 ( n58739, n58740, n58741 );
nand U103222 ( n58740, n58761, n58762 );
nand U103223 ( n58741, n58742, n58743 );
nand U103224 ( n66644, n67620, n67621 );
nand U103225 ( n67621, n67582, n67545 );
nor U103226 ( n67620, n67622, n67623 );
nor U103227 ( n67623, n67545, n67590 );
nand U103228 ( n24809, n25615, n25616 );
nand U103229 ( n25616, n25577, n25540 );
nor U103230 ( n25615, n25617, n25618 );
nor U103231 ( n25618, n25540, n25585 );
nand U103232 ( n57943, n58752, n58753 );
nand U103233 ( n58753, n58714, n58677 );
nor U103234 ( n58752, n58754, n58755 );
nor U103235 ( n58755, n58677, n58722 );
nand U103236 ( n40515, n73496, n73050 );
nand U103237 ( n41668, n76010, n41119 );
nor U103238 ( n39824, n38395, n76404 );
nand U103239 ( n36884, n36953, n36954 );
nand U103240 ( n36954, n76807, n36572 );
nand U103241 ( n36953, n76827, n36955 );
nand U103242 ( n39417, n36802, n36398 );
nand U103243 ( n40518, n73495, n73035 );
xor U103244 ( n36612, n36888, n36481 );
nand U103245 ( n36888, n36889, n36890 );
nand U103246 ( n36889, n76827, n36797 );
nand U103247 ( n36890, n36618, n2035 );
nand U103248 ( n37555, n2179, n36403 );
nor U103249 ( n45366, n44066, n45391 );
nor U103250 ( n33813, n74221, n33635 );
nand U103251 ( n33809, n33810, n33811 );
nor U103252 ( n33810, n33814, n33815 );
nor U103253 ( n33811, n33812, n33813 );
nor U103254 ( n33814, n74230, n33640 );
nor U103255 ( n51814, n49982, n73425 );
nor U103256 ( n33812, n74226, n33636 );
nand U103257 ( n49142, n49143, n49144 );
nand U103258 ( n49144, n569, n40935 );
nand U103259 ( n49143, n76857, n49145 );
nand U103260 ( n36566, n36878, n36879 );
nand U103261 ( n36879, n76808, n36613 );
nand U103262 ( n36878, n76826, n36577 );
nor U103263 ( n33815, n74223, n33639 );
nor U103264 ( n51338, n49989, n73019 );
nand U103265 ( n45643, n45651, n45652 );
nand U103266 ( n45651, n45632, n75208 );
nand U103267 ( n45652, n76663, n45653 );
nand U103268 ( n15826, n45641, n45642 );
nor U103269 ( n45641, n45659, n45660 );
nor U103270 ( n45642, n45643, n45644 );
nor U103271 ( n45659, n75014, n76669 );
nor U103272 ( n46505, n46507, n76330 );
nor U103273 ( n46507, n46508, n46509 );
nand U103274 ( n46508, n46530, n46531 );
nand U103275 ( n46509, n46510, n46511 );
and U103276 ( n45695, n46518, n46519 );
nand U103277 ( n46518, n46525, n46526 );
nand U103278 ( n46519, n46520, n46478 );
nand U103279 ( n46526, n76006, n74919 );
nand U103280 ( n24732, n24740, n24741 );
nand U103281 ( n24740, n24721, n74850 );
nand U103282 ( n24741, n76759, n24742 );
nand U103283 ( n66567, n66575, n66576 );
nand U103284 ( n66575, n66556, n74848 );
nand U103285 ( n66576, n76711, n66577 );
nand U103286 ( n57866, n57874, n57875 );
nand U103287 ( n57874, n57855, n74851 );
nand U103288 ( n57875, n76692, n57876 );
nand U103289 ( n6846, n24730, n24731 );
nor U103290 ( n24730, n24748, n24749 );
nor U103291 ( n24731, n24732, n24733 );
nor U103292 ( n24748, n74999, n76765 );
nand U103293 ( n11336, n66565, n66566 );
nor U103294 ( n66565, n66583, n66584 );
nor U103295 ( n66566, n66567, n66568 );
nor U103296 ( n66583, n75003, n76717 );
nand U103297 ( n13581, n57864, n57865 );
nor U103298 ( n57864, n57882, n57883 );
nor U103299 ( n57865, n57866, n57867 );
nor U103300 ( n57882, n75000, n76698 );
nor U103301 ( n38166, n1892, n38896 );
and U103302 ( n38896, n2138, n38897 );
nand U103303 ( n38897, n38898, n36935 );
nor U103304 ( n67566, n67568, n76870 );
nor U103305 ( n67568, n67569, n67570 );
nand U103306 ( n67569, n67591, n67592 );
nand U103307 ( n67570, n67571, n67572 );
nor U103308 ( n25561, n25563, n76905 );
nor U103309 ( n25563, n25564, n25565 );
nand U103310 ( n25564, n25586, n25587 );
nand U103311 ( n25565, n25566, n25567 );
nor U103312 ( n58698, n58700, n76879 );
nor U103313 ( n58700, n58701, n58702 );
nand U103314 ( n58701, n58723, n58724 );
nand U103315 ( n58702, n58703, n58704 );
and U103316 ( n66619, n67579, n67580 );
nand U103317 ( n67579, n67586, n67587 );
nand U103318 ( n67580, n67581, n67541 );
nand U103319 ( n67587, n75990, n74947 );
and U103320 ( n24784, n25574, n25575 );
nand U103321 ( n25574, n25581, n25582 );
nand U103322 ( n25575, n25576, n25536 );
nand U103323 ( n25582, n76027, n74949 );
and U103324 ( n57918, n58711, n58712 );
nand U103325 ( n58711, n58718, n58719 );
nand U103326 ( n58712, n58713, n58673 );
nand U103327 ( n58719, n75998, n74950 );
nand U103328 ( n62687, n41183, n40801 );
nand U103329 ( n2816, n38113, n38114 );
nor U103330 ( n38113, n38111, n38118 );
nor U103331 ( n38114, n38115, n38116 );
nor U103332 ( n38118, n76809, n74826 );
nor U103333 ( n44817, n44066, n44561 );
nand U103334 ( n16211, n44807, n44808 );
nor U103335 ( n44808, n44809, n44810 );
nor U103336 ( n44807, n44816, n44817 );
nor U103337 ( n44809, n44814, n44815 );
nor U103338 ( n44063, n44066, n43799 );
nand U103339 ( n36961, n39766, n39767 );
nor U103340 ( n39767, n39768, n39769 );
nor U103341 ( n39766, n39771, n39772 );
nor U103342 ( n39769, n76411, n74411 );
nand U103343 ( n71516, n71735, n71736 );
nand U103344 ( n71735, n71739, n71327 );
nand U103345 ( n71736, n71737, n71096 );
nand U103346 ( n71739, n71272, n71740 );
nor U103347 ( n33735, n74260, n33657 );
nand U103348 ( n33731, n33732, n33733 );
nor U103349 ( n33732, n33736, n33737 );
nor U103350 ( n33733, n33734, n33735 );
nor U103351 ( n33736, n74271, n33662 );
nor U103352 ( n37205, n36618, n76802 );
nor U103353 ( n39641, n76415, n74420 );
nand U103354 ( n36613, n39636, n39637 );
nor U103355 ( n39637, n39638, n39639 );
nor U103356 ( n39636, n39641, n39642 );
nor U103357 ( n39639, n76411, n74419 );
nor U103358 ( n64787, n49029, n76242 );
nor U103359 ( n33817, n33818, n33819 );
nor U103360 ( n33818, n74237, n33646 );
nor U103361 ( n33819, n74227, n33645 );
nor U103362 ( n33737, n74262, n33661 );
nand U103363 ( n40967, n64345, n64346 );
nor U103364 ( n64346, n64347, n64348 );
nor U103365 ( n64345, n64350, n64351 );
nor U103366 ( n64348, n76245, n74407 );
nor U103367 ( n64350, n76249, n74413 );
nor U103368 ( n33816, n33820, n33821 );
nor U103369 ( n33820, n74239, n33650 );
nor U103370 ( n33821, n74231, n33649 );
nor U103371 ( n33734, n74267, n33658 );
nor U103372 ( n33741, n74268, n33667 );
nand U103373 ( n33730, n33738, n33739 );
nor U103374 ( n33738, n33742, n33743 );
nor U103375 ( n33739, n33740, n33741 );
nor U103376 ( n33742, n74278, n33672 );
nor U103377 ( n33740, n74276, n33668 );
nand U103378 ( n41595, n730, n40806 );
and U103379 ( n41654, n41658, n41659 );
nand U103380 ( n41658, n76010, n41329 );
nand U103381 ( n41659, n40732, n76378 );
nor U103382 ( n33743, n74272, n33671 );
nand U103383 ( n41004, n41273, n41274 );
nand U103384 ( n41274, n76848, n41178 );
nand U103385 ( n41273, n76844, n41011 );
nor U103386 ( n18238, n17028, n73418 );
nand U103387 ( n36572, n39696, n39697 );
nor U103388 ( n39697, n39698, n39699 );
nor U103389 ( n39696, n39701, n39702 );
nor U103390 ( n39699, n76411, n74421 );
nand U103391 ( n41655, n41660, n41661 );
nand U103392 ( n41661, n41329, n76378 );
nand U103393 ( n41660, n76010, n40732 );
nand U103394 ( n31852, n31863, n31864 );
nand U103395 ( n31863, n31838, n75185 );
nand U103396 ( n31864, n76776, n31865 );
nand U103397 ( n4616, n31850, n31851 );
nor U103398 ( n31850, n31872, n31873 );
nor U103399 ( n31851, n31852, n31853 );
nor U103400 ( n31872, n75069, n76783 );
nor U103401 ( n17752, n16861, n75913 );
nor U103402 ( n33721, n74258, n33635 );
nand U103403 ( n33717, n33718, n33719 );
nor U103404 ( n33718, n33722, n33723 );
nor U103405 ( n33719, n33720, n33721 );
nor U103406 ( n33722, n74269, n33640 );
not U103407 ( n2107, n36907 );
nor U103408 ( n33720, n74264, n33636 );
nor U103409 ( n33723, n74261, n33639 );
nand U103410 ( n41006, n64195, n64196 );
nor U103411 ( n64196, n64197, n64198 );
nor U103412 ( n64195, n64200, n64201 );
nor U103413 ( n64198, n76245, n74415 );
nor U103414 ( n64200, n76249, n74416 );
nand U103415 ( n49023, n49024, n49025 );
nand U103416 ( n49024, n569, n41119 );
nand U103417 ( n49025, n49026, n45754 );
nor U103418 ( n64347, n48794, n76242 );
nand U103419 ( n39319, n2180, n36915 );
nor U103420 ( n32675, n32677, n76896 );
nor U103421 ( n32677, n32678, n32679 );
nand U103422 ( n32678, n32698, n32699 );
nand U103423 ( n32679, n32680, n32681 );
nand U103424 ( n32680, n76772, n31907 );
nand U103425 ( n47237, n47282, n47283 );
nand U103426 ( n47283, n47284, n47285 );
nor U103427 ( n47512, n47515, n47516 );
and U103428 ( n47329, n47433, n47434 );
nand U103429 ( n47434, n47435, n47436 );
nor U103430 ( n47022, n74427, n76005 );
nor U103431 ( n19250, n73020, n17028 );
nor U103432 ( n33725, n33726, n33727 );
nor U103433 ( n33726, n74275, n33646 );
nor U103434 ( n33727, n74265, n33645 );
nor U103435 ( n39698, n38361, n76404 );
nand U103436 ( n37457, n36747, n36907 );
nor U103437 ( n33724, n33728, n33729 );
nor U103438 ( n33728, n74277, n33650 );
nor U103439 ( n33729, n74270, n33649 );
nand U103440 ( n38446, n38447, n38448 );
nand U103441 ( n38448, n76816, n36360 );
nand U103442 ( n38447, n76812, n38449 );
xor U103443 ( n38187, n36935, n38898 );
nor U103444 ( n37197, n36802, n76802 );
nand U103445 ( n49265, n49266, n49267 );
nand U103446 ( n49267, n569, n41150 );
nand U103447 ( n49266, n76857, n49268 );
nor U103448 ( n17486, n16861, n73009 );
nor U103449 ( n38198, n38898, n39030 );
nor U103450 ( n39030, n39021, n1890 );
nand U103451 ( n15816, n45696, n45697 );
nor U103452 ( n45697, n45698, n45699 );
nor U103453 ( n45696, n45713, n45714 );
nand U103454 ( n45698, n45707, n45708 );
nand U103455 ( n45714, n45715, n45716 );
nand U103456 ( n45716, n7434, n42628 );
nand U103457 ( n45715, n76663, n45718 );
nand U103458 ( n36611, n36886, n36887 );
nand U103459 ( n36887, n76807, n36797 );
nand U103460 ( n36886, n76827, n36618 );
nand U103461 ( n6836, n24785, n24786 );
nor U103462 ( n24786, n24787, n24788 );
nor U103463 ( n24785, n24804, n24805 );
nand U103464 ( n24787, n24797, n24798 );
nand U103465 ( n13571, n57919, n57920 );
nor U103466 ( n57920, n57921, n57922 );
nor U103467 ( n57919, n57938, n57939 );
nand U103468 ( n57921, n57931, n57932 );
nand U103469 ( n11326, n66620, n66621 );
nor U103470 ( n66621, n66622, n66623 );
nor U103471 ( n66620, n66639, n66640 );
nand U103472 ( n66622, n66632, n66633 );
nor U103473 ( n18750, n16861, n73422 );
nand U103474 ( n26267, n26312, n26313 );
nand U103475 ( n26313, n26314, n26315 );
nand U103476 ( n59406, n59451, n59452 );
nand U103477 ( n59452, n59453, n59454 );
nor U103478 ( n26532, n26535, n26536 );
nor U103479 ( n59674, n59677, n59678 );
and U103480 ( n26360, n26453, n26454 );
nand U103481 ( n26454, n26455, n26456 );
and U103482 ( n59499, n59592, n59593 );
nand U103483 ( n59593, n59594, n59595 );
nand U103484 ( n68268, n68313, n68314 );
nand U103485 ( n68314, n68315, n68316 );
nor U103486 ( n68533, n68536, n68537 );
and U103487 ( n68361, n68454, n68455 );
nand U103488 ( n68455, n68456, n68457 );
nor U103489 ( n26054, n74439, n76026 );
nor U103490 ( n59195, n74440, n75997 );
nor U103491 ( n68057, n74438, n75989 );
nand U103492 ( n32723, n32739, n32740 );
nand U103493 ( n71410, n72814, n72815 );
nor U103494 ( n72814, n72818, n72819 );
nor U103495 ( n72815, n72816, n72817 );
nor U103496 ( n72819, n73531, n73026 );
nand U103497 ( n38390, n38391, n38392 );
nand U103498 ( n38391, n76816, n36735 );
nand U103499 ( n38392, n1863, n76443 );
nor U103500 ( n72816, n73528, n71105 );
nor U103501 ( n11689, n17014, n76789 );
nand U103502 ( n15821, n45665, n45666 );
nor U103503 ( n45666, n45667, n45668 );
nor U103504 ( n45665, n45690, n45691 );
nand U103505 ( n45668, n45669, n45670 );
nand U103506 ( n39255, n2182, n36907 );
nor U103507 ( n33656, n74302, n33657 );
nand U103508 ( n66615, n66616, n66617 );
nand U103509 ( n66617, n5660, n63167 );
nand U103510 ( n66616, n66619, n76710 );
nand U103511 ( n24780, n24781, n24782 );
nand U103512 ( n24782, n3903, n22085 );
nand U103513 ( n24781, n24784, n76758 );
nand U103514 ( n57914, n57915, n57916 );
nand U103515 ( n57916, n6535, n55195 );
nand U103516 ( n57915, n57918, n76691 );
nand U103517 ( n33652, n33653, n33654 );
nor U103518 ( n33653, n33659, n33660 );
nor U103519 ( n33654, n33655, n33656 );
nor U103520 ( n33659, n74311, n33662 );
nand U103521 ( n11331, n66589, n66590 );
nor U103522 ( n66590, n66591, n66592 );
nor U103523 ( n66589, n66614, n66615 );
nand U103524 ( n66592, n66593, n66594 );
nand U103525 ( n6841, n24754, n24755 );
nor U103526 ( n24755, n24756, n24757 );
nor U103527 ( n24754, n24779, n24780 );
nand U103528 ( n24757, n24758, n24759 );
nand U103529 ( n13576, n57888, n57889 );
nor U103530 ( n57889, n57890, n57891 );
nor U103531 ( n57888, n57913, n57914 );
nand U103532 ( n57891, n57892, n57893 );
nor U103533 ( n33660, n74304, n33661 );
nor U103534 ( n19247, n17028, n75919 );
nor U103535 ( n33655, n74307, n33658 );
nor U103536 ( n33666, n74308, n33667 );
nand U103537 ( n33651, n33663, n33664 );
nor U103538 ( n33663, n33669, n33670 );
nor U103539 ( n33664, n33665, n33666 );
nor U103540 ( n33669, n74317, n33672 );
nor U103541 ( n33665, n74315, n33668 );
nor U103542 ( n51162, n50001, n73021 );
nor U103543 ( n33670, n74312, n33671 );
nand U103544 ( n41329, n64494, n64495 );
nor U103545 ( n64495, n64496, n64497 );
nor U103546 ( n64494, n64499, n64500 );
nor U103547 ( n64497, n76245, n74428 );
nor U103548 ( n64499, n76249, n74430 );
nor U103549 ( n72818, n73529, n71108 );
nor U103550 ( n38215, n1890, n39082 );
and U103551 ( n39082, n2122, n39083 );
nand U103552 ( n39083, n39084, n39085 );
nor U103553 ( n33634, n74299, n33635 );
nand U103554 ( n33630, n33631, n33632 );
nor U103555 ( n33631, n33637, n33638 );
nor U103556 ( n33632, n33633, n33634 );
nor U103557 ( n33637, n74309, n33640 );
nor U103558 ( n33633, n74305, n33636 );
nor U103559 ( n33638, n74303, n33639 );
nand U103560 ( n49574, n49575, n49576 );
nand U103561 ( n49576, n569, n41059 );
nand U103562 ( n49575, n76857, n49577 );
nand U103563 ( n37456, n36512, n36915 );
not U103564 ( n5144, n10763 );
nand U103565 ( n9327, n14797, n14798 );
or U103566 ( n14798, n73525, n10273 );
nor U103567 ( n12224, n13420, n76602 );
nand U103568 ( n12809, n4891, n72970 );
nor U103569 ( n14512, n73980, n14032 );
nand U103570 ( n13472, n13517, n13518 );
nor U103571 ( n13517, n13519, n13520 );
nor U103572 ( n13520, n76602, n73117 );
nor U103573 ( n13519, n13522, n13523 );
nand U103574 ( n12930, n13030, n13032 );
nor U103575 ( n13030, n13033, n13034 );
nor U103576 ( n13034, n76602, n74653 );
nor U103577 ( n13033, n13035, n13037 );
not U103578 ( n4891, n11879 );
nand U103579 ( n13037, n13038, n13039 );
nand U103580 ( n13038, n76603, n74653 );
nand U103581 ( n13523, n13524, n13525 );
nand U103582 ( n13524, n76603, n73117 );
nand U103583 ( n14507, n14508, n14509 );
nor U103584 ( n14508, n14513, n14514 );
nor U103585 ( n14509, n14510, n14512 );
nor U103586 ( n14513, n73992, n14038 );
nand U103587 ( n12693, n76724, n11779 );
nor U103588 ( n14514, n73998, n14037 );
nand U103589 ( n71740, n1222, n71274 );
nor U103590 ( n47855, n73554, n47381 );
nand U103591 ( n47851, n47852, n47853 );
nor U103592 ( n47852, n47857, n47858 );
nor U103593 ( n47853, n47854, n47855 );
nor U103594 ( n47857, n73565, n47386 );
not U103595 ( n7623, n47650 );
nor U103596 ( n47862, n73561, n47391 );
nand U103597 ( n47850, n47859, n47860 );
nor U103598 ( n47859, n47865, n47866 );
nor U103599 ( n47860, n47861, n47862 );
nor U103600 ( n47865, n73574, n47396 );
nor U103601 ( n47854, n73560, n47382 );
nor U103602 ( n11557, n10178, n11594 );
nor U103603 ( n47861, n73571, n47392 );
nor U103604 ( n47858, n73556, n47385 );
nor U103605 ( n45516, n49816, n76834 );
nor U103606 ( n14510, n73985, n14033 );
and U103607 ( n41503, n41508, n41509 );
nand U103608 ( n41508, n41510, n76388 );
nand U103609 ( n41509, n780, n76385 );
nor U103610 ( n14519, n73983, n14044 );
nand U103611 ( n14505, n14515, n14517 );
nor U103612 ( n14515, n14520, n14522 );
nor U103613 ( n14517, n14518, n14519 );
nor U103614 ( n14520, n73995, n14050 );
nor U103615 ( n47866, n73567, n47395 );
nor U103616 ( n11105, n10178, n10785 );
nand U103617 ( n9476, n11093, n11094 );
nor U103618 ( n11094, n11095, n11097 );
nor U103619 ( n11093, n11104, n11105 );
nor U103620 ( n11095, n11102, n11103 );
xor U103621 ( n36695, n36481, n36912 );
nor U103622 ( n36912, n36913, n36914 );
nor U103623 ( n36914, n2180, n36423 );
nor U103624 ( n36913, n36424, n36915 );
nor U103625 ( n14522, n73991, n14049 );
nand U103626 ( n41649, n41804, n41805 );
nand U103627 ( n41804, n76011, n40967 );
nand U103628 ( n41805, n41323, n76379 );
nor U103629 ( n51184, n73419, n49989 );
nand U103630 ( n31904, n31905, n31906 );
nand U103631 ( n31905, n3059, n3558 );
nand U103632 ( n31906, n76776, n31907 );
nand U103633 ( n4611, n31878, n31879 );
nor U103634 ( n31879, n31880, n31881 );
nor U103635 ( n31878, n31903, n31904 );
nand U103636 ( n31881, n31882, n31883 );
xor U103637 ( n36511, n36481, n36904 );
nor U103638 ( n36904, n36905, n36906 );
nor U103639 ( n36906, n2182, n36423 );
nor U103640 ( n36905, n36424, n36907 );
nor U103641 ( n33642, n33643, n33644 );
nor U103642 ( n33643, n74313, n33646 );
nor U103643 ( n33644, n74306, n33645 );
nand U103644 ( n72165, n71143, n71302 );
nand U103645 ( n33371, n76022, n73114 );
nor U103646 ( n14518, n73988, n14045 );
nor U103647 ( n10174, n10178, n9897 );
nor U103648 ( n33641, n33647, n33648 );
nor U103649 ( n33647, n74316, n33650 );
nor U103650 ( n33648, n74310, n33649 );
nor U103651 ( n12864, n12887, n11870 );
nor U103652 ( n12892, n74946, n12809 );
nor U103653 ( n12882, n12840, n12883 );
nand U103654 ( n12883, n12884, n12885 );
nand U103655 ( n12884, n12893, n12857 );
nand U103656 ( n12885, n12864, n76603 );
nor U103657 ( n12844, n12847, n76596 );
nor U103658 ( n12847, n12848, n12849 );
nand U103659 ( n12849, n12850, n12852 );
nand U103660 ( n12848, n12862, n12863 );
nor U103661 ( n26876, n73654, n26412 );
nor U103662 ( n60016, n73653, n59551 );
nor U103663 ( n68875, n73652, n68413 );
nand U103664 ( n26872, n26873, n26874 );
nor U103665 ( n26873, n26878, n26879 );
nor U103666 ( n26874, n26875, n26876 );
nor U103667 ( n26878, n73689, n26417 );
nand U103668 ( n60012, n60013, n60014 );
nor U103669 ( n60013, n60018, n60019 );
nor U103670 ( n60014, n60015, n60016 );
nor U103671 ( n60018, n73688, n59556 );
nand U103672 ( n68871, n68872, n68873 );
nor U103673 ( n68872, n68877, n68878 );
nor U103674 ( n68873, n68874, n68875 );
nor U103675 ( n68877, n73686, n68418 );
not U103676 ( n5835, n68671 );
not U103677 ( n4064, n26670 );
not U103678 ( n6697, n59812 );
nor U103679 ( n47838, n73553, n47359 );
nand U103680 ( n47834, n47835, n47836 );
nor U103681 ( n47835, n47840, n47841 );
nor U103682 ( n47836, n47837, n47838 );
nor U103683 ( n47840, n73562, n47364 );
nor U103684 ( n26883, n73680, n26422 );
nor U103685 ( n60023, n73679, n59561 );
nor U103686 ( n68882, n73675, n68423 );
nand U103687 ( n26871, n26880, n26881 );
nor U103688 ( n26880, n26886, n26887 );
nor U103689 ( n26881, n26882, n26883 );
nor U103690 ( n26886, n73704, n26427 );
nand U103691 ( n60011, n60020, n60021 );
nor U103692 ( n60020, n60026, n60027 );
nor U103693 ( n60021, n60022, n60023 );
nor U103694 ( n60026, n73703, n59566 );
nand U103695 ( n68870, n68879, n68880 );
nor U103696 ( n68879, n68885, n68886 );
nor U103697 ( n68880, n68881, n68882 );
nor U103698 ( n68885, n73702, n68428 );
nor U103699 ( n26875, n73678, n26413 );
nor U103700 ( n60015, n73677, n59552 );
nor U103701 ( n68874, n73674, n68414 );
nor U103702 ( n47837, n73557, n47360 );
nor U103703 ( n26882, n73697, n26423 );
nor U103704 ( n60022, n73696, n59562 );
nor U103705 ( n68881, n73695, n68424 );
nor U103706 ( n26879, n73661, n26416 );
nor U103707 ( n60019, n73660, n59555 );
nor U103708 ( n68878, n73659, n68417 );
nor U103709 ( n47841, n73555, n47363 );
nor U103710 ( n26887, n73691, n26426 );
nor U103711 ( n60027, n73690, n59565 );
nor U103712 ( n68886, n73687, n68427 );
and U103713 ( n41814, n41822, n41823 );
nand U103714 ( n41822, n76011, n41178 );
nand U103715 ( n41823, n41011, n76379 );
xor U103716 ( n71240, n71241, n71242 );
nand U103717 ( n71241, n71245, n71246 );
nand U103718 ( n71242, n71243, n71244 );
nor U103719 ( n16832, n17028, n73009 );
nand U103720 ( n41825, n41832, n41833 );
nand U103721 ( n41833, n40801, n76379 );
nand U103722 ( n41832, n76383, n41183 );
and U103723 ( n41824, n41834, n41835 );
nand U103724 ( n41834, n76383, n40801 );
nand U103725 ( n41835, n41183, n76379 );
nand U103726 ( n12869, n12875, n12877 );
and U103727 ( n12875, n12879, n12818 );
nand U103728 ( n12877, n12864, n12878 );
nand U103729 ( n12878, n4896, n11879 );
nor U103730 ( n14445, n74082, n14032 );
nand U103731 ( n14440, n14442, n14443 );
nor U103732 ( n14442, n14447, n14448 );
nor U103733 ( n14443, n14444, n14445 );
nor U103734 ( n14447, n74101, n14038 );
nand U103735 ( n41813, n41820, n41821 );
nand U103736 ( n41821, n41178, n76379 );
nand U103737 ( n41820, n76011, n41011 );
nor U103738 ( n34087, n74340, n33657 );
nand U103739 ( n34083, n34084, n34085 );
nor U103740 ( n34084, n34088, n34089 );
nor U103741 ( n34085, n34086, n34087 );
nor U103742 ( n34088, n74350, n33662 );
nor U103743 ( n14448, n74111, n14037 );
nor U103744 ( n50690, n49989, n73017 );
not U103745 ( n4892, n12220 );
nor U103746 ( n51347, n50001, n73421 );
nor U103747 ( n34089, n74341, n33661 );
xnor U103748 ( n41174, n41278, n593 );
nand U103749 ( n41278, n41279, n41280 );
nand U103750 ( n41279, n76844, n40801 );
nand U103751 ( n41280, n41183, n41264 );
nor U103752 ( n14444, n74093, n14033 );
nor U103753 ( n26859, n73641, n26390 );
nor U103754 ( n59999, n73642, n59529 );
nor U103755 ( n68858, n73643, n68391 );
nand U103756 ( n26855, n26856, n26857 );
nor U103757 ( n26856, n26861, n26862 );
nor U103758 ( n26857, n26858, n26859 );
nor U103759 ( n26861, n73683, n26395 );
nand U103760 ( n59995, n59996, n59997 );
nor U103761 ( n59996, n60001, n60002 );
nor U103762 ( n59997, n59998, n59999 );
nor U103763 ( n60001, n73682, n59534 );
nand U103764 ( n68854, n68855, n68856 );
nor U103765 ( n68855, n68860, n68861 );
nor U103766 ( n68856, n68857, n68858 );
nor U103767 ( n68860, n73676, n68396 );
nor U103768 ( n14453, n74088, n14044 );
nand U103769 ( n14439, n14449, n14450 );
nor U103770 ( n14449, n14454, n14455 );
nor U103771 ( n14450, n14452, n14453 );
nor U103772 ( n14454, n74103, n14050 );
nor U103773 ( n26858, n73669, n26391 );
nor U103774 ( n59998, n73668, n59530 );
nor U103775 ( n68857, n73665, n68392 );
nor U103776 ( n34086, n74347, n33658 );
nor U103777 ( n49993, n49989, n73008 );
nor U103778 ( n26862, n73658, n26394 );
nor U103779 ( n60002, n73657, n59533 );
nor U103780 ( n68861, n73655, n68395 );
nand U103781 ( n41811, n41826, n41827 );
nand U103782 ( n41827, n41006, n76379 );
nand U103783 ( n41826, n76383, n40972 );
nor U103784 ( n34093, n74348, n33667 );
nand U103785 ( n34082, n34090, n34091 );
nor U103786 ( n34090, n34094, n34095 );
nor U103787 ( n34091, n34092, n34093 );
nor U103788 ( n34094, n74355, n33672 );
nor U103789 ( n18009, n17028, n73015 );
nor U103790 ( n14455, n74100, n14049 );
nor U103791 ( n10273, n11184, n73527 );
nor U103792 ( n34095, n74351, n33671 );
nand U103793 ( n12718, n12697, n12719 );
nor U103794 ( n47843, n47844, n47845 );
nor U103795 ( n47844, n73570, n47370 );
nor U103796 ( n47845, n73559, n47369 );
nor U103797 ( n14452, n74098, n14045 );
nor U103798 ( n34092, n74353, n33668 );
nor U103799 ( n37193, n36403, n76802 );
nor U103800 ( n47842, n47847, n47848 );
nor U103801 ( n47847, n73572, n47374 );
nor U103802 ( n47848, n73563, n47373 );
nor U103803 ( n31944, n31945, n31946 );
nor U103804 ( n31946, n76470, n31948 );
nand U103805 ( n31948, n3514, n31949 );
nand U103806 ( n4606, n31929, n31930 );
nor U103807 ( n31929, n31954, n31955 );
nor U103808 ( n31930, n31931, n31932 );
nor U103809 ( n31954, n75362, n76783 );
nor U103810 ( n14494, n73964, n14004 );
nand U103811 ( n14489, n14490, n14492 );
nor U103812 ( n14490, n14495, n14497 );
nor U103813 ( n14492, n14493, n14494 );
nor U103814 ( n14495, n73986, n14010 );
nand U103815 ( n41810, n41817, n41818 );
nand U103816 ( n41817, n76011, n41006 );
nand U103817 ( n41818, n40972, n76379 );
nor U103818 ( n33295, n74458, n76022 );
nor U103819 ( n50102, n49989, n73412 );
nor U103820 ( n45359, n44113, n45391 );
nor U103821 ( n14497, n73981, n14009 );
nor U103822 ( n12808, n4891, n72970 );
xor U103823 ( n38235, n39085, n39084 );
not U103824 ( n2553, n18558 );
nor U103825 ( n44870, n44113, n44561 );
not U103826 ( n5150, n11184 );
nor U103827 ( n14493, n73979, n14005 );
nor U103828 ( n14499, n14500, n14502 );
nor U103829 ( n14500, n73982, n14018 );
nor U103830 ( n14502, n73978, n14017 );
nor U103831 ( n38246, n39084, n39207 );
and U103832 ( n39207, n2113, n39208 );
nand U103833 ( n39208, n39209, n36907 );
nor U103834 ( n26864, n26865, n26866 );
nor U103835 ( n26865, n73694, n26401 );
nor U103836 ( n26866, n73673, n26400 );
nor U103837 ( n60004, n60005, n60006 );
nor U103838 ( n60005, n73693, n59540 );
nor U103839 ( n60006, n73672, n59539 );
nor U103840 ( n68863, n68864, n68865 );
nor U103841 ( n68864, n73692, n68402 );
nor U103842 ( n68865, n73667, n68401 );
nor U103843 ( n34073, n74338, n33635 );
nand U103844 ( n34069, n34070, n34071 );
nor U103845 ( n34070, n34074, n34075 );
nor U103846 ( n34071, n34072, n34073 );
nor U103847 ( n34074, n74345, n33640 );
nor U103848 ( n34072, n74343, n33636 );
nor U103849 ( n14610, n10260, n21296 );
nor U103850 ( n21296, n73527, n5150 );
nand U103851 ( n47435, n47483, n75934 );
nor U103852 ( n14498, n14503, n14504 );
nor U103853 ( n14503, n73989, n14023 );
nor U103854 ( n14504, n73984, n14022 );
nor U103855 ( n26863, n26868, n26869 );
nor U103856 ( n26868, n73700, n26405 );
nor U103857 ( n26869, n73685, n26404 );
nor U103858 ( n60003, n60008, n60009 );
nor U103859 ( n60008, n73699, n59544 );
nor U103860 ( n60009, n73684, n59543 );
nor U103861 ( n68862, n68867, n68868 );
nor U103862 ( n68867, n73698, n68406 );
nor U103863 ( n68868, n73681, n68405 );
nor U103864 ( n34075, n74339, n33639 );
nor U103865 ( n44110, n44113, n43799 );
or U103866 ( n50419, n49989, n73413 );
xnor U103867 ( n11805, n12705, n12783 );
xor U103868 ( n12783, n74989, n76034 );
nor U103869 ( n12739, n12742, n76596 );
nor U103870 ( n12742, n12743, n12744 );
nand U103871 ( n12744, n12745, n12747 );
nand U103872 ( n12743, n12750, n12752 );
not U103873 ( n2117, n39085 );
xnor U103874 ( n36793, n36891, n2040 );
nand U103875 ( n36891, n36892, n36893 );
nand U103876 ( n36892, n76827, n36398 );
nand U103877 ( n36893, n36802, n2035 );
nand U103878 ( n62786, n62828, n62827 );
nor U103879 ( n62828, n76385, n40806 );
nand U103880 ( n37512, n39085, n36633 );
nor U103881 ( n17013, n17014, n73407 );
nor U103882 ( n14428, n74046, n14004 );
nand U103883 ( n14423, n14424, n14425 );
nor U103884 ( n14424, n14429, n14430 );
nor U103885 ( n14425, n14427, n14428 );
nor U103886 ( n14429, n74097, n14010 );
nor U103887 ( n14430, n74084, n14009 );
nor U103888 ( n34077, n34078, n34079 );
nor U103889 ( n34078, n74352, n33646 );
nor U103890 ( n34079, n74344, n33645 );
or U103891 ( n17884, n17028, n73414 );
nand U103892 ( n68456, n68504, n75937 );
nand U103893 ( n26455, n26503, n75938 );
nand U103894 ( n59594, n59642, n75939 );
xnor U103895 ( n36394, n36901, n2040 );
nand U103896 ( n36901, n36902, n36903 );
nand U103897 ( n36902, n76828, n36702 );
nand U103898 ( n36903, n36403, n2035 );
nor U103899 ( n34076, n34080, n34081 );
nor U103900 ( n34080, n74354, n33650 );
nor U103901 ( n34081, n74349, n33649 );
nor U103902 ( n14427, n74072, n14005 );
nor U103903 ( n14340, n74139, n14032 );
nand U103904 ( n14335, n14337, n14338 );
nor U103905 ( n14337, n14342, n14343 );
nor U103906 ( n14338, n14339, n14340 );
nor U103907 ( n14342, n74156, n14038 );
nor U103908 ( n14433, n14434, n14435 );
nor U103909 ( n14434, n74085, n14018 );
nor U103910 ( n14435, n74071, n14017 );
nand U103911 ( n11775, n11777, n11778 );
nand U103912 ( n11777, n76739, n11780 );
nand U103913 ( n11778, n11779, n76729 );
nand U103914 ( n9111, n11750, n11752 );
nor U103915 ( n11752, n11753, n11754 );
nor U103916 ( n11750, n11774, n11775 );
nand U103917 ( n11753, n11764, n11765 );
nor U103918 ( n14343, n74143, n14037 );
nor U103919 ( n63991, n76249, n74449 );
nand U103920 ( n41178, n63986, n63987 );
nor U103921 ( n63987, n63988, n63989 );
nor U103922 ( n63986, n63991, n63992 );
nor U103923 ( n63989, n76245, n74448 );
nor U103924 ( n14432, n14437, n14438 );
nor U103925 ( n14437, n74099, n14023 );
nor U103926 ( n14438, n74089, n14022 );
nor U103927 ( n52038, n49989, n73424 );
nor U103928 ( n32765, n32767, n76896 );
nor U103929 ( n32767, n32768, n32769 );
nand U103930 ( n32769, n32770, n32771 );
nand U103931 ( n32768, n32772, n32773 );
nand U103932 ( n32773, n76773, n31974 );
nor U103933 ( n14339, n74152, n14033 );
nor U103934 ( n14348, n74153, n14044 );
nand U103935 ( n14334, n14344, n14345 );
nor U103936 ( n14344, n14349, n14350 );
nor U103937 ( n14345, n14347, n14348 );
nor U103938 ( n14349, n74164, n14050 );
nor U103939 ( n64343, n64783, n40935 );
nor U103940 ( n65317, n65925, n41059 );
nor U103941 ( n63663, n64194, n41323 );
nor U103942 ( n62827, n63262, n41183 );
nand U103943 ( n63262, n63664, n63663 );
nor U103944 ( n63664, n40972, n41011 );
nand U103945 ( n64194, n64344, n64343 );
nor U103946 ( n64344, n40732, n41119 );
nand U103947 ( n64783, n65318, n65317 );
nor U103948 ( n65318, n41150, n40765 );
nand U103949 ( n65925, n66005, n66004 );
nor U103950 ( n66005, n40869, n40697 );
and U103951 ( n66349, n66727, n552 );
nor U103952 ( n66727, n41369, n41378 );
and U103953 ( n66179, n66350, n66349 );
nor U103954 ( n66350, n41042, n40789 );
and U103955 ( n66004, n66180, n66179 );
nor U103956 ( n66180, n41203, n40989 );
xnor U103957 ( n40797, n41281, n593 );
nand U103958 ( n41281, n41282, n41283 );
nand U103959 ( n41282, n76844, n41284 );
nand U103960 ( n41283, n40806, n41264 );
nor U103961 ( n14350, n74157, n14049 );
nor U103962 ( n33298, n76021, n74460 );
nand U103963 ( n38482, n38483, n38484 );
nand U103964 ( n38484, n76816, n36467 );
nand U103965 ( n38483, n76812, n38485 );
nor U103966 ( n39579, n76415, n74457 );
nand U103967 ( n36797, n39574, n39575 );
nor U103968 ( n39575, n39576, n39577 );
nor U103969 ( n39574, n39579, n39580 );
nor U103970 ( n39577, n76411, n74456 );
nor U103971 ( n14347, n74162, n14045 );
nand U103972 ( n46733, n7535, n74550 );
nand U103973 ( n46770, n46654, n46808 );
nand U103974 ( n46808, n46694, n46692 );
nor U103975 ( n46752, n46754, n76329 );
nor U103976 ( n46754, n46755, n46756 );
nand U103977 ( n46755, n46771, n46772 );
nand U103978 ( n46756, n46757, n46758 );
nor U103979 ( n46761, n46763, n46764 );
nor U103980 ( n46764, n7535, n74550 );
nor U103981 ( n46763, n76005, n46765 );
nor U103982 ( n46765, n75020, n46733 );
and U103983 ( n45855, n46759, n46760 );
nand U103984 ( n46759, n46766, n46767 );
nand U103985 ( n46760, n46761, n46762 );
nand U103986 ( n46767, n76006, n46734 );
nand U103987 ( n67780, n5749, n74574 );
nand U103988 ( n25777, n3992, n74575 );
nand U103989 ( n58915, n6624, n74576 );
nand U103990 ( n67817, n67701, n67855 );
nand U103991 ( n67855, n67741, n67739 );
nand U103992 ( n25814, n25696, n25852 );
nand U103993 ( n25852, n25736, n25734 );
nand U103994 ( n58952, n58836, n58990 );
nand U103995 ( n58990, n58876, n58874 );
nor U103996 ( n67799, n67801, n76869 );
nor U103997 ( n67801, n67802, n67803 );
nand U103998 ( n67802, n67818, n67819 );
nand U103999 ( n67803, n67804, n67805 );
nor U104000 ( n25796, n25798, n76904 );
nor U104001 ( n25798, n25799, n25800 );
nand U104002 ( n25799, n25815, n25816 );
nand U104003 ( n25800, n25801, n25802 );
nor U104004 ( n58934, n58936, n76878 );
nor U104005 ( n58936, n58937, n58938 );
nand U104006 ( n58937, n58953, n58954 );
nand U104007 ( n58938, n58939, n58940 );
nor U104008 ( n67808, n67810, n67811 );
nor U104009 ( n67811, n5749, n74574 );
nor U104010 ( n67810, n75989, n67812 );
nor U104011 ( n67812, n75017, n67780 );
nor U104012 ( n25805, n25807, n25808 );
nor U104013 ( n25808, n3992, n74575 );
nor U104014 ( n25807, n76026, n25809 );
nor U104015 ( n25809, n75018, n25777 );
nor U104016 ( n58943, n58945, n58946 );
nor U104017 ( n58946, n6624, n74576 );
nor U104018 ( n58945, n75997, n58947 );
nor U104019 ( n58947, n75019, n58915 );
and U104020 ( n66806, n67806, n67807 );
nand U104021 ( n67806, n67813, n67814 );
nand U104022 ( n67807, n67808, n67809 );
nand U104023 ( n67814, n75990, n67781 );
and U104024 ( n24928, n25803, n25804 );
nand U104025 ( n25803, n25810, n25811 );
nand U104026 ( n25804, n25805, n25806 );
nand U104027 ( n25811, n76027, n25778 );
and U104028 ( n58065, n58941, n58942 );
nand U104029 ( n58941, n58948, n58949 );
nand U104030 ( n58942, n58943, n58944 );
nand U104031 ( n58949, n75998, n58916 );
xor U104032 ( n38267, n39209, n36907 );
nor U104033 ( n31943, n31950, n31848 );
and U104034 ( n31950, n74973, n31951 );
and U104035 ( n71897, n71327, n71302 );
nand U104036 ( n47284, n47300, n73065 );
nor U104037 ( n63988, n48566, n76242 );
nand U104038 ( n11178, n73060, n73533 );
nand U104039 ( n14629, n11178, n11184 );
not U104040 ( n5157, n10717 );
nand U104041 ( n10724, n5154, n73533 );
nor U104042 ( n51171, n50001, n73424 );
nor U104043 ( n39576, n38332, n76404 );
nor U104044 ( n18401, n17035, n73020 );
nor U104045 ( n14323, n74128, n14004 );
nand U104046 ( n14318, n14319, n14320 );
nor U104047 ( n14319, n14324, n14325 );
nor U104048 ( n14320, n14322, n14323 );
nor U104049 ( n14324, n74154, n14010 );
xnor U104050 ( n45730, n46581, n46612 );
xor U104051 ( n46612, n74881, n76341 );
nor U104052 ( n46603, n46605, n76330 );
nor U104053 ( n46605, n46606, n46607 );
nand U104054 ( n46607, n46608, n46609 );
nand U104055 ( n46606, n46610, n46611 );
nand U104056 ( n68315, n68331, n73066 );
nand U104057 ( n26314, n26330, n73067 );
nand U104058 ( n59453, n59469, n73068 );
not U104059 ( n5152, n10722 );
xnor U104060 ( n66656, n67628, n67659 );
xor U104061 ( n67659, n74916, n76197 );
xnor U104062 ( n24821, n25623, n25654 );
xor U104063 ( n25654, n74917, n76521 );
xnor U104064 ( n57955, n58760, n58794 );
xor U104065 ( n58794, n74918, n76263 );
nor U104066 ( n67650, n67652, n76870 );
nor U104067 ( n67652, n67653, n67654 );
nand U104068 ( n67654, n67655, n67656 );
nand U104069 ( n67653, n67657, n67658 );
nor U104070 ( n25645, n25647, n76905 );
nor U104071 ( n25647, n25648, n25649 );
nand U104072 ( n25649, n25650, n25651 );
nand U104073 ( n25648, n25652, n25653 );
nor U104074 ( n58785, n58787, n76879 );
nor U104075 ( n58787, n58788, n58789 );
nand U104076 ( n58789, n58790, n58791 );
nand U104077 ( n58788, n58792, n58793 );
nand U104078 ( n10714, n14629, n73533 );
nor U104079 ( n14325, n74140, n14009 );
nor U104080 ( n18904, n17035, n75919 );
nand U104081 ( n36396, n36899, n36900 );
nand U104082 ( n36900, n76807, n36702 );
nand U104083 ( n36899, n76827, n36403 );
nor U104084 ( n14322, n74149, n14005 );
nand U104085 ( n41177, n41253, n41254 );
nand U104086 ( n41254, n76848, n40801 );
nand U104087 ( n41253, n76845, n41183 );
nand U104088 ( n39184, n2183, n39260 );
nor U104089 ( n14328, n14329, n14330 );
nor U104090 ( n14329, n74161, n14018 );
nor U104091 ( n14330, n74150, n14017 );
nand U104092 ( n13522, n13588, n13589 );
nor U104093 ( n14327, n14332, n14333 );
nor U104094 ( n14332, n74163, n14023 );
nor U104095 ( n14333, n74155, n14022 );
nand U104096 ( n13588, n76603, n73116 );
nand U104097 ( n71763, n71302, n71096 );
nor U104098 ( n19550, n17028, n73022 );
or U104099 ( n50946, n50001, n73419 );
nand U104100 ( n72108, n71143, n71410 );
nand U104101 ( n46731, n46732, n46655 );
nand U104102 ( n46732, n46733, n76342 );
nor U104103 ( n46714, n46716, n76329 );
nor U104104 ( n46716, n46717, n46718 );
nand U104105 ( n46717, n46735, n46736 );
nand U104106 ( n46718, n46719, n46720 );
nand U104107 ( n46719, n76658, n45815 );
nand U104108 ( n67778, n67779, n67702 );
nand U104109 ( n67779, n67780, n76198 );
nand U104110 ( n25775, n25776, n25697 );
nand U104111 ( n25776, n25777, n76522 );
nand U104112 ( n58913, n58914, n58837 );
nand U104113 ( n58914, n58915, n76264 );
nor U104114 ( n67761, n67763, n76869 );
nor U104115 ( n67763, n67764, n67765 );
nand U104116 ( n67764, n67782, n67783 );
nand U104117 ( n67765, n67766, n67767 );
nor U104118 ( n25758, n25760, n76904 );
nor U104119 ( n25760, n25761, n25762 );
nand U104120 ( n25761, n25779, n25780 );
nand U104121 ( n25762, n25763, n25764 );
nor U104122 ( n58896, n58898, n76878 );
nor U104123 ( n58898, n58899, n58900 );
nand U104124 ( n58899, n58917, n58918 );
nand U104125 ( n58900, n58901, n58902 );
nand U104126 ( n67766, n76706, n66766 );
nand U104127 ( n25763, n76752, n24888 );
nand U104128 ( n58901, n76685, n58025 );
nand U104129 ( n41831, n41836, n41837 );
nand U104130 ( n41837, n41284, n76379 );
nand U104131 ( n41836, n76383, n40806 );
and U104132 ( n41830, n41838, n41839 );
nand U104133 ( n41838, n76383, n41284 );
nand U104134 ( n41839, n40806, n76379 );
nor U104135 ( n51102, n50001, n73019 );
nor U104136 ( n19228, n17028, n73423 );
nor U104137 ( n32840, n32842, n76896 );
nor U104138 ( n32842, n32843, n32844 );
nand U104139 ( n32843, n32868, n32869 );
nand U104140 ( n32844, n32845, n32846 );
nand U104141 ( n32041, n32855, n32856 );
nand U104142 ( n32856, n32817, n32780 );
nor U104143 ( n32855, n32857, n32858 );
nor U104144 ( n32858, n32780, n32825 );
nor U104145 ( n13590, n74476, n76602 );
nor U104146 ( n13518, n13590, n13592 );
and U104147 ( n13592, n13593, n76035 );
nand U104148 ( n13593, n74468, n73116 );
nor U104149 ( n52193, n49989, n73426 );
nand U104150 ( n37424, n37425, n37426 );
nand U104151 ( n37425, n37354, n37353 );
nand U104152 ( n37426, n2139, n37427 );
not U104153 ( n2139, n37413 );
nand U104154 ( n37312, n37313, n37303 );
nand U104155 ( n37313, n37314, n37315 );
nand U104156 ( n37315, n2064, n37302 );
or U104157 ( n37314, n37307, n37297 );
nand U104158 ( n71910, n71327, n71410 );
nand U104159 ( n40800, n41285, n41286 );
nand U104160 ( n41286, n76848, n41284 );
nand U104161 ( n41285, n76844, n40806 );
nor U104162 ( n14243, n74240, n14032 );
nand U104163 ( n14238, n14239, n14240 );
nor U104164 ( n14239, n14244, n14245 );
nor U104165 ( n14240, n14242, n14243 );
nor U104166 ( n14244, n74250, n14038 );
nor U104167 ( n51830, n49989, n73425 );
nor U104168 ( n14245, n74243, n14037 );
nor U104169 ( n38317, n39334, n39441 );
and U104170 ( n39441, n36802, n39442 );
nand U104171 ( n39442, n39443, n1987 );
nor U104172 ( n14242, n74246, n14033 );
nand U104173 ( n31964, n31972, n31973 );
nand U104174 ( n31972, n31953, n74849 );
nand U104175 ( n31973, n76777, n31974 );
nand U104176 ( n4601, n31962, n31963 );
nor U104177 ( n31962, n31980, n31981 );
nor U104178 ( n31963, n31964, n31965 );
nor U104179 ( n31980, n75004, n76783 );
nor U104180 ( n41598, n76387, n41510 );
nor U104181 ( n14250, n74247, n14044 );
nand U104182 ( n14237, n14247, n14248 );
nor U104183 ( n14247, n14252, n14253 );
nor U104184 ( n14248, n14249, n14250 );
nor U104185 ( n14252, n74255, n14050 );
nor U104186 ( n32801, n32803, n76896 );
nor U104187 ( n32803, n32804, n32805 );
nand U104188 ( n32804, n32826, n32827 );
nand U104189 ( n32805, n32806, n32807 );
and U104190 ( n32016, n32814, n32815 );
nand U104191 ( n32814, n32821, n32822 );
nand U104192 ( n32815, n32816, n32776 );
nand U104193 ( n32822, n76022, n74948 );
nand U104194 ( n36398, n39512, n39513 );
nor U104195 ( n39513, n39514, n39515 );
nor U104196 ( n39512, n39517, n39518 );
nor U104197 ( n39515, n76411, n74482 );
nor U104198 ( n39517, n76415, n74483 );
nand U104199 ( n54620, n54621, n54622 );
nand U104200 ( n54622, n569, n40869 );
nand U104201 ( n54621, n76857, n54623 );
nor U104202 ( n14253, n74251, n14049 );
nor U104203 ( n72820, n72824, n72825 );
nor U104204 ( n72821, n72822, n72823 );
nor U104205 ( n72825, n73551, n73026 );
nand U104206 ( n36796, n36867, n36868 );
nand U104207 ( n36868, n76808, n36398 );
nand U104208 ( n36867, n76826, n36802 );
nor U104209 ( n33025, n32947, n33099 );
and U104210 ( n33099, n32984, n32867 );
nor U104211 ( n33005, n33007, n76895 );
nor U104212 ( n33007, n33008, n33009 );
nand U104213 ( n33008, n33027, n33028 );
nand U104214 ( n33009, n33010, n33011 );
nand U104215 ( n33010, n76773, n32120 );
not U104216 ( n2122, n36848 );
nor U104217 ( n72822, n73061, n71105 );
nor U104218 ( n14249, n74253, n14045 );
nor U104219 ( n63676, n76249, n74475 );
nand U104220 ( n40801, n63671, n63672 );
nor U104221 ( n63672, n63673, n63674 );
nor U104222 ( n63671, n63676, n63677 );
nor U104223 ( n63674, n76245, n74474 );
nor U104224 ( n11552, n10237, n11594 );
nand U104225 ( n45852, n45853, n45854 );
nand U104226 ( n45853, n76671, n45856 );
nand U104227 ( n45854, n45855, n76662 );
nand U104228 ( n15791, n45835, n45836 );
nor U104229 ( n45836, n45837, n45838 );
nor U104230 ( n45835, n45851, n45852 );
nand U104231 ( n45838, n45839, n45840 );
nand U104232 ( n66803, n66804, n66805 );
nand U104233 ( n66804, n76719, n66807 );
nand U104234 ( n66805, n66806, n76710 );
nand U104235 ( n24925, n24926, n24927 );
nand U104236 ( n24926, n76767, n24929 );
nand U104237 ( n24927, n24928, n76758 );
nand U104238 ( n58062, n58063, n58064 );
nand U104239 ( n58063, n76700, n58066 );
nand U104240 ( n58064, n58065, n76691 );
nand U104241 ( n11301, n66786, n66787 );
nor U104242 ( n66787, n66788, n66789 );
nor U104243 ( n66786, n66802, n66803 );
nand U104244 ( n66789, n66790, n66791 );
nand U104245 ( n6811, n24908, n24909 );
nor U104246 ( n24909, n24910, n24911 );
nor U104247 ( n24908, n24924, n24925 );
nand U104248 ( n24911, n24912, n24913 );
nand U104249 ( n13546, n58045, n58046 );
nor U104250 ( n58046, n58047, n58048 );
nor U104251 ( n58045, n58061, n58062 );
nand U104252 ( n58048, n58049, n58050 );
nor U104253 ( n11154, n10237, n10785 );
nand U104254 ( n11789, n11803, n11804 );
nand U104255 ( n11803, n11768, n74924 );
nand U104256 ( n11804, n76730, n11805 );
nand U104257 ( n9106, n11787, n11788 );
nor U104258 ( n11787, n11814, n11815 );
nor U104259 ( n11788, n11789, n11790 );
nor U104260 ( n11814, n75238, n76736 );
nor U104261 ( n10233, n10237, n9897 );
nor U104262 ( n72824, n73062, n71108 );
not U104263 ( n289, n45424 );
nor U104264 ( n14128, n74285, n14032 );
nand U104265 ( n14123, n14124, n14125 );
nor U104266 ( n14124, n14129, n14130 );
nor U104267 ( n14125, n14127, n14128 );
nor U104268 ( n14129, n74295, n14038 );
nand U104269 ( n38514, n38515, n38516 );
nand U104270 ( n38516, n76816, n36822 );
nand U104271 ( n38515, n76812, n38517 );
nor U104272 ( n14130, n74297, n14037 );
nand U104273 ( n33513, n33557, n33558 );
nand U104274 ( n33558, n33559, n33560 );
nor U104275 ( n33777, n33780, n33781 );
and U104276 ( n33605, n33698, n33699 );
nand U104277 ( n33699, n33700, n33701 );
nand U104278 ( n39135, n2184, n39085 );
nor U104279 ( n17612, n17028, n73012 );
nor U104280 ( n14225, n74232, n14004 );
nand U104281 ( n14220, n14222, n14223 );
nor U104282 ( n14222, n14227, n14228 );
nor U104283 ( n14223, n14224, n14225 );
nor U104284 ( n14227, n74248, n14010 );
nor U104285 ( n14127, n74290, n14033 );
nand U104286 ( n45721, n45728, n45729 );
nand U104287 ( n45728, n45710, n74740 );
nand U104288 ( n45729, n76662, n45730 );
nand U104289 ( n15811, n45719, n45720 );
nor U104290 ( n45719, n45736, n45737 );
nor U104291 ( n45720, n45721, n45722 );
nor U104292 ( n45736, n75005, n76668 );
nor U104293 ( n50683, n50001, n73017 );
nor U104294 ( n14135, n74288, n14044 );
nand U104295 ( n14122, n14132, n14133 );
nor U104296 ( n14132, n14137, n14138 );
nor U104297 ( n14133, n14134, n14135 );
nor U104298 ( n14137, n74296, n14050 );
nor U104299 ( n14228, n74241, n14009 );
nand U104300 ( n66647, n66654, n66655 );
nand U104301 ( n66654, n66635, n75210 );
nand U104302 ( n66655, n76711, n66656 );
nand U104303 ( n24812, n24819, n24820 );
nand U104304 ( n24819, n24800, n75211 );
nand U104305 ( n24820, n76759, n24821 );
nand U104306 ( n57946, n57953, n57954 );
nand U104307 ( n57953, n57934, n75212 );
nand U104308 ( n57954, n76692, n57955 );
nand U104309 ( n11321, n66645, n66646 );
nor U104310 ( n66645, n66662, n66663 );
nor U104311 ( n66646, n66647, n66648 );
nor U104312 ( n66662, n74993, n76716 );
nand U104313 ( n6831, n24810, n24811 );
nor U104314 ( n24810, n24827, n24828 );
nor U104315 ( n24811, n24812, n24813 );
nor U104316 ( n24827, n74991, n76764 );
nand U104317 ( n13566, n57944, n57945 );
nor U104318 ( n57944, n57961, n57962 );
nor U104319 ( n57945, n57946, n57947 );
nor U104320 ( n57961, n74990, n76697 );
nor U104321 ( n50412, n50001, n73413 );
nor U104322 ( n48570, n548, n63661 );
and U104323 ( n63661, n41011, n63662 );
nand U104324 ( n63662, n63663, n803 );
nor U104325 ( n14138, n74294, n14049 );
nand U104326 ( n16201, n44918, n44919 );
nor U104327 ( n44919, n44920, n44921 );
nor U104328 ( n44918, n44926, n44927 );
nor U104329 ( n44920, n43808, n44923 );
nor U104330 ( n14224, n74244, n14005 );
nor U104331 ( n14230, n14232, n14233 );
nor U104332 ( n14232, n74252, n14018 );
nor U104333 ( n14233, n74245, n14017 );
nor U104334 ( n49492, n49982, n76834 );
nor U104335 ( n38349, n39443, n39570 );
and U104336 ( n39570, n36577, n39571 );
nand U104337 ( n39571, n39572, n1975 );
nor U104338 ( n14134, n74292, n14045 );
nor U104339 ( n32920, n32922, n76895 );
nor U104340 ( n32922, n32923, n32924 );
nand U104341 ( n32923, n32951, n32952 );
nand U104342 ( n32924, n32925, n32926 );
nand U104343 ( n32936, n32901, n32867 );
nor U104344 ( n32937, n32941, n32942 );
nand U104345 ( n32941, n32950, n32904 );
nand U104346 ( n32942, n3148, n32943 );
nand U104347 ( n32950, n3149, n76472 );
nand U104348 ( n32093, n32933, n32934 );
nand U104349 ( n32934, n3162, n32935 );
nor U104350 ( n32933, n32937, n32938 );
not U104351 ( n3162, n32904 );
not U104352 ( n3148, n32940 );
nor U104353 ( n33045, n33047, n76895 );
nor U104354 ( n33047, n33048, n33049 );
nand U104355 ( n33048, n33062, n33063 );
nand U104356 ( n33049, n33050, n33051 );
and U104357 ( n32160, n33052, n33053 );
nand U104358 ( n33052, n33059, n33060 );
nand U104359 ( n33053, n33054, n33026 );
nand U104360 ( n33060, n76022, n33024 );
nor U104361 ( n14229, n14234, n14235 );
nor U104362 ( n14234, n74254, n14023 );
nor U104363 ( n14235, n74249, n14022 );
xnor U104364 ( n11829, n12719, n12804 );
xor U104365 ( n12804, n73279, n76034 );
nor U104366 ( n12790, n12793, n76596 );
nor U104367 ( n12793, n12794, n12795 );
nand U104368 ( n12795, n12797, n12798 );
nand U104369 ( n12794, n12802, n12803 );
not U104370 ( n8235, n50089 );
or U104371 ( n33022, n33024, n33025 );
nor U104372 ( n32938, n76470, n32939 );
nand U104373 ( n32939, n32940, n75050 );
nand U104374 ( n45812, n45813, n45814 );
nand U104375 ( n45813, n45799, n75202 );
nand U104376 ( n45814, n76663, n45815 );
nand U104377 ( n15796, n45809, n45810 );
nor U104378 ( n45809, n45826, n45827 );
nor U104379 ( n45810, n45811, n45812 );
nor U104380 ( n45826, n74958, n76668 );
nand U104381 ( n66763, n66764, n66765 );
nand U104382 ( n66764, n66707, n74687 );
nand U104383 ( n66765, n76711, n66766 );
nand U104384 ( n24885, n24886, n24887 );
nand U104385 ( n24886, n24872, n74689 );
nand U104386 ( n24887, n76759, n24888 );
nand U104387 ( n58022, n58023, n58024 );
nand U104388 ( n58023, n58009, n74690 );
nand U104389 ( n58024, n76692, n58025 );
nand U104390 ( n11306, n66760, n66761 );
nor U104391 ( n66760, n66777, n66778 );
nor U104392 ( n66761, n66762, n66763 );
nor U104393 ( n66777, n74944, n76716 );
nand U104394 ( n6816, n24882, n24883 );
nor U104395 ( n24882, n24899, n24900 );
nor U104396 ( n24883, n24884, n24885 );
nor U104397 ( n24899, n74939, n76764 );
nand U104398 ( n13551, n58019, n58020 );
nor U104399 ( n58019, n58036, n58037 );
nor U104400 ( n58020, n58021, n58022 );
nor U104401 ( n58036, n74938, n76697 );
nor U104402 ( n17183, n17028, n75913 );
nand U104403 ( n41297, n62941, n62942 );
nor U104404 ( n62942, n62943, n62944 );
nor U104405 ( n62941, n62946, n62947 );
nor U104406 ( n62944, n76244, n74499 );
not U104407 ( n2128, n39021 );
nand U104408 ( n38489, n38490, n38491 );
nand U104409 ( n38490, n76816, n36293 );
nand U104410 ( n38491, n1858, n76443 );
not U104411 ( n1858, n38492 );
nand U104412 ( n4591, n32017, n32018 );
nor U104413 ( n32018, n32019, n32020 );
nor U104414 ( n32017, n32036, n32037 );
nand U104415 ( n32019, n32029, n32030 );
nor U104416 ( n18382, n17035, n73420 );
nand U104417 ( n41284, n63263, n63264 );
nor U104418 ( n63264, n63265, n63266 );
nor U104419 ( n63263, n63268, n63269 );
nor U104420 ( n63266, n76245, n74497 );
nor U104421 ( n18858, n17028, n73422 );
nor U104422 ( n46766, n7545, n46768 );
not U104423 ( n7545, n46655 );
nor U104424 ( n46768, n46769, n46770 );
nor U104425 ( n46769, n76005, n74550 );
nor U104426 ( n67813, n5759, n67815 );
not U104427 ( n5759, n67702 );
nor U104428 ( n67815, n67816, n67817 );
nor U104429 ( n67816, n75989, n74574 );
nor U104430 ( n25810, n4002, n25812 );
not U104431 ( n4002, n25697 );
nor U104432 ( n25812, n25813, n25814 );
nor U104433 ( n25813, n76026, n74575 );
nor U104434 ( n58948, n6634, n58950 );
not U104435 ( n6634, n58837 );
nor U104436 ( n58950, n58951, n58952 );
nor U104437 ( n58951, n75997, n74576 );
nor U104438 ( n14110, n74280, n14004 );
nand U104439 ( n14105, n14107, n14108 );
nor U104440 ( n14107, n14112, n14113 );
nor U104441 ( n14108, n14109, n14110 );
nor U104442 ( n14112, n74291, n14010 );
nor U104443 ( n63265, n48331, n76242 );
nor U104444 ( n62943, n48202, n76242 );
nor U104445 ( n14113, n74286, n14009 );
nand U104446 ( n32117, n32118, n32119 );
nand U104447 ( n32118, n32104, n74688 );
nand U104448 ( n32119, n76777, n32120 );
nand U104449 ( n4571, n32114, n32115 );
nor U104450 ( n32114, n32131, n32132 );
nor U104451 ( n32115, n32116, n32117 );
nor U104452 ( n32131, n74945, n76782 );
nor U104453 ( n16885, n73007, n76162 );
nand U104454 ( n36339, n39269, n39270 );
nor U104455 ( n39270, n39271, n39272 );
nor U104456 ( n39269, n39274, n39275 );
nor U104457 ( n39272, n76410, n74523 );
nor U104458 ( n46634, n46636, n76329 );
nor U104459 ( n46636, n46637, n46638 );
nand U104460 ( n46637, n46658, n46659 );
nand U104461 ( n46638, n46639, n46640 );
xnor U104462 ( n45788, n46647, n46648 );
xor U104463 ( n46648, n73159, n76342 );
nand U104464 ( n46647, n46614, n46617 );
nor U104465 ( n67681, n67683, n76869 );
nor U104466 ( n67683, n67684, n67685 );
nand U104467 ( n67684, n67705, n67706 );
nand U104468 ( n67685, n67686, n67687 );
nor U104469 ( n25676, n25678, n76904 );
nor U104470 ( n25678, n25679, n25680 );
nand U104471 ( n25679, n25700, n25701 );
nand U104472 ( n25680, n25681, n25682 );
nor U104473 ( n58816, n58818, n76878 );
nor U104474 ( n58818, n58819, n58820 );
nand U104475 ( n58819, n58840, n58841 );
nand U104476 ( n58820, n58821, n58822 );
xnor U104477 ( n66696, n67694, n67695 );
xor U104478 ( n67695, n74637, n76198 );
nand U104479 ( n67694, n67661, n67664 );
xnor U104480 ( n24861, n25689, n25690 );
xor U104481 ( n25690, n74638, n76522 );
nand U104482 ( n25689, n25656, n25659 );
xnor U104483 ( n57995, n58829, n58830 );
xor U104484 ( n58830, n74639, n76264 );
nand U104485 ( n58829, n58796, n58799 );
nor U104486 ( n14109, n74284, n14005 );
nand U104487 ( n32012, n32013, n32014 );
nand U104488 ( n32014, n3059, n29404 );
nand U104489 ( n32013, n32016, n76776 );
nand U104490 ( n4596, n31986, n31987 );
nor U104491 ( n31987, n31988, n31989 );
nor U104492 ( n31986, n32011, n32012 );
nand U104493 ( n31989, n31990, n31991 );
nand U104494 ( n48113, n76326, n45420 );
nor U104495 ( n14115, n14117, n14118 );
nor U104496 ( n14117, n74287, n14018 );
nor U104497 ( n14118, n74283, n14017 );
nor U104498 ( n14114, n14119, n14120 );
nor U104499 ( n14119, n74293, n14023 );
nor U104500 ( n14120, n74289, n14022 );
not U104501 ( n1398, n50939 );
nor U104502 ( n34121, n74000, n33657 );
nand U104503 ( n34117, n34118, n34119 );
nor U104504 ( n34118, n34123, n34124 );
nor U104505 ( n34119, n34120, n34121 );
nor U104506 ( n34123, n74010, n33662 );
not U104507 ( n3236, n33915 );
nor U104508 ( n34128, n74007, n33667 );
nand U104509 ( n34116, n34125, n34126 );
nor U104510 ( n34125, n34131, n34132 );
nor U104511 ( n34126, n34127, n34128 );
nor U104512 ( n34131, n74018, n33672 );
nor U104513 ( n34120, n74006, n33658 );
nor U104514 ( n34127, n74014, n33668 );
nor U104515 ( n34124, n74002, n33661 );
nor U104516 ( n38380, n39572, n39692 );
and U104517 ( n39692, n36327, n39693 );
nand U104518 ( n39693, n39694, n1967 );
nor U104519 ( n34132, n74011, n33671 );
nand U104520 ( n71774, n71410, n71096 );
nand U104521 ( n37595, n36551, n36848 );
nand U104522 ( n36702, n39445, n39446 );
nor U104523 ( n39446, n39447, n39448 );
nor U104524 ( n39445, n39450, n39451 );
nor U104525 ( n39448, n76411, n74508 );
nor U104526 ( n14030, n74322, n14032 );
nand U104527 ( n14025, n14027, n14028 );
nor U104528 ( n14027, n14034, n14035 );
nor U104529 ( n14028, n14029, n14030 );
nor U104530 ( n14034, n74332, n14038 );
nand U104531 ( n37532, n36305, n36935 );
nor U104532 ( n14035, n74333, n14037 );
xor U104533 ( n45878, n7535, n46807 );
xor U104534 ( n46807, n74550, n76342 );
nor U104535 ( n46792, n46794, n76329 );
nor U104536 ( n46794, n46795, n46796 );
nand U104537 ( n46795, n46809, n46810 );
nand U104538 ( n46796, n46797, n46798 );
xor U104539 ( n66829, n5749, n67854 );
xor U104540 ( n67854, n74574, n76198 );
xor U104541 ( n24953, n3992, n25851 );
xor U104542 ( n25851, n74575, n76522 );
xor U104543 ( n58088, n6624, n58989 );
xor U104544 ( n58989, n74576, n76264 );
nor U104545 ( n67839, n67841, n76869 );
nor U104546 ( n67841, n67842, n67843 );
nand U104547 ( n67842, n67856, n67857 );
nand U104548 ( n67843, n67844, n67845 );
nor U104549 ( n25836, n25838, n76904 );
nor U104550 ( n25838, n25839, n25840 );
nand U104551 ( n25839, n25853, n25854 );
nand U104552 ( n25840, n25841, n25842 );
nor U104553 ( n58974, n58976, n76878 );
nor U104554 ( n58976, n58977, n58978 );
nand U104555 ( n58977, n58991, n58992 );
nand U104556 ( n58978, n58979, n58980 );
nand U104557 ( n9096, n11854, n11855 );
nor U104558 ( n11854, n11883, n11884 );
nor U104559 ( n11855, n11857, n11858 );
nor U104560 ( n11883, n75303, n76736 );
nand U104561 ( n41945, n41946, n41947 );
xor U104562 ( n41946, n76387, n41948 );
xor U104563 ( n41947, n76387, n41510 );
nand U104564 ( n39000, n2188, n36935 );
nor U104565 ( n39271, n38243, n76403 );
nor U104566 ( n14029, n74327, n14033 );
nor U104567 ( n34104, n73987, n33635 );
nand U104568 ( n34100, n34101, n34102 );
nor U104569 ( n34101, n34106, n34107 );
nor U104570 ( n34102, n34103, n34104 );
nor U104571 ( n34106, n74008, n33640 );
nor U104572 ( n14043, n74325, n14044 );
nand U104573 ( n14024, n14039, n14040 );
nor U104574 ( n14039, n14047, n14048 );
nor U104575 ( n14040, n14042, n14043 );
nor U104576 ( n14047, n74334, n14050 );
nor U104577 ( n52047, n50001, n73426 );
nand U104578 ( n38994, n2187, n39021 );
nor U104579 ( n34103, n74003, n33636 );
nor U104580 ( n34107, n74001, n33639 );
nor U104581 ( n14048, n74331, n14049 );
nor U104582 ( n14180, n14184, n14185 );
and U104583 ( n13983, n14082, n14083 );
nand U104584 ( n14083, n14084, n14085 );
nand U104585 ( n13853, n13908, n13909 );
nand U104586 ( n13909, n13910, n13912 );
nand U104587 ( n54751, n54752, n54753 );
or U104588 ( n54752, n54754, n573 );
nand U104589 ( n54753, n76335, n41041 );
nand U104590 ( n1461, n54748, n54749 );
nor U104591 ( n54748, n54758, n54759 );
nor U104592 ( n54749, n54750, n54751 );
nor U104593 ( n54758, n76856, n74217 );
nand U104594 ( n1451, n54862, n54863 );
nor U104595 ( n54862, n54872, n54873 );
nor U104596 ( n54863, n54864, n54865 );
nor U104597 ( n54872, n76856, n73826 );
nor U104598 ( n14042, n74329, n14045 );
nand U104599 ( n1471, n54639, n54640 );
nor U104600 ( n54639, n54650, n54651 );
nor U104601 ( n54640, n54641, n54642 );
nor U104602 ( n54650, n76856, n74281 );
not U104603 ( n2133, n36935 );
nand U104604 ( n1441, n54980, n54981 );
nor U104605 ( n54981, n54982, n54983 );
nor U104606 ( n54980, n54991, n54992 );
and U104607 ( n54982, n41377, n76338 );
nand U104608 ( n1446, n54908, n54909 );
nor U104609 ( n54908, n54918, n54919 );
nor U104610 ( n54909, n54910, n54911 );
nor U104611 ( n54918, n76857, n73827 );
nand U104612 ( n1456, n54807, n54808 );
nor U104613 ( n54807, n54816, n54817 );
nor U104614 ( n54808, n54809, n54810 );
nor U104615 ( n54816, n76856, n73910 );
nand U104616 ( n54809, n54814, n54815 );
nand U104617 ( n54815, n76338, n40984 );
nand U104618 ( n54814, n76335, n75248 );
nand U104619 ( n1466, n54663, n54664 );
nor U104620 ( n54663, n54673, n54674 );
nor U104621 ( n54664, n54665, n54666 );
nor U104622 ( n54673, n76856, n74259 );
nand U104623 ( n38904, n2185, n36848 );
nor U104624 ( n46677, n46679, n76329 );
nor U104625 ( n46679, n46680, n46681 );
nand U104626 ( n46681, n46682, n46683 );
nand U104627 ( n46680, n46684, n46685 );
nand U104628 ( n46689, n46690, n46657 );
nand U104629 ( n46690, n46650, n46692 );
nand U104630 ( n46685, n76658, n45795 );
nor U104631 ( n67724, n67726, n76869 );
nor U104632 ( n67726, n67727, n67728 );
nand U104633 ( n67728, n67729, n67730 );
nand U104634 ( n67727, n67731, n67732 );
nor U104635 ( n25719, n25721, n76904 );
nor U104636 ( n25721, n25722, n25723 );
nand U104637 ( n25723, n25724, n25725 );
nand U104638 ( n25722, n25726, n25727 );
nor U104639 ( n58859, n58861, n76878 );
nor U104640 ( n58861, n58862, n58863 );
nand U104641 ( n58863, n58864, n58865 );
nand U104642 ( n58862, n58866, n58867 );
nand U104643 ( n67736, n67737, n67704 );
nand U104644 ( n67737, n67697, n67739 );
nand U104645 ( n25731, n25732, n25699 );
nand U104646 ( n25732, n25692, n25734 );
nand U104647 ( n58871, n58872, n58839 );
nand U104648 ( n58872, n58832, n58874 );
nand U104649 ( n67732, n76706, n66703 );
nand U104650 ( n25727, n76752, n24868 );
nand U104651 ( n58867, n76685, n58005 );
not U104652 ( n2152, n37354 );
nand U104653 ( n9101, n11822, n11823 );
nor U104654 ( n11822, n11847, n11848 );
nor U104655 ( n11823, n11824, n11825 );
nor U104656 ( n11847, n73392, n76736 );
nand U104657 ( n4581, n32065, n32066 );
nor U104658 ( n32066, n32067, n32068 );
nor U104659 ( n32065, n32088, n32089 );
nand U104660 ( n32068, n32069, n32070 );
nand U104661 ( n32157, n32158, n32159 );
nand U104662 ( n32158, n76785, n32161 );
nand U104663 ( n32159, n32160, n76776 );
nand U104664 ( n4566, n32140, n32141 );
nor U104665 ( n32141, n32142, n32143 );
nor U104666 ( n32140, n32156, n32157 );
nand U104667 ( n32143, n32144, n32145 );
nor U104668 ( n39447, n38294, n76404 );
nor U104669 ( n34109, n34110, n34111 );
nor U104670 ( n34110, n74013, n33646 );
nor U104671 ( n34111, n74004, n33645 );
nor U104672 ( n34108, n34113, n34114 );
nor U104673 ( n34113, n74015, n33650 );
nor U104674 ( n34114, n74009, n33649 );
and U104675 ( n71514, n71098, n71243 );
nand U104676 ( n41090, n62867, n62868 );
nor U104677 ( n62868, n62869, n62870 );
nor U104678 ( n62867, n62872, n62873 );
nor U104679 ( n62870, n76244, n74520 );
not U104680 ( n2145, n36425 );
nand U104681 ( n36512, n39387, n39388 );
nor U104682 ( n39388, n39389, n39390 );
nor U104683 ( n39387, n39392, n39393 );
nor U104684 ( n39390, n76410, n74518 );
nor U104685 ( n32970, n32972, n76895 );
nor U104686 ( n32972, n32973, n32974 );
nand U104687 ( n32974, n32975, n32976 );
nand U104688 ( n32973, n32977, n32978 );
xnor U104689 ( n32100, n32979, n32980 );
xor U104690 ( n32980, n74652, n76471 );
nand U104691 ( n32979, n32981, n32982 );
nor U104692 ( n32981, n3160, n32949 );
nand U104693 ( n71396, n72477, n72478 );
nor U104694 ( n72477, n72481, n72482 );
nor U104695 ( n72478, n72479, n72480 );
nor U104696 ( n72482, n73828, n73026 );
nor U104697 ( n48914, n547, n64341 );
and U104698 ( n64341, n40732, n64342 );
nand U104699 ( n64342, n64343, n799 );
nor U104700 ( n72479, n73821, n71105 );
not U104701 ( n2148, n37600 );
nor U104702 ( n14003, n74319, n14004 );
nand U104703 ( n13998, n13999, n14000 );
nor U104704 ( n13999, n14007, n14008 );
nor U104705 ( n14000, n14002, n14003 );
nor U104706 ( n14007, n74328, n14010 );
nand U104707 ( n37535, n36925, n39021 );
nor U104708 ( n33146, n33148, n76895 );
nor U104709 ( n33148, n33149, n33150 );
nand U104710 ( n33149, n33166, n33167 );
nand U104711 ( n33150, n33151, n33152 );
nand U104712 ( n33157, n33158, n33159 );
nand U104713 ( n33158, n33160, n33161 );
nand U104714 ( n33161, n33162, n32227 );
and U104715 ( n32224, n33177, n33178 );
xor U104716 ( n33178, n74879, n76470 );
nor U104717 ( n33177, n32229, n33179 );
nor U104718 ( n33179, n3152, n74845 );
not U104719 ( n2138, n36446 );
nor U104720 ( n14008, n74323, n14009 );
xor U104721 ( n32183, n33025, n33098 );
xor U104722 ( n33098, n74610, n76471 );
nor U104723 ( n33083, n33085, n76895 );
nor U104724 ( n33085, n33086, n33087 );
nand U104725 ( n33086, n33100, n33101 );
nand U104726 ( n33087, n33088, n33089 );
nor U104727 ( n18206, n17047, n75919 );
nor U104728 ( n14002, n74321, n14005 );
nor U104729 ( n14013, n14014, n14015 );
nor U104730 ( n14014, n74324, n14018 );
nor U104731 ( n14015, n74320, n14017 );
not U104732 ( n36, n11638 );
nor U104733 ( n62869, n40914, n76241 );
nand U104734 ( n33700, n33748, n75940 );
nor U104735 ( n14012, n14019, n14020 );
nor U104736 ( n14019, n74330, n14023 );
nor U104737 ( n14020, n74326, n14022 );
nor U104738 ( n14575, n74362, n14032 );
nand U104739 ( n14570, n14572, n14573 );
nor U104740 ( n14572, n14577, n14578 );
nor U104741 ( n14573, n14574, n14575 );
nor U104742 ( n14577, n74376, n14038 );
nor U104743 ( n39389, n38275, n76404 );
nor U104744 ( n50404, n50089, n73419 );
nor U104745 ( n14578, n74361, n14037 );
nor U104746 ( n37421, n36767, n2169 );
nand U104747 ( n45784, n45785, n45786 );
nand U104748 ( n45786, n7434, n42703 );
nand U104749 ( n45785, n76663, n45788 );
nand U104750 ( n15806, n45760, n45761 );
nor U104751 ( n45761, n45762, n45763 );
nor U104752 ( n45760, n45783, n45784 );
nand U104753 ( n45763, n45764, n45765 );
nand U104754 ( n11316, n66668, n66669 );
nor U104755 ( n66669, n66670, n66671 );
nor U104756 ( n66668, n66691, n66692 );
nand U104757 ( n66671, n66672, n66673 );
nand U104758 ( n6826, n24833, n24834 );
nor U104759 ( n24834, n24835, n24836 );
nor U104760 ( n24833, n24856, n24857 );
nand U104761 ( n24836, n24837, n24838 );
nand U104762 ( n13561, n57967, n57968 );
nor U104763 ( n57968, n57969, n57970 );
nor U104764 ( n57967, n57990, n57991 );
nand U104765 ( n57970, n57971, n57972 );
nor U104766 ( n14574, n74370, n14033 );
nor U104767 ( n72481, n73822, n71108 );
nor U104768 ( n14583, n74368, n14044 );
nand U104769 ( n14569, n14579, n14580 );
nor U104770 ( n14579, n14584, n14585 );
nor U104771 ( n14580, n14582, n14583 );
nor U104772 ( n14584, n74377, n14050 );
nand U104773 ( n36747, n39336, n39337 );
nor U104774 ( n39337, n39338, n39339 );
nor U104775 ( n39336, n39341, n39342 );
nor U104776 ( n39339, n76410, n74544 );
nor U104777 ( n14585, n74375, n14049 );
nand U104778 ( n9466, n11214, n11215 );
nor U104779 ( n11215, n11217, n11218 );
nor U104780 ( n11214, n11224, n11225 );
nor U104781 ( n11217, n9908, n11220 );
nor U104782 ( n14582, n74373, n14045 );
nand U104783 ( n40913, n62734, n62735 );
nor U104784 ( n62735, n62736, n62737 );
nor U104785 ( n62734, n62739, n62740 );
nor U104786 ( n62737, n76244, n74549 );
nand U104787 ( n54651, n54652, n54653 );
nand U104788 ( n54653, n569, n41203 );
nand U104789 ( n54652, n76857, n54654 );
or U104790 ( n50097, n50001, n73412 );
nor U104791 ( n14618, n74016, n14032 );
nand U104792 ( n14613, n14614, n14615 );
nor U104793 ( n14614, n14620, n14622 );
nor U104794 ( n14615, n14617, n14618 );
nor U104795 ( n14620, n74043, n14038 );
not U104796 ( n4969, n14353 );
nor U104797 ( n14627, n74037, n14044 );
nand U104798 ( n14612, n14623, n14624 );
nor U104799 ( n14623, n14630, n14632 );
nor U104800 ( n14624, n14625, n14627 );
nor U104801 ( n14630, n74061, n14050 );
nor U104802 ( n14617, n74035, n14033 );
nand U104803 ( n33167, n33168, n74879 );
nand U104804 ( n33168, n33169, n33143 );
nor U104805 ( n33169, n33175, n33176 );
nor U104806 ( n33175, n3120, n33180 );
nor U104807 ( n14625, n74059, n14045 );
nor U104808 ( n14622, n74019, n14037 );
nor U104809 ( n14632, n74045, n14049 );
nand U104810 ( n54759, n54760, n54761 );
nand U104811 ( n54761, n569, n41042 );
nand U104812 ( n54760, n76857, n54762 );
nor U104813 ( n50678, n50089, n73019 );
xor U104814 ( n45891, n7534, n46836 );
xor U104815 ( n46836, n74524, n76342 );
nor U104816 ( n46827, n46829, n76329 );
nor U104817 ( n46829, n46830, n46831 );
nand U104818 ( n46831, n46832, n46833 );
nand U104819 ( n46830, n46834, n46835 );
xor U104820 ( n66842, n5748, n67883 );
xor U104821 ( n67883, n74546, n76198 );
xor U104822 ( n24966, n3990, n25880 );
xor U104823 ( n25880, n74547, n76522 );
xor U104824 ( n58101, n6623, n59018 );
xor U104825 ( n59018, n74548, n76264 );
nor U104826 ( n67874, n67876, n76869 );
nor U104827 ( n67876, n67877, n67878 );
nand U104828 ( n67878, n67879, n67880 );
nand U104829 ( n67877, n67881, n67882 );
nor U104830 ( n25871, n25873, n76904 );
nor U104831 ( n25873, n25874, n25875 );
nand U104832 ( n25875, n25876, n25877 );
nand U104833 ( n25874, n25878, n25879 );
nor U104834 ( n59009, n59011, n76878 );
nor U104835 ( n59011, n59012, n59013 );
nand U104836 ( n59013, n59014, n59015 );
nand U104837 ( n59012, n59016, n59017 );
nand U104838 ( n46657, n76341, n46691 );
nand U104839 ( n46691, n74550, n73148 );
and U104840 ( n46614, n46652, n46653 );
and U104841 ( n46653, n46654, n46655 );
nor U104842 ( n46652, n46656, n7547 );
nor U104843 ( n46656, n76005, n74585 );
nand U104844 ( n15786, n45857, n45858 );
nor U104845 ( n45858, n45859, n45860 );
nor U104846 ( n45857, n45874, n45875 );
nand U104847 ( n45859, n45868, n45869 );
nand U104848 ( n45875, n45876, n45877 );
nand U104849 ( n45876, n7434, n42808 );
nand U104850 ( n45877, n76663, n45878 );
nand U104851 ( n11296, n66808, n66809 );
nor U104852 ( n66809, n66810, n66811 );
nor U104853 ( n66808, n66825, n66826 );
nand U104854 ( n66810, n66819, n66820 );
nand U104855 ( n66826, n66827, n66828 );
nand U104856 ( n66827, n5660, n63460 );
nand U104857 ( n66828, n76711, n66829 );
nand U104858 ( n6806, n24932, n24933 );
nor U104859 ( n24933, n24934, n24935 );
nor U104860 ( n24932, n24949, n24950 );
nand U104861 ( n24934, n24943, n24944 );
nand U104862 ( n13541, n58067, n58068 );
nor U104863 ( n58068, n58069, n58070 );
nor U104864 ( n58067, n58084, n58085 );
nand U104865 ( n58069, n58078, n58079 );
nand U104866 ( n24950, n24951, n24952 );
nand U104867 ( n24951, n3903, n22240 );
nand U104868 ( n24952, n76759, n24953 );
nand U104869 ( n58085, n58086, n58087 );
nand U104870 ( n58086, n6535, n55352 );
nand U104871 ( n58087, n76692, n58088 );
nor U104872 ( n14597, n74005, n14004 );
nand U104873 ( n14592, n14593, n14594 );
nor U104874 ( n14593, n14599, n14600 );
nor U104875 ( n14594, n14595, n14597 );
nor U104876 ( n14599, n74038, n14010 );
nor U104877 ( n14595, n74026, n14005 );
nor U104878 ( n14600, n74017, n14009 );
nor U104879 ( n39338, n38259, n76403 );
nor U104880 ( n11740, n16861, n76789 );
nand U104881 ( n45792, n45793, n45794 );
nand U104882 ( n45793, n7434, n7955 );
nand U104883 ( n45794, n76663, n45795 );
nand U104884 ( n15801, n45789, n45790 );
nor U104885 ( n45789, n45803, n45804 );
nor U104886 ( n45790, n45791, n45792 );
nor U104887 ( n45803, n73280, n76668 );
nand U104888 ( n66700, n66701, n66702 );
nand U104889 ( n66701, n5660, n63341 );
nand U104890 ( n66702, n76711, n66703 );
nand U104891 ( n24865, n24866, n24867 );
nand U104892 ( n24866, n3903, n22193 );
nand U104893 ( n24867, n76759, n24868 );
nand U104894 ( n58002, n58003, n58004 );
nand U104895 ( n58003, n6535, n55307 );
nand U104896 ( n58004, n76692, n58005 );
nand U104897 ( n11311, n66697, n66698 );
nor U104898 ( n66697, n66711, n66712 );
nor U104899 ( n66698, n66699, n66700 );
nor U104900 ( n66711, n73277, n76716 );
nand U104901 ( n6821, n24862, n24863 );
nor U104902 ( n24862, n24876, n24877 );
nor U104903 ( n24863, n24864, n24865 );
nor U104904 ( n24876, n73276, n76764 );
nand U104905 ( n13556, n57999, n58000 );
nor U104906 ( n57999, n58013, n58014 );
nor U104907 ( n58000, n58001, n58002 );
nor U104908 ( n58013, n73275, n76697 );
nand U104909 ( n67704, n76197, n67738 );
nand U104910 ( n67738, n74574, n73149 );
nand U104911 ( n25699, n76521, n25733 );
nand U104912 ( n25733, n74575, n73150 );
nand U104913 ( n58839, n76263, n58873 );
nand U104914 ( n58873, n74576, n73151 );
and U104915 ( n67661, n67699, n67700 );
and U104916 ( n67700, n67701, n67702 );
nor U104917 ( n67699, n67703, n5760 );
nor U104918 ( n67703, n75989, n74595 );
and U104919 ( n25656, n25694, n25695 );
and U104920 ( n25695, n25696, n25697 );
nor U104921 ( n25694, n25698, n4003 );
nor U104922 ( n25698, n76026, n74596 );
and U104923 ( n58796, n58834, n58835 );
and U104924 ( n58835, n58836, n58837 );
nor U104925 ( n58834, n58838, n6635 );
nor U104926 ( n58838, n75997, n74597 );
nor U104927 ( n62736, n47958, n76241 );
nor U104928 ( n14558, n74357, n14004 );
nand U104929 ( n14553, n14554, n14555 );
nor U104930 ( n14554, n14559, n14560 );
nor U104931 ( n14555, n14557, n14558 );
nor U104932 ( n14559, n74367, n14010 );
not U104933 ( n284, n45420 );
nand U104934 ( n33559, n33575, n73088 );
and U104935 ( n12908, n75785, n75786 );
nand U104936 ( n75785, n11905, n76724 );
nand U104937 ( n75786, n11918, n4848 );
nor U104938 ( n14560, n74359, n14009 );
nand U104939 ( n41134, n62634, n62635 );
nor U104940 ( n62635, n62636, n62637 );
nor U104941 ( n62634, n62639, n62640 );
nor U104942 ( n62637, n76244, n74552 );
nand U104943 ( n32097, n32098, n32099 );
nand U104944 ( n32098, n3059, n29512 );
nand U104945 ( n32099, n76777, n32100 );
nand U104946 ( n4576, n32094, n32095 );
nor U104947 ( n32094, n32108, n32109 );
nor U104948 ( n32095, n32096, n32097 );
nor U104949 ( n32108, n73278, n76782 );
nor U104950 ( n14557, n74364, n14005 );
nor U104951 ( n18391, n17047, n73020 );
nor U104952 ( n14563, n14564, n14565 );
nor U104953 ( n14564, n74365, n14018 );
nor U104954 ( n14565, n74363, n14017 );
nor U104955 ( n14603, n14604, n14605 );
nor U104956 ( n14604, n74052, n14018 );
nor U104957 ( n14605, n74031, n14017 );
nor U104958 ( n14562, n14567, n14568 );
nor U104959 ( n14567, n74374, n14023 );
nor U104960 ( n14568, n74369, n14022 );
nor U104961 ( n14602, n14608, n14609 );
nor U104962 ( n14608, n74060, n14023 );
nor U104963 ( n14609, n74039, n14022 );
nor U104964 ( n18228, n73018, n17035 );
nand U104965 ( n14914, n76592, n11625 );
nand U104966 ( n16196, n44928, n44929 );
nor U104967 ( n44929, n44930, n44931 );
nor U104968 ( n44928, n44937, n44938 );
nor U104969 ( n44930, n44935, n44936 );
nor U104970 ( n32889, n32891, n76896 );
nor U104971 ( n32891, n32892, n32893 );
nand U104972 ( n32893, n32894, n32895 );
nand U104973 ( n32892, n32896, n32897 );
xnor U104974 ( n32053, n32898, n32899 );
xor U104975 ( n32899, n74671, n76471 );
nand U104976 ( n32898, n32861, n32900 );
nand U104977 ( n32900, n3155, n32867 );
nand U104978 ( n72093, n71396, n71143 );
nor U104979 ( n54988, n66752, n67227 );
nor U104980 ( n67227, n41769, n42184 );
nor U104981 ( n46855, n46857, n76329 );
nor U104982 ( n46857, n46858, n46859 );
nand U104983 ( n46858, n46880, n46881 );
nand U104984 ( n46859, n46860, n46861 );
and U104985 ( n45927, n46869, n46870 );
nand U104986 ( n46870, n7537, n74841 );
nor U104987 ( n46869, n46872, n46873 );
nor U104988 ( n46873, n76341, n46874 );
nor U104989 ( n67902, n67904, n76869 );
nor U104990 ( n67904, n67905, n67906 );
nand U104991 ( n67905, n67927, n67928 );
nand U104992 ( n67906, n67907, n67908 );
nor U104993 ( n25899, n25901, n76904 );
nor U104994 ( n25901, n25902, n25903 );
nand U104995 ( n25902, n25924, n25925 );
nand U104996 ( n25903, n25904, n25905 );
nor U104997 ( n59037, n59039, n76878 );
nor U104998 ( n59039, n59040, n59041 );
nand U104999 ( n59040, n59062, n59063 );
nand U105000 ( n59041, n59042, n59043 );
and U105001 ( n66879, n67916, n67917 );
nand U105002 ( n67917, n5750, n74872 );
nor U105003 ( n67916, n67919, n67920 );
nor U105004 ( n67920, n76197, n67921 );
and U105005 ( n25003, n25913, n25914 );
nand U105006 ( n25914, n3993, n74873 );
nor U105007 ( n25913, n25916, n25917 );
nor U105008 ( n25917, n76521, n25918 );
and U105009 ( n58138, n59051, n59052 );
nand U105010 ( n59052, n6625, n74874 );
nor U105011 ( n59051, n59054, n59055 );
nor U105012 ( n59055, n76263, n59056 );
xor U105013 ( n38432, n39821, n36767 );
nor U105014 ( n17736, n17035, n73418 );
nand U105015 ( n54666, n54667, n54668 );
nand U105016 ( n54667, n569, n40989 );
or U105017 ( n54668, n54669, n573 );
nor U105018 ( n17156, n17035, n73414 );
nand U105019 ( n46694, n76006, n74524 );
and U105020 ( n46650, n46693, n46694 );
nand U105021 ( n46693, n76006, n46695 );
nand U105022 ( n32180, n32181, n32182 );
nand U105023 ( n32181, n3059, n29557 );
nand U105024 ( n32182, n76776, n32183 );
nand U105025 ( n4561, n32162, n32163 );
nor U105026 ( n32163, n32164, n32165 );
nor U105027 ( n32162, n32179, n32180 );
nand U105028 ( n32164, n32173, n32174 );
nand U105029 ( n38545, n38546, n38547 );
nand U105030 ( n38547, n76817, n36655 );
nand U105031 ( n38546, n76812, n38548 );
nor U105032 ( n17039, n17035, n73012 );
nand U105033 ( n37507, n36442, n36446 );
xor U105034 ( n36630, n36481, n36845 );
nor U105035 ( n36845, n36846, n36847 );
nor U105036 ( n36847, n2185, n36423 );
nor U105037 ( n36846, n36424, n36848 );
nor U105038 ( n62636, n40748, n76242 );
nand U105039 ( n14084, n14144, n75941 );
nor U105040 ( n51835, n50001, n73425 );
not U105041 ( n3160, n33023 );
nor U105042 ( n49262, n545, n65315 );
and U105043 ( n65315, n41150, n65316 );
nand U105044 ( n65316, n65317, n795 );
and U105045 ( n32903, n32945, n32946 );
nor U105046 ( n32945, n32948, n32949 );
nor U105047 ( n32946, n32947, n3160 );
nor U105048 ( n32948, n76021, n74652 );
and U105049 ( n32861, n32903, n32904 );
nand U105050 ( n48102, n76326, n45416 );
nor U105051 ( n19082, n17035, n73022 );
nor U105052 ( n17464, n17035, n73015 );
nand U105053 ( n25736, n76027, n74547 );
nand U105054 ( n58876, n75998, n74548 );
and U105055 ( n25692, n25735, n25736 );
nand U105056 ( n25735, n76027, n25737 );
and U105057 ( n58832, n58875, n58876 );
nand U105058 ( n58875, n75998, n58877 );
nand U105059 ( n67741, n75990, n74546 );
and U105060 ( n67697, n67740, n67741 );
nand U105061 ( n67740, n75990, n67742 );
nand U105062 ( n11982, n13024, n13025 );
nand U105063 ( n13025, n12969, n12930 );
nor U105064 ( n13024, n13027, n13028 );
nor U105065 ( n13028, n12930, n12979 );
nor U105066 ( n13007, n13009, n76596 );
nor U105067 ( n13009, n13010, n13012 );
nand U105068 ( n13010, n13040, n13042 );
nand U105069 ( n13012, n13013, n13014 );
nand U105070 ( n38521, n38522, n38523 );
nand U105071 ( n38522, n76816, n36594 );
nand U105072 ( n38523, n1854, n76443 );
not U105073 ( n1854, n38524 );
nand U105074 ( n3111, n36768, n36769 );
nor U105075 ( n36768, n36782, n36783 );
nor U105076 ( n36769, n36770, n36771 );
nor U105077 ( n36782, n2159, n76454 );
nand U105078 ( n37480, n37299, n37298 );
nand U105079 ( n54873, n54874, n54875 );
nand U105080 ( n54874, n76857, n54876 );
nand U105081 ( n54875, n569, n41369 );
nand U105082 ( n49371, n569, n40765 );
nand U105083 ( n54628, n569, n40697 );
nand U105084 ( n54911, n54912, n54913 );
or U105085 ( n54913, n573, n54914 );
nand U105086 ( n54912, n569, n41378 );
nand U105087 ( n54810, n54811, n54812 );
or U105088 ( n54812, n54813, n573 );
nand U105089 ( n54811, n569, n40789 );
nand U105090 ( n45883, n45889, n45890 );
nand U105091 ( n45889, n45871, n74772 );
nand U105092 ( n45890, n76663, n45891 );
nand U105093 ( n15781, n45881, n45882 );
nor U105094 ( n45881, n45897, n45898 );
nor U105095 ( n45882, n45883, n45884 );
nor U105096 ( n45897, n74914, n76668 );
nand U105097 ( n66834, n66840, n66841 );
nand U105098 ( n66840, n66822, n75192 );
nand U105099 ( n66841, n76710, n66842 );
nand U105100 ( n24958, n24964, n24965 );
nand U105101 ( n24964, n24946, n75193 );
nand U105102 ( n24965, n76758, n24966 );
nand U105103 ( n58093, n58099, n58100 );
nand U105104 ( n58099, n58081, n75194 );
nand U105105 ( n58100, n76691, n58101 );
nand U105106 ( n11291, n66832, n66833 );
nor U105107 ( n66832, n66848, n66849 );
nor U105108 ( n66833, n66834, n66835 );
nor U105109 ( n66848, n74900, n76716 );
nand U105110 ( n6801, n24956, n24957 );
nor U105111 ( n24956, n24972, n24973 );
nor U105112 ( n24957, n24958, n24959 );
nor U105113 ( n24972, n74899, n76764 );
nand U105114 ( n13536, n58091, n58092 );
nor U105115 ( n58091, n58107, n58108 );
nor U105116 ( n58092, n58093, n58094 );
nor U105117 ( n58107, n74898, n76697 );
nand U105118 ( n54983, n54984, n54985 );
nand U105119 ( n54984, n54988, n45754 );
nand U105120 ( n54985, n54986, n41769 );
nand U105121 ( n54986, n54923, n54915 );
nand U105122 ( n1886, n41151, n41152 );
nor U105123 ( n41151, n41165, n41166 );
nor U105124 ( n41152, n41153, n41154 );
nor U105125 ( n41165, n635, n76108 );
nor U105126 ( n49552, n49989, n76834 );
nor U105127 ( n38602, n40282, n40337 );
nor U105128 ( n40337, n37764, n37288 );
nand U105129 ( n71924, n71327, n71396 );
nor U105130 ( n12957, n12959, n76596 );
nor U105131 ( n12959, n12960, n12962 );
nand U105132 ( n12960, n12980, n12982 );
nand U105133 ( n12962, n12963, n12964 );
and U105134 ( n11952, n12965, n12967 );
nand U105135 ( n12967, n12968, n12925 );
nand U105136 ( n12965, n12974, n12975 );
nor U105137 ( n12968, n12972, n12973 );
xnor U105138 ( n32196, n32867, n33127 );
xor U105139 ( n33127, n74635, n76471 );
nor U105140 ( n33118, n33120, n76895 );
nor U105141 ( n33120, n33121, n33122 );
nand U105142 ( n33122, n33123, n33124 );
nand U105143 ( n33121, n33125, n33126 );
nor U105144 ( n50087, n50089, n73017 );
nand U105145 ( n38838, n2189, n36446 );
not U105146 ( n1262, n51848 );
and U105147 ( n32949, n76472, n32986 );
nand U105148 ( n32986, n74610, n73167 );
nand U105149 ( n33151, n33165, n33160 );
not U105150 ( n1327, n51121 );
nor U105151 ( n18215, n17047, n73022 );
xnor U105152 ( n36929, n36481, n36932 );
nor U105153 ( n36932, n36933, n36934 );
nor U105154 ( n36934, n2188, n36423 );
nor U105155 ( n36933, n36424, n36935 );
nand U105156 ( n13910, n13930, n73090 );
nor U105157 ( n37753, n36684, n37757 );
nand U105158 ( n37757, n2197, n37080 );
nand U105159 ( n37717, n37751, n37752 );
nor U105160 ( n37751, n37777, n76449 );
nor U105161 ( n37752, n37753, n37754 );
and U105162 ( n37777, n37779, n37708 );
nand U105163 ( n37749, n37750, n37717 );
nand U105164 ( n37750, n2079, n37780 );
xnor U105165 ( n37780, n37781, n37782 );
xor U105166 ( n37782, n74220, n37783 );
nand U105167 ( n37715, n37716, n37717 );
nand U105168 ( n37716, n2079, n37718 );
xnor U105169 ( n37718, n37719, n37720 );
xor U105170 ( n37720, n73896, n37721 );
nand U105171 ( n2901, n37746, n37747 );
nor U105172 ( n37746, n36650, n37787 );
nor U105173 ( n37747, n37748, n37749 );
nand U105174 ( n37787, n37788, n37789 );
nand U105175 ( n2911, n37712, n37713 );
nor U105176 ( n37712, n37725, n37726 );
nor U105177 ( n37713, n37714, n37715 );
nor U105178 ( n37725, P4_STATE_REG, n73895 );
nand U105179 ( n36633, n39211, n39212 );
nor U105180 ( n39212, n39213, n39214 );
nor U105181 ( n39211, n39216, n39217 );
nor U105182 ( n39214, n76410, n74598 );
nand U105183 ( n4586, n32042, n32043 );
nor U105184 ( n32042, n32059, n32060 );
nor U105185 ( n32043, n32044, n32045 );
nor U105186 ( n32059, n74994, n76782 );
nand U105187 ( n32044, n32051, n32052 );
nand U105188 ( n32051, n32032, n75209 );
nand U105189 ( n32052, n76777, n32053 );
nand U105190 ( n38771, n2190, n36425 );
and U105191 ( n71171, n72298, n72299 );
nor U105192 ( n72298, n72302, n72303 );
nor U105193 ( n72299, n72300, n72301 );
nor U105194 ( n72303, n74041, n73026 );
nor U105195 ( n72300, n73063, n71105 );
nor U105196 ( n37348, n37349, n37350 );
nand U105197 ( n37349, n37355, n37356 );
nand U105198 ( n37350, n37351, n37352 );
xor U105199 ( n37351, n37353, n37354 );
nand U105200 ( n15776, n45903, n45904 );
nor U105201 ( n45904, n45905, n45906 );
nor U105202 ( n45903, n45923, n45924 );
nand U105203 ( n45905, n45915, n45916 );
nand U105204 ( n1961, n40870, n40871 );
nor U105205 ( n40870, n40882, n40883 );
nor U105206 ( n40871, n40872, n40873 );
nor U105207 ( n40882, n628, n76114 );
nand U105208 ( n11286, n66854, n66855 );
nor U105209 ( n66855, n66856, n66857 );
nor U105210 ( n66854, n66874, n66875 );
nand U105211 ( n66856, n66866, n66867 );
nand U105212 ( n6796, n24978, n24979 );
nor U105213 ( n24979, n24980, n24981 );
nor U105214 ( n24978, n24998, n24999 );
nand U105215 ( n24980, n24990, n24991 );
nand U105216 ( n13531, n58113, n58114 );
nor U105217 ( n58114, n58115, n58116 );
nor U105218 ( n58113, n58133, n58134 );
nand U105219 ( n58115, n58125, n58126 );
xor U105220 ( n38464, n39922, n36672 );
nor U105221 ( n13248, n13140, n13338 );
and U105222 ( n13338, n13195, n13039 );
nor U105223 ( n13223, n13225, n76595 );
nor U105224 ( n13225, n13227, n13228 );
nand U105225 ( n13227, n13250, n13252 );
nand U105226 ( n13228, n13229, n13230 );
nand U105227 ( n13229, n76725, n12080 );
nand U105228 ( n71510, n71098, n71302 );
nor U105229 ( n13128, n13133, n13134 );
nand U105230 ( n13133, n13144, n13087 );
nand U105231 ( n13134, n4888, n13135 );
nand U105232 ( n13144, n4889, n76606 );
nor U105233 ( n13107, n13109, n76595 );
nor U105234 ( n13109, n13110, n13112 );
nand U105235 ( n13110, n13145, n13147 );
nand U105236 ( n13112, n13113, n13114 );
nand U105237 ( n13127, n13083, n13039 );
nand U105238 ( n12047, n13123, n13124 );
nand U105239 ( n13124, n4899, n13125 );
nor U105240 ( n13123, n13128, n13129 );
not U105241 ( n4899, n13087 );
not U105242 ( n4888, n13132 );
not U105243 ( n8239, n50395 );
nor U105244 ( n38773, n36425, n2190 );
nor U105245 ( n39213, n38227, n76404 );
nand U105246 ( n38575, n38576, n38577 );
nand U105247 ( n38577, n76817, n37007 );
nand U105248 ( n38576, n76812, n38578 );
nand U105249 ( n2676, n38564, n38565 );
nor U105250 ( n38565, n38566, n38567 );
nor U105251 ( n38564, n38574, n38575 );
nand U105252 ( n38567, n38568, n38569 );
nand U105253 ( n11893, n11903, n11904 );
nand U105254 ( n11903, n11882, n75207 );
nand U105255 ( n11904, n76729, n11905 );
nand U105256 ( n9091, n11890, n11892 );
nor U105257 ( n11890, n11913, n11914 );
nor U105258 ( n11892, n11893, n11894 );
nor U105259 ( n11913, n75015, n76736 );
nor U105260 ( n72302, n73064, n71108 );
nor U105261 ( n19238, n17035, n73423 );
xnor U105262 ( n41071, n42275, n41383 );
xor U105263 ( n42275, n593, n41382 );
nor U105264 ( n42270, n41071, n42274 );
nand U105265 ( n42274, n814, n41449 );
nand U105266 ( n42266, n42267, n42225 );
nand U105267 ( n42267, n577, n42295 );
nand U105268 ( n42295, n42296, n42297 );
nand U105269 ( n42296, n42300, n42301 );
nand U105270 ( n42223, n42224, n42225 );
nand U105271 ( n42224, n577, n42226 );
xnor U105272 ( n42226, n42227, n42228 );
xor U105273 ( n42228, n73826, n42229 );
nand U105274 ( n42225, n42268, n42269 );
nor U105275 ( n42268, n42292, n76374 );
nor U105276 ( n42269, n42270, n42271 );
and U105277 ( n42292, n42294, n42209 );
nand U105278 ( n1676, n42263, n42264 );
nor U105279 ( n42263, n41037, n42312 );
nor U105280 ( n42264, n42265, n42266 );
nand U105281 ( n42312, n42313, n42314 );
nand U105282 ( n1686, n42220, n42221 );
nor U105283 ( n42220, n42233, n42234 );
nor U105284 ( n42221, n42222, n42223 );
nor U105285 ( n42233, P3_STATE_REG, n73833 );
not U105286 ( n32, n11625 );
nand U105287 ( n11977, n11978, n11979 );
nand U105288 ( n11979, n4790, n8573 );
nand U105289 ( n11978, n76729, n11982 );
nand U105290 ( n9081, n11954, n11955 );
nor U105291 ( n11955, n11957, n11958 );
nor U105292 ( n11954, n11975, n11977 );
nand U105293 ( n11958, n11959, n11960 );
or U105294 ( n17988, n17047, n73018 );
nand U105295 ( n46874, n7900, n46875 );
nand U105296 ( n67921, n6112, n67922 );
nand U105297 ( n25918, n4334, n25919 );
nand U105298 ( n59056, n6967, n59057 );
xnor U105299 ( n66105, n40697, n654 );
xor U105300 ( n37360, n36618, n36797 );
nor U105301 ( n54991, n76856, n73633 );
nor U105302 ( n49376, n76856, n74381 );
nor U105303 ( n49030, n76855, n74401 );
nor U105304 ( n49573, n76856, n74384 );
nor U105305 ( n49141, n76856, n74396 );
nor U105306 ( n54633, n76856, n74336 );
nor U105307 ( n48571, n76855, n74448 );
nor U105308 ( n37347, n37357, n37358 );
nand U105309 ( n37357, n37361, n37362 );
or U105310 ( n37358, n37359, n37360 );
xor U105311 ( n37362, n37299, n37298 );
nor U105312 ( n48680, n76855, n74415 );
nor U105313 ( n48916, n76855, n74428 );
nor U105314 ( n48454, n76855, n74474 );
nor U105315 ( n54619, n76856, n74382 );
nor U105316 ( n49264, n76856, n74378 );
nor U105317 ( n48799, n76855, n74407 );
nor U105318 ( n48332, n76855, n74497 );
nor U105319 ( n48205, n76855, n74499 );
nor U105320 ( n47961, n76855, n74549 );
nor U105321 ( n46552, n76855, n74714 );
nor U105322 ( n45755, n76855, n74809 );
xnor U105323 ( n66291, n40989, n648 );
nor U105324 ( n54617, n544, n66002 );
and U105325 ( n66002, n40869, n66003 );
nand U105326 ( n66003, n66004, n792 );
nor U105327 ( n13129, n76034, n13130 );
nand U105328 ( n13130, n13132, n74920 );
nand U105329 ( n66435, n41369, n40784 );
nor U105330 ( n13272, n13274, n76595 );
nor U105331 ( n13274, n13275, n13277 );
nand U105332 ( n13275, n13293, n13294 );
nand U105333 ( n13277, n13278, n13279 );
and U105334 ( n12135, n13280, n13282 );
nand U105335 ( n13282, n13283, n13249 );
nand U105336 ( n13280, n13289, n13290 );
nor U105337 ( n13283, n13287, n13288 );
nand U105338 ( n9461, n11227, n11228 );
nor U105339 ( n11228, n11229, n11230 );
nor U105340 ( n11227, n11238, n11239 );
nor U105341 ( n11229, n11235, n11237 );
nor U105342 ( n18874, n17035, n73422 );
nand U105343 ( n38537, n38538, n38539 );
nand U105344 ( n38539, n76446, n36654 );
nand U105345 ( n38538, n38540, n76444 );
xnor U105346 ( n63695, n41011, n714 );
nand U105347 ( n3186, n36468, n36469 );
nor U105348 ( n36468, n36490, n36491 );
nor U105349 ( n36469, n36470, n36471 );
nor U105350 ( n36490, n2158, n76455 );
or U105351 ( n13244, n13247, n13248 );
nand U105352 ( n32188, n32194, n32195 );
nand U105353 ( n32194, n32176, n75191 );
nand U105354 ( n32195, n76776, n32196 );
nand U105355 ( n4556, n32186, n32187 );
nor U105356 ( n32186, n32202, n32203 );
nor U105357 ( n32187, n32188, n32189 );
nor U105358 ( n32202, n74901, n76782 );
nand U105359 ( n11948, n11949, n11950 );
nand U105360 ( n11949, n76738, n11953 );
nand U105361 ( n11950, n11952, n76729 );
nand U105362 ( n9086, n11920, n11922 );
nor U105363 ( n11922, n11923, n11924 );
nor U105364 ( n11920, n11947, n11948 );
nand U105365 ( n11923, n11930, n11932 );
not U105366 ( n278, n45416 );
nor U105367 ( n49988, n73410, n49989 );
nand U105368 ( n40747, n62541, n62542 );
nor U105369 ( n62542, n62543, n62544 );
nor U105370 ( n62541, n62546, n62547 );
nor U105371 ( n62544, n76244, n74645 );
nor U105372 ( n18145, n17047, n73420 );
xnor U105373 ( n37359, n36293, n2164 );
nor U105374 ( n13140, n74599, n76603 );
and U105375 ( n13085, n13138, n13139 );
nor U105376 ( n13138, n13142, n13143 );
nor U105377 ( n13139, n13140, n4898 );
nor U105378 ( n13142, n76602, n74625 );
and U105379 ( n13032, n13085, n13087 );
nor U105380 ( n32223, n32224, n32225 );
nor U105381 ( n32225, n76470, n32226 );
nand U105382 ( n32226, n3497, n32227 );
nand U105383 ( n4551, n32208, n32209 );
nor U105384 ( n32208, n32233, n32234 );
nor U105385 ( n32209, n32210, n32211 );
nor U105386 ( n32233, n74885, n76782 );
nand U105387 ( n42192, n577, n73633 );
nand U105388 ( n1696, n42185, n42186 );
nor U105389 ( n42185, n42199, n42200 );
nor U105390 ( n42186, n42187, n42188 );
nor U105391 ( n42200, P3_STATE_REG, n73637 );
nand U105392 ( n14900, n76592, n11620 );
xor U105393 ( n45935, n7538, n46910 );
xor U105394 ( n46910, n73118, n76342 );
nor U105395 ( n46901, n46903, n76329 );
nor U105396 ( n46903, n46904, n46905 );
nand U105397 ( n46905, n46906, n46907 );
nand U105398 ( n46904, n46908, n46909 );
xor U105399 ( n66886, n5752, n67957 );
xor U105400 ( n67957, n73130, n76198 );
xor U105401 ( n25010, n3994, n25954 );
xor U105402 ( n25954, n73131, n76522 );
xor U105403 ( n58145, n6627, n59092 );
xor U105404 ( n59092, n73132, n76264 );
nor U105405 ( n67948, n67950, n76869 );
nor U105406 ( n67950, n67951, n67952 );
nand U105407 ( n67952, n67953, n67954 );
nand U105408 ( n67951, n67955, n67956 );
nor U105409 ( n25945, n25947, n76904 );
nor U105410 ( n25947, n25948, n25949 );
nand U105411 ( n25949, n25950, n25951 );
nand U105412 ( n25948, n25952, n25953 );
nor U105413 ( n59083, n59085, n76878 );
nor U105414 ( n59085, n59086, n59087 );
nand U105415 ( n59087, n59088, n59089 );
nand U105416 ( n59086, n59090, n59091 );
nand U105417 ( n13195, n76603, n74599 );
nand U105418 ( n13035, n13083, n13084 );
nand U105419 ( n13084, n76603, n13052 );
and U105420 ( n13083, n13194, n13195 );
nand U105421 ( n13194, n76603, n13197 );
nor U105422 ( n38512, n1889, n40087 );
and U105423 ( n40087, n36822, n40088 );
nand U105424 ( n40088, n40089, n1925 );
nor U105425 ( n13287, n13248, n74586 );
nand U105426 ( n71790, n71396, n71096 );
nor U105427 ( n32947, n74635, n76021 );
nor U105428 ( n42007, n42009, n42010 );
nor U105429 ( n42010, n624, n41769 );
and U105430 ( n42009, n42011, n838 );
nand U105431 ( n38552, n38553, n38554 );
nand U105432 ( n38553, n76817, n36386 );
nand U105433 ( n38554, n1853, n76444 );
not U105434 ( n1853, n38555 );
xnor U105435 ( n37361, n37600, n2192 );
nand U105436 ( n12077, n12078, n12079 );
nand U105437 ( n12078, n12060, n75201 );
nand U105438 ( n12079, n76729, n12080 );
nand U105439 ( n9061, n12073, n12074 );
nor U105440 ( n12073, n12094, n12095 );
nor U105441 ( n12074, n12075, n12077 );
nor U105442 ( n12094, n74959, n76735 );
nor U105443 ( n62543, n46937, n76241 );
nor U105444 ( n49596, n50001, n76834 );
nand U105445 ( n32984, n76022, n74635 );
nand U105446 ( n32864, n32901, n32902 );
nand U105447 ( n32902, n76022, n32878 );
and U105448 ( n32901, n32983, n32984 );
nand U105449 ( n32983, n76022, n32985 );
nor U105450 ( n17457, n17047, n73015 );
nor U105451 ( n49756, n50089, n73413 );
nor U105452 ( n37520, n37298, n37598 );
not U105453 ( n8218, n17052 );
nand U105454 ( n12042, n12043, n12044 );
nand U105455 ( n12044, n4790, n8637 );
nand U105456 ( n12043, n76729, n12047 );
nand U105457 ( n9071, n12012, n12013 );
nor U105458 ( n12013, n12014, n12015 );
nor U105459 ( n12012, n12040, n12042 );
nand U105460 ( n12015, n12017, n12018 );
nand U105461 ( n42314, n574, n42299 );
xor U105462 ( n36301, n2040, n36443 );
nor U105463 ( n36443, n36444, n36445 );
nor U105464 ( n36445, n2189, n36423 );
nor U105465 ( n36444, n36424, n36446 );
nand U105466 ( n36551, n39146, n39147 );
nor U105467 ( n39147, n39148, n39149 );
nor U105468 ( n39146, n39151, n39152 );
nor U105469 ( n39149, n76410, n74692 );
or U105470 ( n17728, n17047, n73418 );
nor U105471 ( n54649, n66004, n66177 );
and U105472 ( n66177, n41203, n66178 );
nand U105473 ( n66178, n66179, n789 );
nor U105474 ( n16500, n17028, n76789 );
nand U105475 ( n48091, n76326, n45412 );
nor U105476 ( n33192, n33194, n76895 );
nor U105477 ( n33194, n33195, n33196 );
nand U105478 ( n33196, n33197, n33198 );
nand U105479 ( n33195, n33199, n33200 );
nand U105480 ( n33200, n76773, n32247 );
nor U105481 ( n37479, n37295, n37600 );
nand U105482 ( n37688, n2079, n73798 );
nand U105483 ( n2921, n37681, n37682 );
nor U105484 ( n37681, n37695, n37696 );
nor U105485 ( n37682, n37683, n37684 );
nor U105486 ( n37696, n76920, n73800 );
nand U105487 ( n40402, n40440, n40441 );
nand U105488 ( n40441, n40442, n74634 );
nor U105489 ( n40440, n40437, n40443 );
nor U105490 ( n40443, n74634, n40444 );
nand U105491 ( n38729, n40363, n40364 );
nor U105492 ( n40363, n40382, n40383 );
nor U105493 ( n40364, n40365, n40366 );
nand U105494 ( n40382, n40392, n40393 );
nand U105495 ( n40366, n40367, n40368 );
nand U105496 ( n40367, n2093, n40372 );
nand U105497 ( n40368, n2093, n40369 );
nand U105498 ( n40372, n40373, n40374 );
and U105499 ( n38613, n37113, n2092 );
nand U105500 ( n38119, n2087, n38610 );
nand U105501 ( n38610, n38611, n37110 );
nand U105502 ( n38611, n38612, n38613 );
nor U105503 ( n38612, n37114, n37089 );
nand U105504 ( n40383, n40384, n40385 );
nand U105505 ( n40384, n2093, n40389 );
nand U105506 ( n40385, n2093, n40386 );
nand U105507 ( n40389, n40390, n40391 );
and U105508 ( n44850, n44857, n574 );
and U105509 ( n45065, n45077, n574 );
and U105510 ( n42666, n42678, n574 );
and U105511 ( n42327, n42344, n574 );
nand U105512 ( n1611, n45063, n45064 );
nor U105513 ( n45063, n45086, n41007 );
nor U105514 ( n45064, n45065, n45066 );
nor U105515 ( n45086, n587, n74489 );
nand U105516 ( n1621, n44848, n44849 );
nor U105517 ( n44848, n44861, n41450 );
nor U105518 ( n44849, n44850, n44851 );
nor U105519 ( n44861, n587, n74441 );
nand U105520 ( n1661, n42664, n42665 );
nor U105521 ( n42664, n42687, n40692 );
nor U105522 ( n42665, n42666, n42667 );
nor U105523 ( n42687, n587, n73531 );
nand U105524 ( n1671, n42325, n42326 );
nor U105525 ( n42325, n42358, n40985 );
nor U105526 ( n42326, n42327, n42328 );
nor U105527 ( n42358, n587, n73501 );
xnor U105528 ( n12055, n13189, n13190 );
xor U105529 ( n13190, n74625, n76034 );
nand U105530 ( n13189, n13192, n13193 );
nor U105531 ( n13192, n4898, n13143 );
nor U105532 ( n13178, n13180, n76595 );
nor U105533 ( n13180, n13182, n13183 );
nand U105534 ( n13183, n13184, n13185 );
nand U105535 ( n13182, n13187, n13188 );
nand U105536 ( n2671, n38579, n38580 );
nor U105537 ( n38580, n38581, n38582 );
nor U105538 ( n38579, n38588, n38589 );
nand U105539 ( n38581, n38586, n38587 );
nand U105540 ( n38359, n76816, n36955 );
nand U105541 ( n12132, n12133, n12134 );
nand U105542 ( n12133, n76738, n12137 );
nand U105543 ( n12134, n12135, n76729 );
nand U105544 ( n38422, n76816, n36767 );
nand U105545 ( n38454, n76816, n36672 );
nand U105546 ( n9056, n12110, n12112 );
nor U105547 ( n12112, n12113, n12114 );
nor U105548 ( n12110, n12130, n12132 );
nand U105549 ( n12114, n12115, n12117 );
nand U105550 ( n40365, n40375, n40376 );
nand U105551 ( n40375, n2093, n40380 );
nand U105552 ( n40376, n2093, n40377 );
nand U105553 ( n40380, n40381, n74742 );
not U105554 ( n2149, n37298 );
nor U105555 ( n32222, n32228, n31848 );
and U105556 ( n32228, n74879, n32229 );
not U105557 ( n2518, n17981 );
nand U105558 ( n37136, n37298, n37297 );
nor U105559 ( n47043, n47022, n47044 );
nor U105560 ( n47044, n76005, n47045 );
nor U105561 ( n47045, n73099, n47046 );
nor U105562 ( n47031, n47033, n76329 );
nor U105563 ( n47033, n47034, n47035 );
nand U105564 ( n47035, n47036, n47037 );
nand U105565 ( n47034, n47038, n47039 );
nand U105566 ( n47039, n76658, n46024 );
nor U105567 ( n68074, n68057, n68075 );
nor U105568 ( n68075, n75989, n68076 );
nor U105569 ( n68076, n73104, n68077 );
nor U105570 ( n26071, n26054, n26072 );
nor U105571 ( n26072, n76026, n26073 );
nor U105572 ( n26073, n73105, n26074 );
nor U105573 ( n59212, n59195, n59213 );
nor U105574 ( n59213, n75997, n59214 );
nor U105575 ( n59214, n73106, n59215 );
nor U105576 ( n68062, n68064, n76869 );
nor U105577 ( n68064, n68065, n68066 );
nand U105578 ( n68066, n68067, n68068 );
nand U105579 ( n68065, n68069, n68070 );
nor U105580 ( n26059, n26061, n76904 );
nor U105581 ( n26061, n26062, n26063 );
nand U105582 ( n26063, n26064, n26065 );
nand U105583 ( n26062, n26066, n26067 );
nor U105584 ( n59200, n59202, n76878 );
nor U105585 ( n59202, n59203, n59204 );
nand U105586 ( n59204, n59205, n59206 );
nand U105587 ( n59203, n59207, n59208 );
nand U105588 ( n68070, n76705, n66964 );
nand U105589 ( n26067, n76751, n25088 );
nand U105590 ( n59208, n76684, n58223 );
nand U105591 ( n38582, n38583, n38584 );
nand U105592 ( n38584, n76444, n38585 );
nand U105593 ( n38583, n76817, n37022 );
nor U105594 ( n39148, n38211, n76403 );
nor U105595 ( n50327, n50395, n73019 );
nand U105596 ( n43850, n43851, n43852 );
nand U105597 ( n43852, n43853, n577 );
nand U105598 ( n43851, n43867, n575 );
nor U105599 ( n43853, n43854, n43855 );
nand U105600 ( n43425, n43426, n43427 );
nand U105601 ( n43427, n43428, n577 );
nand U105602 ( n43426, n43441, n575 );
nor U105603 ( n43428, n43429, n43430 );
nand U105604 ( n1631, n43847, n43848 );
nor U105605 ( n43847, n43881, n41115 );
nor U105606 ( n43848, n43849, n43850 );
nor U105607 ( n43881, n587, n74389 );
nand U105608 ( n1646, n43422, n43423 );
nor U105609 ( n43422, n43454, n40761 );
nor U105610 ( n43423, n43424, n43425 );
nor U105611 ( n43454, n587, n74041 );
nor U105612 ( n50665, n50395, n73021 );
nand U105613 ( n43660, n43661, n43662 );
nand U105614 ( n43662, n577, n43663 );
nand U105615 ( n43661, n575, n43667 );
xor U105616 ( n43663, n43664, n43665 );
nand U105617 ( n43553, n43554, n43555 );
nand U105618 ( n43555, n577, n43556 );
nand U105619 ( n43554, n575, n43560 );
xor U105620 ( n43556, n43557, n43558 );
nand U105621 ( n45000, n45001, n45002 );
nand U105622 ( n45002, n577, n45003 );
nand U105623 ( n45001, n575, n45012 );
nand U105624 ( n45003, n45004, n45005 );
nand U105625 ( n43224, n43225, n43226 );
nand U105626 ( n43226, n577, n43227 );
nand U105627 ( n43225, n575, n43231 );
xor U105628 ( n43227, n43228, n43229 );
nand U105629 ( n42951, n42952, n42953 );
nand U105630 ( n42953, n577, n42954 );
nand U105631 ( n42952, n575, n42958 );
xor U105632 ( n42954, n42955, n42956 );
nand U105633 ( n42205, n42206, n42207 );
nand U105634 ( n42207, n577, n42208 );
nand U105635 ( n42206, n575, n42213 );
xnor U105636 ( n42208, n42209, n42210 );
nand U105637 ( n1636, n43657, n43658 );
nor U105638 ( n43657, n43670, n40931 );
nor U105639 ( n43658, n43659, n43660 );
nor U105640 ( n43670, n587, n74346 );
nand U105641 ( n1641, n43550, n43551 );
nor U105642 ( n43550, n43562, n41146 );
nor U105643 ( n43551, n43552, n43553 );
nor U105644 ( n43562, n587, n74279 );
nand U105645 ( n1606, n45132, n45133 );
nor U105646 ( n45132, n45271, n41179 );
nor U105647 ( n45133, n45134, n45135 );
nor U105648 ( n45271, n587, n74496 );
nand U105649 ( n1616, n44997, n44998 );
nor U105650 ( n44997, n45020, n40968 );
nor U105651 ( n44998, n44999, n45000 );
nor U105652 ( n45020, n587, n74447 );
nand U105653 ( n1626, n44383, n44384 );
nor U105654 ( n44383, n44396, n40728 );
nor U105655 ( n44384, n44385, n44386 );
nor U105656 ( n44396, n587, n74405 );
nand U105657 ( n1651, n43221, n43222 );
nor U105658 ( n43221, n43234, n41055 );
nor U105659 ( n43222, n43223, n43224 );
nor U105660 ( n43234, n587, n73828 );
nand U105661 ( n1656, n42948, n42949 );
nor U105662 ( n42948, n42961, n40865 );
nor U105663 ( n42949, n42950, n42951 );
nor U105664 ( n42961, n587, n73551 );
nand U105665 ( n1666, n42412, n42413 );
nor U105666 ( n42412, n42434, n41199 );
nor U105667 ( n42413, n42414, n42415 );
nor U105668 ( n42434, n587, n73523 );
nand U105669 ( n1681, n42237, n42238 );
nor U105670 ( n42237, n42262, n40785 );
nor U105671 ( n42238, n42239, n42240 );
nor U105672 ( n42262, n587, n73475 );
nand U105673 ( n1691, n42202, n42203 );
nor U105674 ( n42202, n42218, n42219 );
nor U105675 ( n42203, n42204, n42205 );
nor U105676 ( n42219, P3_STATE_REG, n73823 );
nand U105677 ( n44851, n44852, n44853 );
nand U105678 ( n44853, n577, n44854 );
nand U105679 ( n44852, n575, n44858 );
xor U105680 ( n44854, n44855, n44856 );
not U105681 ( n1452, n50011 );
nand U105682 ( n1911, n41060, n41061 );
nor U105683 ( n41061, n41062, n41063 );
nor U105684 ( n41060, n41069, n41070 );
nor U105685 ( n41062, n41064, n73637 );
nor U105686 ( n38543, n40089, n40176 );
and U105687 ( n40176, n36655, n40177 );
nand U105688 ( n40177, n40178, n1913 );
nor U105689 ( n13397, n13399, n76595 );
nor U105690 ( n13399, n13400, n13402 );
nand U105691 ( n13400, n13422, n13423 );
nand U105692 ( n13402, n13403, n13404 );
nand U105693 ( n13410, n13412, n13413 );
nand U105694 ( n13412, n13414, n13415 );
nand U105695 ( n13415, n13417, n12220 );
and U105696 ( n12215, n13435, n13437 );
xor U105697 ( n13437, n74847, n76034 );
nor U105698 ( n13435, n12224, n13438 );
nor U105699 ( n13438, n4892, n74818 );
nand U105700 ( n41024, n62425, n62426 );
nor U105701 ( n62426, n62427, n62428 );
nor U105702 ( n62425, n62430, n62431 );
nor U105703 ( n62428, n76244, n74714 );
xor U105704 ( n12164, n13248, n13337 );
xor U105705 ( n13337, n74586, n76034 );
nor U105706 ( n13318, n13320, n76595 );
nor U105707 ( n13320, n13322, n13323 );
nand U105708 ( n13322, n13339, n13340 );
nand U105709 ( n13323, n13324, n13325 );
nor U105710 ( n19091, n17047, n73423 );
nand U105711 ( n15771, n45929, n45930 );
nor U105712 ( n45929, n45944, n45945 );
nor U105713 ( n45930, n45931, n45932 );
nor U105714 ( n45944, n73253, n76668 );
nand U105715 ( n11281, n66880, n66881 );
nor U105716 ( n66880, n66895, n66896 );
nor U105717 ( n66881, n66882, n66883 );
nor U105718 ( n66895, n73249, n76716 );
nand U105719 ( n6791, n25004, n25005 );
nor U105720 ( n25004, n25019, n25020 );
nor U105721 ( n25005, n25006, n25007 );
nor U105722 ( n25019, n73248, n76764 );
nand U105723 ( n13526, n58139, n58140 );
nor U105724 ( n58139, n58154, n58155 );
nor U105725 ( n58140, n58141, n58142 );
nor U105726 ( n58154, n73247, n76697 );
nor U105727 ( n54757, n66179, n66347 );
and U105728 ( n66347, n41042, n66348 );
nand U105729 ( n66348, n66349, n787 );
xor U105730 ( n16393, n16703, n73797 );
nand U105731 ( n72189, n71307, n71143 );
nor U105732 ( n47072, n47074, n76329 );
nor U105733 ( n47074, n47075, n47076 );
nand U105734 ( n47075, n47095, n47096 );
nand U105735 ( n47076, n47077, n47078 );
nand U105736 ( n46050, n47087, n47088 );
nand U105737 ( n47088, n47022, n47046 );
nor U105738 ( n47087, n47089, n47090 );
nor U105739 ( n47089, n47046, n47092 );
nor U105740 ( n68103, n68105, n76869 );
nor U105741 ( n68105, n68106, n68107 );
nand U105742 ( n68106, n68126, n68127 );
nand U105743 ( n68107, n68108, n68109 );
nor U105744 ( n26100, n26102, n76904 );
nor U105745 ( n26102, n26103, n26104 );
nand U105746 ( n26103, n26123, n26124 );
nand U105747 ( n26104, n26105, n26106 );
nor U105748 ( n59241, n59243, n76878 );
nor U105749 ( n59243, n59244, n59245 );
nand U105750 ( n59244, n59264, n59265 );
nand U105751 ( n59245, n59246, n59247 );
nand U105752 ( n66990, n68118, n68119 );
nand U105753 ( n68119, n68057, n68077 );
nor U105754 ( n68118, n68120, n68121 );
nor U105755 ( n68120, n68077, n68123 );
nand U105756 ( n25114, n26115, n26116 );
nand U105757 ( n26116, n26054, n26074 );
nor U105758 ( n26115, n26117, n26118 );
nor U105759 ( n26117, n26074, n26120 );
nand U105760 ( n58252, n59256, n59257 );
nand U105761 ( n59257, n59195, n59215 );
nor U105762 ( n59256, n59258, n59259 );
nor U105763 ( n59258, n59215, n59261 );
xor U105764 ( n21629, n73566, n73024 );
nand U105765 ( n13423, n13424, n74847 );
nand U105766 ( n13424, n13425, n13393 );
nor U105767 ( n13425, n13433, n13434 );
nor U105768 ( n13433, n4862, n13439 );
not U105769 ( n2083, n37102 );
nand U105770 ( n38601, n40322, n2083 );
nor U105771 ( n40322, n37300, n37097 );
nand U105772 ( n37110, n76798, n37303 );
nand U105773 ( n2916, n37697, n37698 );
nor U105774 ( n37697, n37710, n37711 );
nor U105775 ( n37698, n37699, n37700 );
nor U105776 ( n37711, n76920, n73801 );
nand U105777 ( n36305, n39032, n39033 );
nor U105778 ( n39033, n39034, n39035 );
nor U105779 ( n39032, n39037, n39038 );
nor U105780 ( n39035, n76410, n74715 );
nand U105781 ( n37935, n37936, n37937 );
nand U105782 ( n37936, n2079, n37942 );
nand U105783 ( n37937, n2078, n37938 );
xor U105784 ( n37942, n37943, n37944 );
nand U105785 ( n37921, n37922, n37923 );
nand U105786 ( n37922, n2079, n37927 );
nand U105787 ( n37923, n2078, n37924 );
xnor U105788 ( n37927, n37928, n37929 );
nand U105789 ( n37907, n37908, n37909 );
nand U105790 ( n37908, n2079, n37914 );
nand U105791 ( n37909, n2078, n37910 );
xor U105792 ( n37914, n37915, n37916 );
nand U105793 ( n37863, n37864, n37865 );
nand U105794 ( n37864, n2079, n37869 );
nand U105795 ( n37865, n2078, n37866 );
xnor U105796 ( n37869, n37870, n37871 );
nand U105797 ( n37835, n37836, n37837 );
nand U105798 ( n37836, n2079, n37842 );
nand U105799 ( n37837, n2078, n37838 );
xnor U105800 ( n37842, n37843, n37844 );
nand U105801 ( n37793, n37794, n37795 );
nand U105802 ( n37794, n2079, n37800 );
nand U105803 ( n37795, n2078, n37796 );
xor U105804 ( n37800, n37801, n37802 );
nand U105805 ( n37734, n37735, n37736 );
nand U105806 ( n37735, n2079, n37741 );
nand U105807 ( n37736, n2078, n37737 );
xor U105808 ( n37741, n37742, n37743 );
nand U105809 ( n2851, n37918, n37919 );
nor U105810 ( n37918, n37931, n36323 );
nor U105811 ( n37919, n37920, n37921 );
nor U105812 ( n37931, n37745, n73448 );
nand U105813 ( n2871, n37860, n37861 );
nor U105814 ( n37860, n37873, n36356 );
nor U105815 ( n37861, n37862, n37863 );
nor U105816 ( n37873, n37745, n73452 );
nand U105817 ( n2846, n37932, n37933 );
nor U105818 ( n37932, n37945, n37081 );
nor U105819 ( n37933, n37934, n37935 );
nor U105820 ( n37945, n37745, n73456 );
nand U105821 ( n2856, n37904, n37905 );
nor U105822 ( n37904, n37917, n36731 );
nor U105823 ( n37905, n37906, n37907 );
nor U105824 ( n37917, n37745, n73446 );
nand U105825 ( n2881, n37832, n37833 );
nor U105826 ( n37832, n37845, n36463 );
nor U105827 ( n37833, n37834, n37835 );
nor U105828 ( n37845, n37745, n73458 );
nand U105829 ( n2896, n37790, n37791 );
nor U105830 ( n37790, n37803, n36590 );
nor U105831 ( n37791, n37792, n37793 );
nor U105832 ( n37803, n37745, n73470 );
nand U105833 ( n2906, n37731, n37732 );
nor U105834 ( n37731, n37744, n36382 );
nor U105835 ( n37732, n37733, n37734 );
nor U105836 ( n37744, n37745, n73484 );
not U105837 ( n1253, n50884 );
nor U105838 ( n45688, n7527, n74919 );
not U105839 ( n7607, n47611 );
nor U105840 ( n45599, n45617, n74986 );
nor U105841 ( n46894, n7529, n46927 );
nor U105842 ( n46745, n45910, n46788 );
nand U105843 ( n46085, n7890, n47175 );
not U105844 ( n7890, n47138 );
nor U105845 ( n46958, n46085, n47011 );
nor U105846 ( n46597, n45824, n46592 );
nand U105847 ( n47445, n47523, n47524 );
nand U105848 ( n47524, n7607, n47525 );
nor U105849 ( n47523, n47526, n47527 );
nor U105850 ( n47526, n47529, n47530 );
nor U105851 ( n46540, n7528, n46499 );
nor U105852 ( n47527, n47528, n74400 );
nor U105853 ( n47528, n7607, n47525 );
and U105854 ( n47292, n47334, n47335 );
nand U105855 ( n47335, n47336, n47337 );
nor U105856 ( n47334, n47338, n47339 );
nor U105857 ( n47339, n47340, n74443 );
nand U105858 ( n46303, n76660, n45547 );
nor U105859 ( n62427, n46549, n76241 );
nand U105860 ( n37977, n37978, n37979 );
nand U105861 ( n37979, n2079, n37980 );
nand U105862 ( n37978, n2078, n38040 );
nand U105863 ( n37980, n37981, n37982 );
nand U105864 ( n37963, n37964, n37965 );
nand U105865 ( n37965, n2079, n37966 );
nand U105866 ( n37964, n2078, n37970 );
xor U105867 ( n37966, n37967, n37968 );
nand U105868 ( n37949, n37950, n37951 );
nand U105869 ( n37951, n2079, n37952 );
nand U105870 ( n37950, n2078, n37956 );
xnor U105871 ( n37952, n37953, n37954 );
nand U105872 ( n37891, n37892, n37893 );
nand U105873 ( n37893, n2079, n37894 );
nand U105874 ( n37892, n2078, n37898 );
xnor U105875 ( n37894, n37895, n37896 );
nand U105876 ( n37877, n37878, n37879 );
nand U105877 ( n37879, n2079, n37880 );
nand U105878 ( n37878, n2078, n37884 );
xor U105879 ( n37880, n37881, n37882 );
nand U105880 ( n37849, n37850, n37851 );
nand U105881 ( n37851, n2079, n37852 );
nand U105882 ( n37850, n2078, n37856 );
xor U105883 ( n37852, n37853, n37854 );
nand U105884 ( n37821, n37822, n37823 );
nand U105885 ( n37823, n2079, n37824 );
nand U105886 ( n37822, n2078, n37828 );
xor U105887 ( n37824, n37825, n37826 );
nand U105888 ( n37807, n37808, n37809 );
nand U105889 ( n37809, n2079, n37810 );
nand U105890 ( n37808, n2078, n37813 );
xnor U105891 ( n37810, n37811, n37812 );
nand U105892 ( n2891, n37804, n37805 );
nor U105893 ( n37804, n37817, n36818 );
nor U105894 ( n37805, n37806, n37807 );
nor U105895 ( n37817, n37745, n73468 );
nand U105896 ( n2831, n37974, n37975 );
nor U105897 ( n37974, n38100, n36798 );
nor U105898 ( n37975, n37976, n37977 );
nor U105899 ( n38100, n37745, n73509 );
nand U105900 ( n2836, n37960, n37961 );
nor U105901 ( n37960, n37973, n36614 );
nor U105902 ( n37961, n37962, n37963 );
nor U105903 ( n37973, n37745, n73492 );
nand U105904 ( n2841, n37946, n37947 );
nor U105905 ( n37946, n37959, n36573 );
nor U105906 ( n37947, n37948, n37949 );
nor U105907 ( n37959, n37745, n73480 );
nand U105908 ( n2861, n37888, n37889 );
nor U105909 ( n37888, n37901, n36533 );
nor U105910 ( n37889, n37890, n37891 );
nor U105911 ( n37901, n37745, n73442 );
nand U105912 ( n2866, n37874, n37875 );
nor U105913 ( n37874, n37887, n36763 );
nor U105914 ( n37875, n37876, n37877 );
nor U105915 ( n37887, n37745, n73440 );
nand U105916 ( n2876, n37846, n37847 );
nor U105917 ( n37846, n37859, n36668 );
nor U105918 ( n37847, n37848, n37849 );
nor U105919 ( n37859, n37745, n73464 );
nand U105920 ( n2886, n37818, n37819 );
nor U105921 ( n37818, n37831, n36288 );
nor U105922 ( n37819, n37820, n37821 );
nor U105923 ( n37831, n37745, n73459 );
nor U105924 ( n50389, n50395, n73421 );
nand U105925 ( n36925, n39087, n39088 );
nor U105926 ( n39088, n39089, n39090 );
nor U105927 ( n39087, n39092, n39093 );
nor U105928 ( n39090, n76410, n74703 );
nand U105929 ( n71307, n72291, n72292 );
nor U105930 ( n72291, n72295, n72296 );
nor U105931 ( n72292, n72293, n72294 );
nor U105932 ( n72296, n74279, n73026 );
not U105933 ( n27, n11620 );
nor U105934 ( n72293, n74266, n71105 );
nand U105935 ( n37789, n2077, n37783 );
nand U105936 ( n32244, n32245, n32246 );
nand U105937 ( n32245, n3059, n3548 );
nand U105938 ( n32246, n76776, n32247 );
nand U105939 ( n4546, n32241, n32242 );
nor U105940 ( n32241, n32256, n32257 );
nor U105941 ( n32242, n32243, n32244 );
nor U105942 ( n32256, n73250, n76782 );
nor U105943 ( n47049, n7540, n47051 );
nor U105944 ( n47051, n47022, n47046 );
nor U105945 ( n68080, n5754, n68082 );
nor U105946 ( n68082, n68057, n68077 );
nor U105947 ( n26077, n3997, n26079 );
nor U105948 ( n26079, n26054, n26074 );
nor U105949 ( n59218, n6629, n59220 );
nor U105950 ( n59220, n59195, n59215 );
nand U105951 ( n47530, n47531, n7608 );
not U105952 ( n7608, n47608 );
nor U105953 ( n17449, n17052, n73018 );
nand U105954 ( n37143, n36425, n37297 );
nor U105955 ( n38573, n40178, n40255 );
and U105956 ( n40255, n37007, n40256 );
nand U105957 ( n40256, n1893, n2098 );
nor U105958 ( n39089, n38195, n76403 );
nand U105959 ( n9066, n12048, n12049 );
nor U105960 ( n12048, n12065, n12067 );
nor U105961 ( n12049, n12050, n12052 );
nor U105962 ( n12065, n73281, n76735 );
and U105963 ( n37976, n38038, n2077 );
and U105964 ( n37962, n37969, n2077 );
and U105965 ( n37948, n37955, n2077 );
and U105966 ( n37934, n37941, n2077 );
and U105967 ( n37906, n37913, n2077 );
and U105968 ( n37890, n37897, n2077 );
and U105969 ( n37876, n37883, n2077 );
and U105970 ( n37848, n37855, n2077 );
and U105971 ( n37834, n37841, n2077 );
and U105972 ( n37820, n37827, n2077 );
and U105973 ( n37792, n37799, n2077 );
and U105974 ( n37733, n37740, n2077 );
and U105975 ( n37699, n37706, n2077 );
nor U105976 ( n39034, n38182, n76403 );
and U105977 ( n45600, n74986, n45617 );
not U105978 ( n4898, n13245 );
nor U105979 ( n72295, n74273, n71108 );
nand U105980 ( n46021, n46022, n46023 );
nand U105981 ( n46022, n76672, n46025 );
nand U105982 ( n46023, n46024, n76662 );
nand U105983 ( n15756, n46004, n46005 );
nor U105984 ( n46005, n46006, n46007 );
nor U105985 ( n46004, n46020, n46021 );
nand U105986 ( n46007, n46008, n46009 );
nand U105987 ( n66961, n66962, n66963 );
nand U105988 ( n66962, n76720, n66965 );
nand U105989 ( n66963, n66964, n76710 );
nand U105990 ( n25085, n25086, n25087 );
nand U105991 ( n25086, n76768, n25089 );
nand U105992 ( n25087, n25088, n76758 );
nand U105993 ( n58220, n58221, n58222 );
nand U105994 ( n58221, n76701, n58224 );
nand U105995 ( n58222, n58223, n76691 );
nand U105996 ( n11266, n66944, n66945 );
nor U105997 ( n66945, n66946, n66947 );
nor U105998 ( n66944, n66960, n66961 );
nand U105999 ( n66947, n66948, n66949 );
nand U106000 ( n6776, n25068, n25069 );
nor U106001 ( n25069, n25070, n25071 );
nor U106002 ( n25068, n25084, n25085 );
nand U106003 ( n25071, n25072, n25073 );
nand U106004 ( n13511, n58203, n58204 );
nor U106005 ( n58204, n58205, n58206 );
nor U106006 ( n58203, n58219, n58220 );
nand U106007 ( n58206, n58207, n58208 );
nor U106008 ( n13068, n13070, n76596 );
nor U106009 ( n13070, n13072, n13073 );
nand U106010 ( n13073, n13074, n13075 );
nand U106011 ( n13072, n13077, n13078 );
xnor U106012 ( n11997, n13079, n13080 );
xor U106013 ( n13080, n74653, n76034 );
nand U106014 ( n13079, n13032, n13082 );
nand U106015 ( n13082, n4895, n13039 );
nor U106016 ( n54871, n66349, n66725 );
and U106017 ( n66725, n41369, n66726 );
nand U106018 ( n66726, n552, n785 );
xor U106019 ( n40242, n40289, n73803 );
nor U106020 ( n36421, n36424, n36425 );
nand U106021 ( n46342, n76661, n45575 );
nor U106022 ( n46945, n46947, n76329 );
nor U106023 ( n46947, n46948, n46949 );
nand U106024 ( n46949, n46950, n46951 );
nand U106025 ( n46948, n46959, n46960 );
nand U106026 ( n46960, n76658, n45960 );
nor U106027 ( n67980, n67982, n76869 );
nor U106028 ( n67982, n67983, n67984 );
nand U106029 ( n67984, n67985, n67986 );
nand U106030 ( n67983, n67994, n67995 );
nor U106031 ( n25977, n25979, n76904 );
nor U106032 ( n25979, n25980, n25981 );
nand U106033 ( n25981, n25982, n25983 );
nand U106034 ( n25980, n25991, n25992 );
nor U106035 ( n59115, n59117, n76878 );
nor U106036 ( n59117, n59118, n59119 );
nand U106037 ( n59119, n59120, n59121 );
nand U106038 ( n59118, n59129, n59130 );
nand U106039 ( n67995, n76706, n66911 );
nand U106040 ( n25992, n76752, n25035 );
nand U106041 ( n59130, n76685, n58170 );
nand U106042 ( n2666, n38594, n38595 );
nor U106043 ( n38595, n38596, n38597 );
nor U106044 ( n38594, n38605, n38606 );
and U106045 ( n38596, n37023, n76438 );
not U106046 ( n8214, n17053 );
nand U106047 ( n12160, n12162, n12163 );
nand U106048 ( n12162, n4790, n8763 );
nand U106049 ( n12163, n76729, n12164 );
nand U106050 ( n9051, n12138, n12139 );
nor U106051 ( n12139, n12140, n12142 );
nor U106052 ( n12138, n12159, n12160 );
nand U106053 ( n12140, n12152, n12153 );
not U106054 ( n272, n45412 );
or U106055 ( n37987, n37967, n37969 );
nor U106056 ( n49624, n50089, n76834 );
nor U106057 ( n42222, n42230, n42194 );
xor U106058 ( n42230, n42231, n42232 );
xor U106059 ( n42232, n73829, n42229 );
nor U106060 ( n17723, n17052, n73420 );
nand U106061 ( n38040, n38041, n38042 );
nand U106062 ( n38041, n1995, n38048 );
nand U106063 ( n38042, n38043, n38044 );
not U106064 ( n1995, n38043 );
or U106065 ( n38047, n37971, n37969 );
nand U106066 ( n40950, n62359, n62360 );
nor U106067 ( n62360, n62361, n62362 );
nor U106068 ( n62359, n62364, n62365 );
nor U106069 ( n62362, n76244, n74761 );
or U106070 ( n17151, n17047, n73414 );
xor U106071 ( n40167, n73948, n40205 );
nand U106072 ( n16186, n44948, n44949 );
nor U106073 ( n44949, n44950, n44951 );
nor U106074 ( n44948, n44956, n44957 );
nor U106075 ( n44950, n43808, n44953 );
nor U106076 ( n32009, n32024, n74948 );
not U106077 ( n3220, n33876 );
nor U106078 ( n31901, n31939, n75010 );
nor U106079 ( n33185, n3142, n33219 );
nor U106080 ( n32882, n32129, n32878 );
nor U106081 ( n33037, n32218, n33079 );
nand U106082 ( n32386, n3487, n33455 );
not U106083 ( n3487, n33419 );
nor U106084 ( n33238, n32386, n33287 );
nand U106085 ( n33710, n33788, n33789 );
nand U106086 ( n33789, n3220, n33790 );
nor U106087 ( n33788, n33791, n33792 );
nor U106088 ( n33791, n33794, n33795 );
nor U106089 ( n33792, n33793, n74412 );
nor U106090 ( n33793, n3220, n33790 );
and U106091 ( n33567, n33610, n33611 );
nand U106092 ( n33611, n33612, n33613 );
nor U106093 ( n33610, n33614, n33615 );
nor U106094 ( n33615, n33616, n74455 );
nand U106095 ( n14887, n76592, n11615 );
nand U106096 ( n15751, n46026, n46027 );
nor U106097 ( n46027, n46028, n46029 );
nor U106098 ( n46026, n46045, n46046 );
nand U106099 ( n46028, n46039, n46040 );
nand U106100 ( n11261, n66966, n66967 );
nor U106101 ( n66967, n66968, n66969 );
nor U106102 ( n66966, n66985, n66986 );
nand U106103 ( n66968, n66979, n66980 );
nand U106104 ( n6771, n25090, n25091 );
nor U106105 ( n25091, n25092, n25093 );
nor U106106 ( n25090, n25109, n25110 );
nand U106107 ( n25092, n25103, n25104 );
nand U106108 ( n13506, n58228, n58229 );
nor U106109 ( n58229, n58230, n58231 );
nor U106110 ( n58228, n58247, n58248 );
nand U106111 ( n58230, n58241, n58242 );
nor U106112 ( n66612, n66627, n74947 );
nor U106113 ( n24777, n24792, n74949 );
nor U106114 ( n57911, n57926, n74950 );
not U106115 ( n5819, n68632 );
not U106116 ( n4050, n26631 );
not U106117 ( n6683, n59773 );
nor U106118 ( n66524, n66542, n75009 );
nor U106119 ( n24689, n24707, n75007 );
nor U106120 ( n57823, n57841, n75008 );
nor U106121 ( n67941, n5743, n67974 );
nor U106122 ( n25938, n3985, n25971 );
nor U106123 ( n59076, n6618, n59109 );
nor U106124 ( n67643, n66775, n67639 );
nor U106125 ( n25638, n24897, n25634 );
nor U106126 ( n58775, n58034, n58771 );
nor U106127 ( n67792, n66861, n67835 );
nor U106128 ( n25789, n24985, n25832 );
nor U106129 ( n58927, n58120, n58970 );
nand U106130 ( n67049, n6102, n68206 );
not U106131 ( n6102, n68169 );
nand U106132 ( n25149, n4324, n26205 );
not U106133 ( n4324, n26168 );
nand U106134 ( n58287, n6957, n59344 );
not U106135 ( n6957, n59307 );
nor U106136 ( n67993, n67049, n68046 );
nor U106137 ( n25990, n25149, n26043 );
nor U106138 ( n59128, n58287, n59184 );
nand U106139 ( n68466, n68544, n68545 );
nand U106140 ( n68545, n5819, n68546 );
nor U106141 ( n68544, n68547, n68548 );
nor U106142 ( n68547, n68550, n68551 );
nand U106143 ( n26465, n26543, n26544 );
nand U106144 ( n26544, n4050, n26545 );
nor U106145 ( n26543, n26546, n26547 );
nor U106146 ( n26546, n26549, n26550 );
nand U106147 ( n59604, n59685, n59686 );
nand U106148 ( n59686, n6683, n59687 );
nor U106149 ( n59685, n59688, n59689 );
nor U106150 ( n59688, n59691, n59692 );
nor U106151 ( n68548, n68549, n74408 );
nor U106152 ( n68549, n5819, n68546 );
nor U106153 ( n26547, n26548, n74409 );
nor U106154 ( n26548, n4050, n26545 );
nor U106155 ( n59689, n59690, n74410 );
nor U106156 ( n59690, n6683, n59687 );
and U106157 ( n68323, n68366, n68367 );
nand U106158 ( n68367, n68368, n68369 );
nor U106159 ( n68366, n68370, n68371 );
nor U106160 ( n68371, n68372, n74452 );
and U106161 ( n26322, n26365, n26366 );
nand U106162 ( n26366, n26367, n26368 );
nor U106163 ( n26365, n26369, n26370 );
nor U106164 ( n26370, n26371, n74453 );
and U106165 ( n59461, n59504, n59505 );
nand U106166 ( n59505, n59506, n59507 );
nor U106167 ( n59504, n59508, n59509 );
nor U106168 ( n59509, n59510, n74454 );
nand U106169 ( n46461, n45618, n45617 );
nor U106170 ( n46442, n46459, n46460 );
nor U106171 ( n46459, n46415, n46463 );
nor U106172 ( n46460, n46413, n46461 );
nand U106173 ( n46463, n45615, n45614 );
nor U106174 ( n13362, n13364, n76595 );
nor U106175 ( n13364, n13365, n13367 );
nand U106176 ( n13367, n13368, n13369 );
nand U106177 ( n13365, n13370, n13372 );
nand U106178 ( n13372, n76725, n12180 );
nand U106179 ( n37295, n38839, n38840 );
nor U106180 ( n38840, n38841, n38842 );
nor U106181 ( n38839, n38845, n38846 );
nor U106182 ( n38842, n76410, n74782 );
nor U106183 ( n47680, n47682, n73071 );
nand U106184 ( n54999, n67264, n67265 );
nor U106185 ( n67264, n67283, n67284 );
nor U106186 ( n67265, n67266, n67267 );
nand U106187 ( n67283, n67293, n67294 );
nand U106188 ( n67267, n67268, n67269 );
nand U106189 ( n67268, n619, n67273 );
nand U106190 ( n67269, n619, n67270 );
nand U106191 ( n67273, n67274, n67275 );
not U106192 ( n817, n70968 );
nand U106193 ( n67261, n70963, n70964 );
nand U106194 ( n70964, n70965, n74537 );
nor U106195 ( n70963, n67262, n70966 );
nor U106196 ( n70966, n74537, n70967 );
or U106197 ( n41479, n54999, n55000 );
nand U106198 ( n36429, n38906, n38907 );
nor U106199 ( n38907, n38908, n38909 );
nor U106200 ( n38906, n38911, n38912 );
nor U106201 ( n38909, n76410, n74777 );
nand U106202 ( n67284, n67285, n67286 );
nand U106203 ( n67285, n619, n67290 );
nand U106204 ( n67286, n619, n67287 );
nand U106205 ( n67290, n67291, n67292 );
nand U106206 ( n36442, n38965, n38966 );
nor U106207 ( n38966, n38967, n38968 );
nor U106208 ( n38965, n38970, n38971 );
nor U106209 ( n38968, n76410, n74775 );
nor U106210 ( n62361, n46220, n76241 );
nand U106211 ( n33795, n33796, n3222 );
not U106212 ( n3222, n33873 );
nand U106213 ( n40713, n62242, n62243 );
nor U106214 ( n62243, n62244, n62245 );
nor U106215 ( n62242, n62247, n62248 );
nor U106216 ( n62245, n76244, n74809 );
nand U106217 ( n67266, n67276, n67277 );
nand U106218 ( n67276, n619, n67281 );
nand U106219 ( n67277, n619, n67278 );
nand U106220 ( n67281, n67282, n74624 );
nand U106221 ( n68551, n68552, n5820 );
nand U106222 ( n26550, n26551, n4052 );
nand U106223 ( n59692, n59693, n6684 );
not U106224 ( n5820, n68629 );
not U106225 ( n4052, n26628 );
not U106226 ( n6684, n59770 );
nand U106227 ( n37985, n37969, n37967 );
nand U106228 ( n37981, n1997, n37988 );
not U106229 ( n1997, n37983 );
nand U106230 ( n37988, n37987, n37989 );
nand U106231 ( n37989, n37985, n74457 );
nand U106232 ( n38045, n37969, n37971 );
nand U106233 ( n38048, n38047, n38049 );
nand U106234 ( n38049, n38045, n74456 );
not U106235 ( n2444, n18164 );
nand U106236 ( n32351, n33361, n33362 );
nand U106237 ( n33362, n33295, n33320 );
nor U106238 ( n33361, n33363, n33364 );
nor U106239 ( n33363, n33320, n33366 );
nor U106240 ( n33346, n33348, n76895 );
nor U106241 ( n33348, n33349, n33350 );
nand U106242 ( n33349, n33374, n33375 );
nand U106243 ( n33350, n33351, n33352 );
nand U106244 ( n33320, n33296, n33367 );
nand U106245 ( n33367, n33368, n33301 );
and U106246 ( n33368, n33370, n33371 );
nand U106247 ( n38597, n38598, n38599 );
nand U106248 ( n38599, n38600, n37764 );
nand U106249 ( n38598, n38602, n76442 );
nand U106250 ( n38600, n38109, n38108 );
nor U106251 ( n46984, n46986, n76329 );
nor U106252 ( n46986, n46987, n46988 );
nand U106253 ( n46988, n46989, n46990 );
nand U106254 ( n46987, n47003, n47004 );
nor U106255 ( n47019, n47021, n7540 );
and U106256 ( n47003, n75787, n75788 );
nand U106257 ( n75787, n46779, n46993 );
nand U106258 ( n75788, n45978, n76657 );
xnor U106259 ( n45978, n47016, n47017 );
xor U106260 ( n47017, n74417, n76341 );
nand U106261 ( n47016, n46963, n47018 );
nand U106262 ( n47018, n47019, n47020 );
nor U106263 ( n68019, n68021, n76869 );
nor U106264 ( n68021, n68022, n68023 );
nand U106265 ( n68023, n68024, n68025 );
nand U106266 ( n68022, n68038, n68039 );
nor U106267 ( n26016, n26018, n76904 );
nor U106268 ( n26018, n26019, n26020 );
nand U106269 ( n26020, n26021, n26022 );
nand U106270 ( n26019, n26035, n26036 );
nor U106271 ( n59157, n59159, n76878 );
nor U106272 ( n59159, n59160, n59161 );
nand U106273 ( n59161, n59162, n59163 );
nand U106274 ( n59160, n59176, n59177 );
nor U106275 ( n68054, n68056, n5754 );
nor U106276 ( n26051, n26053, n3997 );
nor U106277 ( n59192, n59194, n6629 );
and U106278 ( n68038, n75789, n75790 );
nand U106279 ( n75789, n67826, n68028 );
nand U106280 ( n75790, n66929, n76705 );
and U106281 ( n26035, n75791, n75792 );
nand U106282 ( n75791, n25823, n26025 );
nand U106283 ( n75792, n25053, n76751 );
and U106284 ( n59176, n75793, n75794 );
nand U106285 ( n75793, n58961, n59166 );
nand U106286 ( n75794, n58188, n76684 );
xnor U106287 ( n66929, n68051, n68052 );
xor U106288 ( n68052, n74431, n76197 );
nand U106289 ( n68051, n67998, n68053 );
nand U106290 ( n68053, n68054, n68055 );
xnor U106291 ( n25053, n26048, n26049 );
xor U106292 ( n26049, n74432, n76521 );
nand U106293 ( n26048, n25995, n26050 );
nand U106294 ( n26050, n26051, n26052 );
xnor U106295 ( n58188, n59189, n59190 );
xor U106296 ( n59190, n74433, n76263 );
nand U106297 ( n59189, n59133, n59191 );
nand U106298 ( n59191, n59192, n59193 );
and U106299 ( n31902, n75010, n31939 );
nand U106300 ( n13403, n13420, n13414 );
nor U106301 ( n45685, n74919, n7557 );
nand U106302 ( n47596, n47514, n47649 );
nand U106303 ( n47649, n47650, n7605 );
nor U106304 ( n45596, n74986, n45614 );
nor U106305 ( n46897, n46927, n7559 );
nor U106306 ( n46748, n46788, n45921 );
nor U106307 ( n46955, n47011, n7560 );
nor U106308 ( n46600, n46592, n45821 );
nor U106309 ( n47108, n47138, n47178 );
nor U106310 ( n46542, n46499, n7558 );
nand U106311 ( n46323, n7490, n45533 );
nand U106312 ( n47252, n47282, n47298 );
nand U106313 ( n47298, n47299, n47284 );
not U106314 ( n7605, n47515 );
and U106315 ( n47349, n47433, n47481 );
nand U106316 ( n47481, n47482, n47435 );
not U106317 ( n2194, n37353 );
and U106318 ( n66525, n75009, n66542 );
and U106319 ( n24690, n75007, n24707 );
and U106320 ( n57824, n75008, n57841 );
nor U106321 ( n50907, n73426, n50395 );
xnor U106322 ( n32272, n33206, n33241 );
xor U106323 ( n33241, n74855, n76471 );
nor U106324 ( n33225, n33227, n76895 );
nor U106325 ( n33227, n33228, n33229 );
nand U106326 ( n33229, n33230, n33231 );
nand U106327 ( n33228, n33239, n33240 );
nand U106328 ( n32641, n76774, n31877 );
nor U106329 ( n33305, n33307, n76895 );
nor U106330 ( n33307, n33308, n33309 );
nand U106331 ( n33309, n33310, n33311 );
nand U106332 ( n33308, n33312, n33313 );
nor U106333 ( n33317, n33295, n33318 );
nor U106334 ( n33318, n76021, n33319 );
nor U106335 ( n33319, n74460, n33320 );
nand U106336 ( n33313, n76772, n32325 );
nor U106337 ( n38841, n76403, n38128 );
nand U106338 ( n25401, n76754, n24663 );
nand U106339 ( n58538, n76687, n57799 );
nand U106340 ( n67406, n76708, n66500 );
nor U106341 ( n38908, n38147, n76403 );
nor U106342 ( n38967, n38163, n76403 );
nor U106343 ( n18183, n73022, n17052 );
and U106344 ( n37076, n37092, n37093 );
nor U106345 ( n37092, n37099, n37100 );
nor U106346 ( n37093, n37094, n37095 );
nor U106347 ( n37099, n37101, n37102 );
nor U106348 ( n37095, n37096, n37097 );
and U106349 ( n37096, n2039, n37098 );
nor U106350 ( n18879, n17047, n73422 );
nand U106351 ( n11985, n11994, n11995 );
nand U106352 ( n11994, n11963, n74737 );
nand U106353 ( n11995, n76729, n11997 );
nand U106354 ( n9076, n11983, n11984 );
nor U106355 ( n11983, n12004, n12005 );
nor U106356 ( n11984, n11985, n11987 );
nor U106357 ( n12004, n75006, n76735 );
nor U106358 ( n62244, n45750, n76241 );
nand U106359 ( n45952, n45958, n45959 );
nand U106360 ( n45958, n45940, n75197 );
nand U106361 ( n45959, n76662, n45960 );
nand U106362 ( n15766, n45950, n45951 );
nor U106363 ( n45950, n45966, n45967 );
nor U106364 ( n45951, n45952, n45953 );
nor U106365 ( n45966, n74868, n76668 );
nand U106366 ( n66903, n66909, n66910 );
nand U106367 ( n66909, n66891, n75196 );
nand U106368 ( n66910, n76710, n66911 );
nand U106369 ( n25027, n25033, n25034 );
nand U106370 ( n25033, n25015, n75198 );
nand U106371 ( n25034, n76758, n25035 );
nand U106372 ( n58162, n58168, n58169 );
nand U106373 ( n58168, n58150, n75199 );
nand U106374 ( n58169, n76691, n58170 );
nand U106375 ( n11276, n66901, n66902 );
nor U106376 ( n66901, n66917, n66918 );
nor U106377 ( n66902, n66903, n66904 );
nor U106378 ( n66917, n74840, n76716 );
nor U106379 ( n46530, n46537, n46538 );
nor U106380 ( n46537, n46415, n46541 );
nor U106381 ( n46538, n46413, n46539 );
or U106382 ( n46541, n45686, n45685 );
or U106383 ( n46539, n45689, n45688 );
nand U106384 ( n6786, n25025, n25026 );
nor U106385 ( n25025, n25041, n25042 );
nor U106386 ( n25026, n25027, n25028 );
nor U106387 ( n25041, n74838, n76764 );
nand U106388 ( n13521, n58160, n58161 );
nor U106389 ( n58160, n58176, n58177 );
nor U106390 ( n58161, n58162, n58163 );
nor U106391 ( n58176, n74837, n76697 );
nand U106392 ( n45571, n45572, n45573 );
nand U106393 ( n45573, n76347, n45574 );
nand U106394 ( n45572, n76671, n45575 );
nor U106395 ( n18148, n17053, n75919 );
nand U106396 ( n46343, n7490, n45574 );
nand U106397 ( n48066, n76326, n45404 );
nor U106398 ( n46521, n73220, n76005 );
not U106399 ( n2377, n18892 );
nor U106400 ( n33316, n33321, n33322 );
nor U106401 ( n33322, n74460, n76470 );
nor U106402 ( n33321, n3153, n74458 );
and U106403 ( n45597, n74986, n45614 );
nand U106404 ( n32759, n31940, n31939 );
nor U106405 ( n32741, n32757, n32758 );
nor U106406 ( n32757, n32714, n32761 );
nor U106407 ( n32758, n32712, n32759 );
nand U106408 ( n32761, n31937, n31936 );
nand U106409 ( n67524, n66543, n66542 );
nand U106410 ( n25519, n24708, n24707 );
nand U106411 ( n58656, n57842, n57841 );
nor U106412 ( n67506, n67522, n67523 );
nor U106413 ( n67522, n67479, n67526 );
nor U106414 ( n67523, n67477, n67524 );
nand U106415 ( n67526, n66540, n66539 );
nor U106416 ( n25501, n25517, n25518 );
nor U106417 ( n25517, n25474, n25521 );
nor U106418 ( n25518, n25472, n25519 );
nand U106419 ( n25521, n24705, n24704 );
nor U106420 ( n58638, n58654, n58655 );
nor U106421 ( n58654, n58611, n58658 );
nor U106422 ( n58655, n58609, n58656 );
nand U106423 ( n58658, n57839, n57838 );
nor U106424 ( n12969, n74774, n76602 );
not U106425 ( n1284, n50873 );
nor U106426 ( n32817, n73232, n76021 );
nor U106427 ( n25577, n73224, n76026 );
nor U106428 ( n58714, n73225, n75997 );
nor U106429 ( n33945, n33947, n73077 );
nor U106430 ( n67582, n73223, n75989 );
xor U106431 ( n11780, n12695, n75051 );
nand U106432 ( n12695, n4882, n12697 );
not U106433 ( n4953, n14304 );
nor U106434 ( n13445, n4884, n13488 );
nor U106435 ( n13263, n12208, n13313 );
nand U106436 ( n12427, n5237, n13784 );
not U106437 ( n5237, n13738 );
nor U106438 ( n12859, n4883, n12952 );
nor U106439 ( n13512, n12427, n13578 );
nor U106440 ( n13059, n12092, n13052 );
nand U106441 ( n14097, n14194, n14195 );
nand U106442 ( n14195, n4953, n14197 );
nor U106443 ( n14194, n14198, n14199 );
nor U106444 ( n14198, n14202, n14203 );
xnor U106445 ( n16599, n16602, n16603 );
nor U106446 ( n14199, n14200, n74429 );
nor U106447 ( n14200, n4953, n14197 );
nand U106448 ( n12800, n12859, n12839 );
and U106449 ( n13920, n13965, n13967 );
nand U106450 ( n13967, n13968, n13969 );
nor U106451 ( n13965, n13970, n13972 );
nor U106452 ( n13972, n13973, n74461 );
nand U106453 ( n12745, n76728, n11820 );
nor U106454 ( n47336, n7582, n75934 );
not U106455 ( n7582, n47521 );
nor U106456 ( n68701, n68703, n73076 );
nor U106457 ( n26700, n26702, n73075 );
nor U106458 ( n59842, n59844, n73074 );
nor U106459 ( n17142, n17052, n73418 );
not U106460 ( n780, n41948 );
nor U106461 ( n16575, n17035, n76789 );
nand U106462 ( n46472, n76661, n45664 );
nand U106463 ( n12170, n12178, n12179 );
nand U106464 ( n12178, n12155, n74785 );
nand U106465 ( n12179, n76729, n12180 );
nand U106466 ( n9046, n12168, n12169 );
nor U106467 ( n12168, n12188, n12189 );
nor U106468 ( n12169, n12170, n12172 );
nor U106469 ( n12188, n74915, n76735 );
nand U106470 ( n14203, n14204, n4954 );
not U106471 ( n4954, n14300 );
xor U106472 ( n38592, n37022, n37764 );
nand U106473 ( n40834, n62298, n62299 );
nor U106474 ( n62299, n62300, n62301 );
nor U106475 ( n62298, n62303, n62304 );
nor U106476 ( n62301, n76244, n74821 );
nand U106477 ( n12909, n76728, n11919 );
xnor U106478 ( n32290, n33245, n33292 );
xor U106479 ( n33292, n73160, n76471 );
nor U106480 ( n33260, n33262, n76895 );
nor U106481 ( n33262, n33263, n33264 );
nand U106482 ( n33264, n33265, n33266 );
nand U106483 ( n33263, n33279, n33280 );
and U106484 ( n33279, n75795, n75796 );
nand U106485 ( n75795, n33070, n33269 );
nand U106486 ( n75796, n32290, n76772 );
and U106487 ( n33323, n33302, n75797 );
or U106488 ( n75797, n33295, n33320 );
nand U106489 ( n4526, n32327, n32328 );
nor U106490 ( n32328, n32329, n32330 );
nor U106491 ( n32327, n32346, n32347 );
nand U106492 ( n32329, n32340, n32341 );
nand U106493 ( n45526, n45527, n45528 );
or U106494 ( n45528, n45529, n43367 );
nand U106495 ( n45527, n76347, n45533 );
nand U106496 ( n40852, n61591, n61592 );
nor U106497 ( n61592, n61593, n61594 );
nor U106498 ( n61591, n61597, n61598 );
nor U106499 ( n61594, n76244, n74862 );
xor U106500 ( n16142, n74105, n16270 );
nor U106501 ( n32006, n74948, n32034 );
nand U106502 ( n33861, n33779, n33914 );
nand U106503 ( n33914, n33915, n3219 );
nor U106504 ( n31898, n75010, n31936 );
nor U106505 ( n33188, n33219, n3173 );
nor U106506 ( n32885, n32878, n32126 );
nor U106507 ( n33040, n33079, n32215 );
nor U106508 ( n33235, n33287, n3174 );
nor U106509 ( n33387, n33419, n33458 );
nand U106510 ( n33527, n33557, n33573 );
nand U106511 ( n33573, n33574, n33559 );
not U106512 ( n3219, n33780 );
and U106513 ( n33625, n33698, n33746 );
nand U106514 ( n33746, n33747, n33700 );
nand U106515 ( n12797, n76728, n11853 );
nor U106516 ( n47539, n74400, n47618 );
nand U106517 ( n13057, n11974, n4881 );
nor U106518 ( n13040, n13053, n13054 );
nor U106519 ( n13053, n13060, n13062 );
nor U106520 ( n13054, n13055, n13057 );
nand U106521 ( n13062, n11972, n4907 );
nor U106522 ( n66609, n74947, n66637 );
nor U106523 ( n24774, n74949, n24802 );
nor U106524 ( n57908, n74950, n57936 );
nand U106525 ( n68617, n68535, n68670 );
nand U106526 ( n68670, n68671, n5818 );
nand U106527 ( n26616, n26534, n26669 );
nand U106528 ( n26669, n26670, n4049 );
nand U106529 ( n59758, n59676, n59811 );
nand U106530 ( n59811, n59812, n6682 );
nor U106531 ( n66521, n75009, n66539 );
nor U106532 ( n24686, n75007, n24704 );
nor U106533 ( n57820, n75008, n57838 );
nor U106534 ( n67944, n67974, n5772 );
nor U106535 ( n25941, n25971, n4013 );
nor U106536 ( n59079, n59109, n6645 );
nor U106537 ( n67646, n67639, n66772 );
nor U106538 ( n25641, n25634, n24894 );
nor U106539 ( n58778, n58771, n58031 );
nor U106540 ( n67795, n67835, n66872 );
nor U106541 ( n25792, n25832, n24996 );
nor U106542 ( n58930, n58970, n58131 );
nor U106543 ( n67990, n68046, n5773 );
nor U106544 ( n25987, n26043, n4014 );
nor U106545 ( n59125, n59184, n6647 );
nor U106546 ( n68139, n68169, n68209 );
nor U106547 ( n26136, n26168, n26208 );
nor U106548 ( n59277, n59307, n59347 );
nand U106549 ( n68283, n68313, n68329 );
nand U106550 ( n68329, n68330, n68315 );
nand U106551 ( n26282, n26312, n26328 );
nand U106552 ( n26328, n26329, n26314 );
nand U106553 ( n59421, n59451, n59467 );
nand U106554 ( n59467, n59468, n59453 );
not U106555 ( n5818, n68536 );
not U106556 ( n4049, n26535 );
not U106557 ( n6682, n59677 );
and U106558 ( n68381, n68454, n68502 );
nand U106559 ( n68502, n68503, n68456 );
and U106560 ( n26380, n26453, n26501 );
nand U106561 ( n26501, n26502, n26455 );
and U106562 ( n59519, n59592, n59640 );
nand U106563 ( n59640, n59641, n59594 );
nand U106564 ( n71313, n72071, n72072 );
nor U106565 ( n72071, n72075, n72076 );
nor U106566 ( n72072, n72073, n72074 );
nor U106567 ( n72076, n74346, n73026 );
nand U106568 ( n32264, n32270, n32271 );
nand U106569 ( n32270, n32252, n75195 );
nand U106570 ( n32271, n76776, n32272 );
nand U106571 ( n4541, n32262, n32263 );
nor U106572 ( n32262, n32278, n32279 );
nor U106573 ( n32263, n32264, n32265 );
nor U106574 ( n32278, n74839, n76782 );
nor U106575 ( n50621, n50395, n76834 );
nand U106576 ( n32322, n32323, n32324 );
nand U106577 ( n32323, n76786, n32326 );
nand U106578 ( n32324, n32325, n76776 );
nand U106579 ( n4531, n32305, n32306 );
nor U106580 ( n32306, n32307, n32308 );
nor U106581 ( n32305, n32321, n32322 );
nand U106582 ( n32308, n32309, n32310 );
nor U106583 ( n72073, n73069, n71105 );
nor U106584 ( n47111, n47113, n76328 );
nor U106585 ( n47113, n47114, n47115 );
nand U106586 ( n47115, n47116, n47117 );
nand U106587 ( n47114, n47118, n47119 );
nand U106588 ( n47119, n76657, n46057 );
nor U106589 ( n68142, n68144, n76868 );
nor U106590 ( n68144, n68145, n68146 );
nand U106591 ( n68146, n68147, n68148 );
nand U106592 ( n68145, n68149, n68150 );
nor U106593 ( n26141, n26143, n76903 );
nor U106594 ( n26143, n26144, n26145 );
nand U106595 ( n26145, n26146, n26147 );
nand U106596 ( n26144, n26148, n26149 );
nor U106597 ( n59280, n59282, n76877 );
nor U106598 ( n59282, n59283, n59284 );
nand U106599 ( n59284, n59285, n59286 );
nand U106600 ( n59283, n59287, n59288 );
nand U106601 ( n68150, n76705, n67021 );
nand U106602 ( n26149, n76751, n25121 );
nand U106603 ( n59288, n76684, n58259 );
nor U106604 ( n50022, n50331, n73421 );
nand U106605 ( n31873, n31874, n31875 );
nand U106606 ( n31875, n76481, n31876 );
nand U106607 ( n31874, n76785, n31877 );
nand U106608 ( n24659, n24660, n24661 );
nand U106609 ( n24661, n76527, n24662 );
nand U106610 ( n24660, n76767, n24663 );
nand U106611 ( n57795, n57796, n57797 );
nand U106612 ( n57797, n76269, n57798 );
nand U106613 ( n57796, n76700, n57799 );
nand U106614 ( n66496, n66497, n66498 );
nand U106615 ( n66498, n76203, n66499 );
nand U106616 ( n66497, n76719, n66500 );
not U106617 ( n22, n11615 );
not U106618 ( n8213, n17440 );
nor U106619 ( n62300, n40715, n76241 );
nand U106620 ( n46595, n45703, n7527 );
nor U106621 ( n46582, n46593, n46594 );
nor U106622 ( n46593, n46415, n46598 );
nor U106623 ( n46594, n46413, n46595 );
nand U106624 ( n46598, n45712, n7557 );
nand U106625 ( n9041, n12195, n12197 );
nor U106626 ( n12195, n12229, n12230 );
nor U106627 ( n12197, n12198, n12199 );
nor U106628 ( n12229, n74905, n76735 );
nor U106629 ( n12214, n12215, n12217 );
nor U106630 ( n12217, n76034, n12219 );
nand U106631 ( n12219, n5247, n12220 );
nand U106632 ( n32642, n3103, n31876 );
nand U106633 ( n71689, n71307, n71096 );
nand U106634 ( n25402, n3947, n24662 );
nand U106635 ( n58539, n6579, n57798 );
nand U106636 ( n67407, n5704, n66499 );
nand U106637 ( n47617, n47618, n74400 );
xor U106638 ( n15348, n15482, n74301 );
and U106639 ( n31899, n75010, n31936 );
nand U106640 ( n9451, n11258, n11259 );
nor U106641 ( n11259, n11260, n11262 );
nor U106642 ( n11258, n11268, n11269 );
nor U106643 ( n11260, n9908, n11264 );
and U106644 ( n66522, n75009, n66539 );
and U106645 ( n24687, n75007, n24704 );
and U106646 ( n57821, n75008, n57838 );
nor U106647 ( n72075, n73070, n71108 );
nand U106648 ( n45610, n45611, n45612 );
nand U106649 ( n45612, n45613, n76346 );
nand U106650 ( n45611, n45616, n76670 );
and U106651 ( n45613, n45614, n45615 );
and U106652 ( n45616, n45617, n45618 );
xor U106653 ( n38508, n74198, n40095 );
nor U106654 ( n40095, n74123, n40142 );
not U106655 ( n618, n61073 );
nor U106656 ( n33612, n3195, n75940 );
not U106657 ( n3195, n33786 );
nor U106658 ( n61593, n76241, n45491 );
nor U106659 ( n26367, n4030, n75938 );
not U106660 ( n4030, n26541 );
nor U106661 ( n59506, n6663, n75939 );
not U106662 ( n6663, n59683 );
nor U106663 ( n68368, n5794, n75937 );
not U106664 ( n5794, n68542 );
nor U106665 ( n33390, n33392, n76894 );
nor U106666 ( n33392, n33393, n33394 );
nand U106667 ( n33394, n33395, n33396 );
nand U106668 ( n33393, n33397, n33398 );
nand U106669 ( n33398, n76772, n32358 );
nor U106670 ( n14408, n14410, n73079 );
and U106671 ( n32010, n74948, n32024 );
nand U106672 ( n45975, n45976, n45977 );
nand U106673 ( n45976, n42977, n45841 );
nand U106674 ( n45977, n76662, n45978 );
nand U106675 ( n15761, n45972, n45973 );
nor U106676 ( n45972, n45987, n45988 );
nor U106677 ( n45973, n45974, n45975 );
nor U106678 ( n45987, n74860, n76668 );
nand U106679 ( n66926, n66927, n66928 );
nand U106680 ( n66927, n63615, n66792 );
nand U106681 ( n66928, n76710, n66929 );
nand U106682 ( n25050, n25051, n25052 );
nand U106683 ( n25051, n22395, n24914 );
nand U106684 ( n25052, n76758, n25053 );
nand U106685 ( n58185, n58186, n58187 );
nand U106686 ( n58186, n55507, n58051 );
nand U106687 ( n58187, n76691, n58188 );
nand U106688 ( n11271, n66923, n66924 );
nor U106689 ( n66923, n66938, n66939 );
nor U106690 ( n66924, n66925, n66926 );
nor U106691 ( n66938, n74830, n76716 );
nand U106692 ( n6781, n25047, n25048 );
nor U106693 ( n25047, n25062, n25063 );
nor U106694 ( n25048, n25049, n25050 );
nor U106695 ( n25062, n74828, n76764 );
nand U106696 ( n13516, n58182, n58183 );
nor U106697 ( n58182, n58197, n58198 );
nor U106698 ( n58183, n58184, n58185 );
nor U106699 ( n58197, n74827, n76697 );
and U106700 ( n66613, n74947, n66627 );
and U106701 ( n24778, n74949, n24792 );
and U106702 ( n57912, n74950, n57926 );
nand U106703 ( n40401, n40437, n2094 );
nand U106704 ( n32770, n76775, n31985 );
nand U106705 ( n25530, n76755, n24753 );
nand U106706 ( n67535, n76709, n66588 );
nand U106707 ( n58667, n76688, n57887 );
nand U106708 ( n11815, n11817, n11818 );
nand U106709 ( n11818, n76608, n11819 );
nand U106710 ( n11817, n76738, n11820 );
not U106711 ( n8240, n50331 );
not U106712 ( n2199, n40445 );
nand U106713 ( n14285, n14183, n14352 );
nand U106714 ( n14352, n14353, n4952 );
nor U106715 ( n13449, n13488, n4910 );
nor U106716 ( n13267, n13313, n12204 );
nor U106717 ( n12854, n12952, n4909 );
nor U106718 ( n13508, n13578, n4911 );
nor U106719 ( n13064, n13052, n12088 );
nor U106720 ( n13700, n13738, n13788 );
nand U106721 ( n13870, n13908, n13928 );
nand U106722 ( n13928, n13929, n13910 );
not U106723 ( n4952, n14184 );
and U106724 ( n13992, n14082, n14142 );
nand U106725 ( n14142, n14143, n14084 );
and U106726 ( n11889, n12858, n12800 );
nand U106727 ( n12858, n74946, n12860 );
nand U106728 ( n12860, n12859, n12857 );
nor U106729 ( n38847, n76406, n36425 );
nor U106730 ( n12213, n12222, n12223 );
and U106731 ( n12222, n74847, n12224 );
nor U106732 ( n38774, n76406, n37600 );
nand U106733 ( n32622, n3103, n31834 );
xor U106734 ( n15873, n16002, n74225 );
nand U106735 ( n67387, n5704, n66457 );
nand U106736 ( n25382, n3947, n24620 );
nand U106737 ( n58519, n6579, n57752 );
or U106738 ( n49759, n50001, n73008 );
nand U106739 ( n71491, n71143, n71313 );
nor U106740 ( n39276, n76406, n36907 );
nand U106741 ( n45660, n45661, n45662 );
nand U106742 ( n45662, n76347, n45663 );
nand U106743 ( n45661, n76671, n45664 );
nor U106744 ( n38976, n76406, n36935 );
nor U106745 ( n13454, n13457, n76595 );
nor U106746 ( n13457, n13458, n13459 );
nand U106747 ( n13459, n13460, n13462 );
nand U106748 ( n13458, n13463, n13464 );
nand U106749 ( n13464, n76725, n12247 );
and U106750 ( n13143, n76606, n13198 );
nand U106751 ( n13198, n74586, n73158 );
xor U106752 ( n39683, n39755, n74391 );
nand U106753 ( n31827, n31828, n31829 );
or U106754 ( n31829, n31830, n30094 );
nand U106755 ( n31828, n76481, n31834 );
nand U106756 ( n24613, n24614, n24615 );
or U106757 ( n24615, n24616, n22773 );
nand U106758 ( n24614, n76527, n24620 );
nand U106759 ( n57745, n57746, n57747 );
or U106760 ( n57747, n57748, n55887 );
nand U106761 ( n57746, n76269, n57752 );
nand U106762 ( n66450, n66451, n66452 );
or U106763 ( n66452, n66453, n64111 );
nand U106764 ( n66451, n76203, n66457 );
xor U106765 ( n40078, n40128, n74257 );
nand U106766 ( n12964, n76728, n11953 );
nand U106767 ( n11914, n11915, n11917 );
nand U106768 ( n11917, n76608, n11918 );
nand U106769 ( n11915, n76738, n11919 );
nor U106770 ( n39153, n76406, n39085 );
nand U106771 ( n12747, n4848, n11819 );
nand U106772 ( n12799, n12839, n12854 );
nor U106773 ( n39039, n76406, n39021 );
nor U106774 ( n38913, n76406, n36446 );
nor U106775 ( n39350, n76406, n36915 );
nor U106776 ( n39094, n76406, n36848 );
not U106777 ( n265, n45404 );
nand U106778 ( n46473, n7490, n45663 );
nand U106779 ( n36575, n76806, n36577 );
nand U106780 ( n36616, n76806, n36618 );
nand U106781 ( n36400, n36401, n36402 );
nand U106782 ( n36402, n2893, n36292 );
nand U106783 ( n36401, n76806, n36403 );
xor U106784 ( n15619, n74300, n15745 );
nor U106785 ( n50077, n50331, n73021 );
nand U106786 ( n36800, n76806, n36802 );
xor U106787 ( n39990, n74298, n40035 );
xor U106788 ( n11763, n12723, n75051 );
nand U106789 ( n12723, n12697, n4908 );
nand U106790 ( n46054, n46055, n46056 );
nand U106791 ( n46055, n43032, n45841 );
nand U106792 ( n46056, n76662, n46057 );
nand U106793 ( n15746, n46051, n46052 );
nor U106794 ( n46051, n46066, n46067 );
nor U106795 ( n46052, n46053, n46054 );
nor U106796 ( n46066, n74811, n76667 );
nand U106797 ( n32881, n32025, n32024 );
nor U106798 ( n32868, n32879, n32880 );
nor U106799 ( n32879, n32714, n32884 );
nor U106800 ( n32880, n32712, n32881 );
nand U106801 ( n32884, n32035, n32034 );
nand U106802 ( n67018, n67019, n67020 );
nand U106803 ( n67019, n63731, n66792 );
nand U106804 ( n67020, n76710, n67021 );
nand U106805 ( n25118, n25119, n25120 );
nand U106806 ( n25119, n22450, n24914 );
nand U106807 ( n25120, n76758, n25121 );
nand U106808 ( n58256, n58257, n58258 );
nand U106809 ( n58257, n55565, n58051 );
nand U106810 ( n58258, n76691, n58259 );
nand U106811 ( n11256, n67015, n67016 );
nor U106812 ( n67015, n67030, n67031 );
nor U106813 ( n67016, n67017, n67018 );
nor U106814 ( n67030, n74790, n76715 );
nand U106815 ( n6766, n25115, n25116 );
nor U106816 ( n25115, n25130, n25131 );
nor U106817 ( n25116, n25117, n25118 );
nor U106818 ( n25130, n74789, n76763 );
nand U106819 ( n13501, n58253, n58254 );
nor U106820 ( n58253, n58268, n58269 );
nor U106821 ( n58254, n58255, n58256 );
nor U106822 ( n58268, n74788, n76696 );
nand U106823 ( n67642, n66628, n66627 );
nand U106824 ( n25637, n24793, n24792 );
nand U106825 ( n58774, n57927, n57926 );
nand U106826 ( n45667, n45682, n45683 );
nand U106827 ( n45683, n45684, n76346 );
nand U106828 ( n45682, n45687, n76670 );
nor U106829 ( n45684, n45685, n45686 );
nor U106830 ( n45687, n45688, n45689 );
nor U106831 ( n67629, n67640, n67641 );
nor U106832 ( n67640, n67479, n67645 );
nor U106833 ( n67641, n67477, n67642 );
nand U106834 ( n67645, n66638, n66637 );
nor U106835 ( n25624, n25635, n25636 );
nor U106836 ( n25635, n25474, n25640 );
nor U106837 ( n25636, n25472, n25637 );
nand U106838 ( n25640, n24803, n24802 );
nor U106839 ( n58761, n58772, n58773 );
nor U106840 ( n58772, n58611, n58777 );
nor U106841 ( n58773, n58609, n58774 );
nand U106842 ( n58777, n57937, n57936 );
nand U106843 ( n36765, n76805, n36767 );
nand U106844 ( n36820, n76805, n36822 );
nand U106845 ( n14873, n76592, n11610 );
nand U106846 ( n36592, n76806, n36594 );
nand U106847 ( n36670, n76806, n36672 );
nand U106848 ( n36290, n76805, n36293 );
nand U106849 ( n36733, n76806, n36735 );
nand U106850 ( n36384, n76806, n36386 );
nand U106851 ( n36652, n76806, n36655 );
nand U106852 ( n37083, n76806, n36955 );
nand U106853 ( n36325, n76805, n36327 );
nand U106854 ( n11848, n11849, n11850 );
nand U106855 ( n11850, n76608, n11852 );
nand U106856 ( n11849, n76738, n11853 );
nor U106857 ( n33804, n74412, n33883 );
nor U106858 ( n39218, n76406, n39260 );
nor U106859 ( n16801, n17052, n73015 );
xor U106860 ( n39913, n39955, n74335 );
nand U106861 ( n36535, n76806, n36537 );
nand U106862 ( n36358, n76806, n36360 );
nand U106863 ( n36465, n76806, n36467 );
nand U106864 ( n16181, n44958, n44959 );
nor U106865 ( n44959, n44960, n44961 );
nor U106866 ( n44958, n44967, n44968 );
nor U106867 ( n44960, n44965, n44966 );
nor U106868 ( n68560, n74408, n68639 );
nor U106869 ( n26559, n74409, n26638 );
nor U106870 ( n59701, n74410, n59780 );
nor U106871 ( n17034, n75913, n17035 );
not U106872 ( n2193, n37299 );
nand U106873 ( n40694, n578, n40697 );
xnor U106874 ( n37956, n37957, n37958 );
xor U106875 ( n37958, n74419, n37955 );
nand U106876 ( n31932, n31933, n31934 );
nand U106877 ( n31934, n31935, n76480 );
nand U106878 ( n31933, n31938, n76784 );
and U106879 ( n31935, n31936, n31937 );
and U106880 ( n31938, n31939, n31940 );
nand U106881 ( n40987, n578, n40989 );
and U106882 ( n71931, n71327, n71313 );
nand U106883 ( n24700, n24701, n24702 );
nand U106884 ( n24702, n24703, n76526 );
nand U106885 ( n24701, n24706, n76766 );
and U106886 ( n24703, n24704, n24705 );
nand U106887 ( n66535, n66536, n66537 );
nand U106888 ( n66537, n66538, n76202 );
nand U106889 ( n66536, n66541, n76718 );
and U106890 ( n66538, n66539, n66540 );
nand U106891 ( n57834, n57835, n57836 );
nand U106892 ( n57836, n57837, n76268 );
nand U106893 ( n57835, n57840, n76699 );
and U106894 ( n57837, n57838, n57839 );
and U106895 ( n24706, n24707, n24708 );
and U106896 ( n66541, n66542, n66543 );
and U106897 ( n57840, n57841, n57842 );
nand U106898 ( n41009, n578, n41011 );
nand U106899 ( n41201, n578, n41203 );
nand U106900 ( n9650, n67262, n817 );
nand U106901 ( n41117, n578, n41119 );
nand U106902 ( n40933, n578, n40935 );
nand U106903 ( n40763, n578, n40765 );
nand U106904 ( n41057, n578, n41059 );
xor U106905 ( n39808, n74390, n39856 );
nand U106906 ( n41452, n578, n41323 );
nand U106907 ( n40970, n578, n40972 );
nand U106908 ( n40803, n40804, n40805 );
nand U106909 ( n40805, n1777, n40696 );
nand U106910 ( n40804, n578, n40806 );
nand U106911 ( n41181, n578, n41183 );
nand U106912 ( n41148, n578, n41150 );
nand U106913 ( n40867, n578, n40869 );
nand U106914 ( n40730, n578, n40732 );
nand U106915 ( n12798, n4848, n11852 );
nor U106916 ( n13968, n4928, n75941 );
not U106917 ( n4928, n14192 );
nand U106918 ( n32287, n32288, n32289 );
nand U106919 ( n32288, n29716, n32146 );
nand U106920 ( n32289, n76776, n32290 );
nand U106921 ( n4536, n32284, n32285 );
nor U106922 ( n32284, n32299, n32300 );
nor U106923 ( n32285, n32286, n32287 );
nor U106924 ( n32299, n74829, n76782 );
nand U106925 ( n33882, n33883, n74412 );
nand U106926 ( n68638, n68639, n74408 );
nand U106927 ( n26637, n26638, n74409 );
nand U106928 ( n59779, n59780, n74410 );
nand U106929 ( n32355, n32356, n32357 );
nand U106930 ( n32356, n29771, n32146 );
nand U106931 ( n32357, n76776, n32358 );
nand U106932 ( n4521, n32352, n32353 );
nor U106933 ( n32352, n32367, n32368 );
nor U106934 ( n32353, n32354, n32355 );
nor U106935 ( n32367, n74791, n76781 );
nand U106936 ( n36944, n37087, n37088 );
nor U106937 ( n37088, n2088, n37089 );
nor U106938 ( n37087, n37090, n37091 );
nor U106939 ( n37090, n37076, n2090 );
nand U106940 ( n48055, n76326, n45400 );
nor U106941 ( n47142, n47144, n76328 );
nor U106942 ( n47144, n47145, n47146 );
nand U106943 ( n47145, n47161, n47162 );
nand U106944 ( n47146, n47147, n47148 );
nand U106945 ( n47147, n76657, n46079 );
nor U106946 ( n68173, n68175, n76868 );
nor U106947 ( n68175, n68176, n68177 );
nand U106948 ( n68176, n68192, n68193 );
nand U106949 ( n68177, n68178, n68179 );
nor U106950 ( n26172, n26174, n76903 );
nor U106951 ( n26174, n26175, n26176 );
nand U106952 ( n26175, n26191, n26192 );
nand U106953 ( n26176, n26177, n26178 );
nor U106954 ( n59311, n59313, n76877 );
nor U106955 ( n59313, n59314, n59315 );
nand U106956 ( n59314, n59330, n59331 );
nand U106957 ( n59315, n59316, n59317 );
nand U106958 ( n68178, n76705, n67043 );
nand U106959 ( n26177, n76751, n25143 );
nand U106960 ( n59316, n76684, n58281 );
nor U106961 ( n16612, n17047, n76788 );
nor U106962 ( n38116, n37298, n38108 );
nor U106963 ( n33426, n33428, n76894 );
nor U106964 ( n33428, n33429, n33430 );
nand U106965 ( n33429, n33441, n33442 );
nand U106966 ( n33430, n33431, n33432 );
xnor U106967 ( n32380, n33439, n33440 );
xor U106968 ( n33440, n73115, n76471 );
nand U106969 ( n33439, n33405, n33299 );
nand U106970 ( n40787, n578, n40789 );
xor U106971 ( n38440, n72933, n39927 );
nor U106972 ( n39927, n72932, n39970 );
nor U106973 ( n40004, n40049, n72930 );
nand U106974 ( n41039, n578, n41042 );
not U106975 ( n76258, n61177 );
nand U106976 ( n61177, n67257, n61072 );
nor U106977 ( n67257, n41445, n61073 );
and U106978 ( n61072, n67258, n55000 );
nor U106979 ( n67258, n67263, n54999 );
nor U106980 ( n67263, n67300, n67301 );
nor U106981 ( n67300, n829, n41466 );
nand U106982 ( n31981, n31982, n31983 );
nand U106983 ( n31983, n76481, n31984 );
nand U106984 ( n31982, n76785, n31985 );
nand U106985 ( n24749, n24750, n24751 );
nand U106986 ( n24751, n76527, n24752 );
nand U106987 ( n24750, n76767, n24753 );
nand U106988 ( n57883, n57884, n57885 );
nand U106989 ( n57885, n76269, n57886 );
nand U106990 ( n57884, n76700, n57887 );
nand U106991 ( n66584, n66585, n66586 );
nand U106992 ( n66586, n76203, n66587 );
nand U106993 ( n66585, n76719, n66588 );
nand U106994 ( n32087, n75050, n32965 );
or U106995 ( n32965, n32129, n74652 );
nand U106996 ( n45782, n73159, n46672 );
or U106997 ( n46672, n45824, n74585 );
nand U106998 ( n12039, n74920, n13163 );
or U106999 ( n13163, n12092, n74625 );
nand U107000 ( n66690, n74637, n67719 );
or U107001 ( n67719, n66775, n74595 );
nand U107002 ( n24855, n74638, n25714 );
or U107003 ( n25714, n24897, n74596 );
nand U107004 ( n57989, n74639, n58854 );
or U107005 ( n58854, n58034, n74597 );
nand U107006 ( n9036, n12239, n12240 );
nor U107007 ( n12239, n12258, n12259 );
nor U107008 ( n12240, n12242, n12243 );
nor U107009 ( n12258, n73254, n76735 );
not U107010 ( n2368, n17928 );
nand U107011 ( n12243, n12244, n12245 );
nand U107012 ( n12244, n4790, n5295 );
nand U107013 ( n12245, n76729, n12247 );
nor U107014 ( n38107, n37354, n38108 );
nor U107015 ( n50580, n50031, n73426 );
nor U107016 ( n14214, n74429, n14313 );
and U107017 ( n71311, n72064, n72065 );
nor U107018 ( n72064, n72068, n72069 );
nor U107019 ( n72065, n72066, n72067 );
nor U107020 ( n72069, n74389, n73026 );
nor U107021 ( n65806, n72931, n65930 );
nor U107022 ( n66010, n66096, n72929 );
nor U107023 ( n66185, n74170, n66278 );
nor U107024 ( n16788, n17053, n73418 );
nor U107025 ( n17377, n17440, n73420 );
nor U107026 ( n13597, n13599, n76595 );
nor U107027 ( n13599, n13600, n13602 );
nand U107028 ( n13600, n13622, n13623 );
nand U107029 ( n13602, n13603, n13604 );
nor U107030 ( n13609, n13590, n13610 );
nor U107031 ( n13610, n76602, n13612 );
nor U107032 ( n13612, n74468, n13613 );
nand U107033 ( n13603, n76725, n12344 );
nand U107034 ( n32771, n3103, n31984 );
nand U107035 ( n36653, n36654, n36292 );
nor U107036 ( n13655, n13658, n76595 );
nor U107037 ( n13658, n13659, n13660 );
nand U107038 ( n13659, n13684, n13685 );
nand U107039 ( n13660, n13662, n13663 );
nand U107040 ( n12377, n13674, n13675 );
nand U107041 ( n13675, n13590, n13613 );
nor U107042 ( n13674, n13677, n13678 );
nor U107043 ( n13677, n13613, n13680 );
nand U107044 ( n25531, n3947, n24752 );
nand U107045 ( n67536, n5704, n66587 );
nand U107046 ( n58668, n6579, n57886 );
nor U107047 ( n72066, n74385, n71105 );
nand U107048 ( n11957, n11968, n11969 );
nand U107049 ( n11969, n11970, n76607 );
nand U107050 ( n11968, n11973, n76737 );
and U107051 ( n11970, n4907, n11972 );
and U107052 ( n11973, n4881, n11974 );
nand U107053 ( n36385, n36292, n75247 );
or U107054 ( n50069, n50031, n73021 );
and U107055 ( n45702, n7527, n45703 );
xor U107056 ( n38345, n72947, n39578 );
nor U107057 ( n39826, n72938, n39871 );
nor U107058 ( n39700, n72941, n39770 );
nor U107059 ( n39578, n72944, n39640 );
xor U107060 ( n39561, n73495, n39626 );
and U107061 ( n11888, n12853, n12799 );
nand U107062 ( n12853, n74946, n12855 );
nand U107063 ( n12855, n12854, n12857 );
xor U107064 ( n14778, n14923, n74395 );
nand U107065 ( n11754, n11755, n11757 );
or U107066 ( n11757, n11758, n9425 );
nand U107067 ( n11755, n76608, n11763 );
nor U107068 ( n47182, n47184, n76328 );
nor U107069 ( n47184, n47185, n47186 );
nand U107070 ( n47186, n47187, n47188 );
nand U107071 ( n47185, n47195, n47196 );
nor U107072 ( n47203, n7544, n73178 );
nand U107073 ( n47196, n76657, n46113 );
nor U107074 ( n68213, n68215, n76868 );
nor U107075 ( n68215, n68216, n68217 );
nand U107076 ( n68217, n68218, n68219 );
nand U107077 ( n68216, n68226, n68227 );
nor U107078 ( n26212, n26214, n76903 );
nor U107079 ( n26214, n26215, n26216 );
nand U107080 ( n26216, n26217, n26218 );
nand U107081 ( n26215, n26225, n26226 );
nor U107082 ( n59351, n59353, n76877 );
nor U107083 ( n59353, n59354, n59355 );
nand U107084 ( n59355, n59356, n59357 );
nand U107085 ( n59354, n59364, n59365 );
nor U107086 ( n68234, n5758, n73187 );
nor U107087 ( n26233, n4000, n73188 );
nor U107088 ( n59372, n6633, n73189 );
nand U107089 ( n68227, n76706, n67077 );
nand U107090 ( n26226, n76752, n25179 );
nand U107091 ( n59365, n76685, n58315 );
nand U107092 ( n14312, n14313, n74429 );
nor U107093 ( n72068, n74387, n71108 );
not U107094 ( n2198, n37091 );
nor U107095 ( n40451, n73496, n40450 );
nor U107096 ( n40449, n40450, n40451 );
nand U107097 ( n71798, n71313, n71096 );
and U107098 ( n32007, n74948, n32034 );
nor U107099 ( n40324, n37097, n37303 );
xor U107100 ( n15084, n74392, n15214 );
and U107101 ( n66610, n74947, n66637 );
and U107102 ( n24775, n74949, n24802 );
and U107103 ( n57909, n74950, n57936 );
nand U107104 ( n32894, n76775, n32064 );
nand U107105 ( n67655, n76709, n66667 );
nand U107106 ( n25650, n76755, n24832 );
nand U107107 ( n58790, n76688, n57966 );
nor U107108 ( n17710, n17440, n75919 );
nand U107109 ( n13074, n76728, n12010 );
nand U107110 ( n46608, n76660, n45741 );
nor U107111 ( n33462, n33464, n76894 );
nor U107112 ( n33464, n33465, n33466 );
nand U107113 ( n33466, n33467, n33468 );
nand U107114 ( n33465, n33475, n33476 );
nand U107115 ( n32414, n33477, n33478 );
nand U107116 ( n33477, n33480, n33370 );
nand U107117 ( n33478, n33479, n3144 );
nand U107118 ( n33480, n33371, n33405 );
not U107119 ( n3144, n33370 );
nand U107120 ( n9768, n67262, n620 );
nand U107121 ( n12982, n4848, n11929 );
nor U107122 ( n50368, n50031, n73424 );
xor U107123 ( n49373, n72935, n65806 );
nor U107124 ( n17434, n17440, n73020 );
nand U107125 ( n36264, n37102, n37097 );
and U107126 ( n13617, n13589, n75798 );
or U107127 ( n75798, n13590, n13613 );
and U107128 ( n47206, n47157, n75799 );
or U107129 ( n75799, n76341, n47204 );
and U107130 ( n68237, n68188, n75800 );
or U107131 ( n75800, n76197, n68235 );
and U107132 ( n26236, n26187, n75801 );
or U107133 ( n75801, n76521, n26234 );
and U107134 ( n59375, n59326, n75802 );
or U107135 ( n75802, n76263, n59373 );
nor U107136 ( n36675, n36677, n73800 );
nor U107137 ( n36677, n36678, n36679 );
nand U107138 ( n36678, n36681, n76920 );
nand U107139 ( n36679, n2003, n36680 );
not U107140 ( n76428, n38617 );
nand U107141 ( n38617, n38727, n38728 );
nor U107142 ( n38727, n37113, n38729 );
xor U107143 ( n48679, n72946, n63990 );
nor U107144 ( n64789, n72937, n65323 );
nor U107145 ( n64349, n72939, n64498 );
nor U107146 ( n63990, n72943, n64199 );
nor U107147 ( n37137, n37299, n37300 );
nor U107148 ( n38318, n76811, n74482 );
nor U107149 ( n38216, n76811, n74692 );
nor U107150 ( n38295, n76811, n74508 );
nor U107151 ( n38396, n76811, n74402 );
nor U107152 ( n38365, n76811, n74421 );
nor U107153 ( n38263, n76811, n74544 );
nor U107154 ( n38248, n76811, n74523 );
xor U107155 ( n54645, n74256, n66185 );
nand U107156 ( n33036, n32130, n32129 );
nor U107157 ( n33027, n33034, n33035 );
nor U107158 ( n33034, n32714, n33039 );
nor U107159 ( n33035, n32712, n33036 );
nand U107160 ( n33039, n32127, n32126 );
nand U107161 ( n46744, n45825, n45824 );
nor U107162 ( n46735, n46742, n46743 );
nor U107163 ( n46742, n46415, n46747 );
nor U107164 ( n46743, n46413, n46744 );
nand U107165 ( n46747, n45822, n45821 );
nand U107166 ( n67791, n66776, n66775 );
nand U107167 ( n13262, n12093, n12092 );
nor U107168 ( n13250, n13259, n13260 );
nor U107169 ( n13259, n13060, n13265 );
nor U107170 ( n13260, n13055, n13262 );
nand U107171 ( n13265, n12089, n12088 );
nand U107172 ( n25788, n24898, n24897 );
nand U107173 ( n58926, n58035, n58034 );
nor U107174 ( n67782, n67789, n67790 );
nor U107175 ( n67789, n67479, n67794 );
nor U107176 ( n67790, n67477, n67791 );
nand U107177 ( n67794, n66773, n66772 );
nor U107178 ( n25779, n25786, n25787 );
nor U107179 ( n25786, n25474, n25791 );
nor U107180 ( n25787, n25472, n25788 );
nand U107181 ( n25791, n24895, n24894 );
nor U107182 ( n58917, n58924, n58925 );
nor U107183 ( n58924, n58611, n58929 );
nor U107184 ( n58925, n58609, n58926 );
nand U107185 ( n58929, n58032, n58031 );
nand U107186 ( n46075, n46076, n46077 );
nand U107187 ( n46077, n46062, n74554 );
nand U107188 ( n46076, n76662, n46079 );
nand U107189 ( n15741, n46072, n46073 );
nor U107190 ( n46072, n46087, n46088 );
nor U107191 ( n46073, n46074, n46075 );
nor U107192 ( n46087, n74769, n76667 );
nand U107193 ( n67039, n67040, n67041 );
nand U107194 ( n67041, n67026, n74558 );
nand U107195 ( n67040, n76710, n67043 );
nand U107196 ( n25139, n25140, n25141 );
nand U107197 ( n25141, n25126, n74559 );
nand U107198 ( n25140, n76758, n25143 );
nand U107199 ( n58277, n58278, n58279 );
nand U107200 ( n58279, n58264, n74560 );
nand U107201 ( n58278, n76691, n58281 );
nand U107202 ( n11251, n67036, n67037 );
nor U107203 ( n67036, n67051, n67052 );
nor U107204 ( n67037, n67038, n67039 );
nor U107205 ( n67051, n74745, n76715 );
nand U107206 ( n6761, n25136, n25137 );
nor U107207 ( n25136, n25151, n25152 );
nor U107208 ( n25137, n25138, n25139 );
nor U107209 ( n25151, n74744, n76763 );
nand U107210 ( n13496, n58274, n58275 );
nor U107211 ( n58274, n58289, n58290 );
nor U107212 ( n58275, n58276, n58277 );
nor U107213 ( n58289, n74743, n76696 );
nand U107214 ( n48044, n76326, n45396 );
nand U107215 ( n32376, n32377, n32378 );
nand U107216 ( n32378, n32363, n74557 );
nand U107217 ( n32377, n76776, n32380 );
nand U107218 ( n4516, n32373, n32374 );
nor U107219 ( n32373, n32388, n32389 );
nor U107220 ( n32374, n32375, n32376 );
nor U107221 ( n32388, n74746, n76781 );
not U107222 ( n17, n11610 );
xor U107223 ( n32113, n32129, n74652 );
xor U107224 ( n12072, n12092, n74625 );
and U107225 ( n32023, n32024, n32025 );
xor U107226 ( n45808, n45824, n74585 );
xor U107227 ( n66716, n66775, n74595 );
xor U107228 ( n24881, n24897, n74596 );
xor U107229 ( n58018, n58034, n74597 );
and U107230 ( n66626, n66627, n66628 );
and U107231 ( n24791, n24792, n24793 );
and U107232 ( n57925, n57926, n57927 );
nor U107233 ( n38605, n76809, n73799 );
nor U107234 ( n38333, n76810, n74456 );
nor U107235 ( n38413, n76809, n74398 );
nor U107236 ( n38350, n76810, n74419 );
nor U107237 ( n38588, n76809, n73802 );
nor U107238 ( n38481, n76809, n74371 );
nor U107239 ( n38428, n76810, n74393 );
nor U107240 ( n38445, n76810, n74356 );
nor U107241 ( n38460, n76810, n74360 );
nor U107242 ( n38513, n76809, n74234 );
nor U107243 ( n38528, n76809, n74165 );
nor U107244 ( n38496, n76810, n74314 );
nor U107245 ( n38558, n76809, n73997 );
nor U107246 ( n38574, n76809, n73897 );
nor U107247 ( n38544, n76809, n74218 );
nor U107248 ( n38382, n76810, n74411 );
nor U107249 ( n38183, n76810, n74715 );
nor U107250 ( n38131, n76809, n74782 );
nor U107251 ( n38280, n76810, n74518 );
nor U107252 ( n38231, n76810, n74598 );
nor U107253 ( n38200, n76810, n74703 );
nor U107254 ( n38168, n76810, n74775 );
nor U107255 ( n38152, n76809, n74777 );
nand U107256 ( n9446, n11270, n11272 );
nor U107257 ( n11272, n11273, n11274 );
nor U107258 ( n11270, n11282, n11283 );
nor U107259 ( n11273, n11279, n11280 );
nor U107260 ( n50637, n73425, n50331 );
nor U107261 ( n39340, n74459, n39391 );
nor U107262 ( n39215, n74485, n39273 );
nor U107263 ( n39449, n72953, n39516 );
xnor U107264 ( n12278, n13472, n13515 );
xor U107265 ( n13515, n74823, n76034 );
nor U107266 ( n13495, n13498, n76595 );
nor U107267 ( n13498, n13499, n13500 );
nand U107268 ( n13500, n13502, n13503 );
nand U107269 ( n13499, n13513, n13514 );
nand U107270 ( n12340, n12342, n12343 );
nand U107271 ( n12342, n76739, n12345 );
nand U107272 ( n12343, n12344, n76729 );
nand U107273 ( n9021, n12319, n12320 );
nor U107274 ( n12320, n12322, n12323 );
nor U107275 ( n12319, n12339, n12340 );
nand U107276 ( n12323, n12324, n12325 );
nand U107277 ( n9016, n12347, n12348 );
nor U107278 ( n12348, n12349, n12350 );
nor U107279 ( n12347, n12370, n12372 );
nand U107280 ( n12349, n12363, n12364 );
nand U107281 ( n15736, n46094, n46095 );
nor U107282 ( n46095, n46096, n46097 );
nor U107283 ( n46094, n46109, n46110 );
nand U107284 ( n46097, n46098, n46099 );
nand U107285 ( n46110, n46111, n46112 );
nand U107286 ( n46111, n46114, n76670 );
nand U107287 ( n46112, n76662, n46113 );
nand U107288 ( n11246, n67058, n67059 );
nor U107289 ( n67059, n67060, n67061 );
nor U107290 ( n67058, n67073, n67074 );
nand U107291 ( n67061, n67062, n67063 );
nand U107292 ( n67074, n67075, n67076 );
nand U107293 ( n67075, n67078, n76718 );
nand U107294 ( n67076, n76710, n67077 );
nand U107295 ( n6756, n25160, n25161 );
nor U107296 ( n25161, n25162, n25163 );
nor U107297 ( n25160, n25175, n25176 );
nand U107298 ( n25163, n25164, n25165 );
nand U107299 ( n13491, n58296, n58297 );
nor U107300 ( n58297, n58298, n58299 );
nor U107301 ( n58296, n58311, n58312 );
nand U107302 ( n58299, n58300, n58301 );
nand U107303 ( n25176, n25177, n25178 );
nand U107304 ( n25177, n25180, n76766 );
nand U107305 ( n25178, n76758, n25179 );
nand U107306 ( n58312, n58313, n58314 );
nand U107307 ( n58313, n58316, n76699 );
nand U107308 ( n58314, n76691, n58315 );
not U107309 ( n259, n45400 );
xor U107310 ( n13652, n74418, n14375 );
xor U107311 ( n38377, n72945, n39700 );
nand U107312 ( n32060, n32061, n32062 );
nand U107313 ( n32062, n76481, n32063 );
nand U107314 ( n32061, n76785, n32064 );
nor U107315 ( n16648, n17052, n76788 );
nand U107316 ( n32169, n74610, n33113 );
or U107317 ( n33113, n32218, n74635 );
nand U107318 ( n47207, n47204, n73178 );
nand U107319 ( n68238, n68235, n73187 );
nand U107320 ( n26237, n26234, n73188 );
nand U107321 ( n59376, n59373, n73189 );
nand U107322 ( n66663, n66664, n66665 );
nand U107323 ( n66665, n76202, n66666 );
nand U107324 ( n66664, n76719, n66667 );
nand U107325 ( n45864, n74550, n46822 );
or U107326 ( n46822, n45910, n74524 );
nand U107327 ( n24828, n24829, n24830 );
nand U107328 ( n24830, n76526, n24831 );
nand U107329 ( n24829, n76767, n24832 );
nand U107330 ( n57962, n57963, n57964 );
nand U107331 ( n57964, n76268, n57965 );
nand U107332 ( n57963, n76700, n57966 );
nand U107333 ( n12147, n74586, n13355 );
or U107334 ( n13355, n12208, n74599 );
nand U107335 ( n66815, n74574, n67869 );
or U107336 ( n67869, n66861, n74546 );
xor U107337 ( n38476, n72934, n40004 );
nand U107338 ( n24939, n74575, n25866 );
or U107339 ( n25866, n24985, n74547 );
nand U107340 ( n58074, n74576, n59004 );
or U107341 ( n59004, n58120, n74548 );
nand U107342 ( n14859, n76592, n11605 );
nand U107343 ( n45737, n45738, n45739 );
nand U107344 ( n45739, n76346, n45740 );
nand U107345 ( n45738, n76671, n45741 );
nand U107346 ( n12005, n12007, n12008 );
nand U107347 ( n12008, n76608, n12009 );
nand U107348 ( n12007, n76738, n12010 );
and U107349 ( n38728, n40403, n37114 );
nor U107350 ( n40403, n40407, n37108 );
nor U107351 ( n40407, n40408, n40409 );
xor U107352 ( n40408, n37102, n37097 );
nor U107353 ( n28740, n22674, n74058 );
nor U107354 ( n62045, n55787, n74057 );
nand U107355 ( n23095, n23160, n23161 );
nand U107356 ( n23161, n76540, n73394 );
nand U107357 ( n56216, n56281, n56282 );
nand U107358 ( n56282, n76282, n73393 );
nand U107359 ( n28730, n28738, n28739 );
nor U107360 ( n28738, n28742, n28743 );
nor U107361 ( n28739, n28740, n28741 );
nor U107362 ( n28743, n28673, n74120 );
nand U107363 ( n62035, n62043, n62044 );
nor U107364 ( n62043, n62047, n62048 );
nor U107365 ( n62044, n62045, n62046 );
nor U107366 ( n62048, n61978, n74119 );
or U107367 ( n23093, n23095, n75803 );
and U107368 ( n75803, n76541, n75205 );
or U107369 ( n56214, n56216, n75804 );
and U107370 ( n75804, n76283, n75203 );
nand U107371 ( n7336, n23084, n23085 );
nor U107372 ( n23084, n23147, n23148 );
nor U107373 ( n23085, n23086, n23087 );
nor U107374 ( n23147, n23151, n23152 );
nand U107375 ( n14071, n56205, n56206 );
nor U107376 ( n56205, n56268, n56269 );
nor U107377 ( n56206, n56207, n56208 );
nor U107378 ( n56268, n56272, n56273 );
nor U107379 ( n70645, n63953, n74056 );
nand U107380 ( n64585, n64648, n64649 );
nand U107381 ( n64649, n76216, n73390 );
nand U107382 ( n70635, n70643, n70644 );
nor U107383 ( n70643, n70647, n70648 );
nor U107384 ( n70644, n70645, n70646 );
nor U107385 ( n70648, n70578, n74118 );
nand U107386 ( n11826, n64574, n64575 );
nor U107387 ( n64574, n64637, n64638 );
nor U107388 ( n64575, n64576, n64577 );
nor U107389 ( n64637, n75304, n64640 );
or U107390 ( n64583, n64585, n75805 );
and U107391 ( n75805, n76217, n75204 );
nor U107392 ( n35919, n29997, n74304 );
nand U107393 ( n30426, n30489, n30490 );
nand U107394 ( n30490, n76483, n73395 );
nand U107395 ( n35909, n35917, n35918 );
nor U107396 ( n35917, n35921, n35922 );
nor U107397 ( n35918, n35919, n35920 );
nor U107398 ( n35922, n35852, n74317 );
or U107399 ( n30424, n30426, n75806 );
and U107400 ( n75806, n76484, n75206 );
nand U107401 ( n5091, n30415, n30416 );
nor U107402 ( n30415, n30478, n30479 );
nor U107403 ( n30416, n30417, n30418 );
nor U107404 ( n30478, n75311, n30481 );
nor U107405 ( n28770, n22674, n73908 );
nor U107406 ( n62075, n55787, n73909 );
nand U107407 ( n28760, n28768, n28769 );
nor U107408 ( n28768, n28772, n28773 );
nor U107409 ( n28769, n28770, n28771 );
nor U107410 ( n28773, n28673, n73946 );
nand U107411 ( n62065, n62073, n62074 );
nor U107412 ( n62073, n62077, n62078 );
nor U107413 ( n62074, n62075, n62076 );
nor U107414 ( n62078, n61978, n73947 );
nor U107415 ( n70675, n63953, n73907 );
nand U107416 ( n70665, n70673, n70674 );
nor U107417 ( n70673, n70677, n70678 );
nor U107418 ( n70674, n70675, n70676 );
nor U107419 ( n70678, n70578, n73945 );
nor U107420 ( n35949, n29997, n74262 );
nand U107421 ( n35939, n35947, n35948 );
nor U107422 ( n35947, n35951, n35952 );
nor U107423 ( n35948, n35949, n35950 );
nor U107424 ( n35952, n35852, n74278 );
xor U107425 ( n38408, n72940, n39826 );
nor U107426 ( n28734, n28661, n74096 );
nand U107427 ( n28731, n28732, n28733 );
nor U107428 ( n28732, n28736, n28737 );
nor U107429 ( n28733, n28734, n28735 );
nor U107430 ( n28736, n28665, n74076 );
nor U107431 ( n62039, n61966, n74095 );
nand U107432 ( n62036, n62037, n62038 );
nor U107433 ( n62037, n62041, n62042 );
nor U107434 ( n62038, n62039, n62040 );
nor U107435 ( n62041, n61970, n74075 );
nor U107436 ( n70639, n70566, n74094 );
nand U107437 ( n70636, n70637, n70638 );
nor U107438 ( n70637, n70641, n70642 );
nor U107439 ( n70638, n70639, n70640 );
nor U107440 ( n70641, n70570, n74073 );
nor U107441 ( n35913, n35840, n74312 );
nand U107442 ( n32411, n32412, n32413 );
nand U107443 ( n32412, n32415, n76784 );
nand U107444 ( n32413, n76776, n32414 );
nand U107445 ( n35910, n35911, n35912 );
nor U107446 ( n35911, n35915, n35916 );
nor U107447 ( n35912, n35913, n35914 );
nor U107448 ( n35915, n35844, n74307 );
nand U107449 ( n4511, n32395, n32396 );
nor U107450 ( n32396, n32397, n32398 );
nor U107451 ( n32395, n32410, n32411 );
nand U107452 ( n32398, n32399, n32400 );
nor U107453 ( n28764, n28661, n73934 );
nor U107454 ( n62069, n61966, n73935 );
nand U107455 ( n28761, n28762, n28763 );
nor U107456 ( n28762, n28766, n28767 );
nor U107457 ( n28763, n28764, n28765 );
nor U107458 ( n28766, n28665, n73920 );
nand U107459 ( n62066, n62067, n62068 );
nor U107460 ( n62067, n62071, n62072 );
nor U107461 ( n62068, n62069, n62070 );
nor U107462 ( n62071, n61970, n73921 );
nand U107463 ( n61986, n56587, n73504 );
nand U107464 ( n28681, n23465, n73503 );
nor U107465 ( n28749, n28681, n74055 );
nor U107466 ( n62054, n61986, n74054 );
nand U107467 ( n28745, n28746, n28747 );
nor U107468 ( n28746, n28750, n28751 );
nor U107469 ( n28747, n28748, n28749 );
nor U107470 ( n28750, n28686, n74068 );
nand U107471 ( n62050, n62051, n62052 );
nor U107472 ( n62051, n62055, n62056 );
nor U107473 ( n62052, n62053, n62054 );
nor U107474 ( n62055, n61991, n74067 );
nor U107475 ( n70669, n70566, n73933 );
nand U107476 ( n70666, n70667, n70668 );
nor U107477 ( n70667, n70671, n70672 );
nor U107478 ( n70668, n70669, n70670 );
nor U107479 ( n70671, n70570, n73918 );
nand U107480 ( n70586, n64974, n73502 );
nor U107481 ( n35943, n35840, n74272 );
nor U107482 ( n70654, n70586, n74053 );
nand U107483 ( n35940, n35941, n35942 );
nor U107484 ( n35941, n35945, n35946 );
nor U107485 ( n35942, n35943, n35944 );
nor U107486 ( n35945, n35844, n74267 );
nor U107487 ( n49719, n50030, n73424 );
nand U107488 ( n70650, n70651, n70652 );
nor U107489 ( n70651, n70655, n70656 );
nor U107490 ( n70652, n70653, n70654 );
nor U107491 ( n70655, n70591, n74065 );
nand U107492 ( n35860, n30772, n73524 );
nor U107493 ( n35928, n35860, n74303 );
nand U107494 ( n35924, n35925, n35926 );
nor U107495 ( n35925, n35929, n35930 );
nor U107496 ( n35926, n35927, n35928 );
nor U107497 ( n35929, n35865, n74305 );
nor U107498 ( n28779, n28681, n73905 );
nor U107499 ( n62084, n61986, n73906 );
nand U107500 ( n28775, n28776, n28777 );
nor U107501 ( n28776, n28780, n28781 );
nor U107502 ( n28777, n28778, n28779 );
nor U107503 ( n28780, n28686, n73914 );
nand U107504 ( n62080, n62081, n62082 );
nor U107505 ( n62081, n62085, n62086 );
nor U107506 ( n62082, n62083, n62084 );
nor U107507 ( n62085, n61991, n73915 );
nor U107508 ( n70684, n70586, n73904 );
nand U107509 ( n32085, n75050, n32967 );
or U107510 ( n32967, n32126, n74652 );
nand U107511 ( n70680, n70681, n70682 );
nor U107512 ( n70681, n70685, n70686 );
nor U107513 ( n70682, n70683, n70684 );
nor U107514 ( n70685, n70591, n73912 );
nor U107515 ( n35958, n35860, n74261 );
nand U107516 ( n35954, n35955, n35956 );
nor U107517 ( n35955, n35959, n35960 );
nor U107518 ( n35956, n35957, n35958 );
nor U107519 ( n35959, n35865, n74264 );
nand U107520 ( n12037, n74920, n13165 );
or U107521 ( n13165, n12088, n74625 );
nand U107522 ( n45780, n73159, n46674 );
or U107523 ( n46674, n45821, n74585 );
nand U107524 ( n66688, n74637, n67721 );
or U107525 ( n67721, n66772, n74595 );
nand U107526 ( n24853, n74638, n25716 );
or U107527 ( n25716, n24894, n74596 );
nand U107528 ( n57987, n74639, n58856 );
or U107529 ( n58856, n58031, n74597 );
nand U107530 ( n11924, n11925, n11927 );
nand U107531 ( n11927, n4790, n5303 );
nand U107532 ( n11925, n76608, n11929 );
nor U107533 ( n28705, n28664, n73605 );
nor U107534 ( n62010, n61969, n73604 );
nand U107535 ( n28699, n28700, n28701 );
nor U107536 ( n28701, n28702, n28703 );
nor U107537 ( n28700, n28704, n28705 );
nor U107538 ( n28702, n28661, n73627 );
nand U107539 ( n62004, n62005, n62006 );
nor U107540 ( n62006, n62007, n62008 );
nor U107541 ( n62005, n62009, n62010 );
nor U107542 ( n62007, n61966, n73626 );
nor U107543 ( n39502, n73035, n39501 );
nor U107544 ( n39500, n39501, n39502 );
nor U107545 ( n70610, n70569, n73588 );
nand U107546 ( n70604, n70605, n70606 );
nor U107547 ( n70606, n70607, n70608 );
nor U107548 ( n70605, n70609, n70610 );
nor U107549 ( n70607, n70566, n73610 );
nor U107550 ( n35884, n35843, n73953 );
nand U107551 ( n35878, n35879, n35880 );
nor U107552 ( n35880, n35881, n35882 );
nor U107553 ( n35879, n35883, n35884 );
nor U107554 ( n35881, n35840, n73962 );
nor U107555 ( n28741, n28670, n74078 );
nor U107556 ( n62046, n61975, n74077 );
nor U107557 ( n70646, n70575, n74074 );
nor U107558 ( n35920, n35849, n74308 );
nor U107559 ( n28737, n28664, n74051 );
nor U107560 ( n62042, n61969, n74050 );
nor U107561 ( n28771, n28670, n73922 );
nor U107562 ( n62076, n61975, n73923 );
nor U107563 ( n70642, n70569, n74049 );
nor U107564 ( n35916, n35843, n74302 );
nor U107565 ( n70676, n70575, n73919 );
nor U107566 ( n50605, n50031, n73425 );
nor U107567 ( n35950, n35849, n74268 );
nor U107568 ( n28767, n28664, n73902 );
nor U107569 ( n62072, n61969, n73903 );
nor U107570 ( n33162, n76470, n74845 );
nor U107571 ( n70672, n70569, n73901 );
nor U107572 ( n35946, n35843, n74260 );
nand U107573 ( n28685, n23469, n73503 );
nand U107574 ( n61990, n56591, n73504 );
nor U107575 ( n28719, n28685, n73569 );
nor U107576 ( n62024, n61990, n73568 );
nand U107577 ( n28713, n28714, n28715 );
nor U107578 ( n28715, n28716, n28717 );
nor U107579 ( n28714, n28718, n28719 );
nor U107580 ( n28717, n28681, n73607 );
nand U107581 ( n62018, n62019, n62020 );
nor U107582 ( n62020, n62021, n62022 );
nor U107583 ( n62019, n62023, n62024 );
nor U107584 ( n62022, n61986, n73606 );
nand U107585 ( n70590, n64978, n73502 );
nor U107586 ( n70624, n70590, n73564 );
nor U107587 ( n28752, n28756, n28757 );
nor U107588 ( n28756, n28695, n74110 );
nor U107589 ( n28757, n28694, n74070 );
nor U107590 ( n62057, n62061, n62062 );
nor U107591 ( n62061, n62000, n74109 );
nor U107592 ( n62062, n61999, n74069 );
nand U107593 ( n70618, n70619, n70620 );
nor U107594 ( n70620, n70621, n70622 );
nor U107595 ( n70619, n70623, n70624 );
nor U107596 ( n70622, n70586, n73589 );
nand U107597 ( n35864, n30776, n73524 );
nor U107598 ( n35898, n35864, n73949 );
nand U107599 ( n35892, n35893, n35894 );
nor U107600 ( n35894, n35895, n35896 );
nor U107601 ( n35893, n35897, n35898 );
nor U107602 ( n35896, n35860, n73954 );
nor U107603 ( n28800, n22674, n74178 );
nor U107604 ( n62105, n55787, n74179 );
nor U107605 ( n70657, n70661, n70662 );
nor U107606 ( n70661, n70600, n74108 );
nor U107607 ( n70662, n70599, n74066 );
nand U107608 ( n28790, n28798, n28799 );
nor U107609 ( n28798, n28802, n28803 );
nor U107610 ( n28799, n28800, n28801 );
nor U107611 ( n28803, n28673, n74215 );
nand U107612 ( n62095, n62103, n62104 );
nor U107613 ( n62103, n62107, n62108 );
nor U107614 ( n62104, n62105, n62106 );
nor U107615 ( n62108, n61978, n74216 );
nor U107616 ( n28751, n28685, n74029 );
nor U107617 ( n62056, n61990, n74028 );
nor U107618 ( n35931, n35935, n35936 );
nor U107619 ( n35935, n35874, n74313 );
nor U107620 ( n35936, n35873, n74306 );
nor U107621 ( n70705, n63953, n74177 );
nand U107622 ( n70695, n70703, n70704 );
nor U107623 ( n70703, n70707, n70708 );
nor U107624 ( n70704, n70705, n70706 );
nor U107625 ( n70708, n70578, n74214 );
nor U107626 ( n35979, n29997, n74341 );
nor U107627 ( n70656, n70590, n74027 );
nand U107628 ( n35969, n35977, n35978 );
nor U107629 ( n35977, n35981, n35982 );
nor U107630 ( n35978, n35979, n35980 );
nor U107631 ( n35982, n35852, n74355 );
nor U107632 ( n35930, n35864, n74299 );
nor U107633 ( n28782, n28786, n28787 );
nor U107634 ( n28786, n28695, n73937 );
nor U107635 ( n28787, n28694, n73916 );
nor U107636 ( n62087, n62091, n62092 );
nor U107637 ( n62091, n62000, n73938 );
nor U107638 ( n62092, n61999, n73917 );
nor U107639 ( n70687, n70691, n70692 );
nor U107640 ( n70691, n70600, n73936 );
nor U107641 ( n70692, n70599, n73913 );
nor U107642 ( n28781, n28685, n73899 );
nor U107643 ( n28709, n28670, n73614 );
nand U107644 ( n28698, n28706, n28707 );
nor U107645 ( n28706, n28710, n28711 );
nor U107646 ( n28707, n28708, n28709 );
nor U107647 ( n28710, n28674, n73623 );
nor U107648 ( n62086, n61990, n73900 );
nor U107649 ( n62014, n61975, n73613 );
nor U107650 ( n35961, n35965, n35966 );
nor U107651 ( n35965, n35874, n74275 );
nor U107652 ( n35966, n35873, n74265 );
nand U107653 ( n62003, n62011, n62012 );
nor U107654 ( n62011, n62015, n62016 );
nor U107655 ( n62012, n62013, n62014 );
nor U107656 ( n62015, n61979, n73622 );
nor U107657 ( n70686, n70590, n73898 );
nor U107658 ( n70614, n70575, n73592 );
nand U107659 ( n70603, n70611, n70612 );
nor U107660 ( n70611, n70615, n70616 );
nor U107661 ( n70612, n70613, n70614 );
nor U107662 ( n70615, n70579, n73602 );
nor U107663 ( n35960, n35864, n74258 );
nor U107664 ( n35888, n35849, n73956 );
nor U107665 ( n61968, n61969, n73653 );
nor U107666 ( n28663, n28664, n73654 );
nand U107667 ( n35877, n35885, n35886 );
nor U107668 ( n35885, n35889, n35890 );
nor U107669 ( n35886, n35887, n35888 );
nor U107670 ( n35889, n35853, n73960 );
nand U107671 ( n61960, n61961, n61962 );
nor U107672 ( n61962, n61963, n61964 );
nor U107673 ( n61961, n61967, n61968 );
nor U107674 ( n61963, n61966, n73690 );
nand U107675 ( n28655, n28656, n28657 );
nor U107676 ( n28657, n28658, n28659 );
nor U107677 ( n28656, n28662, n28663 );
nor U107678 ( n28658, n28661, n73691 );
nor U107679 ( n70568, n70569, n73652 );
nand U107680 ( n70560, n70561, n70562 );
nor U107681 ( n70562, n70563, n70564 );
nor U107682 ( n70561, n70567, n70568 );
nor U107683 ( n70563, n70566, n73687 );
nor U107684 ( n35842, n35843, n74000 );
nand U107685 ( n35834, n35835, n35836 );
nor U107686 ( n35836, n35837, n35838 );
nor U107687 ( n35835, n35841, n35842 );
nor U107688 ( n35837, n35840, n74011 );
nor U107689 ( n28794, n28661, n74203 );
nor U107690 ( n62099, n61966, n74204 );
nand U107691 ( n28791, n28792, n28793 );
nor U107692 ( n28792, n28796, n28797 );
nor U107693 ( n28793, n28794, n28795 );
nor U107694 ( n28796, n28665, n74190 );
nand U107695 ( n62096, n62097, n62098 );
nor U107696 ( n62097, n62101, n62102 );
nor U107697 ( n62098, n62099, n62100 );
nor U107698 ( n62101, n61970, n74191 );
nor U107699 ( n70699, n70566, n74202 );
nand U107700 ( n70696, n70697, n70698 );
nor U107701 ( n70697, n70701, n70702 );
nor U107702 ( n70698, n70699, n70700 );
nor U107703 ( n70701, n70570, n74189 );
nor U107704 ( n35973, n35840, n74351 );
nand U107705 ( n35970, n35971, n35972 );
nor U107706 ( n35971, n35975, n35976 );
nor U107707 ( n35972, n35973, n35974 );
nor U107708 ( n35975, n35844, n74347 );
nand U107709 ( n7331, n23153, n23154 );
nor U107710 ( n23153, n23163, n23164 );
nor U107711 ( n23154, n23155, n23156 );
nor U107712 ( n23163, n23199, n23152 );
nand U107713 ( n33051, n76774, n32161 );
nand U107714 ( n14066, n56274, n56275 );
nor U107715 ( n56274, n56284, n56285 );
nor U107716 ( n56275, n56276, n56277 );
nor U107717 ( n56284, n56320, n56273 );
nor U107718 ( n28809, n28681, n74172 );
nor U107719 ( n62114, n61986, n74173 );
nand U107720 ( n28805, n28806, n28807 );
nor U107721 ( n28806, n28810, n28811 );
nor U107722 ( n28807, n28808, n28809 );
nor U107723 ( n28810, n28686, n74182 );
nand U107724 ( n62110, n62111, n62112 );
nor U107725 ( n62111, n62115, n62116 );
nor U107726 ( n62112, n62113, n62114 );
nor U107727 ( n62115, n61991, n74183 );
nand U107728 ( n11821, n64641, n64642 );
nor U107729 ( n64641, n64682, n64683 );
nor U107730 ( n64642, n64643, n64644 );
nor U107731 ( n64682, n75305, n64640 );
nor U107732 ( n70714, n70586, n74171 );
nand U107733 ( n70710, n70711, n70712 );
nor U107734 ( n70711, n70715, n70716 );
nor U107735 ( n70712, n70713, n70714 );
nor U107736 ( n70715, n70591, n74180 );
nand U107737 ( n5086, n30482, n30483 );
nor U107738 ( n30482, n30523, n30524 );
nor U107739 ( n30483, n30484, n30485 );
nor U107740 ( n30523, n75316, n30481 );
nor U107741 ( n35988, n35860, n74339 );
nand U107742 ( n35984, n35985, n35986 );
nor U107743 ( n35985, n35989, n35990 );
nor U107744 ( n35986, n35987, n35988 );
nor U107745 ( n35989, n35865, n74343 );
nand U107746 ( n13279, n76727, n12137 );
nand U107747 ( n46758, n76660, n45856 );
nand U107748 ( n45707, n45711, n76346 );
and U107749 ( n45711, n7557, n45712 );
nand U107750 ( n32895, n3103, n32063 );
nor U107751 ( n28753, n28754, n28755 );
nor U107752 ( n28755, n27016, n74087 );
nor U107753 ( n28754, n28691, n74117 );
nor U107754 ( n62058, n62059, n62060 );
nor U107755 ( n62060, n60157, n74086 );
nor U107756 ( n62059, n61996, n74116 );
nor U107757 ( n49502, n50331, n76834 );
nor U107758 ( n28720, n28724, n28725 );
nor U107759 ( n28724, n28695, n73609 );
nor U107760 ( n28725, n28694, n73598 );
nor U107761 ( n62025, n62029, n62030 );
nor U107762 ( n62029, n62000, n73608 );
nor U107763 ( n62030, n61999, n73597 );
nand U107764 ( n67805, n76708, n66807 );
nand U107765 ( n25802, n76754, n24929 );
nand U107766 ( n58940, n76687, n58066 );
nor U107767 ( n61989, n61990, n73642 );
nor U107768 ( n28684, n28685, n73641 );
nand U107769 ( n61981, n61982, n61983 );
nor U107770 ( n61983, n61984, n61985 );
nor U107771 ( n61982, n61988, n61989 );
nor U107772 ( n61985, n61986, n73657 );
nand U107773 ( n28676, n28677, n28678 );
nor U107774 ( n28678, n28679, n28680 );
nor U107775 ( n28677, n28683, n28684 );
nor U107776 ( n28680, n28681, n73658 );
nor U107777 ( n70658, n70659, n70660 );
nor U107778 ( n70660, n69013, n74083 );
nor U107779 ( n70659, n70596, n74115 );
nor U107780 ( n35932, n35933, n35934 );
nor U107781 ( n35934, n34259, n74310 );
nor U107782 ( n35933, n35870, n74316 );
nor U107783 ( n70625, n70629, n70630 );
nor U107784 ( n70629, n70600, n73590 );
nor U107785 ( n70630, n70599, n73583 );
nand U107786 ( n40664, n41471, n41466 );
nor U107787 ( n35899, n35903, n35904 );
nor U107788 ( n35903, n35874, n73955 );
nor U107789 ( n35904, n35873, n73951 );
nor U107790 ( n70589, n70590, n73643 );
nand U107791 ( n70581, n70582, n70583 );
nor U107792 ( n70583, n70584, n70585 );
nor U107793 ( n70582, n70588, n70589 );
nor U107794 ( n70585, n70586, n73655 );
nor U107795 ( n35863, n35864, n73987 );
nand U107796 ( n35855, n35856, n35857 );
nor U107797 ( n35857, n35858, n35859 );
nor U107798 ( n35856, n35862, n35863 );
nor U107799 ( n35859, n35860, n74001 );
nor U107800 ( n28783, n28784, n28785 );
nor U107801 ( n28785, n27016, n73928 );
nor U107802 ( n28784, n28691, n73943 );
nor U107803 ( n62088, n62089, n62090 );
nor U107804 ( n62090, n60157, n73929 );
nor U107805 ( n62089, n61996, n73944 );
nor U107806 ( n67498, n76197, n74962 );
nor U107807 ( n46434, n76341, n74930 );
nor U107808 ( n25493, n76521, n74960 );
nor U107809 ( n58630, n76263, n74963 );
nand U107810 ( n67656, n5704, n66666 );
nand U107811 ( n25651, n3947, n24831 );
nand U107812 ( n58791, n6579, n57965 );
nor U107813 ( n70688, n70689, n70690 );
nor U107814 ( n70690, n69013, n73927 );
nor U107815 ( n70689, n70596, n73942 );
nor U107816 ( n35962, n35963, n35964 );
nor U107817 ( n35964, n34259, n74270 );
nor U107818 ( n35963, n35870, n74277 );
nor U107819 ( n32733, n76470, n74961 );
xor U107820 ( n46122, n47233, n47204 );
nor U107821 ( n47226, n47228, n76328 );
nor U107822 ( n47228, n47229, n47230 );
nand U107823 ( n47229, n47246, n47247 );
nand U107824 ( n47230, n47231, n47232 );
not U107825 ( n4248, n22737 );
xor U107826 ( n67086, n68264, n68235 );
xor U107827 ( n25188, n26263, n26234 );
xor U107828 ( n58324, n59402, n59373 );
nor U107829 ( n28703, n28660, n73630 );
not U107830 ( n6880, n55853 );
nor U107831 ( n62008, n61965, n73629 );
nor U107832 ( n68257, n68259, n76868 );
nor U107833 ( n68259, n68260, n68261 );
nand U107834 ( n68260, n68277, n68278 );
nand U107835 ( n68261, n68262, n68263 );
nor U107836 ( n26256, n26258, n76903 );
nor U107837 ( n26258, n26259, n26260 );
nand U107838 ( n26259, n26276, n26277 );
nand U107839 ( n26260, n26261, n26262 );
nor U107840 ( n59395, n59397, n76877 );
nor U107841 ( n59397, n59398, n59399 );
nand U107842 ( n59398, n59415, n59416 );
nand U107843 ( n59399, n59400, n59401 );
nor U107844 ( n61974, n61975, n73679 );
nor U107845 ( n28669, n28670, n73680 );
nand U107846 ( n61959, n61971, n61972 );
nor U107847 ( n61971, n61976, n61977 );
nor U107848 ( n61972, n61973, n61974 );
nor U107849 ( n61976, n61979, n73696 );
nand U107850 ( n28654, n28666, n28667 );
nor U107851 ( n28666, n28671, n28672 );
nor U107852 ( n28667, n28668, n28669 );
nor U107853 ( n28671, n28674, n73697 );
not U107854 ( n6025, n64077 );
nor U107855 ( n70608, n70565, n73612 );
not U107856 ( n3410, n30060 );
nor U107857 ( n70574, n70575, n73675 );
nor U107858 ( n35882, n35839, n73963 );
nand U107859 ( n70559, n70571, n70572 );
nor U107860 ( n70571, n70576, n70577 );
nor U107861 ( n70572, n70573, n70574 );
nor U107862 ( n70576, n70579, n73695 );
nor U107863 ( n35848, n35849, n74007 );
nand U107864 ( n35833, n35845, n35846 );
nor U107865 ( n35845, n35850, n35851 );
nor U107866 ( n35846, n35847, n35848 );
nor U107867 ( n35850, n35853, n74014 );
nor U107868 ( n28797, n28664, n74175 );
nand U107869 ( n13075, n4848, n12009 );
nor U107870 ( n62102, n61969, n74176 );
nor U107871 ( n70702, n70569, n74174 );
nor U107872 ( n35976, n35843, n74340 );
nor U107873 ( n28801, n28670, n74193 );
nor U107874 ( n62106, n61975, n74194 );
nor U107875 ( n28742, n28674, n74114 );
nor U107876 ( n62047, n61979, n74113 );
nor U107877 ( n70706, n70575, n74192 );
nor U107878 ( n35980, n35849, n74348 );
nor U107879 ( n61992, n61997, n61998 );
nor U107880 ( n61997, n62000, n73693 );
nor U107881 ( n61998, n61999, n73672 );
nor U107882 ( n28687, n28692, n28693 );
nor U107883 ( n28692, n28695, n73694 );
nor U107884 ( n28693, n28694, n73673 );
nor U107885 ( n70647, n70579, n74112 );
nand U107886 ( n46609, n7490, n45740 );
nor U107887 ( n35921, n35853, n74315 );
nor U107888 ( n70592, n70597, n70598 );
nor U107889 ( n70597, n70600, n73692 );
nor U107890 ( n70598, n70599, n73667 );
nor U107891 ( n35866, n35871, n35872 );
nor U107892 ( n35871, n35874, n74013 );
nor U107893 ( n35872, n35873, n74004 );
nor U107894 ( n28772, n28674, n73940 );
nor U107895 ( n62077, n61979, n73941 );
nor U107896 ( n70677, n70579, n73939 );
nor U107897 ( n35951, n35853, n74276 );
nand U107898 ( n28686, n23470, n73503 );
nand U107899 ( n61991, n56592, n73504 );
xnor U107900 ( n12300, n13584, n13585 );
xor U107901 ( n13585, n73117, n76034 );
nand U107902 ( n13584, n13518, n13587 );
nand U107903 ( n13587, n4893, n13525 );
nor U107904 ( n13544, n13547, n76595 );
nor U107905 ( n13547, n13548, n13549 );
nand U107906 ( n13549, n13550, n13552 );
nand U107907 ( n13548, n13568, n13569 );
and U107908 ( n13568, n75807, n75808 );
nand U107909 ( n75807, n12828, n13555 );
nand U107910 ( n75808, n12300, n76724 );
xor U107911 ( n49136, n72942, n64789 );
nand U107912 ( n70591, n64979, n73502 );
nand U107913 ( n35865, n30777, n73524 );
nor U107914 ( n61964, n61965, n73688 );
nor U107915 ( n28659, n28660, n73689 );
nor U107916 ( n70564, n70565, n73686 );
nor U107917 ( n35838, n35839, n74010 );
nor U107918 ( n28811, n28685, n74168 );
nor U107919 ( n62116, n61990, n74169 );
nor U107920 ( n70716, n70590, n74167 );
nor U107921 ( n35990, n35864, n74338 );
nor U107922 ( n28812, n28816, n28817 );
nor U107923 ( n28816, n28695, n74206 );
nor U107924 ( n28817, n28694, n74184 );
nor U107925 ( n62117, n62121, n62122 );
nor U107926 ( n62121, n62000, n74207 );
nor U107927 ( n62122, n61999, n74185 );
nor U107928 ( n28827, n28664, n73753 );
nor U107929 ( n62132, n61969, n73754 );
nand U107930 ( n28821, n28822, n28823 );
nor U107931 ( n28823, n28824, n28825 );
nor U107932 ( n28822, n28826, n28827 );
nor U107933 ( n28824, n28661, n73783 );
nand U107934 ( n62126, n62127, n62128 );
nor U107935 ( n62128, n62129, n62130 );
nor U107936 ( n62127, n62131, n62132 );
nor U107937 ( n62129, n61966, n73784 );
nor U107938 ( n70717, n70721, n70722 );
nor U107939 ( n70721, n70600, n74205 );
nor U107940 ( n70722, n70599, n74181 );
nor U107941 ( n70732, n70569, n73752 );
nand U107942 ( n70726, n70727, n70728 );
nor U107943 ( n70728, n70729, n70730 );
nor U107944 ( n70727, n70731, n70732 );
nor U107945 ( n70729, n70566, n73782 );
nor U107946 ( n35991, n35995, n35996 );
nor U107947 ( n35995, n35874, n74352 );
nor U107948 ( n35996, n35873, n74344 );
nor U107949 ( n36006, n35843, n74102 );
nand U107950 ( n36000, n36001, n36002 );
nor U107951 ( n36002, n36003, n36004 );
nor U107952 ( n36001, n36005, n36006 );
nor U107953 ( n36003, n35840, n74131 );
nand U107954 ( n28682, n23466, n73503 );
nand U107955 ( n61987, n56588, n73504 );
nor U107956 ( n28716, n28682, n73620 );
nor U107957 ( n62021, n61987, n73619 );
nor U107958 ( n28841, n28685, n73750 );
nor U107959 ( n62146, n61990, n73751 );
nand U107960 ( n28835, n28836, n28837 );
nor U107961 ( n28837, n28838, n28839 );
nor U107962 ( n28836, n28840, n28841 );
nor U107963 ( n28839, n28681, n73756 );
nand U107964 ( n62140, n62141, n62142 );
nor U107965 ( n62142, n62143, n62144 );
nor U107966 ( n62141, n62145, n62146 );
nor U107967 ( n62144, n61986, n73757 );
nor U107968 ( n28735, n28660, n74092 );
nor U107969 ( n62040, n61965, n74091 );
nand U107970 ( n70587, n64975, n73502 );
nor U107971 ( n70621, n70587, n73596 );
nor U107972 ( n70746, n70590, n73749 );
nand U107973 ( n70740, n70741, n70742 );
nor U107974 ( n70742, n70743, n70744 );
nor U107975 ( n70741, n70745, n70746 );
nor U107976 ( n70744, n70586, n73755 );
nand U107977 ( n35861, n30773, n73524 );
nor U107978 ( n35895, n35861, n73959 );
nor U107979 ( n36020, n35864, n74063 );
nand U107980 ( n36014, n36015, n36016 );
nor U107981 ( n36016, n36017, n36018 );
nor U107982 ( n36015, n36019, n36020 );
nor U107983 ( n36018, n35860, n74104 );
nor U107984 ( n70640, n70565, n74090 );
nor U107985 ( n35914, n35839, n74311 );
nor U107986 ( n28765, n28660, n73931 );
nor U107987 ( n62070, n61965, n73932 );
nor U107988 ( n70670, n70565, n73930 );
nor U107989 ( n35944, n35839, n74271 );
nand U107990 ( n28673, n4248, n23494 );
nand U107991 ( n61978, n6880, n56616 );
nor U107992 ( n28711, n28673, n73632 );
nor U107993 ( n62016, n61978, n73631 );
nand U107994 ( n70578, n6025, n65003 );
nor U107995 ( n70616, n70578, n73621 );
nand U107996 ( n35852, n3410, n30801 );
nor U107997 ( n17950, n73423, n17440 );
nor U107998 ( n35890, n35852, n73965 );
nor U107999 ( n28813, n28814, n28815 );
nor U108000 ( n28815, n27016, n74196 );
nor U108001 ( n28814, n28691, n74212 );
nor U108002 ( n62118, n62119, n62120 );
nor U108003 ( n62120, n60157, n74197 );
nor U108004 ( n62119, n61996, n74213 );
nor U108005 ( n28831, n28670, n73771 );
nor U108006 ( n62136, n61975, n73772 );
nand U108007 ( n28820, n28828, n28829 );
nor U108008 ( n28828, n28832, n28833 );
nor U108009 ( n28829, n28830, n28831 );
nor U108010 ( n28832, n28674, n73789 );
nand U108011 ( n62125, n62133, n62134 );
nor U108012 ( n62133, n62137, n62138 );
nor U108013 ( n62134, n62135, n62136 );
nor U108014 ( n62137, n61979, n73790 );
nor U108015 ( n70718, n70719, n70720 );
nor U108016 ( n70720, n69013, n74195 );
nor U108017 ( n70719, n70596, n74211 );
nor U108018 ( n35992, n35993, n35994 );
nor U108019 ( n35994, n34259, n74349 );
nor U108020 ( n35993, n35870, n74354 );
nor U108021 ( n70736, n70575, n73768 );
nand U108022 ( n70725, n70733, n70734 );
nor U108023 ( n70733, n70737, n70738 );
nor U108024 ( n70734, n70735, n70736 );
nor U108025 ( n70737, n70579, n73788 );
nor U108026 ( n36010, n35849, n74125 );
nand U108027 ( n35999, n36007, n36008 );
nor U108028 ( n36007, n36011, n36012 );
nor U108029 ( n36008, n36009, n36010 );
nor U108030 ( n36011, n35853, n74136 );
nand U108031 ( n68055, n75990, n72950 );
nand U108032 ( n47020, n76006, n72948 );
nand U108033 ( n26052, n76027, n72951 );
nand U108034 ( n59193, n75998, n72952 );
nor U108035 ( n28795, n28660, n74200 );
nor U108036 ( n62100, n61965, n74201 );
nor U108037 ( n70700, n70565, n74199 );
nand U108038 ( n36943, n37112, n2092 );
nor U108039 ( n37112, n37113, n37114 );
nor U108040 ( n35974, n35839, n74350 );
nor U108041 ( n62871, n74462, n62945 );
nor U108042 ( n63267, n72954, n63675 );
not U108043 ( n4250, n22736 );
not U108044 ( n6883, n55852 );
not U108045 ( n6028, n64076 );
not U108046 ( n3413, n30059 );
nor U108047 ( n28842, n28846, n28847 );
nor U108048 ( n28846, n28695, n73786 );
nor U108049 ( n28847, n28694, n73765 );
nor U108050 ( n62147, n62151, n62152 );
nor U108051 ( n62151, n62000, n73787 );
nor U108052 ( n62152, n61999, n73766 );
nor U108053 ( n28721, n28722, n28723 );
nor U108054 ( n28723, n27016, n73616 );
nor U108055 ( n28722, n28691, n73625 );
nor U108056 ( n62026, n62027, n62028 );
nor U108057 ( n62028, n60157, n73615 );
nor U108058 ( n62027, n61996, n73624 );
nor U108059 ( n61984, n61987, n73682 );
nor U108060 ( n28679, n28682, n73683 );
nor U108061 ( n70747, n70751, n70752 );
nor U108062 ( n70751, n70600, n73785 );
nor U108063 ( n70752, n70599, n73762 );
nor U108064 ( n70626, n70627, n70628 );
nor U108065 ( n70628, n69013, n73594 );
nor U108066 ( n70627, n70596, n73603 );
nor U108067 ( n36021, n36025, n36026 );
nor U108068 ( n36025, n35874, n74134 );
nor U108069 ( n36026, n35873, n74122 );
nor U108070 ( n70584, n70587, n73676 );
nor U108071 ( n35900, n35901, n35902 );
nor U108072 ( n35902, n34259, n73957 );
nor U108073 ( n35901, n35870, n73961 );
nor U108074 ( n35858, n35861, n74008 );
and U108075 ( n24607, n75809, n28638 );
nand U108076 ( n75809, n28629, n28913 );
and U108077 ( n57739, n75810, n61943 );
nand U108078 ( n75810, n61934, n62218 );
nor U108079 ( n28748, n28682, n74081 );
nor U108080 ( n62053, n61987, n74080 );
not U108081 ( n4255, n28914 );
not U108082 ( n6888, n62219 );
nor U108083 ( n28629, n28645, n28641 );
nor U108084 ( n61934, n61950, n61946 );
not U108085 ( n4230, n28912 );
not U108086 ( n6863, n62217 );
nor U108087 ( n28718, n28686, n73601 );
nor U108088 ( n62023, n61991, n73600 );
and U108089 ( n66415, n75811, n70543 );
nand U108090 ( n75811, n70534, n70818 );
nor U108091 ( n70653, n70587, n74079 );
not U108092 ( n6033, n70819 );
nor U108093 ( n70534, n70550, n70546 );
not U108094 ( n6008, n70817 );
and U108095 ( n31823, n75812, n35817 );
nand U108096 ( n75812, n35808, n36092 );
nor U108097 ( n70623, n70591, n73585 );
nor U108098 ( n35927, n35861, n74309 );
not U108099 ( n3418, n36093 );
nor U108100 ( n35808, n35824, n35820 );
not U108101 ( n3393, n36091 );
nor U108102 ( n35897, n35865, n73952 );
nor U108103 ( n28778, n28682, n73925 );
nor U108104 ( n62083, n61987, n73926 );
nor U108105 ( n61977, n61978, n73703 );
nor U108106 ( n28672, n28673, n73704 );
nor U108107 ( n70683, n70587, n73924 );
nor U108108 ( n70577, n70578, n73702 );
nor U108109 ( n35957, n35861, n74269 );
nor U108110 ( n28802, n28674, n74209 );
nor U108111 ( n62107, n61979, n74210 );
nor U108112 ( n35851, n35852, n74018 );
nor U108113 ( n28825, n28660, n73780 );
nor U108114 ( n62130, n61965, n73781 );
nor U108115 ( n70707, n70579, n74208 );
nor U108116 ( n35981, n35853, n74353 );
nor U108117 ( n70730, n70565, n73779 );
nor U108118 ( n36004, n35839, n74129 );
nor U108119 ( n28857, n28664, n73835 );
nor U108120 ( n62162, n61969, n73836 );
nand U108121 ( n28851, n28852, n28853 );
nor U108122 ( n28853, n28854, n28855 );
nor U108123 ( n28852, n28856, n28857 );
nor U108124 ( n28854, n28661, n73865 );
nand U108125 ( n62156, n62157, n62158 );
nor U108126 ( n62158, n62159, n62160 );
nor U108127 ( n62157, n62161, n62162 );
nor U108128 ( n62159, n61966, n73866 );
nand U108129 ( n71031, n71098, n71313 );
nor U108130 ( n70762, n70569, n73834 );
nand U108131 ( n70756, n70757, n70758 );
nor U108132 ( n70758, n70759, n70760 );
nor U108133 ( n70757, n70761, n70762 );
nor U108134 ( n70759, n70566, n73864 );
nor U108135 ( n36036, n35843, n74222 );
nand U108136 ( n36030, n36031, n36032 );
nor U108137 ( n36032, n36033, n36034 );
nor U108138 ( n36031, n36035, n36036 );
nor U108139 ( n36033, n35840, n74235 );
nor U108140 ( n41464, n41465, n41466 );
and U108141 ( n41465, n833, n41467 );
and U108142 ( n41444, n41461, n41462 );
nor U108143 ( n41461, n41468, n41469 );
nor U108144 ( n41462, n41463, n41464 );
nor U108145 ( n41468, n41470, n41471 );
nor U108146 ( n61993, n61994, n61995 );
nor U108147 ( n61995, n60157, n73684 );
nor U108148 ( n61994, n61996, n73699 );
nor U108149 ( n28688, n28689, n28690 );
nor U108150 ( n28690, n27016, n73685 );
nor U108151 ( n28689, n28691, n73700 );
xnor U108152 ( n32430, n33509, n33484 );
nor U108153 ( n33502, n33504, n76894 );
nor U108154 ( n33504, n33505, n33506 );
nand U108155 ( n33505, n33522, n33523 );
nand U108156 ( n33506, n33507, n33508 );
nor U108157 ( n70593, n70594, n70595 );
nor U108158 ( n70595, n69013, n73681 );
nor U108159 ( n70594, n70596, n73698 );
nor U108160 ( n35867, n35868, n35869 );
nor U108161 ( n35869, n34259, n74009 );
nor U108162 ( n35868, n35870, n74015 );
nor U108163 ( n61988, n61991, n73668 );
nor U108164 ( n28683, n28686, n73669 );
xor U108165 ( n49513, n49514, n49515 );
nor U108166 ( n70588, n70591, n73665 );
nor U108167 ( n35862, n35865, n74003 );
nor U108168 ( n28871, n28685, n73831 );
nor U108169 ( n62176, n61990, n73832 );
nand U108170 ( n28865, n28866, n28867 );
nor U108171 ( n28867, n28868, n28869 );
nor U108172 ( n28866, n28870, n28871 );
nor U108173 ( n28869, n28681, n73838 );
nand U108174 ( n62170, n62171, n62172 );
nor U108175 ( n62172, n62173, n62174 );
nor U108176 ( n62171, n62175, n62176 );
nor U108177 ( n62174, n61986, n73839 );
nor U108178 ( n70776, n70590, n73830 );
nand U108179 ( n70770, n70771, n70772 );
nor U108180 ( n70772, n70773, n70774 );
nor U108181 ( n70771, n70775, n70776 );
nor U108182 ( n70774, n70586, n73837 );
nor U108183 ( n36050, n35864, n74221 );
nand U108184 ( n36044, n36045, n36046 );
nor U108185 ( n36046, n36047, n36048 );
nor U108186 ( n36045, n36049, n36050 );
nor U108187 ( n36048, n35860, n74223 );
nor U108188 ( n28808, n28682, n74187 );
nor U108189 ( n62113, n61987, n74188 );
nor U108190 ( n70713, n70587, n74186 );
nor U108191 ( n35987, n35861, n74345 );
nor U108192 ( n28704, n28665, n73618 );
nor U108193 ( n62009, n61970, n73617 );
nor U108194 ( n70609, n70570, n73595 );
nor U108195 ( n28861, n28670, n73853 );
nor U108196 ( n62166, n61975, n73854 );
nor U108197 ( n35883, n35844, n73958 );
nand U108198 ( n28850, n28858, n28859 );
nor U108199 ( n28858, n28862, n28863 );
nor U108200 ( n28859, n28860, n28861 );
nor U108201 ( n28862, n28674, n73872 );
nand U108202 ( n62155, n62163, n62164 );
nor U108203 ( n62163, n62167, n62168 );
nor U108204 ( n62164, n62165, n62166 );
nor U108205 ( n62167, n61979, n73873 );
nand U108206 ( n12268, n12275, n12277 );
nand U108207 ( n12275, n12253, n75200 );
nand U108208 ( n12277, n76729, n12278 );
nand U108209 ( n9031, n12265, n12267 );
nor U108210 ( n12265, n12285, n12287 );
nor U108211 ( n12267, n12268, n12269 );
nor U108212 ( n12285, n74869, n76735 );
nor U108213 ( n70766, n70575, n73850 );
nand U108214 ( n70755, n70763, n70764 );
nor U108215 ( n70763, n70767, n70768 );
nor U108216 ( n70764, n70765, n70766 );
nor U108217 ( n70767, n70579, n73871 );
nor U108218 ( n36040, n35849, n74229 );
nand U108219 ( n36029, n36037, n36038 );
nor U108220 ( n36037, n36041, n36042 );
nor U108221 ( n36038, n36039, n36040 );
nor U108222 ( n36041, n35853, n74238 );
nand U108223 ( n40406, n40437, n2199 );
nand U108224 ( n7326, n23200, n23201 );
nor U108225 ( n23200, n23210, n23211 );
nor U108226 ( n23201, n23202, n23203 );
nor U108227 ( n23210, n23248, n23152 );
nand U108228 ( n11816, n64684, n64685 );
nor U108229 ( n64684, n64727, n64728 );
nor U108230 ( n64685, n64686, n64687 );
nor U108231 ( n64727, n75306, n64640 );
nand U108232 ( n14061, n56321, n56322 );
nor U108233 ( n56321, n56331, n56332 );
nor U108234 ( n56322, n56323, n56324 );
nor U108235 ( n56331, n56369, n56273 );
nor U108236 ( n62638, n74492, n62738 );
nand U108237 ( n5081, n30525, n30526 );
nor U108238 ( n30525, n30568, n30569 );
nor U108239 ( n30526, n30527, n30528 );
nor U108240 ( n30568, n75317, n30481 );
nor U108241 ( n28838, n28682, n73774 );
nor U108242 ( n62143, n61987, n73775 );
nor U108243 ( n70743, n70587, n73773 );
nor U108244 ( n36017, n35861, n74126 );
nand U108245 ( n33184, n32219, n32218 );
nor U108246 ( n33166, n33182, n33183 );
nor U108247 ( n33182, n32714, n33187 );
nor U108248 ( n33183, n32712, n33184 );
nand U108249 ( n33187, n32216, n32215 );
nor U108250 ( n28872, n28876, n28877 );
nor U108251 ( n28876, n28695, n73869 );
nor U108252 ( n28877, n28694, n73847 );
nor U108253 ( n62177, n62181, n62182 );
nor U108254 ( n62181, n62000, n73870 );
nor U108255 ( n62182, n61999, n73848 );
nand U108256 ( n46893, n45911, n45910 );
nor U108257 ( n46880, n46891, n46892 );
nor U108258 ( n46891, n46415, n46896 );
nor U108259 ( n46892, n46413, n46893 );
nand U108260 ( n46896, n45922, n45921 );
nor U108261 ( n70777, n70781, n70782 );
nor U108262 ( n70781, n70600, n73868 );
nor U108263 ( n70782, n70599, n73844 );
nor U108264 ( n36051, n36055, n36056 );
nor U108265 ( n36055, n35874, n74237 );
nor U108266 ( n36056, n35873, n74227 );
nand U108267 ( n67940, n66862, n66861 );
nand U108268 ( n25937, n24986, n24985 );
nand U108269 ( n59075, n58121, n58120 );
nor U108270 ( n67927, n67938, n67939 );
nor U108271 ( n67938, n67479, n67943 );
nor U108272 ( n67939, n67477, n67940 );
nand U108273 ( n67943, n66873, n66872 );
nor U108274 ( n25924, n25935, n25936 );
nor U108275 ( n25935, n25474, n25940 );
nor U108276 ( n25936, n25472, n25937 );
nand U108277 ( n25940, n24997, n24996 );
nor U108278 ( n59062, n59073, n59074 );
nor U108279 ( n59073, n58611, n59078 );
nor U108280 ( n59074, n58609, n59075 );
nand U108281 ( n59078, n58132, n58131 );
nand U108282 ( n13444, n12209, n12208 );
nor U108283 ( n13422, n13442, n13443 );
nor U108284 ( n13442, n13060, n13448 );
nor U108285 ( n13443, n13055, n13444 );
nand U108286 ( n13448, n12205, n12204 );
nor U108287 ( n28833, n28673, n73795 );
nor U108288 ( n62138, n61978, n73796 );
nor U108289 ( n61967, n61970, n73677 );
nor U108290 ( n28662, n28665, n73678 );
nor U108291 ( n70738, n70578, n73794 );
nand U108292 ( n23211, n23212, n23213 );
nand U108293 ( n23212, n164, n22814 );
or U108294 ( n23213, n73394, n23160 );
nand U108295 ( n56332, n56333, n56334 );
nand U108296 ( n56333, n437, n55928 );
or U108297 ( n56334, n73393, n56281 );
nor U108298 ( n36012, n35852, n74142 );
nor U108299 ( n70567, n70570, n73674 );
nor U108300 ( n28855, n28660, n73862 );
nor U108301 ( n62160, n61965, n73863 );
nor U108302 ( n35841, n35844, n74006 );
nor U108303 ( n70760, n70565, n73861 );
nor U108304 ( n36034, n35839, n74233 );
nor U108305 ( n28843, n28844, n28845 );
nor U108306 ( n28845, n27016, n73777 );
nor U108307 ( n28844, n28691, n73792 );
nor U108308 ( n62148, n62149, n62150 );
nor U108309 ( n62150, n60157, n73778 );
nor U108310 ( n62149, n61996, n73793 );
nor U108311 ( n70748, n70749, n70750 );
nor U108312 ( n70750, n69013, n73776 );
nor U108313 ( n70749, n70596, n73791 );
nor U108314 ( n36022, n36023, n36024 );
nor U108315 ( n36024, n34259, n74127 );
nor U108316 ( n36023, n35870, n74137 );
nor U108317 ( n28840, n28686, n73763 );
nor U108318 ( n62145, n61991, n73764 );
nor U108319 ( n70745, n70591, n73761 );
nor U108320 ( n36019, n35865, n74121 );
not U108321 ( n2400, n17917 );
xor U108322 ( n9425, n74964, n11759 );
nor U108323 ( n11759, n11760, n74924 );
not U108324 ( n4760, n8480 );
nor U108325 ( n12167, n74512, n12184 );
nor U108326 ( n12328, n74450, n12375 );
nor U108327 ( n12282, n5310, n12284 );
nor U108328 ( n12104, n5309, n12103 );
nor U108329 ( n12387, n73107, n12437 );
nor U108330 ( n11802, n74880, n11830 );
not U108331 ( n5307, n12032 );
nor U108332 ( n12563, n73072, n12573 );
nor U108333 ( n12445, n73097, n12489 );
nor U108334 ( n11993, n74677, n12045 );
nor U108335 ( n11928, n74737, n11980 );
nor U108336 ( n11865, n74808, n11902 );
nor U108337 ( n12513, n73087, n12537 );
or U108338 ( n12184, n12238, n12187 );
nand U108339 ( n9866, n8652, n8653 );
nor U108340 ( n8652, n8669, n8670 );
nor U108341 ( n8653, n8654, n8655 );
nor U108342 ( n8669, n74997, n8414 );
nand U108343 ( n9756, n9363, n9364 );
nor U108344 ( n9364, n9365, n9367 );
nor U108345 ( n9363, n9384, n9385 );
nand U108346 ( n9365, n9375, n9377 );
not U108347 ( n253, n45396 );
nand U108348 ( n9796, n9105, n9107 );
nor U108349 ( n9105, n9119, n9120 );
nor U108350 ( n9107, n9108, n9109 );
nand U108351 ( n9120, n9122, n9123 );
nand U108352 ( n8720, n8722, n8723 );
nand U108353 ( n8723, n8724, n76742 );
nand U108354 ( n8722, n8708, n8725 );
nor U108355 ( n8724, n5274, n8708 );
nand U108356 ( n8592, n8593, n8594 );
nand U108357 ( n8594, n8595, n76742 );
nand U108358 ( n8593, n8573, n8597 );
nor U108359 ( n8595, n5272, n8573 );
nand U108360 ( n9856, n8717, n8718 );
nor U108361 ( n8717, n8733, n8734 );
nor U108362 ( n8718, n8719, n8720 );
nor U108363 ( n8733, n75201, n8414 );
nand U108364 ( n9876, n8588, n8589 );
nor U108365 ( n8588, n8607, n8608 );
nor U108366 ( n8589, n8590, n8592 );
nor U108367 ( n8607, n75235, n8414 );
nand U108368 ( n9826, n8910, n8912 );
nor U108369 ( n8912, n8913, n8914 );
nor U108370 ( n8910, n8923, n8924 );
nand U108371 ( n8913, n8920, n8789 );
nand U108372 ( n9786, n9169, n9170 );
nor U108373 ( n9170, n9172, n9173 );
nor U108374 ( n9169, n9183, n9184 );
nand U108375 ( n9172, n9179, n8789 );
nand U108376 ( n9816, n8974, n8975 );
nor U108377 ( n8975, n8977, n8978 );
nor U108378 ( n8974, n8988, n8989 );
nand U108379 ( n8977, n8984, n8789 );
nand U108380 ( n9846, n8778, n8779 );
nor U108381 ( n8779, n8780, n8782 );
nor U108382 ( n8778, n8794, n8795 );
nand U108383 ( n8780, n8788, n8789 );
nor U108384 ( n28830, n22674, n73759 );
nor U108385 ( n62135, n55787, n73760 );
nor U108386 ( n70735, n63953, n73758 );
nor U108387 ( n36009, n29997, n74107 );
xor U108388 ( n38313, n72956, n39449 );
nor U108389 ( n28868, n28682, n73856 );
nor U108390 ( n62173, n61987, n73857 );
nor U108391 ( n70773, n70587, n73855 );
nor U108392 ( n36047, n35861, n74230 );
nor U108393 ( n28863, n28673, n73878 );
nor U108394 ( n62168, n61978, n73879 );
nor U108395 ( n28826, n28665, n73769 );
nor U108396 ( n62131, n61970, n73770 );
nor U108397 ( n70768, n70578, n73877 );
nor U108398 ( n36042, n35852, n74242 );
nor U108399 ( n70731, n70570, n73767 );
not U108400 ( n7405, n43338 );
nor U108401 ( n45880, n74515, n45894 );
nor U108402 ( n46011, n74451, n46049 );
nor U108403 ( n36005, n35844, n74124 );
nor U108404 ( n45963, n7965, n45965 );
nor U108405 ( n45834, n7964, n45833 );
nor U108406 ( n46058, n73108, n46093 );
not U108407 ( n7962, n45776 );
nor U108408 ( n46194, n73073, n46202 );
nor U108409 ( n46100, n73098, n46135 );
nor U108410 ( n45727, n74680, n45787 );
nor U108411 ( n45560, n74891, n45606 );
nor U108412 ( n45694, n74740, n45717 );
nor U108413 ( n45640, n74810, n45650 );
nor U108414 ( n46154, n73089, n46174 );
xor U108415 ( n43367, n74967, n45530 );
nor U108416 ( n45530, n45531, n74931 );
or U108417 ( n45894, n45928, n45896 );
nand U108418 ( n16601, n42715, n42716 );
nor U108419 ( n42715, n42729, n42730 );
nor U108420 ( n42716, n42717, n42718 );
nor U108421 ( n42729, n74998, n42500 );
nor U108422 ( n50588, n50030, n73425 );
nand U108423 ( n14845, n76592, n11600 );
xor U108424 ( n54614, n72936, n66010 );
xor U108425 ( n32207, n32218, n74635 );
nand U108426 ( n16491, n43316, n43317 );
nor U108427 ( n43317, n43318, n43319 );
nor U108428 ( n43316, n43333, n43334 );
nand U108429 ( n43318, n43326, n43327 );
nand U108430 ( n16531, n43096, n43097 );
nor U108431 ( n43096, n43107, n43108 );
nor U108432 ( n43097, n43098, n43099 );
nand U108433 ( n43108, n43109, n43110 );
xor U108434 ( n12194, n12208, n74599 );
xor U108435 ( n45902, n45910, n74524 );
nand U108436 ( n16561, n42926, n42927 );
nor U108437 ( n42927, n42928, n42929 );
nor U108438 ( n42926, n42936, n42937 );
nand U108439 ( n42928, n42934, n42829 );
nand U108440 ( n16521, n43147, n43148 );
nor U108441 ( n43148, n43149, n43150 );
nor U108442 ( n43147, n43158, n43159 );
nand U108443 ( n43149, n43155, n42829 );
nor U108444 ( n28873, n28874, n28875 );
nor U108445 ( n28875, n27016, n73859 );
nor U108446 ( n28874, n28691, n73875 );
nor U108447 ( n62178, n62179, n62180 );
nor U108448 ( n62180, n60157, n73860 );
nor U108449 ( n62179, n61996, n73876 );
nand U108450 ( n16551, n42991, n42992 );
nor U108451 ( n42992, n42993, n42994 );
nor U108452 ( n42991, n43002, n43003 );
nand U108453 ( n42993, n42999, n42829 );
nand U108454 ( n16581, n42820, n42821 );
nor U108455 ( n42821, n42822, n42823 );
nor U108456 ( n42820, n42833, n42834 );
nand U108457 ( n42822, n42828, n42829 );
xor U108458 ( n66853, n66861, n74546 );
xor U108459 ( n24977, n24985, n74547 );
xor U108460 ( n58112, n58120, n74548 );
nor U108461 ( n70778, n70779, n70780 );
nor U108462 ( n70780, n69013, n73858 );
nor U108463 ( n70779, n70596, n73874 );
nor U108464 ( n36052, n36053, n36054 );
nor U108465 ( n36054, n34259, n74231 );
nor U108466 ( n36053, n35870, n74239 );
nor U108467 ( n28870, n28686, n73845 );
nor U108468 ( n62175, n61991, n73846 );
nor U108469 ( n70775, n70591, n73843 );
nor U108470 ( n36049, n35865, n74226 );
nand U108471 ( n32116, n32123, n32124 );
nand U108472 ( n32124, n32125, n76480 );
nand U108473 ( n32123, n32128, n76785 );
and U108474 ( n32125, n32126, n32127 );
and U108475 ( n32128, n32129, n32130 );
nand U108476 ( n12075, n12084, n12085 );
nand U108477 ( n12085, n12087, n76607 );
nand U108478 ( n12084, n12090, n76737 );
and U108479 ( n12087, n12088, n12089 );
and U108480 ( n12090, n12092, n12093 );
nand U108481 ( n45811, n45818, n45819 );
nand U108482 ( n45819, n45820, n76346 );
nand U108483 ( n45818, n45823, n76671 );
and U108484 ( n45820, n45821, n45822 );
and U108485 ( n45823, n45824, n45825 );
nor U108486 ( n28708, n22674, n73635 );
nor U108487 ( n62013, n55787, n73634 );
nor U108488 ( n70613, n63953, n73628 );
nor U108489 ( n35887, n29997, n73969 );
nand U108490 ( n66762, n66769, n66770 );
nand U108491 ( n66770, n66771, n76202 );
nand U108492 ( n66769, n66774, n76719 );
and U108493 ( n66771, n66772, n66773 );
nand U108494 ( n24884, n24891, n24892 );
nand U108495 ( n24892, n24893, n76526 );
nand U108496 ( n24891, n24896, n76767 );
and U108497 ( n24893, n24894, n24895 );
nand U108498 ( n58021, n58028, n58029 );
nand U108499 ( n58029, n58030, n76268 );
nand U108500 ( n58028, n58033, n76700 );
and U108501 ( n58030, n58031, n58032 );
and U108502 ( n66774, n66775, n66776 );
and U108503 ( n24896, n24897, n24898 );
and U108504 ( n58033, n58034, n58035 );
nand U108505 ( n16171, n44977, n44978 );
nor U108506 ( n44978, n44979, n44980 );
nor U108507 ( n44977, n44983, n44984 );
nor U108508 ( n44979, n43808, n44982 );
xor U108509 ( n48911, n72949, n64349 );
nand U108510 ( n71496, n71327, n71144 );
nand U108511 ( n71135, n71143, n71144 );
nand U108512 ( n13971, n57222, n57223 );
nor U108513 ( n57222, n57231, n57232 );
nor U108514 ( n57223, n57224, n57225 );
nor U108515 ( n57232, n56468, n57007 );
nand U108516 ( n7236, n24100, n24101 );
nor U108517 ( n24100, n24109, n24110 );
nor U108518 ( n24101, n24102, n24103 );
nor U108519 ( n24110, n23344, n23883 );
nand U108520 ( n4991, n31394, n31395 );
nor U108521 ( n31394, n31403, n31404 );
nor U108522 ( n31395, n31396, n31397 );
nor U108523 ( n31404, n75321, n31181 );
nand U108524 ( n11726, n65644, n65645 );
nor U108525 ( n65644, n65653, n65654 );
nor U108526 ( n65645, n65646, n65647 );
nor U108527 ( n65654, n75310, n65435 );
nand U108528 ( n5011, n31228, n31229 );
nor U108529 ( n31228, n31237, n31238 );
nor U108530 ( n31229, n31230, n31231 );
nor U108531 ( n31238, n75311, n31181 );
nand U108532 ( n5001, n31313, n31314 );
nor U108533 ( n31313, n31322, n31323 );
nor U108534 ( n31314, n31315, n31316 );
nor U108535 ( n31323, n75317, n31181 );
nand U108536 ( n7246, n24019, n24020 );
nor U108537 ( n24019, n24028, n24029 );
nor U108538 ( n24020, n24021, n24022 );
nor U108539 ( n24029, n23248, n23883 );
nand U108540 ( n13991, n57060, n57061 );
nor U108541 ( n57060, n57069, n57070 );
nor U108542 ( n57061, n57062, n57063 );
nor U108543 ( n57070, n56272, n57007 );
nand U108544 ( n13981, n57141, n57142 );
nor U108545 ( n57141, n57150, n57151 );
nor U108546 ( n57142, n57143, n57144 );
nor U108547 ( n57151, n56369, n57007 );
nand U108548 ( n7256, n23938, n23939 );
nor U108549 ( n23938, n23947, n23948 );
nor U108550 ( n23939, n23940, n23941 );
nor U108551 ( n23948, n23151, n23883 );
nand U108552 ( n13951, n57374, n57375 );
nor U108553 ( n57374, n57383, n57384 );
nor U108554 ( n57375, n57376, n57377 );
nor U108555 ( n57384, n6649, n56217 );
nand U108556 ( n13941, n57395, n57396 );
nor U108557 ( n57395, n57404, n57405 );
nor U108558 ( n57396, n57397, n57398 );
nor U108559 ( n57405, n6664, n56217 );
nand U108560 ( n13931, n57415, n57416 );
nor U108561 ( n57415, n57424, n57425 );
nor U108562 ( n57416, n57417, n57418 );
nor U108563 ( n57425, n6685, n56217 );
nand U108564 ( n7226, n24181, n24182 );
nor U108565 ( n24181, n24190, n24191 );
nor U108566 ( n24182, n24183, n24184 );
nor U108567 ( n24191, n23441, n23883 );
nand U108568 ( n7216, n24249, n24250 );
nor U108569 ( n24249, n24258, n24259 );
nor U108570 ( n24250, n24251, n24252 );
nor U108571 ( n24259, n4017, n23096 );
nand U108572 ( n7206, n24272, n24273 );
nor U108573 ( n24272, n24281, n24282 );
nor U108574 ( n24273, n24274, n24275 );
nor U108575 ( n24282, n4032, n23096 );
nand U108576 ( n7196, n24292, n24293 );
nor U108577 ( n24292, n24301, n24302 );
nor U108578 ( n24293, n24294, n24295 );
nor U108579 ( n24302, n4053, n23096 );
xor U108580 ( n32112, n32126, n74652 );
nand U108581 ( n11746, n65482, n65483 );
nor U108582 ( n65482, n65491, n65492 );
nor U108583 ( n65483, n65484, n65485 );
nor U108584 ( n65492, n75304, n65435 );
nand U108585 ( n11736, n65563, n65564 );
nor U108586 ( n65563, n65572, n65573 );
nor U108587 ( n65564, n65565, n65566 );
nor U108588 ( n65573, n75306, n65435 );
nand U108589 ( n13961, n57303, n57304 );
nor U108590 ( n57303, n57312, n57313 );
nor U108591 ( n57304, n57305, n57306 );
nor U108592 ( n57313, n56563, n57007 );
nand U108593 ( n4981, n31475, n31476 );
nor U108594 ( n31475, n31484, n31485 );
nor U108595 ( n31476, n31477, n31478 );
nor U108596 ( n31485, n75320, n31181 );
nand U108597 ( n4971, n31543, n31544 );
nor U108598 ( n31543, n31552, n31553 );
nor U108599 ( n31544, n31545, n31546 );
nor U108600 ( n31552, n75314, n31181 );
nand U108601 ( n4961, n31564, n31565 );
nor U108602 ( n31564, n31573, n31574 );
nor U108603 ( n31565, n31566, n31567 );
nor U108604 ( n31573, n75313, n31181 );
nand U108605 ( n4951, n31588, n31589 );
nor U108606 ( n31588, n31597, n31598 );
nor U108607 ( n31589, n31590, n31591 );
nor U108608 ( n31597, n75296, n31181 );
nand U108609 ( n11716, n65725, n65726 );
nor U108610 ( n65725, n65734, n65735 );
nor U108611 ( n65726, n65727, n65728 );
nor U108612 ( n65735, n75309, n65435 );
nand U108613 ( n11706, n65833, n65834 );
nor U108614 ( n65833, n65842, n65843 );
nor U108615 ( n65834, n65835, n65836 );
nor U108616 ( n65842, n75290, n65435 );
nand U108617 ( n11696, n65854, n65855 );
nor U108618 ( n65854, n65863, n65864 );
nor U108619 ( n65855, n65856, n65857 );
nor U108620 ( n65863, n75293, n65435 );
nand U108621 ( n11686, n65874, n65875 );
nor U108622 ( n65874, n65883, n65884 );
nor U108623 ( n65875, n65876, n65877 );
nor U108624 ( n65883, n75292, n65435 );
xor U108625 ( n12070, n12088, n74625 );
nand U108626 ( n32029, n32033, n76480 );
and U108627 ( n32033, n32034, n32035 );
nand U108628 ( n38556, n76446, n75247 );
xor U108629 ( n33509, n76471, n73197 );
xor U108630 ( n45807, n45821, n74585 );
xor U108631 ( n32429, n33469, n33509 );
nor U108632 ( n61973, n55787, n73660 );
nor U108633 ( n28668, n22674, n73661 );
nor U108634 ( n28856, n28665, n73851 );
nor U108635 ( n62161, n61970, n73852 );
nor U108636 ( n70573, n63953, n73659 );
nand U108637 ( n66632, n66636, n76202 );
and U108638 ( n66636, n66637, n66638 );
nand U108639 ( n24797, n24801, n76526 );
and U108640 ( n24801, n24802, n24803 );
nand U108641 ( n57931, n57935, n76268 );
and U108642 ( n57935, n57936, n57937 );
xor U108643 ( n66715, n66772, n74595 );
xor U108644 ( n24880, n24894, n74596 );
xor U108645 ( n58017, n58031, n74597 );
nor U108646 ( n35847, n29997, n74002 );
nor U108647 ( n70761, n70570, n73849 );
nor U108648 ( n36035, n35844, n74228 );
xor U108649 ( n48449, n72955, n63267 );
not U108650 ( n4229, n28551 );
not U108651 ( n6862, n61856 );
not U108652 ( n6007, n70456 );
not U108653 ( n3392, n35730 );
and U108654 ( n68264, n68188, n68279 );
nand U108655 ( n68279, n75990, n73187 );
and U108656 ( n47233, n47157, n47248 );
nand U108657 ( n47248, n76006, n73178 );
and U108658 ( n26263, n26187, n26278 );
nand U108659 ( n26278, n76027, n73188 );
and U108660 ( n59402, n59326, n59417 );
nand U108661 ( n59417, n75998, n73189 );
nor U108662 ( n13284, n74586, n76603 );
nand U108663 ( n31969, n32583, n32584 );
nand U108664 ( n32583, n32589, n74591 );
nand U108665 ( n32584, n3077, n32585 );
nand U108666 ( n32585, n32586, n32587 );
not U108667 ( n3058, n31869 );
or U108668 ( n32170, n32172, n75813 );
and U108669 ( n75813, n31841, n75191 );
nand U108670 ( n31960, n31891, n31968 );
nand U108671 ( n31968, n3055, n31894 );
nand U108672 ( n66572, n67348, n67349 );
nand U108673 ( n67348, n67354, n74593 );
nand U108674 ( n67349, n5678, n67350 );
nand U108675 ( n67350, n67351, n67352 );
nand U108676 ( n45648, n46287, n46288 );
nand U108677 ( n46287, n46293, n74648 );
nand U108678 ( n46288, n7463, n46289 );
nand U108679 ( n46289, n46290, n46291 );
nand U108680 ( n24737, n25341, n25342 );
nand U108681 ( n25341, n25347, n74592 );
nand U108682 ( n25342, n3920, n25343 );
nand U108683 ( n25343, n25344, n25345 );
nand U108684 ( n57871, n58480, n58481 );
nand U108685 ( n58480, n58486, n74594 );
nand U108686 ( n58481, n6553, n58482 );
nand U108687 ( n58482, n58483, n58484 );
nor U108688 ( n54382, n54341, n73538 );
nand U108689 ( n54376, n54377, n54378 );
nor U108690 ( n54378, n54379, n54380 );
nor U108691 ( n54377, n54381, n54382 );
nor U108692 ( n54379, n54338, n73548 );
not U108693 ( n7433, n45567 );
not U108694 ( n3902, n24655 );
not U108695 ( n6534, n57791 );
not U108696 ( n5659, n66492 );
or U108697 ( n66816, n66818, n75814 );
and U108698 ( n75814, n66464, n75192 );
or U108699 ( n45865, n45867, n75815 );
and U108700 ( n75815, n45540, n74772 );
or U108701 ( n24940, n24942, n75816 );
and U108702 ( n75816, n24627, n75193 );
or U108703 ( n58075, n58077, n75817 );
and U108704 ( n75817, n57759, n75194 );
nand U108705 ( n32255, n32238, n32268 );
nand U108706 ( n32268, n3055, n32240 );
xnor U108707 ( n67085, n68220, n68264 );
xnor U108708 ( n46121, n47189, n47233 );
or U108709 ( n32253, n32255, n75818 );
and U108710 ( n75818, n31841, n75195 );
xnor U108711 ( n25187, n26219, n26263 );
xnor U108712 ( n58323, n59358, n59402 );
nand U108713 ( n24728, n24679, n24736 );
nand U108714 ( n24736, n3899, n24682 );
nand U108715 ( n66563, n66514, n66571 );
nand U108716 ( n66571, n5657, n66517 );
nand U108717 ( n57862, n57813, n57870 );
nand U108718 ( n57870, n6532, n57816 );
and U108719 ( n32238, n31969, n32269 );
nand U108720 ( n32269, n76779, n32232 );
nand U108721 ( n45706, n45678, n45725 );
nand U108722 ( n45725, n7430, n45681 );
nand U108723 ( n32107, n32078, n32135 );
nand U108724 ( n32135, n3055, n32081 );
or U108725 ( n32105, n32107, n75819 );
and U108726 ( n75819, n31841, n74688 );
not U108727 ( n818, n41460 );
nand U108728 ( n45943, n45913, n45956 );
nand U108729 ( n45956, n7430, n45928 );
nand U108730 ( n66894, n66864, n66907 );
nand U108731 ( n66907, n5657, n66878 );
nand U108732 ( n25018, n24988, n25031 );
nand U108733 ( n25031, n3899, n25002 );
nand U108734 ( n58153, n58123, n58166 );
nand U108735 ( n58166, n6532, n58137 );
and U108736 ( n66864, n66572, n66908 );
nand U108737 ( n66908, n76713, n66870 );
and U108738 ( n45913, n45648, n45957 );
nand U108739 ( n45957, n76665, n45919 );
and U108740 ( n24988, n24737, n25032 );
nand U108741 ( n25032, n76761, n24994 );
and U108742 ( n58123, n57871, n58167 );
nand U108743 ( n58167, n76694, n58129 );
or U108744 ( n66892, n66894, n75820 );
and U108745 ( n75820, n66464, n75196 );
or U108746 ( n45941, n45943, n75821 );
and U108747 ( n75821, n45540, n75197 );
or U108748 ( n25016, n25018, n75822 );
and U108749 ( n75822, n24627, n75198 );
or U108750 ( n58151, n58153, n75823 );
and U108751 ( n75823, n57759, n75199 );
nand U108752 ( n45639, n45589, n45647 );
nand U108753 ( n45647, n7430, n45592 );
nand U108754 ( n66710, n66681, n66781 );
nand U108755 ( n66781, n5657, n66684 );
nand U108756 ( n24875, n24846, n24903 );
nand U108757 ( n24903, n3899, n24849 );
nand U108758 ( n58012, n57980, n58040 );
nand U108759 ( n58040, n6532, n57983 );
or U108760 ( n66708, n66710, n75824 );
and U108761 ( n75824, n66464, n74687 );
or U108762 ( n24873, n24875, n75825 );
and U108763 ( n75825, n24627, n74689 );
or U108764 ( n58010, n58012, n75826 );
and U108765 ( n75826, n57759, n74690 );
nand U108766 ( n32028, n31999, n32048 );
nand U108767 ( n32048, n3055, n32002 );
nor U108768 ( n28887, n28664, n73713 );
nor U108769 ( n62192, n61969, n73712 );
nand U108770 ( n28881, n28882, n28883 );
nor U108771 ( n28883, n28884, n28885 );
nor U108772 ( n28882, n28886, n28887 );
nor U108773 ( n28884, n28661, n73739 );
nand U108774 ( n62186, n62187, n62188 );
nor U108775 ( n62188, n62189, n62190 );
nor U108776 ( n62187, n62191, n62192 );
nor U108777 ( n62189, n61966, n73738 );
or U108778 ( n32318, n32320, n75827 );
and U108779 ( n75827, n31841, n74615 );
nor U108780 ( n67223, n829, n842 );
nand U108781 ( n45802, n45773, n45830 );
nand U108782 ( n45830, n7430, n45776 );
or U108783 ( n45800, n45802, n75828 );
and U108784 ( n75828, n45540, n75202 );
nor U108785 ( n70792, n70569, n73710 );
nand U108786 ( n66631, n66602, n66651 );
nand U108787 ( n66651, n5657, n66605 );
nand U108788 ( n24796, n24767, n24816 );
nand U108789 ( n24816, n3899, n24770 );
nand U108790 ( n57930, n57901, n57950 );
nand U108791 ( n57950, n6532, n57904 );
nand U108792 ( n70786, n70787, n70788 );
nor U108793 ( n70788, n70789, n70790 );
nor U108794 ( n70787, n70791, n70792 );
nor U108795 ( n70789, n70566, n73737 );
nor U108796 ( n36066, n35843, n74023 );
nand U108797 ( n36060, n36061, n36062 );
nor U108798 ( n36062, n36063, n36064 );
nor U108799 ( n36061, n36065, n36066 );
nor U108800 ( n36063, n35840, n74042 );
or U108801 ( n66957, n66959, n75829 );
and U108802 ( n75829, n66464, n74616 );
or U108803 ( n46017, n46019, n75830 );
and U108804 ( n75830, n45540, n74607 );
or U108805 ( n25081, n25083, n75831 );
and U108806 ( n75831, n24627, n74617 );
or U108807 ( n58216, n58218, n75832 );
and U108808 ( n75832, n57759, n74618 );
nand U108809 ( n54362, n44136, n73497 );
nor U108810 ( n54396, n54362, n73534 );
nand U108811 ( n54390, n54391, n54392 );
nor U108812 ( n54392, n54393, n54394 );
nor U108813 ( n54391, n54395, n54396 );
nor U108814 ( n54394, n54358, n73539 );
nand U108815 ( n32532, n76779, n74699 );
nand U108816 ( n4491, n32483, n32484 );
nor U108817 ( n32483, n32498, n32499 );
nor U108818 ( n32484, n32485, n32486 );
nor U108819 ( n32498, n73194, n76781 );
nand U108820 ( n32495, n32496, n32497 );
nand U108821 ( n32497, n76780, n74478 );
nor U108822 ( n28901, n28685, n73671 );
nor U108823 ( n62206, n61990, n73670 );
nand U108824 ( n28895, n28896, n28897 );
nor U108825 ( n28897, n28898, n28899 );
nor U108826 ( n28896, n28900, n28901 );
nor U108827 ( n28899, n28681, n73716 );
nand U108828 ( n62200, n62201, n62202 );
nor U108829 ( n62202, n62203, n62204 );
nor U108830 ( n62201, n62205, n62206 );
nor U108831 ( n62204, n61986, n73715 );
nor U108832 ( n70806, n70590, n73666 );
nor U108833 ( n36080, n35864, n74012 );
nand U108834 ( n67188, n76713, n74700 );
nand U108835 ( n25290, n76761, n74701 );
nand U108836 ( n58426, n76694, n74702 );
nand U108837 ( n46236, n76665, n74717 );
nand U108838 ( n70800, n70801, n70802 );
nor U108839 ( n70802, n70803, n70804 );
nor U108840 ( n70801, n70805, n70806 );
nor U108841 ( n70804, n70586, n73714 );
nand U108842 ( n36074, n36075, n36076 );
nor U108843 ( n36076, n36077, n36078 );
nor U108844 ( n36075, n36079, n36080 );
nor U108845 ( n36078, n35860, n74024 );
nand U108846 ( n11226, n67139, n67140 );
nor U108847 ( n67139, n67154, n67155 );
nor U108848 ( n67140, n67141, n67142 );
nor U108849 ( n67154, n73193, n76715 );
nand U108850 ( n6736, n25241, n25242 );
nor U108851 ( n25241, n25256, n25257 );
nor U108852 ( n25242, n25243, n25244 );
nor U108853 ( n25256, n74694, n76763 );
nand U108854 ( n13471, n58377, n58378 );
nor U108855 ( n58377, n58392, n58393 );
nor U108856 ( n58378, n58379, n58380 );
nor U108857 ( n58392, n74693, n76696 );
nand U108858 ( n15716, n46175, n46176 );
nor U108859 ( n46175, n46190, n46191 );
nor U108860 ( n46176, n46177, n46178 );
nor U108861 ( n46190, n74726, n76667 );
nand U108862 ( n67151, n67152, n67153 );
nand U108863 ( n67153, n76714, n74479 );
nand U108864 ( n25253, n25254, n25255 );
nand U108865 ( n25255, n76762, n74480 );
nand U108866 ( n58389, n58390, n58391 );
nand U108867 ( n58391, n76695, n74481 );
nand U108868 ( n46187, n46188, n46189 );
nand U108869 ( n46189, n76666, n74473 );
nand U108870 ( n71144, n72840, n72841 );
nor U108871 ( n72840, n72844, n72845 );
nor U108872 ( n72841, n72842, n72843 );
nor U108873 ( n72845, n74405, n73026 );
nor U108874 ( n54386, n54347, n73541 );
nand U108875 ( n54375, n54383, n54384 );
nor U108876 ( n54383, n54387, n54388 );
nor U108877 ( n54384, n54385, n54386 );
nor U108878 ( n54387, n54351, n73546 );
nor U108879 ( n54477, n43268, n74132 );
nand U108880 ( n54467, n54475, n54476 );
nor U108881 ( n54475, n54479, n54480 );
nor U108882 ( n54476, n54477, n54478 );
nor U108883 ( n54480, n54350, n74160 );
nor U108884 ( n72842, n73095, n71105 );
xnor U108885 ( n67106, n68268, n68311 );
xor U108886 ( n68311, n74695, n76197 );
xnor U108887 ( n25208, n26267, n26310 );
xor U108888 ( n26310, n74697, n76521 );
xnor U108889 ( n58344, n59406, n59449 );
xor U108890 ( n59449, n74698, n76263 );
nor U108891 ( n68304, n68306, n76868 );
nor U108892 ( n68306, n68307, n68308 );
nand U108893 ( n68307, n68325, n68326 );
nand U108894 ( n68308, n68309, n68310 );
nor U108895 ( n26303, n26305, n76903 );
nor U108896 ( n26305, n26306, n26307 );
nand U108897 ( n26306, n26324, n26325 );
nand U108898 ( n26307, n26308, n26309 );
nor U108899 ( n59442, n59444, n76877 );
nor U108900 ( n59444, n59445, n59446 );
nand U108901 ( n59445, n59463, n59464 );
nand U108902 ( n59446, n59447, n59448 );
xnor U108903 ( n46142, n47237, n47280 );
xor U108904 ( n47280, n74659, n76341 );
xnor U108905 ( n32450, n33513, n33555 );
xor U108906 ( n33555, n74696, n76470 );
nor U108907 ( n28891, n28670, n73721 );
nor U108908 ( n62196, n61975, n73720 );
nand U108909 ( n28880, n28888, n28889 );
nor U108910 ( n28888, n28892, n28893 );
nor U108911 ( n28889, n28890, n28891 );
nor U108912 ( n28892, n28674, n73733 );
nand U108913 ( n62185, n62193, n62194 );
nor U108914 ( n62193, n62197, n62198 );
nor U108915 ( n62194, n62195, n62196 );
nor U108916 ( n62197, n61979, n73732 );
nor U108917 ( n33548, n33550, n76894 );
nor U108918 ( n33550, n33551, n33552 );
nand U108919 ( n33551, n33569, n33570 );
nand U108920 ( n33552, n33553, n33554 );
nor U108921 ( n47273, n47275, n76328 );
nor U108922 ( n47275, n47276, n47277 );
nand U108923 ( n47276, n47294, n47295 );
nand U108924 ( n47277, n47278, n47279 );
nor U108925 ( n70796, n70575, n73719 );
nand U108926 ( n70785, n70793, n70794 );
nor U108927 ( n70793, n70797, n70798 );
nor U108928 ( n70794, n70795, n70796 );
nor U108929 ( n70797, n70579, n73731 );
nor U108930 ( n36070, n35849, n74030 );
nand U108931 ( n36059, n36067, n36068 );
nor U108932 ( n36067, n36071, n36072 );
nor U108933 ( n36068, n36069, n36070 );
nor U108934 ( n36071, n35853, n74036 );
nor U108935 ( n54564, n54341, n73576 );
nand U108936 ( n54558, n54559, n54560 );
nor U108937 ( n54560, n54561, n54562 );
nor U108938 ( n54559, n54563, n54564 );
nor U108939 ( n54561, n54338, n73591 );
not U108940 ( n4896, n11877 );
nor U108941 ( n54471, n54338, n74148 );
nand U108942 ( n54468, n54469, n54470 );
nor U108943 ( n54469, n54473, n54474 );
nor U108944 ( n54470, n54471, n54472 );
nor U108945 ( n54473, n54342, n74144 );
nand U108946 ( n54358, n44132, n73497 );
nor U108947 ( n54486, n54358, n74130 );
nand U108948 ( n54482, n54483, n54484 );
nor U108949 ( n54483, n54487, n54488 );
nor U108950 ( n54484, n54485, n54486 );
nor U108951 ( n54487, n54363, n74135 );
nor U108952 ( n54397, n54401, n54402 );
nor U108953 ( n54401, n54372, n73540 );
nor U108954 ( n54402, n54371, n73536 );
nand U108955 ( n9766, n9304, n9305 );
nor U108956 ( n9304, n9322, n9323 );
nor U108957 ( n9305, n9307, n9308 );
nand U108958 ( n9323, n9324, n9325 );
nor U108959 ( n28902, n28906, n28907 );
nor U108960 ( n28906, n28695, n73718 );
nor U108961 ( n28907, n28694, n73706 );
nor U108962 ( n62207, n62211, n62212 );
nor U108963 ( n62211, n62000, n73717 );
nor U108964 ( n62212, n61999, n73705 );
nand U108965 ( n4506, n32423, n32424 );
nor U108966 ( n32423, n32438, n32439 );
nor U108967 ( n32424, n32425, n32426 );
nor U108968 ( n32438, n74750, n76781 );
nand U108969 ( n32435, n32436, n32437 );
nand U108970 ( n32437, n76780, n73102 );
nor U108971 ( n70807, n70811, n70812 );
nor U108972 ( n70811, n70600, n73711 );
nor U108973 ( n70812, n70599, n73701 );
nand U108974 ( n32506, n32512, n32513 );
nand U108975 ( n32513, n32494, n74478 );
or U108976 ( n32512, n74478, n32496 );
nor U108977 ( n36081, n36085, n36086 );
nor U108978 ( n36085, n35874, n74025 );
nor U108979 ( n36086, n35873, n74021 );
nand U108980 ( n4486, n32504, n32505 );
nor U108981 ( n32504, n32516, n32517 );
nor U108982 ( n32505, n32506, n32507 );
nor U108983 ( n32516, n74643, n76781 );
nand U108984 ( n11241, n67079, n67080 );
nor U108985 ( n67079, n67094, n67095 );
nor U108986 ( n67080, n67081, n67082 );
nor U108987 ( n67094, n74749, n76715 );
nand U108988 ( n15731, n46115, n46116 );
nor U108989 ( n46115, n46130, n46131 );
nor U108990 ( n46116, n46117, n46118 );
nor U108991 ( n46130, n75965, n76667 );
nand U108992 ( n6751, n25181, n25182 );
nor U108993 ( n25181, n25196, n25197 );
nor U108994 ( n25182, n25183, n25184 );
nor U108995 ( n25196, n74748, n76763 );
nand U108996 ( n13486, n58317, n58318 );
nor U108997 ( n58317, n58332, n58333 );
nor U108998 ( n58318, n58319, n58320 );
nor U108999 ( n58332, n74747, n76696 );
nand U109000 ( n67091, n67092, n67093 );
nand U109001 ( n67093, n76714, n73100 );
nand U109002 ( n46127, n46128, n46129 );
nand U109003 ( n46129, n76666, n73098 );
nand U109004 ( n25193, n25194, n25195 );
nand U109005 ( n25195, n76762, n73103 );
nand U109006 ( n58329, n58330, n58331 );
nand U109007 ( n58331, n76695, n73101 );
nand U109008 ( n32364, n32365, n32366 );
nand U109009 ( n32366, n76780, n74557 );
nor U109010 ( n54578, n54362, n73558 );
nand U109011 ( n54572, n54573, n54574 );
nor U109012 ( n54574, n54575, n54576 );
nor U109013 ( n54573, n54577, n54578 );
nor U109014 ( n54576, n54358, n73577 );
nand U109015 ( n67162, n67168, n67169 );
nand U109016 ( n67169, n67150, n74479 );
or U109017 ( n67168, n74479, n67152 );
nand U109018 ( n25264, n25270, n25271 );
nand U109019 ( n25271, n25252, n74480 );
or U109020 ( n25270, n74480, n25254 );
nand U109021 ( n58400, n58406, n58407 );
nand U109022 ( n58407, n58388, n74481 );
or U109023 ( n58406, n74481, n58390 );
nand U109024 ( n46198, n46204, n46205 );
nand U109025 ( n46205, n46186, n74473 );
or U109026 ( n46204, n74473, n46188 );
nand U109027 ( n11221, n67160, n67161 );
nor U109028 ( n67160, n67172, n67173 );
nor U109029 ( n67161, n67162, n67163 );
nor U109030 ( n67172, n74642, n76715 );
nand U109031 ( n6731, n25262, n25263 );
nor U109032 ( n25262, n25274, n25275 );
nor U109033 ( n25263, n25264, n25265 );
nor U109034 ( n25274, n74641, n76763 );
nand U109035 ( n13466, n58398, n58399 );
nor U109036 ( n58398, n58410, n58411 );
nor U109037 ( n58399, n58400, n58401 );
nor U109038 ( n58410, n74640, n76696 );
nand U109039 ( n15711, n46196, n46197 );
nor U109040 ( n46196, n46208, n46209 );
nor U109041 ( n46197, n46198, n46199 );
nor U109042 ( n46208, n74672, n76667 );
nand U109043 ( n67027, n67028, n67029 );
nand U109044 ( n67029, n76714, n74558 );
nand U109045 ( n46063, n46064, n46065 );
nand U109046 ( n46065, n76666, n74554 );
nand U109047 ( n25127, n25128, n25129 );
nand U109048 ( n25129, n76762, n74559 );
nand U109049 ( n58265, n58266, n58267 );
nand U109050 ( n58267, n76695, n74560 );
not U109051 ( n7813, n43331 );
nor U109052 ( n54380, n54337, n73549 );
nand U109053 ( n11899, n12673, n12674 );
nand U109054 ( n12673, n12680, n74649 );
nand U109055 ( n12674, n4819, n12675 );
nand U109056 ( n12675, n12677, n12678 );
nor U109057 ( n21399, n21358, n73980 );
nand U109058 ( n11864, n11842, n11898 );
nand U109059 ( n11898, n4787, n11845 );
nand U109060 ( n21393, n21394, n21395 );
nor U109061 ( n21395, n21396, n21397 );
nor U109062 ( n21394, n21398, n21399 );
nor U109063 ( n21396, n21355, n73991 );
not U109064 ( n4789, n11810 );
not U109065 ( n5754, n68003 );
not U109066 ( n7540, n46968 );
not U109067 ( n3997, n26000 );
not U109068 ( n6629, n59138 );
nor U109069 ( n28885, n28660, n73742 );
nor U109070 ( n62190, n61965, n73741 );
nand U109071 ( n8528, n8529, n8530 );
nand U109072 ( n8530, n8532, n76742 );
nand U109073 ( n8529, n8515, n8533 );
nor U109074 ( n8532, n5270, n8515 );
nand U109075 ( n9886, n8524, n8525 );
nor U109076 ( n8524, n8540, n8542 );
nor U109077 ( n8525, n8527, n8528 );
nor U109078 ( n8540, n75207, n8414 );
nor U109079 ( n54507, n43268, n73640 );
nor U109080 ( n70790, n70565, n73740 );
nand U109081 ( n54497, n54505, n54506 );
nor U109082 ( n54505, n54509, n54510 );
nor U109083 ( n54506, n54507, n54508 );
nor U109084 ( n54510, n54350, n73664 );
nand U109085 ( n9806, n9039, n9040 );
nor U109086 ( n9040, n9042, n9043 );
nor U109087 ( n9039, n9050, n9052 );
nand U109088 ( n9042, n9049, n8789 );
nand U109089 ( n9776, n9234, n9235 );
nor U109090 ( n9235, n9237, n9238 );
nor U109091 ( n9234, n9245, n9247 );
nand U109092 ( n9237, n9244, n8789 );
nor U109093 ( n36064, n35839, n74044 );
nor U109094 ( n54568, n54347, n73580 );
nand U109095 ( n54557, n54565, n54566 );
nor U109096 ( n54565, n54569, n54570 );
nor U109097 ( n54566, n54567, n54568 );
nor U109098 ( n54569, n54351, n73586 );
nand U109099 ( n26901, n28638, n28639 );
nand U109100 ( n28639, n4227, n28640 );
nand U109101 ( n28640, n28641, n28642 );
not U109102 ( n4227, n28645 );
nand U109103 ( n60041, n61943, n61944 );
nand U109104 ( n61944, n6859, n61945 );
nand U109105 ( n61945, n61946, n61947 );
not U109106 ( n6859, n61950 );
nand U109107 ( n16501, n43269, n43270 );
nor U109108 ( n43269, n43283, n43284 );
nor U109109 ( n43270, n43271, n43272 );
nand U109110 ( n43284, n43285, n43286 );
nand U109111 ( n68900, n70543, n70544 );
nand U109112 ( n70544, n6004, n70545 );
nand U109113 ( n70545, n70546, n70547 );
not U109114 ( n6004, n70550 );
nand U109115 ( n34146, n35817, n35818 );
nand U109116 ( n35818, n3389, n35819 );
nand U109117 ( n35819, n35820, n35821 );
not U109118 ( n3389, n35824 );
nand U109119 ( n11967, n11942, n11990 );
nand U109120 ( n11990, n4787, n11945 );
nand U109121 ( n12257, n12235, n12273 );
nand U109122 ( n12273, n4787, n12238 );
and U109123 ( n12235, n11899, n12274 );
nand U109124 ( n12274, n76732, n12228 );
or U109125 ( n12254, n12257, n75833 );
and U109126 ( n75833, n11772, n75200 );
nor U109127 ( n28860, n22674, n73841 );
nand U109128 ( n12064, n12028, n12099 );
nand U109129 ( n12099, n4787, n12032 );
or U109130 ( n12062, n12064, n75834 );
and U109131 ( n75834, n11772, n75201 );
nor U109132 ( n62165, n55787, n73842 );
nor U109133 ( n70765, n63953, n73840 );
or U109134 ( n12335, n12338, n75835 );
and U109135 ( n75835, n11772, n74644 );
nor U109136 ( n36039, n29997, n74224 );
nor U109137 ( n54501, n54338, n73651 );
nand U109138 ( n54498, n54499, n54500 );
nor U109139 ( n54499, n54503, n54504 );
nor U109140 ( n54500, n54501, n54502 );
nor U109141 ( n54503, n54342, n73646 );
nand U109142 ( n21379, n10265, n73525 );
nor U109143 ( n54516, n54358, n73639 );
nor U109144 ( n21413, n21379, n73964 );
nand U109145 ( n54512, n54513, n54514 );
nor U109146 ( n54513, n54517, n54518 );
nor U109147 ( n54514, n54515, n54516 );
nor U109148 ( n54517, n54363, n73644 );
nand U109149 ( n21407, n21408, n21409 );
nor U109150 ( n21409, n21410, n21411 );
nor U109151 ( n21408, n21412, n21413 );
nor U109152 ( n21411, n21375, n73981 );
nor U109153 ( n54478, n54347, n74145 );
nand U109154 ( n32389, n32390, n32391 );
nand U109155 ( n32390, n3544, n32146 );
or U109156 ( n32391, n74557, n32365 );
nand U109157 ( n32457, n32458, n32459 );
nand U109158 ( n32458, n29871, n32146 );
or U109159 ( n32459, n73102, n32436 );
nor U109160 ( n54579, n54583, n54584 );
nor U109161 ( n54583, n54372, n73578 );
nor U109162 ( n54584, n54371, n73573 );
nand U109163 ( n42643, n42644, n42645 );
nand U109164 ( n42645, n42646, n76675 );
nand U109165 ( n42644, n42628, n42647 );
nor U109166 ( n42646, n7927, n42628 );
nand U109167 ( n42774, n42775, n42776 );
nand U109168 ( n42776, n42777, n76675 );
nand U109169 ( n42775, n42764, n42778 );
nor U109170 ( n42777, n7929, n42764 );
nand U109171 ( n42592, n42593, n42594 );
nand U109172 ( n42594, n42595, n76675 );
nand U109173 ( n42593, n42582, n42596 );
nor U109174 ( n42595, n7925, n42582 );
nand U109175 ( n67052, n67053, n67054 );
nand U109176 ( n67053, n6159, n66792 );
or U109177 ( n67054, n74558, n67028 );
nand U109178 ( n67113, n67114, n67115 );
nand U109179 ( n67114, n63827, n66792 );
or U109180 ( n67115, n73100, n67092 );
nand U109181 ( n46088, n46089, n46090 );
nand U109182 ( n46089, n7947, n45841 );
or U109183 ( n46090, n74554, n46064 );
nand U109184 ( n46149, n46150, n46151 );
nand U109185 ( n46150, n43128, n45841 );
or U109186 ( n46151, n73098, n46128 );
nand U109187 ( n25215, n25216, n25217 );
nand U109188 ( n25216, n22548, n24914 );
or U109189 ( n25217, n73103, n25194 );
nand U109190 ( n25152, n25153, n25154 );
nand U109191 ( n25153, n4382, n24914 );
or U109192 ( n25154, n74559, n25128 );
nand U109193 ( n58351, n58352, n58353 );
nand U109194 ( n58352, n55661, n58051 );
or U109195 ( n58353, n73101, n58330 );
nand U109196 ( n58290, n58291, n58292 );
nand U109197 ( n58291, n7014, n58051 );
or U109198 ( n58292, n74560, n58266 );
nand U109199 ( n16591, n42771, n42772 );
nor U109200 ( n42771, n42784, n42785 );
nor U109201 ( n42772, n42773, n42774 );
nor U109202 ( n42784, n75202, n42500 );
nand U109203 ( n16621, n42589, n42590 );
nor U109204 ( n42589, n42602, n42603 );
nor U109205 ( n42590, n42591, n42592 );
nor U109206 ( n42602, n75208, n42500 );
nand U109207 ( n16611, n42640, n42641 );
nor U109208 ( n42640, n42655, n42656 );
nor U109209 ( n42641, n42642, n42643 );
nor U109210 ( n42655, n75236, n42500 );
nor U109211 ( n54474, n54341, n74133 );
nand U109212 ( n16541, n43043, n43044 );
nor U109213 ( n43044, n43045, n43046 );
nor U109214 ( n43043, n43052, n43053 );
nand U109215 ( n43045, n43051, n42829 );
nand U109216 ( n16511, n43199, n43200 );
nor U109217 ( n43200, n43201, n43202 );
nor U109218 ( n43199, n43208, n43209 );
nand U109219 ( n43201, n43207, n42829 );
nand U109220 ( n9901, n8419, n8420 );
nor U109221 ( n8419, n8440, n8442 );
nor U109222 ( n8420, n8422, n8423 );
nor U109223 ( n8440, n74924, n8414 );
nand U109224 ( n16636, n42504, n42505 );
nor U109225 ( n42504, n42519, n42520 );
nor U109226 ( n42505, n42506, n42507 );
nor U109227 ( n42519, n74931, n42500 );
nor U109228 ( n21494, n9303, n74361 );
nor U109229 ( n21403, n21364, n73983 );
nand U109230 ( n21484, n21492, n21493 );
nor U109231 ( n21492, n21496, n21497 );
nor U109232 ( n21493, n21494, n21495 );
nor U109233 ( n21497, n21367, n74377 );
nand U109234 ( n21392, n21400, n21401 );
nor U109235 ( n21400, n21404, n21405 );
nor U109236 ( n21401, n21402, n21403 );
nor U109237 ( n21404, n21368, n73988 );
not U109238 ( n12, n11605 );
nand U109239 ( n12600, n76732, n74718 );
nand U109240 ( n8981, n12539, n12540 );
nor U109241 ( n12539, n12558, n12559 );
nor U109242 ( n12540, n12542, n12543 );
nor U109243 ( n12558, n74727, n76734 );
nand U109244 ( n12554, n12555, n12557 );
nand U109245 ( n12557, n76733, n74484 );
nand U109246 ( n9373, n8438, n9374 );
nand U109247 ( n9374, n76745, n75226 );
nor U109248 ( n54562, n54337, n73593 );
nand U109249 ( n7266, n23808, n23809 );
nor U109250 ( n23808, n23820, n23821 );
nor U109251 ( n23809, n23810, n23811 );
nand U109252 ( n23821, n23822, n23823 );
nand U109253 ( n14001, n56933, n56934 );
nor U109254 ( n56933, n56945, n56946 );
nor U109255 ( n56934, n56935, n56936 );
nand U109256 ( n56946, n56947, n56948 );
nor U109257 ( n23636, n74878, n76539 );
nor U109258 ( n23725, n74820, n76539 );
nor U109259 ( n23547, n74923, n76539 );
nor U109260 ( n56758, n74877, n76281 );
nor U109261 ( n56669, n74922, n76281 );
nor U109262 ( n56847, n74819, n76281 );
nor U109263 ( n23814, n74780, n76539 );
nor U109264 ( n56939, n74779, n76281 );
nand U109265 ( n7286, n23630, n23631 );
nor U109266 ( n23630, n23641, n23642 );
nor U109267 ( n23631, n23632, n23633 );
nor U109268 ( n23641, n24, n23152 );
nand U109269 ( n7276, n23719, n23720 );
nor U109270 ( n23719, n23730, n23731 );
nor U109271 ( n23720, n23721, n23722 );
nor U109272 ( n23730, n14, n23152 );
nand U109273 ( n7296, n23541, n23542 );
nor U109274 ( n23541, n23552, n23553 );
nor U109275 ( n23542, n23543, n23544 );
nor U109276 ( n23552, n34, n23152 );
nand U109277 ( n14021, n56752, n56753 );
nor U109278 ( n56752, n56763, n56764 );
nor U109279 ( n56753, n56754, n56755 );
nor U109280 ( n56763, n274, n56273 );
nand U109281 ( n14031, n56663, n56664 );
nor U109282 ( n56663, n56674, n56675 );
nor U109283 ( n56664, n56665, n56666 );
nor U109284 ( n56674, n287, n56273 );
nand U109285 ( n14011, n56841, n56842 );
nor U109286 ( n56841, n56852, n56853 );
nor U109287 ( n56842, n56843, n56844 );
nor U109288 ( n56852, n262, n56273 );
nor U109289 ( n23303, n75037, n76539 );
nor U109290 ( n56427, n75036, n76281 );
nor U109291 ( n31111, n74778, n76482 );
nand U109292 ( n7316, n23297, n23298 );
nor U109293 ( n23297, n23308, n23309 );
nor U109294 ( n23298, n23299, n23300 );
nor U109295 ( n23308, n23344, n23152 );
nor U109296 ( n54489, n54493, n54494 );
nor U109297 ( n54493, n54372, n74151 );
nor U109298 ( n54494, n54371, n74138 );
nand U109299 ( n7306, n23394, n23395 );
nor U109300 ( n23394, n23437, n23438 );
nor U109301 ( n23395, n23396, n23397 );
nor U109302 ( n23437, n23441, n23152 );
nand U109303 ( n5021, n31105, n31106 );
nor U109304 ( n31105, n31117, n31118 );
nor U109305 ( n31106, n31107, n31108 );
nor U109306 ( n31117, n75411, n30480 );
nand U109307 ( n11756, n65359, n65360 );
nor U109308 ( n65359, n65371, n65372 );
nor U109309 ( n65360, n65361, n65362 );
nor U109310 ( n65371, n75412, n64639 );
nor U109311 ( n21581, n21358, n74082 );
nand U109312 ( n21575, n21576, n21577 );
nor U109313 ( n21577, n21578, n21579 );
nor U109314 ( n21576, n21580, n21581 );
nor U109315 ( n21578, n21355, n74100 );
nor U109316 ( n30941, n74876, n76482 );
nor U109317 ( n56522, n74971, n76281 );
nor U109318 ( n23400, n74972, n76539 );
nor U109319 ( n65365, n74776, n76215 );
nand U109320 ( n14051, n56421, n56422 );
nor U109321 ( n56421, n56432, n56433 );
nor U109322 ( n56422, n56423, n56424 );
nor U109323 ( n56432, n56468, n56273 );
nor U109324 ( n65058, n74921, n76215 );
nor U109325 ( n65143, n74875, n76215 );
nor U109326 ( n65228, n74814, n76215 );
nor U109327 ( n31026, n74817, n76482 );
nand U109328 ( n14041, n56516, n56517 );
nor U109329 ( n56516, n56559, n56560 );
nor U109330 ( n56517, n56518, n56519 );
nor U109331 ( n56559, n56563, n56273 );
nand U109332 ( n5041, n30935, n30936 );
nor U109333 ( n30935, n30976, n30977 );
nor U109334 ( n30936, n30937, n30938 );
nor U109335 ( n30976, n75313, n30481 );
nand U109336 ( n11786, n65052, n65053 );
nor U109337 ( n65052, n65093, n65094 );
nor U109338 ( n65053, n65054, n65055 );
nor U109339 ( n65093, n75290, n64640 );
nand U109340 ( n11776, n65137, n65138 );
nor U109341 ( n65137, n65178, n65179 );
nor U109342 ( n65138, n65139, n65140 );
nor U109343 ( n65178, n75293, n64640 );
nand U109344 ( n11766, n65222, n65223 );
nor U109345 ( n65222, n65263, n65264 );
nor U109346 ( n65223, n65224, n65225 );
nor U109347 ( n65263, n75292, n64640 );
nand U109348 ( n5031, n31020, n31021 );
nor U109349 ( n31020, n31061, n31062 );
nor U109350 ( n31021, n31022, n31023 );
nor U109351 ( n31061, n75296, n30481 );
nor U109352 ( n30856, n74927, n76482 );
nand U109353 ( n5051, n30850, n30851 );
nor U109354 ( n30850, n30891, n30892 );
nor U109355 ( n30851, n30852, n30853 );
nor U109356 ( n30891, n75314, n30481 );
nor U109357 ( n64827, n75028, n76215 );
nor U109358 ( n64916, n74968, n76215 );
nand U109359 ( n11806, n64821, n64822 );
nor U109360 ( n64821, n64864, n64865 );
nor U109361 ( n64822, n64823, n64824 );
nor U109362 ( n64864, n75310, n64640 );
nand U109363 ( n11796, n64910, n64911 );
nor U109364 ( n64910, n64953, n64954 );
nor U109365 ( n64911, n64912, n64913 );
nor U109366 ( n64953, n75309, n64640 );
nor U109367 ( n54488, n54362, n74106 );
nand U109368 ( n5071, n30615, n30616 );
nor U109369 ( n30615, n30658, n30659 );
nor U109370 ( n30616, n30617, n30618 );
nor U109371 ( n30658, n75321, n30481 );
nand U109372 ( n5061, n30704, n30705 );
nor U109373 ( n30704, n30747, n30748 );
nor U109374 ( n30705, n30706, n30707 );
nor U109375 ( n30747, n75320, n30481 );
nor U109376 ( n30621, n75041, n76482 );
nor U109377 ( n30710, n74984, n76482 );
nor U109378 ( n21488, n21355, n74375 );
nor U109379 ( n49530, n50031, n76834 );
nand U109380 ( n21485, n21486, n21487 );
nor U109381 ( n21486, n21490, n21491 );
nor U109382 ( n21487, n21488, n21489 );
nor U109383 ( n21490, n21359, n74370 );
nand U109384 ( n54359, n44133, n73497 );
nor U109385 ( n54393, n54359, n73545 );
nand U109386 ( n21375, n10260, n73525 );
nor U109387 ( n21503, n21375, n74359 );
nand U109388 ( n21499, n21500, n21501 );
nor U109389 ( n21500, n21504, n21505 );
nor U109390 ( n21501, n21502, n21503 );
nor U109391 ( n21504, n21380, n74364 );
nor U109392 ( n21414, n21418, n21419 );
nor U109393 ( n21418, n21389, n73982 );
nor U109394 ( n21419, n21388, n73978 );
nor U109395 ( n28898, n28682, n73730 );
nor U109396 ( n62203, n61987, n73729 );
nor U109397 ( n70803, n70587, n73728 );
nor U109398 ( n36077, n35861, n74034 );
nor U109399 ( n21595, n21379, n74046 );
nand U109400 ( n21589, n21590, n21591 );
nor U109401 ( n21591, n21592, n21593 );
nor U109402 ( n21590, n21594, n21595 );
nor U109403 ( n21593, n21375, n74084 );
nand U109404 ( n43324, n42512, n43325 );
nand U109405 ( n43325, n76678, n75225 );
nand U109406 ( n54350, n7813, n44161 );
nor U109407 ( n54388, n54350, n73550 );
not U109408 ( n5158, n9382 );
nor U109409 ( n21397, n21354, n73992 );
nor U109410 ( n54508, n54347, n73647 );
nor U109411 ( n54447, n43268, n73882 );
nand U109412 ( n54437, n54445, n54446 );
nor U109413 ( n54445, n54449, n54450 );
nor U109414 ( n54446, n54447, n54448 );
nor U109415 ( n54450, n54350, n73894 );
nor U109416 ( n54504, n54341, n73638 );
nand U109417 ( n8996, n12464, n12465 );
nor U109418 ( n12464, n12483, n12484 );
nor U109419 ( n12465, n12467, n12468 );
nor U109420 ( n12483, n75967, n76734 );
nand U109421 ( n12479, n12480, n12482 );
nand U109422 ( n12482, n76733, n73097 );
nor U109423 ( n40326, n2083, n2069 );
nor U109424 ( n28893, n28673, n73745 );
nor U109425 ( n62198, n61978, n73744 );
nand U109426 ( n12568, n12575, n12577 );
nand U109427 ( n12577, n12553, n74484 );
or U109428 ( n12575, n74484, n12555 );
nand U109429 ( n8976, n12565, n12567 );
nor U109430 ( n12565, n12580, n12582 );
nor U109431 ( n12567, n12568, n12569 );
nor U109432 ( n12580, n74673, n76734 );
nor U109433 ( n54490, n54491, n54492 );
nor U109434 ( n54492, n48005, n74146 );
nor U109435 ( n54491, n54368, n74159 );
nand U109436 ( n9011, n12378, n12379 );
nor U109437 ( n12378, n12397, n12398 );
nor U109438 ( n12379, n12380, n12382 );
nor U109439 ( n12397, n74812, n76734 );
nand U109440 ( n12393, n12394, n12395 );
nand U109441 ( n12395, n76733, n74577 );
nor U109442 ( n70798, n70578, n73743 );
not U109443 ( n8212, n17129 );
nor U109444 ( n21524, n9303, n74143 );
nor U109445 ( n36072, n35852, n74047 );
nand U109446 ( n21514, n21522, n21523 );
nor U109447 ( n21522, n21526, n21527 );
nor U109448 ( n21523, n21524, n21525 );
nor U109449 ( n21527, n21367, n74164 );
nor U109450 ( n28890, n22674, n73748 );
nor U109451 ( n62195, n55787, n73747 );
nor U109452 ( n21585, n21364, n74088 );
nand U109453 ( n21574, n21582, n21583 );
nor U109454 ( n21582, n21586, n21587 );
nor U109455 ( n21583, n21584, n21585 );
nor U109456 ( n21586, n21368, n74098 );
nor U109457 ( n54417, n43268, n73968 );
nor U109458 ( n70795, n63953, n73746 );
nand U109459 ( n54407, n54415, n54416 );
nor U109460 ( n54415, n54419, n54420 );
nor U109461 ( n54416, n54417, n54418 );
nor U109462 ( n54420, n54350, n73996 );
nor U109463 ( n36069, n29997, n74048 );
nor U109464 ( n54519, n54523, n54524 );
nor U109465 ( n54523, n54372, n73656 );
nor U109466 ( n54524, n54371, n73645 );
nand U109467 ( n9264, n9279, n9280 );
nor U109468 ( n9279, n4765, n9290 );
nand U109469 ( n9280, n9282, n76744 );
not U109470 ( n4765, n8789 );
nand U109471 ( n9771, n9262, n9263 );
nor U109472 ( n9262, n9294, n9295 );
nor U109473 ( n9263, n9264, n9265 );
nand U109474 ( n9294, n9299, n9300 );
nor U109475 ( n54441, n54338, n73890 );
nor U109476 ( n54518, n54362, n73636 );
nand U109477 ( n54438, n54439, n54440 );
nor U109478 ( n54439, n54443, n54444 );
nor U109479 ( n54440, n54441, n54442 );
nor U109480 ( n54443, n54342, n73885 );
nand U109481 ( n9836, n8845, n8847 );
nor U109482 ( n8845, n8859, n8860 );
nor U109483 ( n8847, n8848, n8849 );
nand U109484 ( n8860, n8862, n8863 );
nand U109485 ( n36287, n37079, n37078 );
nor U109486 ( n37079, n37080, n36943 );
nor U109487 ( n54398, n54399, n54400 );
nor U109488 ( n54400, n48005, n73542 );
nor U109489 ( n54399, n54368, n73547 );
nand U109490 ( n9072, n9073, n9074 );
nand U109491 ( n9073, n9084, n76890 );
nand U109492 ( n9074, n9075, n76743 );
nor U109493 ( n9084, n5460, n9085 );
nand U109494 ( n9137, n9138, n9139 );
nand U109495 ( n9138, n9149, n76890 );
nand U109496 ( n9139, n9140, n76743 );
nor U109497 ( n9149, n5462, n9150 );
nand U109498 ( n8875, n8877, n8878 );
nand U109499 ( n8877, n8888, n76889 );
nand U109500 ( n8878, n8879, n76743 );
nor U109501 ( n8888, n5457, n8889 );
nand U109502 ( n9801, n9068, n9069 );
nor U109503 ( n9068, n9094, n9095 );
nor U109504 ( n9069, n9070, n9072 );
nand U109505 ( n9094, n9099, n9100 );
nand U109506 ( n9791, n9133, n9134 );
nor U109507 ( n9133, n9157, n9158 );
nor U109508 ( n9134, n9135, n9137 );
nand U109509 ( n9157, n9162, n9163 );
nand U109510 ( n9831, n8872, n8873 );
nor U109511 ( n8872, n8899, n8900 );
nor U109512 ( n8873, n8874, n8875 );
nand U109513 ( n8899, n8904, n8905 );
nor U109514 ( n21518, n21355, n74157 );
nor U109515 ( n54456, n54358, n73881 );
nand U109516 ( n21515, n21516, n21517 );
nor U109517 ( n21516, n21520, n21521 );
nor U109518 ( n21517, n21518, n21519 );
nor U109519 ( n21520, n21359, n74152 );
nand U109520 ( n54452, n54453, n54454 );
nor U109521 ( n54453, n54457, n54458 );
nor U109522 ( n54454, n54455, n54456 );
nor U109523 ( n54457, n54363, n73883 );
nor U109524 ( n28903, n28904, n28905 );
nor U109525 ( n28905, n27016, n73724 );
nor U109526 ( n28904, n28691, n73736 );
nor U109527 ( n62208, n62209, n62210 );
nor U109528 ( n62210, n60157, n73723 );
nor U109529 ( n62209, n61996, n73735 );
nor U109530 ( n21533, n21375, n74140 );
nand U109531 ( n21529, n21530, n21531 );
nor U109532 ( n21530, n21534, n21535 );
nor U109533 ( n21531, n21532, n21533 );
nor U109534 ( n21534, n21380, n74149 );
nand U109535 ( n8395, n8397, n8398 );
nand U109536 ( n8397, n8403, n8404 );
nand U109537 ( n8398, n8399, n76743 );
nor U109538 ( n8403, n73392, n75238 );
nand U109539 ( n9906, n8392, n8393 );
nor U109540 ( n8392, n8412, n8413 );
nor U109541 ( n8393, n8394, n8395 );
nor U109542 ( n8413, n74964, n8414 );
nor U109543 ( n54411, n54338, n73977 );
nand U109544 ( n54408, n54409, n54410 );
nor U109545 ( n54409, n54413, n54414 );
nor U109546 ( n54410, n54411, n54412 );
nor U109547 ( n54413, n54342, n73972 );
nand U109548 ( n9781, n9199, n9200 );
nor U109549 ( n9199, n9224, n9225 );
nor U109550 ( n9200, n9202, n9203 );
nand U109551 ( n9224, n9229, n9230 );
nor U109552 ( n70808, n70809, n70810 );
nor U109553 ( n70810, n69013, n73722 );
nor U109554 ( n70809, n70596, n73734 );
nand U109555 ( n54363, n44137, n73497 );
nor U109556 ( n54395, n54363, n73537 );
nor U109557 ( n54575, n54359, n73584 );
nor U109558 ( n36082, n36083, n36084 );
nor U109559 ( n36084, n34259, n74032 );
nor U109560 ( n36083, n35870, n74040 );
nor U109561 ( n21596, n21600, n21601 );
nor U109562 ( n21600, n21389, n74085 );
nor U109563 ( n21601, n21388, n74071 );
nand U109564 ( n9871, n8618, n8619 );
nor U109565 ( n8618, n8647, n8648 );
nor U109566 ( n8619, n8620, n8622 );
nor U109567 ( n8647, n74737, n8414 );
nand U109568 ( n8745, n8755, n8757 );
nand U109569 ( n8755, n8767, n76889 );
nand U109570 ( n8757, n8758, n76742 );
nor U109571 ( n8767, n5454, n8768 );
nand U109572 ( n8553, n8565, n8567 );
nand U109573 ( n8565, n8577, n76889 );
nand U109574 ( n8567, n8568, n76742 );
nor U109575 ( n8577, n5450, n8578 );
nand U109576 ( n8620, n8629, n8630 );
nand U109577 ( n8629, n8640, n76889 );
nand U109578 ( n8630, n8632, n76742 );
nor U109579 ( n8640, n5452, n8642 );
nand U109580 ( n9851, n8743, n8744 );
nor U109581 ( n8743, n8773, n8774 );
nor U109582 ( n8744, n8745, n8747 );
nor U109583 ( n8773, n74956, n8414 );
nand U109584 ( n9881, n8550, n8552 );
nor U109585 ( n8550, n8583, n8584 );
nor U109586 ( n8552, n8553, n8554 );
nor U109587 ( n8583, n74808, n8414 );
nor U109588 ( n72844, n73096, n71108 );
nor U109589 ( n28900, n28686, n73709 );
nor U109590 ( n62205, n61991, n73708 );
nand U109591 ( n9761, n9334, n9335 );
nor U109592 ( n9334, n9355, n9357 );
nor U109593 ( n9335, n9337, n9338 );
nand U109594 ( n9355, n9360, n9362 );
nor U109595 ( n70805, n70591, n73707 );
nor U109596 ( n36079, n35865, n74022 );
nor U109597 ( n54426, n54358, n73967 );
nand U109598 ( n54422, n54423, n54424 );
nor U109599 ( n54423, n54427, n54428 );
nor U109600 ( n54424, n54425, n54426 );
nor U109601 ( n54427, n54363, n73970 );
nand U109602 ( n9821, n8938, n8939 );
nor U109603 ( n8938, n8962, n8963 );
nor U109604 ( n8939, n8940, n8942 );
nand U109605 ( n8962, n8967, n8968 );
nand U109606 ( n9811, n9004, n9005 );
nor U109607 ( n9004, n9029, n9030 );
nor U109608 ( n9005, n9007, n9008 );
nand U109609 ( n9029, n9034, n9035 );
nand U109610 ( n9841, n8810, n8812 );
nor U109611 ( n8810, n8835, n8837 );
nor U109612 ( n8812, n8813, n8814 );
nand U109613 ( n8835, n8840, n8842 );
nand U109614 ( n12430, n12432, n12433 );
nand U109615 ( n12432, n5292, n12118 );
or U109616 ( n12433, n74577, n12394 );
nand U109617 ( n12507, n12508, n12509 );
nand U109618 ( n12508, n9145, n12118 );
or U109619 ( n12509, n73097, n12480 );
nor U109620 ( n54479, n54351, n74158 );
nand U109621 ( n9891, n8487, n8488 );
nor U109622 ( n8487, n8519, n8520 );
nor U109623 ( n8488, n8489, n8490 );
nor U109624 ( n8519, n74880, n8414 );
nand U109625 ( n9861, n8679, n8680 );
nor U109626 ( n8679, n8712, n8713 );
nor U109627 ( n8680, n8682, n8683 );
nor U109628 ( n8712, n74677, n8414 );
nor U109629 ( n54570, n54350, n73599 );
nor U109630 ( n21579, n21354, n74101 );
nor U109631 ( n54520, n54521, n54522 );
nor U109632 ( n54522, n48005, n73649 );
nor U109633 ( n54521, n54368, n73663 );
nor U109634 ( n54534, n54341, n73806 );
nand U109635 ( n54528, n54529, n54530 );
nor U109636 ( n54530, n54531, n54532 );
nor U109637 ( n54529, n54533, n54534 );
nor U109638 ( n54531, n54338, n73816 );
xnor U109639 ( n12385, n13525, n13715 );
xor U109640 ( n13715, n73116, n76034 );
nor U109641 ( n13704, n13707, n76594 );
nor U109642 ( n13707, n13708, n13709 );
nand U109643 ( n13709, n13710, n13712 );
nand U109644 ( n13708, n13713, n13714 );
nand U109645 ( n31842, n31856, n31857 );
nor U109646 ( n31856, n3063, n31859 );
nand U109647 ( n31857, n76779, n31858 );
nor U109648 ( n31859, n31860, n31861 );
nand U109649 ( n43069, n43070, n43071 );
nand U109650 ( n43070, n43079, n76862 );
nand U109651 ( n43071, n43072, n76677 );
nor U109652 ( n43079, n8114, n43080 );
nand U109653 ( n16536, n43066, n43067 );
nor U109654 ( n43066, n43087, n43088 );
nor U109655 ( n43067, n43068, n43069 );
nand U109656 ( n43087, n43091, n43092 );
nand U109657 ( n24628, n24642, n24643 );
nor U109658 ( n24642, n3907, n24645 );
nand U109659 ( n24643, n76761, n24644 );
nor U109660 ( n24645, n24646, n24647 );
nand U109661 ( n57760, n57778, n57779 );
nor U109662 ( n57778, n6539, n57781 );
nand U109663 ( n57779, n76694, n57780 );
nor U109664 ( n57781, n57782, n57783 );
nand U109665 ( n66465, n66479, n66480 );
nor U109666 ( n66479, n5664, n66482 );
nand U109667 ( n66480, n76713, n66481 );
nor U109668 ( n66482, n66483, n66484 );
nand U109669 ( n21376, n10262, n73525 );
nor U109670 ( n21410, n21376, n73986 );
nor U109671 ( n21495, n21364, n74368 );
nor U109672 ( n16685, n17053, n76788 );
nand U109673 ( n43237, n43249, n43250 );
nor U109674 ( n43249, n7410, n43258 );
nand U109675 ( n43250, n43251, n76677 );
not U109676 ( n7410, n42829 );
nor U109677 ( n54580, n54581, n54582 );
nor U109678 ( n54582, n48005, n73581 );
nor U109679 ( n54581, n54368, n73587 );
nand U109680 ( n16506, n43235, n43236 );
nor U109681 ( n43235, n43261, n43262 );
nor U109682 ( n43236, n43237, n43238 );
nand U109683 ( n43261, n43265, n43266 );
nor U109684 ( n21491, n21358, n74362 );
nand U109685 ( n16571, n42874, n42875 );
nor U109686 ( n42874, n42885, n42886 );
nor U109687 ( n42875, n42876, n42877 );
nand U109688 ( n42886, n42887, n42888 );
nor U109689 ( n54448, n54347, n73886 );
nand U109690 ( n32178, n74610, n33115 );
or U109691 ( n33115, n32215, n74635 );
nor U109692 ( n54472, n54337, n74147 );
nor U109693 ( n54444, n54341, n73880 );
nand U109694 ( n12158, n74586, n13358 );
or U109695 ( n13358, n12204, n74599 );
nand U109696 ( n45873, n74550, n46824 );
or U109697 ( n46824, n45921, n74524 );
nand U109698 ( n45541, n45554, n45555 );
nor U109699 ( n45554, n7438, n45557 );
nand U109700 ( n45555, n76665, n45556 );
nor U109701 ( n45557, n45558, n45559 );
nand U109702 ( n43121, n43122, n43123 );
nand U109703 ( n43122, n43131, n76863 );
nand U109704 ( n43123, n43124, n76676 );
nor U109705 ( n43131, n8115, n43132 );
nand U109706 ( n42898, n42899, n42900 );
nand U109707 ( n42899, n42908, n76862 );
nand U109708 ( n42900, n42901, n76676 );
nor U109709 ( n42908, n8110, n42909 );
nand U109710 ( n16526, n43118, n43119 );
nor U109711 ( n43118, n43137, n43138 );
nor U109712 ( n43119, n43120, n43121 );
nand U109713 ( n43137, n43141, n43142 );
nand U109714 ( n16566, n42895, n42896 );
nor U109715 ( n42895, n42917, n42918 );
nor U109716 ( n42896, n42897, n42898 );
nand U109717 ( n42917, n42921, n42922 );
and U109718 ( n32000, n31979, n76778 );
nor U109719 ( n54577, n54363, n73575 );
nand U109720 ( n21367, n5158, n10297 );
nor U109721 ( n17665, n17440, n76788 );
nor U109722 ( n21405, n21367, n73995 );
nand U109723 ( n42485, n42486, n42487 );
nand U109724 ( n42486, n42491, n42492 );
nand U109725 ( n42487, n42488, n76676 );
nor U109726 ( n42491, n73391, n75237 );
nand U109727 ( n16641, n42482, n42483 );
nor U109728 ( n42482, n42498, n42499 );
nor U109729 ( n42483, n42484, n42485 );
nor U109730 ( n42499, n74967, n42500 );
nor U109731 ( n54548, n54362, n73805 );
nand U109732 ( n54542, n54543, n54544 );
nor U109733 ( n54544, n54545, n54546 );
nor U109734 ( n54543, n54547, n54548 );
nor U109735 ( n54546, n54358, n73807 );
and U109736 ( n66603, n66582, n76712 );
and U109737 ( n24768, n24747, n76760 );
and U109738 ( n57902, n57881, n76693 );
and U109739 ( n45774, n45735, n76664 );
nand U109740 ( n66824, n74574, n67871 );
or U109741 ( n67871, n66872, n74546 );
nand U109742 ( n24948, n74575, n25868 );
or U109743 ( n25868, n24996, n74547 );
nand U109744 ( n58083, n74576, n59006 );
or U109745 ( n59006, n58131, n74548 );
not U109746 ( n7815, n43330 );
nor U109747 ( n21464, n9303, n74297 );
nor U109748 ( n54418, n54347, n73973 );
nor U109749 ( n54381, n54342, n73543 );
nand U109750 ( n21454, n21462, n21463 );
nor U109751 ( n21462, n21466, n21467 );
nor U109752 ( n21463, n21464, n21465 );
nor U109753 ( n21467, n21367, n74296 );
nor U109754 ( n17068, n17129, n73020 );
nand U109755 ( n42612, n42622, n42623 );
nand U109756 ( n42622, n42631, n76862 );
nand U109757 ( n42623, n42624, n76675 );
nor U109758 ( n42631, n8104, n42632 );
nand U109759 ( n16606, n42688, n42689 );
nor U109760 ( n42688, n42711, n42712 );
nor U109761 ( n42689, n42690, n42691 );
nor U109762 ( n42711, n74740, n42500 );
nand U109763 ( n42794, n42802, n42803 );
nand U109764 ( n42802, n42811, n76862 );
nand U109765 ( n42803, n42804, n76675 );
nor U109766 ( n42811, n8108, n42812 );
nand U109767 ( n42690, n42697, n42698 );
nand U109768 ( n42697, n42706, n76862 );
nand U109769 ( n42698, n42699, n76675 );
nor U109770 ( n42706, n8105, n42707 );
nand U109771 ( n16586, n42792, n42793 );
nor U109772 ( n42792, n42816, n42817 );
nor U109773 ( n42793, n42794, n42795 );
nor U109774 ( n42816, n74957, n42500 );
nand U109775 ( n16616, n42610, n42611 );
nor U109776 ( n42610, n42636, n42637 );
nor U109777 ( n42611, n42612, n42613 );
nor U109778 ( n42636, n74810, n42500 );
and U109779 ( n31892, n31871, n76778 );
and U109780 ( n45679, n45658, n76664 );
and U109781 ( n32079, n32058, n76778 );
nor U109782 ( n54414, n54341, n73966 );
nand U109783 ( n16496, n43293, n43294 );
nor U109784 ( n43293, n43310, n43311 );
nor U109785 ( n43294, n43295, n43296 );
nand U109786 ( n43310, n43314, n43315 );
and U109787 ( n66515, n66494, n76712 );
and U109788 ( n24680, n24657, n76760 );
and U109789 ( n57814, n57793, n76693 );
nor U109790 ( n21507, n21508, n21509 );
nor U109791 ( n21509, n14797, n74369 );
nor U109792 ( n21508, n21385, n74374 );
and U109793 ( n66682, n66661, n76712 );
and U109794 ( n24847, n24826, n76760 );
and U109795 ( n57981, n57960, n76693 );
nor U109796 ( n21506, n21510, n21511 );
nor U109797 ( n21510, n21389, n74365 );
nor U109798 ( n21511, n21388, n74363 );
and U109799 ( n45590, n45569, n76664 );
nor U109800 ( n54538, n54347, n73812 );
nor U109801 ( n28886, n28665, n73727 );
nor U109802 ( n62191, n61970, n73726 );
nand U109803 ( n54527, n54535, n54536 );
nor U109804 ( n54535, n54539, n54540 );
nor U109805 ( n54536, n54537, n54538 );
nor U109806 ( n54539, n54351, n73818 );
nor U109807 ( n21434, n9303, n74333 );
nor U109808 ( n21505, n21379, n74357 );
nor U109809 ( n70791, n70570, n73725 );
nand U109810 ( n21424, n21432, n21433 );
nor U109811 ( n21432, n21436, n21437 );
nor U109812 ( n21433, n21434, n21435 );
nor U109813 ( n21437, n21367, n74334 );
nor U109814 ( n36065, n35844, n74033 );
nand U109815 ( n16556, n42962, n42963 );
nor U109816 ( n42962, n42981, n42982 );
nor U109817 ( n42963, n42964, n42965 );
nand U109818 ( n42981, n42985, n42986 );
nand U109819 ( n16546, n43015, n43016 );
nor U109820 ( n43015, n43035, n43036 );
nor U109821 ( n43016, n43017, n43018 );
nand U109822 ( n43035, n43039, n43040 );
nand U109823 ( n16576, n42846, n42847 );
nor U109824 ( n42846, n42866, n42867 );
nor U109825 ( n42847, n42848, n42849 );
nand U109826 ( n42866, n42870, n42871 );
nand U109827 ( n16516, n43171, n43172 );
nor U109828 ( n43171, n43191, n43192 );
nor U109829 ( n43172, n43173, n43174 );
nand U109830 ( n43191, n43195, n43196 );
nor U109831 ( n54459, n54463, n54464 );
nor U109832 ( n54463, n54372, n73891 );
nor U109833 ( n54464, n54371, n73884 );
nor U109834 ( n54509, n54351, n73662 );
nor U109835 ( n54458, n54362, n73867 );
nand U109836 ( n16631, n42529, n42530 );
nor U109837 ( n42529, n42555, n42556 );
nor U109838 ( n42530, n42531, n42532 );
nor U109839 ( n42555, n75077, n42500 );
nand U109840 ( n16626, n42559, n42560 );
nor U109841 ( n42559, n42585, n42586 );
nor U109842 ( n42560, n42561, n42562 );
nor U109843 ( n42585, n74891, n42500 );
nand U109844 ( n16596, n42741, n42742 );
nor U109845 ( n42741, n42767, n42768 );
nor U109846 ( n42742, n42743, n42744 );
nor U109847 ( n42767, n74680, n42500 );
nor U109848 ( n21458, n21355, n74294 );
nand U109849 ( n21455, n21456, n21457 );
nor U109850 ( n21456, n21460, n21461 );
nor U109851 ( n21457, n21458, n21459 );
nor U109852 ( n21460, n21359, n74290 );
nor U109853 ( n54429, n54433, n54434 );
nor U109854 ( n54433, n54372, n73990 );
nor U109855 ( n54434, n54371, n73971 );
nor U109856 ( n21415, n21416, n21417 );
nor U109857 ( n21417, n14797, n73984 );
nor U109858 ( n21416, n21385, n73989 );
nor U109859 ( n21473, n21375, n74286 );
not U109860 ( n2075, n38120 );
nand U109861 ( n21469, n21470, n21471 );
nor U109862 ( n21470, n21474, n21475 );
nor U109863 ( n21471, n21472, n21473 );
nor U109864 ( n21474, n21380, n74284 );
nor U109865 ( n54428, n54362, n73950 );
nor U109866 ( n21428, n21355, n74331 );
nand U109867 ( n21425, n21426, n21427 );
nor U109868 ( n21426, n21430, n21431 );
nor U109869 ( n21427, n21428, n21429 );
nor U109870 ( n21430, n21359, n74327 );
nor U109871 ( n21592, n21376, n74097 );
nor U109872 ( n37708, n73799, n73023 );
nand U109873 ( n33197, n76774, n32261 );
nor U109874 ( n21525, n21364, n74153 );
nor U109875 ( n54549, n54553, n54554 );
nor U109876 ( n54553, n54372, n73817 );
nor U109877 ( n54554, n54371, n73810 );
nor U109878 ( n21443, n21375, n74323 );
nand U109879 ( n21439, n21440, n21441 );
nor U109880 ( n21440, n21444, n21445 );
nor U109881 ( n21441, n21442, n21443 );
nor U109882 ( n21444, n21380, n74321 );
nand U109883 ( n13460, n76727, n12264 );
and U109884 ( n71661, n71144, n71096 );
nor U109885 ( n21521, n21358, n74139 );
nand U109886 ( n46906, n76660, n45949 );
nor U109887 ( n37704, n73798, n73023 );
nand U109888 ( n67953, n76708, n66900 );
nand U109889 ( n25950, n76754, n25024 );
nand U109890 ( n59088, n76687, n58159 );
nand U109891 ( n21380, n10267, n73525 );
nor U109892 ( n21412, n21380, n73979 );
nor U109893 ( n21587, n21367, n74103 );
nor U109894 ( n54532, n54337, n73815 );
nor U109895 ( n54460, n54461, n54462 );
nor U109896 ( n54462, n48005, n73888 );
nor U109897 ( n54461, n54368, n73893 );
nor U109898 ( n21537, n21538, n21539 );
nor U109899 ( n21539, n14797, n74155 );
nor U109900 ( n21538, n21385, n74163 );
nor U109901 ( n21536, n21540, n21541 );
nor U109902 ( n21540, n21389, n74161 );
nor U109903 ( n21541, n21388, n74150 );
nor U109904 ( n54485, n54359, n74141 );
nor U109905 ( n54563, n54342, n73582 );
nor U109906 ( n21551, n21358, n74240 );
nand U109907 ( n32032, n32054, n32055 );
or U109908 ( n32055, n31861, n32002 );
nand U109909 ( n32054, n76779, n3567 );
nand U109910 ( n21545, n21546, n21547 );
nor U109911 ( n21547, n21548, n21549 );
nor U109912 ( n21546, n21550, n21551 );
nor U109913 ( n21548, n21355, n74251 );
nor U109914 ( n21535, n21379, n74128 );
nand U109915 ( n66635, n66657, n66658 );
or U109916 ( n66658, n66484, n66605 );
nand U109917 ( n66657, n76713, n6182 );
nand U109918 ( n24800, n24822, n24823 );
or U109919 ( n24823, n24647, n24770 );
nand U109920 ( n24822, n76761, n4404 );
nand U109921 ( n57934, n57956, n57957 );
or U109922 ( n57957, n57783, n57904 );
nand U109923 ( n57956, n76694, n7037 );
nor U109924 ( n54502, n54337, n73650 );
nor U109925 ( n54430, n54431, n54432 );
nor U109926 ( n54432, n48005, n73975 );
nor U109927 ( n54431, n54368, n73994 );
nand U109928 ( n32104, n32121, n32122 );
or U109929 ( n32122, n31861, n32081 );
nand U109930 ( n32121, n76779, n3568 );
nand U109931 ( n45710, n45731, n45732 );
or U109932 ( n45732, n45559, n45681 );
nand U109933 ( n45731, n76665, n7970 );
nand U109934 ( n66707, n66767, n66768 );
or U109935 ( n66768, n66484, n66684 );
nand U109936 ( n66767, n76713, n6183 );
nand U109937 ( n24872, n24889, n24890 );
or U109938 ( n24890, n24647, n24849 );
nand U109939 ( n24889, n76761, n4405 );
nand U109940 ( n58009, n58026, n58027 );
or U109941 ( n58027, n57783, n57983 );
nand U109942 ( n58026, n76694, n7038 );
xor U109943 ( n17049, n17050, n17051 );
nor U109944 ( n17050, n73015, n17053 );
nor U109945 ( n17051, n73414, n17052 );
nor U109946 ( n21597, n21598, n21599 );
nor U109947 ( n21599, n14797, n74089 );
nor U109948 ( n21598, n21385, n74099 );
nand U109949 ( n32153, n32154, n32155 );
nand U109950 ( n32155, n76779, n32138 );
or U109951 ( n50052, n50030, n73426 );
nand U109952 ( n45632, n45654, n45655 );
or U109953 ( n45655, n45559, n45592 );
nand U109954 ( n45654, n76665, n7969 );
nand U109955 ( n66799, n66800, n66801 );
nand U109956 ( n66801, n76713, n66784 );
nand U109957 ( n45848, n45849, n45850 );
nand U109958 ( n45850, n76665, n45833 );
nand U109959 ( n24921, n24922, n24923 );
nand U109960 ( n24923, n76761, n24906 );
nand U109961 ( n58058, n58059, n58060 );
nand U109962 ( n58060, n76694, n58043 );
nand U109963 ( n31953, n31975, n31976 );
or U109964 ( n31976, n31861, n31894 );
nand U109965 ( n31975, n76779, n3565 );
nand U109966 ( n66863, n66864, n66865 );
nand U109967 ( n66865, n76713, n66847 );
nand U109968 ( n45912, n45913, n45914 );
nand U109969 ( n45914, n76665, n45896 );
nand U109970 ( n24987, n24988, n24989 );
nand U109971 ( n24989, n76761, n24971 );
nand U109972 ( n58122, n58123, n58124 );
nand U109973 ( n58124, n76694, n58106 );
nand U109974 ( n32296, n32297, n32298 );
nand U109975 ( n32298, n76780, n32277 );
nor U109976 ( n21565, n21379, n74232 );
nand U109977 ( n21559, n21560, n21561 );
nor U109978 ( n21561, n21562, n21563 );
nor U109979 ( n21560, n21564, n21565 );
nor U109980 ( n21563, n21375, n74241 );
nand U109981 ( n31848, n32572, n32573 );
nand U109982 ( n24721, n24743, n24744 );
or U109983 ( n24744, n24647, n24682 );
nand U109984 ( n24743, n76761, n4403 );
nand U109985 ( n66556, n66578, n66579 );
or U109986 ( n66579, n66484, n66517 );
nand U109987 ( n66578, n76713, n6180 );
nand U109988 ( n57855, n57877, n57878 );
or U109989 ( n57878, n57783, n57816 );
nand U109990 ( n57877, n76694, n7035 );
nand U109991 ( n4471, n32554, n32555 );
nor U109992 ( n32554, n32563, n32564 );
nor U109993 ( n32555, n32556, n32557 );
nor U109994 ( n32564, n73164, n76781 );
nand U109995 ( n66935, n66936, n66937 );
nand U109996 ( n66937, n76714, n66916 );
nand U109997 ( n45984, n45985, n45986 );
nand U109998 ( n45986, n76666, n45965 );
nand U109999 ( n25059, n25060, n25061 );
nand U110000 ( n25061, n76762, n25040 );
nand U110001 ( n58194, n58195, n58196 );
nand U110002 ( n58196, n76695, n58175 );
nor U110003 ( n21489, n21354, n74376 );
nand U110004 ( n13294, n4848, n12119 );
nor U110005 ( n21496, n21368, n74373 );
nor U110006 ( n54449, n54351, n73892 );
nand U110007 ( n33063, n3103, n32147 );
nand U110008 ( n11773, n11794, n11795 );
nor U110009 ( n11794, n4794, n11798 );
nand U110010 ( n11795, n76732, n11797 );
nor U110011 ( n11798, n11799, n11800 );
nor U110012 ( n21594, n21380, n74072 );
nor U110013 ( n21555, n21364, n74247 );
nand U110014 ( n21544, n21552, n21553 );
nor U110015 ( n21552, n21556, n21557 );
nor U110016 ( n21553, n21554, n21555 );
nor U110017 ( n21556, n21368, n74253 );
and U110018 ( n12029, n12003, n76731 );
nand U110019 ( n46772, n7490, n45842 );
not U110020 ( n5160, n9380 );
nor U110021 ( n54515, n54359, n73648 );
nor U110022 ( n21398, n21359, n73985 );
nand U110023 ( n67819, n5704, n66793 );
nand U110024 ( n25816, n3947, n24915 );
nand U110025 ( n58954, n6579, n58052 );
and U110026 ( n11943, n11912, n76731 );
nor U110027 ( n54419, n54351, n73993 );
nand U110028 ( n33266, n76774, n32304 );
nand U110029 ( n13552, n76727, n12318 );
nand U110030 ( n46990, n76660, n45992 );
nand U110031 ( n11839, n11840, n11842 );
nor U110032 ( n11840, n11843, n11844 );
nor U110033 ( n11844, n11809, n11800 );
and U110034 ( n11843, n11813, n76731 );
nand U110035 ( n26022, n76754, n25067 );
nand U110036 ( n59163, n76687, n58202 );
nand U110037 ( n68025, n76708, n66943 );
nor U110038 ( n21465, n21364, n74288 );
nor U110039 ( n32283, n33236, n33185 );
and U110040 ( n33236, n74855, n33237 );
nand U110041 ( n33237, n33234, n33238 );
nor U110042 ( n21461, n21358, n74285 );
nor U110043 ( n12292, n13509, n13445 );
and U110044 ( n13509, n74823, n13510 );
nand U110045 ( n13510, n13507, n13512 );
nor U110046 ( n45971, n46956, n46894 );
and U110047 ( n46956, n74822, n46957 );
nand U110048 ( n46957, n46954, n46958 );
nor U110049 ( n54545, n54359, n73813 );
nor U110050 ( n21566, n21570, n21571 );
nor U110051 ( n21570, n21389, n74252 );
nor U110052 ( n21571, n21388, n74245 );
nor U110053 ( n21435, n21364, n74325 );
nor U110054 ( n66922, n67991, n67941 );
and U110055 ( n67991, n74852, n67992 );
nand U110056 ( n67992, n67989, n67993 );
nor U110057 ( n25046, n25988, n25938 );
and U110058 ( n25988, n74853, n25989 );
nand U110059 ( n25989, n25986, n25990 );
nor U110060 ( n58181, n59126, n59076 );
and U110061 ( n59126, n74854, n59127 );
nand U110062 ( n59127, n59124, n59128 );
nor U110063 ( n21431, n21358, n74322 );
nand U110064 ( n12297, n12298, n12299 );
nand U110065 ( n12298, n8957, n12118 );
nand U110066 ( n12299, n76729, n12300 );
nand U110067 ( n9026, n12293, n12294 );
nor U110068 ( n12293, n12312, n12313 );
nor U110069 ( n12294, n12295, n12297 );
nor U110070 ( n12312, n74861, n76735 );
nor U110071 ( n54540, n54350, n73820 );
nor U110072 ( n21549, n21354, n74250 );
nor U110073 ( n33055, n74610, n76021 );
nor U110074 ( n21502, n21376, n74367 );
nor U110075 ( n21477, n21478, n21479 );
nor U110076 ( n21479, n14797, n74289 );
nor U110077 ( n21478, n21385, n74293 );
nor U110078 ( n54442, n54337, n73889 );
nor U110079 ( n21476, n21480, n21481 );
nor U110080 ( n21480, n21389, n74287 );
nor U110081 ( n21481, n21388, n74283 );
nor U110082 ( n21475, n21379, n74280 );
nor U110083 ( n21526, n21368, n74162 );
nand U110084 ( n24634, n25330, n25331 );
nand U110085 ( n66471, n67337, n67338 );
nand U110086 ( n57766, n58469, n58470 );
nor U110087 ( n21519, n21354, n74156 );
nand U110088 ( n11206, n67319, n67320 );
nor U110089 ( n67319, n67328, n67329 );
nor U110090 ( n67320, n67321, n67322 );
nor U110091 ( n67329, n73163, n76715 );
nand U110092 ( n6716, n25312, n25313 );
nor U110093 ( n25312, n25321, n25322 );
nor U110094 ( n25313, n25314, n25315 );
nor U110095 ( n25322, n72958, n76763 );
nand U110096 ( n13451, n58451, n58452 );
nor U110097 ( n58451, n58460, n58461 );
nor U110098 ( n58452, n58453, n58454 );
nor U110099 ( n58461, n72959, n76696 );
nor U110100 ( n21447, n21448, n21449 );
nor U110101 ( n21449, n14797, n74326 );
nor U110102 ( n21448, n21385, n74330 );
nor U110103 ( n54412, n54337, n73976 );
nor U110104 ( n21446, n21450, n21451 );
nor U110105 ( n21450, n21389, n74324 );
nor U110106 ( n21451, n21388, n74320 );
nor U110107 ( n21445, n21379, n74319 );
nor U110108 ( n21580, n21359, n74093 );
nand U110109 ( n11963, n11998, n11999 );
or U110110 ( n11999, n11800, n11945 );
nand U110111 ( n11998, n76732, n5315 );
nor U110112 ( n54550, n54551, n54552 );
nor U110113 ( n54552, n48005, n73814 );
nor U110114 ( n54551, n54368, n73819 );
nor U110115 ( n54547, n54363, n73809 );
nand U110116 ( n11882, n11907, n11908 );
or U110117 ( n11908, n11800, n11845 );
nand U110118 ( n11907, n76732, n5314 );
nor U110119 ( n54385, n43268, n73552 );
nand U110120 ( n12127, n12128, n12129 );
nand U110121 ( n12129, n76732, n12103 );
nand U110122 ( n45629, n46276, n46277 );
nand U110123 ( n15696, n46258, n46259 );
nor U110124 ( n46258, n46267, n46268 );
nor U110125 ( n46259, n46260, n46261 );
nor U110126 ( n46268, n72962, n76667 );
nor U110127 ( n21532, n21376, n74154 );
nand U110128 ( n12308, n12309, n12310 );
nand U110129 ( n12310, n76733, n12284 );
nor U110130 ( n54455, n54359, n73887 );
nor U110131 ( n39091, n74578, n39150 );
nor U110132 ( n38969, n74627, n39036 );
nor U110133 ( n38844, n74708, n38910 );
nor U110134 ( n62429, n74567, n62545 );
nor U110135 ( n54425, n54359, n73974 );
nand U110136 ( n4481, n32522, n32523 );
nor U110137 ( n32522, n32533, n32534 );
nor U110138 ( n32523, n32524, n32525 );
nor U110139 ( n32533, n73169, n76781 );
nand U110140 ( n11216, n67178, n67179 );
nor U110141 ( n67178, n67189, n67190 );
nor U110142 ( n67179, n67180, n67181 );
nor U110143 ( n67189, n73168, n76715 );
nand U110144 ( n6726, n25280, n25281 );
nor U110145 ( n25280, n25291, n25292 );
nor U110146 ( n25281, n25282, n25283 );
nor U110147 ( n25291, n72961, n76763 );
nand U110148 ( n13461, n58416, n58417 );
nor U110149 ( n58416, n58427, n58428 );
nor U110150 ( n58417, n58418, n58419 );
nor U110151 ( n58427, n72960, n76696 );
nand U110152 ( n15706, n46226, n46227 );
nor U110153 ( n46226, n46237, n46238 );
nor U110154 ( n46227, n46228, n46229 );
nor U110155 ( n46237, n72964, n76667 );
nor U110156 ( n21562, n21376, n74248 );
nand U110157 ( n13135, n76603, n74920 );
nor U110158 ( n21466, n21368, n74292 );
nor U110159 ( n21557, n21367, n74255 );
nor U110160 ( n21459, n21354, n74295 );
nor U110161 ( n54533, n54342, n73811 );
nand U110162 ( n45408, n61286, n830 );
nor U110163 ( n61286, n782, n61287 );
nor U110164 ( n61287, n76390, n61288 );
not U110165 ( n782, n41510 );
nor U110166 ( n13793, n13795, n76594 );
nor U110167 ( n13795, n13797, n13798 );
nand U110168 ( n13797, n13814, n13815 );
nand U110169 ( n13798, n13799, n13800 );
nand U110170 ( n13799, n76724, n12462 );
nand U110171 ( n13812, n13763, n76603 );
nor U110172 ( n54567, n43268, n73611 );
nor U110173 ( n21436, n21368, n74329 );
nor U110174 ( n21429, n21354, n74332 );
nand U110175 ( n7186, n24312, n24313 );
nor U110176 ( n24313, n24314, n24315 );
nor U110177 ( n24312, n24317, n24318 );
nor U110178 ( n24315, n4069, n23096 );
nand U110179 ( n13921, n57435, n57436 );
nor U110180 ( n57436, n57437, n57438 );
nor U110181 ( n57435, n57440, n57441 );
nor U110182 ( n57438, n6702, n56217 );
nand U110183 ( n4941, n31608, n31609 );
nor U110184 ( n31609, n31610, n31611 );
nor U110185 ( n31608, n31613, n31614 );
nor U110186 ( n31610, n75288, n31181 );
nand U110187 ( n11676, n65894, n65895 );
nor U110188 ( n65895, n65896, n65897 );
nor U110189 ( n65894, n65899, n65900 );
nor U110190 ( n65896, n75287, n65435 );
nand U110191 ( n4496, n32463, n32464 );
nor U110192 ( n32463, n32477, n32478 );
nor U110193 ( n32464, n32465, n32466 );
nor U110194 ( n32477, n74712, n76781 );
nand U110195 ( n11231, n67119, n67120 );
nor U110196 ( n67119, n67133, n67134 );
nor U110197 ( n67120, n67121, n67122 );
nor U110198 ( n67133, n74711, n76715 );
nand U110199 ( n15721, n46155, n46156 );
nor U110200 ( n46155, n46169, n46170 );
nor U110201 ( n46156, n46157, n46158 );
nor U110202 ( n46169, n74728, n76667 );
nand U110203 ( n6741, n25221, n25222 );
nor U110204 ( n25221, n25235, n25236 );
nor U110205 ( n25222, n25223, n25224 );
nor U110206 ( n25235, n74710, n76763 );
nand U110207 ( n13476, n58357, n58358 );
nor U110208 ( n58357, n58371, n58372 );
nor U110209 ( n58358, n58359, n58360 );
nor U110210 ( n58371, n74709, n76696 );
nor U110211 ( n21567, n21568, n21569 );
nor U110212 ( n21569, n14797, n74249 );
nor U110213 ( n21568, n21385, n74254 );
nor U110214 ( n62302, n74674, n62363 );
nor U110215 ( n61596, n74736, n62246 );
nor U110216 ( n21402, n9303, n73998 );
nor U110217 ( n21472, n21376, n74291 );
nand U110218 ( n33383, n32345, n3142 );
nor U110219 ( n33374, n33381, n33382 );
nor U110220 ( n33381, n32714, n33385 );
nor U110221 ( n33382, n32712, n33383 );
nand U110222 ( n33385, n32343, n3173 );
nor U110223 ( n21564, n21380, n74244 );
nand U110224 ( n41312, n41456, n41457 );
nor U110225 ( n41457, n41458, n604 );
nor U110226 ( n41456, n41459, n41460 );
nor U110227 ( n41459, n41444, n41443 );
nand U110228 ( n47104, n46044, n7529 );
nor U110229 ( n47095, n47102, n47103 );
nor U110230 ( n47102, n46415, n47106 );
nor U110231 ( n47103, n46413, n47104 );
nand U110232 ( n47106, n46042, n7559 );
nand U110233 ( n13996, n57002, n57003 );
nor U110234 ( n57002, n57009, n57010 );
nor U110235 ( n57003, n57004, n57005 );
and U110236 ( n57010, n56055, n437 );
nand U110237 ( n7261, n23878, n23879 );
nor U110238 ( n23878, n23885, n23886 );
nor U110239 ( n23879, n23880, n23881 );
and U110240 ( n23886, n22937, n164 );
nand U110241 ( n5016, n31171, n31172 );
nor U110242 ( n31171, n31179, n31180 );
nor U110243 ( n31172, n31173, n31174 );
nor U110244 ( n31180, n75363, n31181 );
nand U110245 ( n11751, n65425, n65426 );
nor U110246 ( n65425, n65433, n65434 );
nor U110247 ( n65426, n65427, n65428 );
nor U110248 ( n65434, n75364, n65435 );
nand U110249 ( n12223, n12659, n12660 );
nor U110250 ( n23981, n76539, n23984 );
nand U110251 ( n23984, n4528, n74733 );
nor U110252 ( n24062, n76539, n24065 );
nand U110253 ( n24065, n4527, n74679 );
nor U110254 ( n57103, n76281, n57106 );
nand U110255 ( n57106, n7160, n74732 );
nor U110256 ( n57184, n76281, n57187 );
nand U110257 ( n57187, n7159, n74678 );
nor U110258 ( n57265, n76281, n57268 );
nand U110259 ( n57268, n7158, n75249 );
nor U110260 ( n57366, n76281, n57369 );
nand U110261 ( n57369, n7157, n74583 );
nor U110262 ( n57387, n76281, n57390 );
nand U110263 ( n57390, n7155, n74542 );
nor U110264 ( n57408, n76281, n57411 );
nand U110265 ( n57411, n7154, n74509 );
nor U110266 ( n24143, n76539, n24146 );
nand U110267 ( n24146, n4525, n75251 );
nor U110268 ( n24241, n76539, n24244 );
nand U110269 ( n24244, n4524, n74584 );
nor U110270 ( n24262, n76539, n24265 );
nand U110271 ( n24265, n4523, n74543 );
nor U110272 ( n24285, n76539, n24288 );
nand U110273 ( n24288, n4522, n74510 );
nand U110274 ( n68135, n66984, n5743 );
nand U110275 ( n26132, n25108, n3985 );
nand U110276 ( n59273, n58246, n6618 );
nand U110277 ( n7251, n23979, n23980 );
nor U110278 ( n23979, n23987, n23988 );
nor U110279 ( n23980, n23981, n23982 );
nor U110280 ( n23988, n23199, n23883 );
nand U110281 ( n7241, n24060, n24061 );
nor U110282 ( n24060, n24068, n24069 );
nor U110283 ( n24061, n24062, n24063 );
nor U110284 ( n24069, n23296, n23883 );
nand U110285 ( n7221, n24239, n24240 );
nor U110286 ( n24239, n24247, n24248 );
nor U110287 ( n24240, n24241, n24242 );
nor U110288 ( n24248, n3987, n23096 );
nand U110289 ( n7211, n24260, n24261 );
nor U110290 ( n24260, n24268, n24269 );
nor U110291 ( n24261, n24262, n24263 );
nor U110292 ( n24269, n4023, n23096 );
nand U110293 ( n7201, n24283, n24284 );
nor U110294 ( n24283, n24290, n24291 );
nor U110295 ( n24284, n24285, n24286 );
nor U110296 ( n24291, n4042, n23096 );
nor U110297 ( n68126, n68133, n68134 );
nor U110298 ( n68133, n67479, n68137 );
nor U110299 ( n68134, n67477, n68135 );
nand U110300 ( n68137, n66982, n5772 );
nor U110301 ( n26123, n26130, n26131 );
nor U110302 ( n26130, n25474, n26134 );
nor U110303 ( n26131, n25472, n26132 );
nand U110304 ( n26134, n25106, n4013 );
nor U110305 ( n59264, n59271, n59272 );
nor U110306 ( n59271, n58611, n59275 );
nor U110307 ( n59272, n58609, n59273 );
nand U110308 ( n59275, n58244, n6645 );
nor U110309 ( n31275, n76482, n31278 );
nand U110310 ( n31278, n3640, n74731 );
nor U110311 ( n31356, n76482, n31359 );
nand U110312 ( n31359, n3639, n74676 );
nor U110313 ( n65525, n76215, n65528 );
nand U110314 ( n65528, n6268, n74730 );
nor U110315 ( n65606, n76215, n65609 );
nand U110316 ( n65609, n6267, n74675 );
nor U110317 ( n31437, n76482, n31440 );
nand U110318 ( n31440, n3638, n75252 );
nor U110319 ( n31535, n76482, n31538 );
nand U110320 ( n31538, n3637, n74582 );
nor U110321 ( n31556, n76482, n31559 );
nand U110322 ( n31559, n3635, n74540 );
nor U110323 ( n31581, n76482, n31584 );
nand U110324 ( n31584, n3634, n73135 );
nor U110325 ( n65687, n76215, n65690 );
nand U110326 ( n65690, n6265, n75250 );
nor U110327 ( n65785, n76215, n65788 );
nand U110328 ( n65788, n6264, n74581 );
nor U110329 ( n65846, n76215, n65849 );
nand U110330 ( n65849, n6263, n74539 );
nor U110331 ( n65867, n76215, n65870 );
nand U110332 ( n65870, n6262, n74507 );
nand U110333 ( n4996, n31354, n31355 );
nor U110334 ( n31354, n31362, n31363 );
nor U110335 ( n31355, n31356, n31357 );
nor U110336 ( n31363, n75318, n31181 );
nand U110337 ( n13986, n57101, n57102 );
nor U110338 ( n57101, n57109, n57110 );
nor U110339 ( n57102, n57103, n57104 );
nor U110340 ( n57110, n56320, n57007 );
nand U110341 ( n13976, n57182, n57183 );
nor U110342 ( n57182, n57190, n57191 );
nor U110343 ( n57183, n57184, n57185 );
nor U110344 ( n57191, n56420, n57007 );
nand U110345 ( n13966, n57263, n57264 );
nor U110346 ( n57263, n57271, n57272 );
nor U110347 ( n57264, n57265, n57266 );
nor U110348 ( n57272, n56515, n57007 );
nand U110349 ( n13956, n57364, n57365 );
nor U110350 ( n57364, n57372, n57373 );
nor U110351 ( n57365, n57366, n57367 );
nor U110352 ( n57373, n6619, n56217 );
nand U110353 ( n13946, n57385, n57386 );
nor U110354 ( n57385, n57393, n57394 );
nor U110355 ( n57386, n57387, n57388 );
nor U110356 ( n57394, n6655, n56217 );
nand U110357 ( n13936, n57406, n57407 );
nor U110358 ( n57406, n57413, n57414 );
nor U110359 ( n57407, n57408, n57409 );
nor U110360 ( n57414, n6674, n56217 );
nand U110361 ( n13926, n57426, n57427 );
nor U110362 ( n57426, n57432, n57433 );
nor U110363 ( n57427, n57428, n57429 );
nor U110364 ( n57432, n255, n57007 );
nand U110365 ( n7231, n24141, n24142 );
nor U110366 ( n24141, n24149, n24150 );
nor U110367 ( n24142, n24143, n24144 );
nor U110368 ( n24150, n23391, n23883 );
nand U110369 ( n7191, n24303, n24304 );
nor U110370 ( n24303, n24309, n24310 );
nor U110371 ( n24304, n24305, n24306 );
nor U110372 ( n24309, n9, n23883 );
nand U110373 ( n8961, n12628, n12629 );
nor U110374 ( n12628, n12639, n12640 );
nor U110375 ( n12629, n12630, n12632 );
nor U110376 ( n12640, n72963, n76734 );
nand U110377 ( n5006, n31273, n31274 );
nor U110378 ( n31273, n31281, n31282 );
nor U110379 ( n31274, n31275, n31276 );
nor U110380 ( n31282, n75316, n31181 );
nand U110381 ( n11741, n65523, n65524 );
nor U110382 ( n65523, n65531, n65532 );
nor U110383 ( n65524, n65525, n65526 );
nor U110384 ( n65532, n75305, n65435 );
nand U110385 ( n11731, n65604, n65605 );
nor U110386 ( n65604, n65612, n65613 );
nor U110387 ( n65605, n65606, n65607 );
nor U110388 ( n65613, n75307, n65435 );
nand U110389 ( n4986, n31435, n31436 );
nor U110390 ( n31435, n31443, n31444 );
nor U110391 ( n31436, n31437, n31438 );
nor U110392 ( n31444, n75319, n31181 );
nand U110393 ( n4976, n31533, n31534 );
nor U110394 ( n31533, n31541, n31542 );
nor U110395 ( n31534, n31535, n31536 );
nor U110396 ( n31541, n75315, n31181 );
nand U110397 ( n4966, n31554, n31555 );
nor U110398 ( n31554, n31562, n31563 );
nor U110399 ( n31555, n31556, n31557 );
nor U110400 ( n31562, n75312, n31181 );
nand U110401 ( n4956, n31579, n31580 );
nor U110402 ( n31579, n31586, n31587 );
nor U110403 ( n31580, n31581, n31582 );
nor U110404 ( n31586, n75298, n31181 );
nand U110405 ( n4946, n31599, n31600 );
nor U110406 ( n31599, n31605, n31606 );
nor U110407 ( n31600, n31601, n31602 );
nor U110408 ( n31605, n75297, n31181 );
nand U110409 ( n11681, n65885, n65886 );
nor U110410 ( n65885, n65891, n65892 );
nor U110411 ( n65886, n65887, n65888 );
nor U110412 ( n65891, n75295, n65435 );
nand U110413 ( n13695, n12369, n4884 );
nor U110414 ( n13684, n13693, n13694 );
nor U110415 ( n13693, n13060, n13698 );
nor U110416 ( n13694, n13055, n13695 );
nand U110417 ( n13698, n12367, n4910 );
nand U110418 ( n11721, n65685, n65686 );
nor U110419 ( n65685, n65693, n65694 );
nor U110420 ( n65686, n65687, n65688 );
nor U110421 ( n65694, n75308, n65435 );
nand U110422 ( n11711, n65783, n65784 );
nor U110423 ( n65783, n65791, n65792 );
nor U110424 ( n65784, n65785, n65786 );
nor U110425 ( n65791, n75294, n65435 );
nand U110426 ( n11701, n65844, n65845 );
nor U110427 ( n65844, n65852, n65853 );
nor U110428 ( n65845, n65846, n65847 );
nor U110429 ( n65852, n75291, n65435 );
nand U110430 ( n11691, n65865, n65866 );
nor U110431 ( n65865, n65872, n65873 );
nor U110432 ( n65866, n65867, n65868 );
nor U110433 ( n65872, n75289, n65435 );
nor U110434 ( n21442, n21376, n74328 );
nand U110435 ( n8971, n12588, n12589 );
nor U110436 ( n12588, n12602, n12603 );
nor U110437 ( n12589, n12590, n12592 );
nor U110438 ( n12602, n72965, n76734 );
nand U110439 ( n32239, n76779, n32201 );
nand U110440 ( n31883, n31884, n74912 );
nand U110441 ( n31884, n31885, n31886 );
nand U110442 ( n31885, n3055, n31868 );
nand U110443 ( n31886, n31887, n76778 );
nand U110444 ( n32070, n32071, n74752 );
nand U110445 ( n32071, n32072, n32073 );
nand U110446 ( n32072, n3055, n32056 );
nand U110447 ( n32073, n32074, n76778 );
nor U110448 ( n49558, n50030, n76834 );
nand U110449 ( n66506, n66507, n74913 );
nand U110450 ( n66507, n66508, n66509 );
nand U110451 ( n66508, n5657, n66491 );
nand U110452 ( n66509, n66510, n76712 );
nand U110453 ( n24671, n24672, n74910 );
nand U110454 ( n24672, n24673, n24674 );
nand U110455 ( n24673, n3899, n24654 );
nand U110456 ( n24674, n24675, n76760 );
nand U110457 ( n57805, n57806, n74911 );
nand U110458 ( n57806, n57807, n57808 );
nand U110459 ( n57807, n6532, n57790 );
nand U110460 ( n57808, n57809, n76693 );
nand U110461 ( n66673, n66674, n74751 );
nand U110462 ( n66674, n66675, n66676 );
nand U110463 ( n66675, n5657, n66659 );
nand U110464 ( n66676, n66677, n76712 );
nand U110465 ( n57972, n57973, n74754 );
nand U110466 ( n57973, n57974, n57975 );
nand U110467 ( n57974, n6532, n57958 );
nand U110468 ( n57975, n57976, n76693 );
nand U110469 ( n31991, n31992, n75044 );
nand U110470 ( n31992, n31993, n31994 );
nand U110471 ( n31993, n3055, n31977 );
nand U110472 ( n31994, n31995, n76778 );
nand U110473 ( n45581, n45582, n75077 );
nand U110474 ( n45582, n45583, n45584 );
nand U110475 ( n45583, n7430, n45566 );
nand U110476 ( n45584, n45585, n76664 );
nand U110477 ( n24838, n24839, n74753 );
nand U110478 ( n24839, n24840, n24841 );
nand U110479 ( n24840, n3899, n24824 );
nand U110480 ( n24841, n24842, n76760 );
nor U110481 ( n38111, n38119, n38120 );
nand U110482 ( n45670, n45671, n74810 );
nand U110483 ( n45671, n45672, n45673 );
nand U110484 ( n45672, n7430, n45656 );
nand U110485 ( n45673, n45674, n76664 );
nand U110486 ( n66594, n66595, n75045 );
nand U110487 ( n66595, n66596, n66597 );
nand U110488 ( n66596, n5657, n66580 );
nand U110489 ( n66597, n66598, n76712 );
nand U110490 ( n45765, n45766, n74998 );
nand U110491 ( n45766, n45767, n45768 );
nand U110492 ( n45767, n7430, n45733 );
nand U110493 ( n45768, n45769, n76664 );
nand U110494 ( n24759, n24760, n75043 );
nand U110495 ( n24760, n24761, n24762 );
nand U110496 ( n24761, n3899, n24745 );
nand U110497 ( n24762, n24763, n76760 );
nand U110498 ( n57893, n57894, n75046 );
nand U110499 ( n57894, n57895, n57896 );
nand U110500 ( n57895, n6532, n57879 );
nand U110501 ( n57896, n57897, n76693 );
nor U110502 ( n54345, n43268, n73556 );
nor U110503 ( n21584, n9303, n74111 );
nand U110504 ( n54331, n54343, n54344 );
nor U110505 ( n54343, n54348, n54349 );
nor U110506 ( n54344, n54345, n54346 );
nor U110507 ( n54349, n54350, n73574 );
nor U110508 ( n21550, n21359, n74246 );
nor U110509 ( n54335, n54338, n73567 );
nand U110510 ( n54332, n54333, n54334 );
nor U110511 ( n54333, n54339, n54340 );
nor U110512 ( n54334, n54335, n54336 );
nor U110513 ( n54339, n54342, n73560 );
nand U110514 ( n8986, n12514, n12515 );
nor U110515 ( n12514, n12532, n12533 );
nor U110516 ( n12515, n12517, n12518 );
nor U110517 ( n12532, n74729, n76734 );
not U110518 ( n7794, n54228 );
nand U110519 ( n9001, n12438, n12439 );
nor U110520 ( n12438, n12457, n12458 );
nor U110521 ( n12439, n12440, n12442 );
nor U110522 ( n12457, n73222, n76734 );
nor U110523 ( n54357, n54358, n73555 );
nand U110524 ( n54353, n54354, n54355 );
nor U110525 ( n54354, n54360, n54361 );
nor U110526 ( n54355, n54356, n54357 );
nor U110527 ( n54360, n54363, n73557 );
nand U110528 ( n32211, n32212, n32213 );
nand U110529 ( n32213, n32214, n76480 );
nand U110530 ( n32212, n32217, n76785 );
and U110531 ( n32214, n32215, n32216 );
and U110532 ( n32217, n32218, n32219 );
and U110533 ( n32363, n32379, n76778 );
nor U110534 ( n32379, n73112, n32339 );
and U110535 ( n32434, n32454, n76778 );
nor U110536 ( n32454, n74503, n32409 );
nand U110537 ( n12199, n12200, n12202 );
nand U110538 ( n12202, n12203, n76607 );
nand U110539 ( n12200, n12207, n76737 );
and U110540 ( n12203, n12204, n12205 );
and U110541 ( n12207, n12208, n12209 );
nand U110542 ( n40710, n40711, n40712 );
nand U110543 ( n40712, n583, n40713 );
nand U110544 ( n40711, n1787, n40714 );
not U110545 ( n1787, n40715 );
nand U110546 ( n40744, n40745, n40746 );
nand U110547 ( n40746, n583, n40747 );
nand U110548 ( n40745, n1782, n40714 );
not U110549 ( n1782, n40748 );
nand U110550 ( n40910, n40911, n40912 );
nand U110551 ( n40912, n583, n40913 );
nand U110552 ( n40911, n1779, n40714 );
not U110553 ( n1779, n40914 );
and U110554 ( n67026, n67042, n76712 );
nor U110555 ( n67042, n73110, n66978 );
and U110556 ( n67090, n67110, n76712 );
nor U110557 ( n67110, n74502, n67072 );
and U110558 ( n46062, n46078, n76664 );
nor U110559 ( n46078, n73108, n46038 );
and U110560 ( n46126, n46146, n76664 );
nor U110561 ( n46146, n74500, n46108 );
and U110562 ( n25126, n25142, n76760 );
nor U110563 ( n25142, n73113, n25102 );
and U110564 ( n25192, n25212, n76760 );
nor U110565 ( n25212, n74504, n25174 );
and U110566 ( n58264, n58280, n76693 );
nor U110567 ( n58280, n73111, n58240 );
and U110568 ( n58328, n58348, n76693 );
nor U110569 ( n58348, n74505, n58310 );
nand U110570 ( n32453, n32434, n73102 );
nand U110571 ( n67109, n67090, n73100 );
nand U110572 ( n25211, n25192, n73103 );
nand U110573 ( n58347, n58328, n73101 );
nand U110574 ( n46145, n46126, n73098 );
nor U110575 ( n54346, n54347, n73561 );
nor U110576 ( n54340, n54341, n73554 );
not U110577 ( n7, n11600 );
nand U110578 ( n12237, n76732, n12187 );
nor U110579 ( n54537, n43268, n73808 );
nor U110580 ( n21362, n9303, n74019 );
nand U110581 ( n21348, n21360, n21361 );
nor U110582 ( n21360, n21365, n21366 );
nor U110583 ( n21361, n21362, n21363 );
nor U110584 ( n21366, n21367, n74061 );
nand U110585 ( n11835, n11837, n76731 );
nor U110586 ( n11837, n11813, n11838 );
nand U110587 ( n12018, n12019, n74997 );
nand U110588 ( n12019, n12020, n12022 );
nand U110589 ( n12020, n4787, n12000 );
nand U110590 ( n12022, n12023, n76731 );
nand U110591 ( n11932, n11933, n74808 );
nand U110592 ( n11933, n11934, n11935 );
nand U110593 ( n11934, n4787, n11909 );
nand U110594 ( n11935, n11937, n76731 );
or U110595 ( n16804, n17047, n73012 );
nor U110596 ( n54364, n54369, n54370 );
nor U110597 ( n54369, n54372, n73570 );
nor U110598 ( n54370, n54371, n73559 );
nor U110599 ( n54361, n54362, n73553 );
nand U110600 ( n32943, n76022, n75050 );
nor U110601 ( n21352, n21355, n74045 );
nand U110602 ( n21349, n21350, n21351 );
nor U110603 ( n21350, n21356, n21357 );
nor U110604 ( n21351, n21352, n21353 );
nor U110605 ( n21356, n21359, n74035 );
not U110606 ( n5139, n21230 );
nor U110607 ( n21374, n21375, n74017 );
nand U110608 ( n21370, n21371, n21372 );
nor U110609 ( n21371, n21377, n21378 );
nor U110610 ( n21372, n21373, n21374 );
nor U110611 ( n21377, n21380, n74026 );
nor U110612 ( n54365, n54366, n54367 );
nor U110613 ( n54367, n48005, n73563 );
nor U110614 ( n54366, n54368, n73572 );
and U110615 ( n71325, n71665, n71666 );
nor U110616 ( n71665, n71669, n71670 );
nor U110617 ( n71666, n71667, n71668 );
nor U110618 ( n71670, n74441, n73026 );
and U110619 ( n12392, n12418, n76731 );
nor U110620 ( n12418, n73107, n12362 );
and U110621 ( n12478, n12503, n76731 );
nor U110622 ( n12503, n74506, n12455 );
nor U110623 ( n71667, n74434, n71105 );
xnor U110624 ( n12419, n13759, n13760 );
xor U110625 ( n13760, n74735, n76035 );
nand U110626 ( n13759, n13717, n13720 );
nor U110627 ( n13743, n13745, n76594 );
nor U110628 ( n13745, n13747, n13748 );
nand U110629 ( n13747, n13767, n13768 );
nand U110630 ( n13748, n13749, n13750 );
nand U110631 ( n9436, n11294, n11295 );
nor U110632 ( n11295, n11297, n11298 );
nor U110633 ( n11294, n11302, n11303 );
nor U110634 ( n11297, n9908, n11300 );
nand U110635 ( n12414, n12415, n12417 );
nand U110636 ( n12415, n76729, n12419 );
nand U110637 ( n12417, n12392, n74577 );
nand U110638 ( n12493, n12500, n12502 );
nand U110639 ( n12500, n76608, n12504 );
nand U110640 ( n12502, n12478, n73097 );
nor U110641 ( n21554, n9303, n74243 );
xor U110642 ( n32206, n32215, n74635 );
xor U110643 ( n12193, n12204, n74599 );
nor U110644 ( n54348, n54351, n73571 );
xor U110645 ( n45901, n45921, n74524 );
xor U110646 ( n66852, n66872, n74546 );
xor U110647 ( n24976, n24996, n74547 );
xor U110648 ( n58111, n58131, n74548 );
xor U110649 ( n50027, n75836, n75837 );
nor U110650 ( n75836, n50031, n73421 );
nor U110651 ( n75837, n50030, n73021 );
nor U110652 ( n21363, n21364, n74037 );
nor U110653 ( n21357, n21358, n74016 );
nor U110654 ( n54336, n54337, n73565 );
nor U110655 ( n21382, n21383, n21384 );
nor U110656 ( n21384, n14797, n74039 );
nor U110657 ( n21383, n21385, n74060 );
nor U110658 ( n21381, n21386, n21387 );
nor U110659 ( n21386, n21389, n74052 );
nor U110660 ( n21387, n21388, n74031 );
nor U110661 ( n21378, n21379, n74005 );
nand U110662 ( n41040, n41041, n40696 );
nand U110663 ( n32257, n32258, n32259 );
nand U110664 ( n32259, n76480, n32260 );
nand U110665 ( n32258, n76785, n32261 );
nand U110666 ( n45945, n45946, n45947 );
nand U110667 ( n45947, n76346, n45948 );
nand U110668 ( n45946, n76671, n45949 );
nand U110669 ( n12259, n12260, n12262 );
nand U110670 ( n12262, n76607, n12263 );
nand U110671 ( n12260, n76738, n12264 );
nand U110672 ( n66896, n66897, n66898 );
nand U110673 ( n66898, n76202, n66899 );
nand U110674 ( n66897, n76719, n66900 );
nand U110675 ( n25020, n25021, n25022 );
nand U110676 ( n25022, n76526, n25023 );
nand U110677 ( n25021, n76767, n25024 );
nand U110678 ( n58155, n58156, n58157 );
nand U110679 ( n58157, n76268, n58158 );
nand U110680 ( n58156, n76700, n58159 );
nand U110681 ( n40788, n40696, n75248 );
nor U110682 ( n17122, n17129, n75919 );
nor U110683 ( n54356, n54359, n73562 );
nor U110684 ( n71669, n74436, n71108 );
nand U110685 ( n4476, n32539, n32540 );
nor U110686 ( n32539, n32548, n32549 );
nor U110687 ( n32540, n32541, n32542 );
nor U110688 ( n32548, n74699, n31969 );
nor U110689 ( n21365, n21368, n74059 );
nor U110690 ( n21353, n21354, n74043 );
nand U110691 ( n11211, n67195, n67196 );
nor U110692 ( n67195, n67204, n67205 );
nor U110693 ( n67196, n67197, n67198 );
nor U110694 ( n67204, n74700, n66572 );
nand U110695 ( n15701, n46243, n46244 );
nor U110696 ( n46243, n46252, n46253 );
nor U110697 ( n46244, n46245, n46246 );
nor U110698 ( n46252, n74717, n45648 );
nand U110699 ( n6721, n25297, n25298 );
nor U110700 ( n25297, n25306, n25307 );
nor U110701 ( n25298, n25299, n25300 );
nor U110702 ( n25306, n74701, n24737 );
nand U110703 ( n13456, n58436, n58437 );
nor U110704 ( n58436, n58445, n58446 );
nor U110705 ( n58437, n58438, n58439 );
nor U110706 ( n58445, n74702, n57871 );
nand U110707 ( n32144, n76480, n32147 );
nand U110708 ( n12115, n76607, n12119 );
nand U110709 ( n45839, n76346, n45842 );
nand U110710 ( n32300, n32301, n32302 );
nand U110711 ( n32302, n76480, n32303 );
nand U110712 ( n32301, n76786, n32304 );
nand U110713 ( n12313, n12314, n12315 );
nand U110714 ( n12315, n76607, n12317 );
nand U110715 ( n12314, n76739, n12318 );
nand U110716 ( n66790, n76202, n66793 );
nand U110717 ( n45988, n45989, n45990 );
nand U110718 ( n45990, n76346, n45991 );
nand U110719 ( n45989, n76672, n45992 );
nand U110720 ( n24912, n76526, n24915 );
nand U110721 ( n58049, n76268, n58052 );
nand U110722 ( n66939, n66940, n66941 );
nand U110723 ( n66941, n76202, n66942 );
nand U110724 ( n66940, n76720, n66943 );
nand U110725 ( n25063, n25064, n25065 );
nand U110726 ( n25065, n76526, n25066 );
nand U110727 ( n25064, n76768, n25067 );
nand U110728 ( n58198, n58199, n58200 );
nand U110729 ( n58200, n76268, n58201 );
nand U110730 ( n58199, n76701, n58202 );
nand U110731 ( n13290, n76603, n13247 );
nand U110732 ( n12975, n76603, n74886 );
nor U110733 ( n21373, n21376, n74038 );
nor U110734 ( n17623, n17077, n73423 );
nand U110735 ( n13604, n76727, n12345 );
xor U110736 ( n45203, n45204, n45205 );
xor U110737 ( n45205, n74475, n847 );
nand U110738 ( n45204, n45206, n45207 );
nand U110739 ( n45207, n850, n45077 );
nand U110740 ( n44393, n45218, n45219 );
nand U110741 ( n45219, n45220, n45221 );
nand U110742 ( n45218, n45228, n862 );
nand U110743 ( n45221, n45222, n45223 );
nand U110744 ( n42959, n45245, n45246 );
nand U110745 ( n45246, n894, n42678 );
nor U110746 ( n45245, n45247, n45248 );
nor U110747 ( n45248, n45249, n74337 );
nand U110748 ( n42431, n45251, n45252 );
nand U110749 ( n45252, n904, n42344 );
nor U110750 ( n45251, n45253, n45254 );
nor U110751 ( n45254, n45255, n74263 );
nand U110752 ( n45085, n45017, n45019 );
nor U110753 ( n45259, n45260, n45261 );
nor U110754 ( n45261, n73829, n45262 );
nor U110755 ( n45260, n45263, n45264 );
nand U110756 ( n45262, n42257, n42229 );
nand U110757 ( n45264, n42257, n42231 );
nand U110758 ( n43880, n45231, n45232 );
nand U110759 ( n45232, n45233, n45234 );
nand U110760 ( n45231, n45241, n873 );
nand U110761 ( n45234, n45235, n45236 );
nor U110762 ( n45206, n45208, n45209 );
nor U110763 ( n45209, n45210, n74449 );
nor U110764 ( n45208, n45211, n45085 );
nor U110765 ( n45210, n850, n45077 );
nand U110766 ( n8966, n12609, n12610 );
nor U110767 ( n12609, n12620, n12622 );
nor U110768 ( n12610, n12612, n12613 );
nor U110769 ( n12620, n74718, n11899 );
nand U110770 ( n33310, n76774, n32326 );
nand U110771 ( n12458, n12459, n12460 );
nand U110772 ( n12459, n12463, n76737 );
nand U110773 ( n12460, n76730, n12462 );
nand U110774 ( n47036, n76660, n46025 );
nand U110775 ( n68067, n76708, n66965 );
nand U110776 ( n26064, n76754, n25089 );
nand U110777 ( n59205, n76687, n58224 );
nand U110778 ( n71326, n72886, n72887 );
nor U110779 ( n72886, n72895, n72896 );
nor U110780 ( n72887, n72888, n72889 );
nor U110781 ( n72896, n74447, n73026 );
nor U110782 ( n17115, n17077, n75919 );
nor U110783 ( n1071, n76638, n74623 );
nor U110784 ( n996, n76638, n74624 );
nor U110785 ( n50359, n50034, n73425 );
not U110786 ( n917, n45201 );
nand U110787 ( n44390, n45153, n45154 );
nand U110788 ( n45154, n45155, n45156 );
nand U110789 ( n45153, n45163, n863 );
nand U110790 ( n45156, n45157, n45158 );
nand U110791 ( n42955, n45179, n45180 );
nand U110792 ( n45180, n895, n42678 );
nor U110793 ( n45179, n45181, n45182 );
nor U110794 ( n45182, n45183, n74336 );
nand U110795 ( n43557, n45166, n45167 );
nand U110796 ( n45167, n45168, n45169 );
nand U110797 ( n45166, n45176, n877 );
nand U110798 ( n45169, n45170, n45171 );
nand U110799 ( n42423, n45186, n45187 );
nand U110800 ( n45187, n905, n42344 );
nor U110801 ( n45186, n45188, n45189 );
nor U110802 ( n45189, n45190, n74259 );
nand U110803 ( n45076, n45009, n45011 );
nand U110804 ( n42212, n917, n73827 );
nand U110805 ( n45139, n45141, n45142 );
nand U110806 ( n45142, n852, n45077 );
nor U110807 ( n45141, n45143, n45144 );
nor U110808 ( n45144, n45145, n74448 );
nor U110809 ( n45194, n45195, n45196 );
nor U110810 ( n45196, n73826, n45197 );
nor U110811 ( n45195, n45198, n45199 );
nand U110812 ( n45197, n42247, n42229 );
nand U110813 ( n42227, n42211, n45200 );
nand U110814 ( n45200, n42209, n42212 );
nand U110815 ( n33454, n32387, n32386 );
nand U110816 ( n13783, n12428, n12427 );
nand U110817 ( n47174, n46086, n46085 );
nand U110818 ( n68205, n67050, n67049 );
nand U110819 ( n26204, n25150, n25149 );
nand U110820 ( n59343, n58288, n58287 );
nor U110821 ( n13417, n76034, n74818 );
nand U110822 ( n13462, n4848, n12263 );
nand U110823 ( n33198, n3103, n32260 );
nand U110824 ( n46907, n7490, n45948 );
nand U110825 ( n33395, n76774, n32372 );
nand U110826 ( n67954, n5704, n66899 );
nand U110827 ( n25951, n3947, n25023 );
nand U110828 ( n59089, n6579, n58158 );
nand U110829 ( n47116, n76660, n46071 );
xnor U110830 ( n37898, n37899, n37900 );
xor U110831 ( n37900, n74398, n37897 );
nand U110832 ( n68147, n76708, n67035 );
nand U110833 ( n26146, n76754, n25135 );
nand U110834 ( n59285, n76687, n58273 );
nand U110835 ( n13710, n76727, n12403 );
nand U110836 ( n45081, n45082, n45019 );
nand U110837 ( n45082, n857, n45018 );
nor U110838 ( n45078, n45079, n45080 );
nor U110839 ( n45079, n45083, n45084 );
nor U110840 ( n45080, n853, n45081 );
nand U110841 ( n45084, n45085, n45018 );
not U110842 ( n857, n45017 );
nor U110843 ( n50045, n50034, n73426 );
xor U110844 ( n12473, n13848, n13763 );
nor U110845 ( n13839, n13842, n76594 );
nor U110846 ( n13842, n13843, n13844 );
nand U110847 ( n13843, n13864, n13865 );
nand U110848 ( n13844, n13845, n13847 );
not U110849 ( n422, n61735 );
not U110850 ( n149, n28430 );
not U110851 ( n187, n35607 );
not U110852 ( n458, n70335 );
nand U110853 ( n34240, n35688, n35689 );
nand U110854 ( n35689, n3410, n35685 );
nor U110855 ( n35688, n35690, n35691 );
nor U110856 ( n35691, n31612, n34130 );
nand U110857 ( n26995, n28509, n28510 );
nand U110858 ( n28510, n4248, n28506 );
nor U110859 ( n28509, n28511, n28512 );
nor U110860 ( n28512, n24316, n26885 );
nand U110861 ( n68994, n70414, n70415 );
nand U110862 ( n70415, n6025, n70411 );
nor U110863 ( n70414, n70416, n70417 );
nor U110864 ( n70417, n65898, n68884 );
nand U110865 ( n60138, n61814, n61815 );
nand U110866 ( n61815, n6880, n61811 );
nor U110867 ( n61814, n61816, n61817 );
nor U110868 ( n61817, n57439, n60025 );
nand U110869 ( n35610, n35644, n35645 );
nor U110870 ( n35644, n29190, n35700 );
nor U110871 ( n35645, n35646, n35647 );
nand U110872 ( n35700, n35701, n35702 );
nand U110873 ( n28433, n28465, n28466 );
nor U110874 ( n28465, n21873, n28521 );
nor U110875 ( n28466, n28467, n28468 );
nand U110876 ( n28521, n28522, n28523 );
nand U110877 ( n70338, n70370, n70371 );
nor U110878 ( n70370, n62908, n70426 );
nor U110879 ( n70371, n70372, n70373 );
nand U110880 ( n70426, n70427, n70428 );
nand U110881 ( n61738, n61770, n61771 );
nor U110882 ( n61770, n54964, n61826 );
nor U110883 ( n61771, n61772, n61773 );
nand U110884 ( n61826, n61827, n61828 );
nor U110885 ( n35669, n35672, n35673 );
nor U110886 ( n35673, n73138, n35668 );
nor U110887 ( n35672, n34708, n35674 );
nand U110888 ( n35674, n35675, n35676 );
nor U110889 ( n28490, n28493, n28494 );
nor U110890 ( n28494, n73136, n28489 );
nor U110891 ( n28493, n27463, n28495 );
nand U110892 ( n28495, n28496, n28497 );
nor U110893 ( n70395, n70398, n70399 );
nor U110894 ( n70399, n73139, n70394 );
nor U110895 ( n70398, n69452, n70400 );
nand U110896 ( n70400, n70401, n70402 );
nor U110897 ( n61795, n61798, n61799 );
nor U110898 ( n61799, n73137, n61794 );
nor U110899 ( n61798, n60612, n61800 );
nand U110900 ( n61800, n61801, n61802 );
nor U110901 ( n35608, n35611, n74591 );
nor U110902 ( n35611, n34166, n187 );
nor U110903 ( n28431, n28434, n74592 );
nor U110904 ( n28434, n26921, n149 );
nor U110905 ( n70336, n70339, n74593 );
nor U110906 ( n70339, n68920, n458 );
nor U110907 ( n61736, n61739, n74594 );
nor U110908 ( n61739, n60061, n422 );
nand U110909 ( n35676, n35677, n35678 );
nand U110910 ( n35677, n35679, n35680 );
nand U110911 ( n35679, n34240, n34191 );
nand U110912 ( n35680, n35681, n34233 );
nand U110913 ( n28497, n28498, n28499 );
nand U110914 ( n28498, n28500, n28501 );
nand U110915 ( n28500, n26995, n26946 );
nand U110916 ( n28501, n28502, n26988 );
nand U110917 ( n70402, n70403, n70404 );
nand U110918 ( n70403, n70405, n70406 );
nand U110919 ( n70405, n68994, n68945 );
nand U110920 ( n70406, n70407, n68987 );
nand U110921 ( n61802, n61803, n61804 );
nand U110922 ( n61803, n61805, n61806 );
nand U110923 ( n61805, n60138, n60086 );
nand U110924 ( n61806, n61807, n60131 );
nand U110925 ( n35665, n35666, n35667 );
nand U110926 ( n35667, n35668, n73138 );
nand U110927 ( n35666, n35669, n35670 );
or U110928 ( n35670, n35671, n74513 );
nand U110929 ( n28486, n28487, n28488 );
nand U110930 ( n28488, n28489, n73136 );
nand U110931 ( n28487, n28490, n28491 );
or U110932 ( n28491, n28492, n74516 );
nand U110933 ( n70391, n70392, n70393 );
nand U110934 ( n70393, n70394, n73139 );
nand U110935 ( n70392, n70395, n70396 );
or U110936 ( n70396, n70397, n74514 );
nand U110937 ( n61791, n61792, n61793 );
nand U110938 ( n61793, n61794, n73137 );
nand U110939 ( n61792, n61795, n61796 );
or U110940 ( n61796, n61797, n74517 );
or U110941 ( n35681, n34240, n74561 );
or U110942 ( n28502, n26995, n74555 );
or U110943 ( n70407, n68994, n74562 );
or U110944 ( n61807, n60138, n74556 );
nand U110945 ( n3611, n35599, n35600 );
nor U110946 ( n35600, n35601, n35602 );
nor U110947 ( n35599, n35608, n35609 );
nand U110948 ( n35602, n30099, n35603 );
nand U110949 ( n5856, n28422, n28423 );
nor U110950 ( n28423, n28424, n28425 );
nor U110951 ( n28422, n28431, n28432 );
nand U110952 ( n28425, n22778, n28426 );
nand U110953 ( n10346, n70327, n70328 );
nor U110954 ( n70328, n70329, n70330 );
nor U110955 ( n70327, n70336, n70337 );
nand U110956 ( n70330, n64116, n70331 );
nand U110957 ( n12591, n61727, n61728 );
nor U110958 ( n61728, n61729, n61730 );
nor U110959 ( n61727, n61736, n61737 );
nand U110960 ( n61730, n55892, n61731 );
nor U110961 ( n54108, n54111, n74648 );
nor U110962 ( n54111, n47900, n492 );
not U110963 ( n492, n54107 );
nand U110964 ( n47986, n54186, n54187 );
nand U110965 ( n54187, n7813, n54183 );
nor U110966 ( n54186, n54188, n54189 );
nor U110967 ( n54189, n44990, n47864 );
nand U110968 ( n54110, n54142, n54143 );
nor U110969 ( n54142, n42399, n54198 );
nor U110970 ( n54143, n54144, n54145 );
nand U110971 ( n54198, n54199, n54200 );
nor U110972 ( n54167, n54170, n54171 );
nor U110973 ( n54171, n74525, n54166 );
nor U110974 ( n54170, n48514, n54172 );
nand U110975 ( n54172, n54173, n54174 );
nand U110976 ( n54174, n54175, n54176 );
nand U110977 ( n54175, n54177, n54178 );
nand U110978 ( n54177, n47986, n47926 );
nand U110979 ( n54178, n54179, n47979 );
nand U110980 ( n54163, n54164, n54165 );
nand U110981 ( n54165, n54166, n74525 );
nand U110982 ( n54164, n54167, n54168 );
or U110983 ( n54168, n54169, n73133 );
or U110984 ( n54179, n47986, n73140 );
nand U110985 ( n14836, n54099, n54100 );
nor U110986 ( n54100, n54101, n54102 );
nor U110987 ( n54099, n54108, n54109 );
nand U110988 ( n54102, n43372, n54103 );
nand U110989 ( n32566, n32582, n3232 );
nor U110990 ( n32582, n3063, n74591 );
nand U110991 ( n46270, n46286, n7618 );
nor U110992 ( n46286, n7438, n74648 );
nand U110993 ( n25324, n25340, n4059 );
nor U110994 ( n25340, n3907, n74592 );
nand U110995 ( n67331, n67347, n5830 );
nor U110996 ( n67347, n5664, n74593 );
nand U110997 ( n58463, n58479, n6692 );
nor U110998 ( n58479, n6539, n74594 );
nor U110999 ( n32282, n33232, n33188 );
and U111000 ( n33232, n74855, n33233 );
nand U111001 ( n33233, n33234, n33235 );
nor U111002 ( n12290, n13504, n13449 );
and U111003 ( n13504, n74823, n13505 );
nand U111004 ( n13505, n13507, n13508 );
nor U111005 ( n45970, n46952, n46897 );
and U111006 ( n46952, n74822, n46953 );
nand U111007 ( n46953, n46954, n46955 );
nor U111008 ( n66921, n67987, n67944 );
and U111009 ( n67987, n74852, n67988 );
nand U111010 ( n67988, n67989, n67990 );
nor U111011 ( n25045, n25984, n25941 );
and U111012 ( n25984, n74853, n25985 );
nand U111013 ( n25985, n25986, n25987 );
nor U111014 ( n58180, n59122, n59079 );
and U111015 ( n59122, n74854, n59123 );
nand U111016 ( n59123, n59124, n59125 );
buf U111017 ( n76921, n76923 );
nand U111018 ( n32340, n32344, n76784 );
and U111019 ( n32344, n3142, n32345 );
nor U111020 ( n45071, n854, n45072 );
not U111021 ( n854, n45074 );
nand U111022 ( n45072, n45073, n45011 );
nand U111023 ( n45073, n858, n45010 );
not U111024 ( n858, n45009 );
nand U111025 ( n66979, n66983, n76718 );
and U111026 ( n66983, n5743, n66984 );
nand U111027 ( n46039, n46043, n76670 );
and U111028 ( n46043, n7529, n46044 );
nand U111029 ( n25103, n25107, n76766 );
and U111030 ( n25107, n3985, n25108 );
nand U111031 ( n58241, n58245, n76699 );
and U111032 ( n58245, n6618, n58246 );
nor U111033 ( n61176, n41471, n67217 );
nor U111034 ( n41463, n41908, n834 );
nand U111035 ( n42247, n915, n73910 );
not U111036 ( n915, n42251 );
and U111037 ( n71028, n71098, n71144 );
nand U111038 ( n42257, n915, n73911 );
nand U111039 ( n47996, n54203, n54204 );
nor U111040 ( n54204, n54205, n54206 );
nor U111041 ( n54203, n54213, n54214 );
nor U111042 ( n54206, n54207, n73511 );
nand U111043 ( n34250, n35705, n35706 );
nor U111044 ( n35706, n35707, n35708 );
nor U111045 ( n35705, n35715, n35716 );
nor U111046 ( n35708, n35709, n73526 );
nand U111047 ( n27005, n28526, n28527 );
nor U111048 ( n28527, n28528, n28529 );
nor U111049 ( n28526, n28536, n28537 );
nor U111050 ( n28529, n28530, n73516 );
nand U111051 ( n69004, n70431, n70432 );
nor U111052 ( n70432, n70433, n70434 );
nor U111053 ( n70431, n70441, n70442 );
nor U111054 ( n70434, n70435, n73515 );
nand U111055 ( n60148, n61831, n61832 );
nor U111056 ( n61832, n61833, n61834 );
nor U111057 ( n61831, n61841, n61842 );
nor U111058 ( n61834, n61835, n73517 );
nand U111059 ( n54173, n54169, n73133 );
nand U111060 ( n35675, n35671, n74513 );
nand U111061 ( n28496, n28492, n74516 );
nand U111062 ( n70401, n70397, n74514 );
nand U111063 ( n61801, n61797, n74517 );
nor U111064 ( n61744, n61745, n61746 );
nand U111065 ( n61746, n6514, n54949 );
nor U111066 ( n54116, n54117, n54118 );
nand U111067 ( n54118, n7414, n42384 );
nor U111068 ( n28439, n28440, n28441 );
nand U111069 ( n28441, n3882, n21858 );
nor U111070 ( n35618, n35619, n35620 );
nand U111071 ( n35620, n3038, n29171 );
nor U111072 ( n70344, n70345, n70346 );
nand U111073 ( n70346, n5639, n62893 );
nand U111074 ( n12586, n61742, n61743 );
nor U111075 ( n61742, n61749, n61750 );
nor U111076 ( n61743, n55891, n61744 );
nor U111077 ( n61749, n61752, n73180 );
nand U111078 ( n14831, n54114, n54115 );
nor U111079 ( n54114, n54121, n54122 );
nor U111080 ( n54115, n43371, n54116 );
nor U111081 ( n54121, n54124, n74686 );
nand U111082 ( n5851, n28437, n28438 );
nor U111083 ( n28437, n28444, n28445 );
nor U111084 ( n28438, n22777, n28439 );
nor U111085 ( n28444, n28447, n73181 );
nand U111086 ( n3606, n35616, n35617 );
nor U111087 ( n35616, n35623, n35624 );
nor U111088 ( n35617, n30098, n35618 );
nor U111089 ( n35623, n35626, n73182 );
nand U111090 ( n10341, n70342, n70343 );
nor U111091 ( n70342, n70349, n70350 );
nor U111092 ( n70343, n64115, n70344 );
nor U111093 ( n70349, n70352, n73183 );
nand U111094 ( n32368, n32369, n32370 );
nand U111095 ( n32370, n76481, n32371 );
nand U111096 ( n32369, n76786, n32372 );
nand U111097 ( n67031, n67032, n67033 );
nand U111098 ( n67033, n76203, n67034 );
nand U111099 ( n67032, n76720, n67035 );
nand U111100 ( n46067, n46068, n46069 );
nand U111101 ( n46069, n76347, n46070 );
nand U111102 ( n46068, n76672, n46071 );
nand U111103 ( n25131, n25132, n25133 );
nand U111104 ( n25133, n76527, n25134 );
nand U111105 ( n25132, n76768, n25135 );
nand U111106 ( n58269, n58270, n58271 );
nand U111107 ( n58271, n76269, n58272 );
nand U111108 ( n58270, n76701, n58273 );
nand U111109 ( n12643, n12672, n4964 );
nor U111110 ( n12672, n4794, n74649 );
nor U111111 ( n41448, n41449, n617 );
or U111112 ( n17413, n17077, n73022 );
nor U111113 ( n27748, n75427, n76512 );
nor U111114 ( n27849, n73427, n76512 );
nor U111115 ( n54074, n54078, n54079 );
nand U111116 ( n54078, n73046, n73499 );
nand U111117 ( n54079, n73028, n73473 );
nand U111118 ( n27751, n76516, n796 );
nand U111119 ( n27750, n796, n31913 );
or U111120 ( n31913, n31914, n21769 );
nand U111121 ( n12363, n12368, n76737 );
and U111122 ( n12368, n4884, n12369 );
nand U111123 ( n12420, n12425, n76737 );
and U111124 ( n12425, n12427, n12428 );
nand U111125 ( n8559, n9428, n9429 );
nor U111126 ( n9429, n4767, n9430 );
nor U111127 ( n9428, n8263, n9433 );
not U111128 ( n4767, n9432 );
nor U111129 ( n61750, n422, n54967 );
nor U111130 ( n28445, n149, n21876 );
nor U111131 ( n35624, n187, n29193 );
nor U111132 ( n70350, n458, n62911 );
nor U111133 ( n54122, n492, n42402 );
nand U111134 ( n42617, n43369, n43370 );
nor U111135 ( n43370, n7412, n43371 );
nor U111136 ( n43369, n42323, n43373 );
not U111137 ( n7412, n43372 );
not U111138 ( n220, n21124 );
nand U111139 ( n21127, n21159, n21160 );
nor U111140 ( n21159, n8315, n21215 );
nor U111141 ( n21160, n21161, n21162 );
nand U111142 ( n21215, n21216, n21217 );
nor U111143 ( n21125, n21128, n74649 );
nor U111144 ( n21128, n14674, n220 );
nor U111145 ( n21184, n21186, n21187 );
nor U111146 ( n21187, n73134, n21188 );
nor U111147 ( n21186, n21189, n21190 );
and U111148 ( n21189, n73134, n21188 );
nand U111149 ( n14767, n21203, n21204 );
nand U111150 ( n21204, n5158, n21199 );
nor U111151 ( n21203, n21205, n21206 );
nor U111152 ( n21206, n11310, n14629 );
nand U111153 ( n21190, n21191, n21192 );
or U111154 ( n21191, n21195, n21194 );
nand U111155 ( n21192, n21193, n73141 );
nand U111156 ( n21193, n21194, n21195 );
nand U111157 ( n21180, n21181, n21182 );
nand U111158 ( n21182, n21183, n74538 );
nand U111159 ( n21181, n21184, n21185 );
or U111160 ( n21185, n21183, n74538 );
nand U111161 ( n8101, n21116, n21117 );
nor U111162 ( n21117, n21118, n21119 );
nor U111163 ( n21116, n21125, n21126 );
nand U111164 ( n21119, n9432, n21120 );
nor U111165 ( n49605, n50034, n76834 );
nand U111166 ( n12398, n12399, n12400 );
nand U111167 ( n12400, n76608, n12402 );
nand U111168 ( n12399, n76739, n12403 );
not U111169 ( n185, n35619 );
not U111170 ( n148, n28440 );
not U111171 ( n457, n70345 );
not U111172 ( n420, n61745 );
not U111173 ( n490, n54117 );
nor U111174 ( n35707, n73059, n35714 );
nand U111175 ( n35714, n35693, n73526 );
nor U111176 ( n28528, n73055, n28535 );
nand U111177 ( n28535, n28514, n73516 );
nor U111178 ( n70433, n73053, n70440 );
nand U111179 ( n70440, n70419, n73515 );
nor U111180 ( n61833, n73054, n61840 );
nand U111181 ( n61840, n61819, n73517 );
nor U111182 ( n54075, n54076, n54077 );
nand U111183 ( n54076, n73062, n73822 );
nand U111184 ( n54077, n73057, n73529 );
nor U111185 ( n54205, n73052, n54212 );
nand U111186 ( n54212, n54191, n73511 );
nand U111187 ( n54085, n73070, n74387 );
nand U111188 ( n54084, n73096, n74436 );
and U111189 ( n31833, n32572, n3143 );
nor U111190 ( n32581, n75258, n76781 );
nor U111191 ( n46285, n75259, n76667 );
nor U111192 ( n25339, n75260, n76763 );
nor U111193 ( n67346, n75257, n76715 );
nor U111194 ( n58478, n75261, n76696 );
and U111195 ( n24619, n25330, n3987 );
and U111196 ( n45532, n46276, n7530 );
and U111197 ( n66456, n67337, n5744 );
and U111198 ( n57751, n58469, n6619 );
nand U111199 ( n54091, n73125, n74494 );
nor U111200 ( n35601, n35605, n35606 );
nor U111201 ( n35605, n29162, n34234 );
nand U111202 ( n35606, n35607, n74591 );
nor U111203 ( n28424, n28428, n28429 );
nor U111204 ( n28428, n21849, n26989 );
nand U111205 ( n28429, n28430, n74592 );
nor U111206 ( n70329, n70333, n70334 );
nor U111207 ( n70333, n62884, n68988 );
nand U111208 ( n70334, n70335, n74593 );
nor U111209 ( n61729, n61733, n61734 );
nor U111210 ( n61733, n54940, n60132 );
nand U111211 ( n61734, n61735, n74594 );
nor U111212 ( n54101, n54105, n54106 );
nor U111213 ( n54105, n42375, n47980 );
nand U111214 ( n54106, n54107, n74648 );
and U111215 ( n61752, n61731, n61735 );
and U111216 ( n28447, n28426, n28430 );
and U111217 ( n35626, n35603, n35607 );
and U111218 ( n70352, n70331, n70335 );
and U111219 ( n54124, n54103, n54107 );
nor U111220 ( n66874, n74884, n76716 );
nor U111221 ( n45783, n74995, n76668 );
nor U111222 ( n45851, n74951, n76668 );
nor U111223 ( n45923, n74904, n76668 );
nor U111224 ( n24856, n74970, n76764 );
nor U111225 ( n24924, n74926, n76764 );
nor U111226 ( n24998, n74883, n76764 );
nor U111227 ( n57990, n74969, n76697 );
nor U111228 ( n58061, n74925, n76697 );
nor U111229 ( n58133, n74882, n76697 );
nor U111230 ( n32156, n74929, n76782 );
nor U111231 ( n66802, n74928, n76716 );
nor U111232 ( n32088, n74988, n76782 );
nor U111233 ( n66691, n74987, n76716 );
nor U111234 ( n32179, n73264, n76782 );
nor U111235 ( n32321, n73235, n76782 );
nor U111236 ( n32456, n72967, n76781 );
nor U111237 ( n66825, n73263, n76716 );
nor U111238 ( n66960, n73236, n76716 );
nor U111239 ( n67112, n72966, n76715 );
nor U111240 ( n45874, n73267, n76668 );
nor U111241 ( n46020, n73239, n76668 );
nor U111242 ( n46148, n73206, n76667 );
nor U111243 ( n24949, n73262, n76764 );
nor U111244 ( n25084, n73234, n76764 );
nor U111245 ( n25214, n73199, n76763 );
nor U111246 ( n58084, n73261, n76697 );
nor U111247 ( n58219, n73233, n76697 );
nor U111248 ( n58350, n73198, n76696 );
nor U111249 ( n32346, n74801, n76781 );
nor U111250 ( n32410, n73217, n76781 );
nor U111251 ( n45070, n45074, n45075 );
nand U111252 ( n45075, n45076, n45010 );
nor U111253 ( n66985, n74800, n76715 );
nor U111254 ( n67073, n73216, n76715 );
nor U111255 ( n46045, n74815, n76667 );
nor U111256 ( n46109, n73221, n76667 );
nor U111257 ( n25109, n74799, n76763 );
nor U111258 ( n25175, n73215, n76763 );
nor U111259 ( n58247, n74798, n76696 );
nor U111260 ( n58311, n73214, n76696 );
nor U111261 ( n45690, n73308, n76669 );
nor U111262 ( n24779, n73294, n76765 );
nor U111263 ( n57913, n73295, n76698 );
nor U111264 ( n24691, n73317, n76765 );
nor U111265 ( n57825, n73316, n76698 );
nor U111266 ( n45601, n73391, n76669 );
nor U111267 ( n32011, n73297, n76783 );
nand U111268 ( n5211, n30191, n30192 );
nand U111269 ( n30192, n3072, n30193 );
nor U111270 ( n30191, n30194, n30195 );
nor U111271 ( n30194, n30199, n30200 );
nand U111272 ( n5201, n30214, n30215 );
nand U111273 ( n30215, n3072, n30216 );
nor U111274 ( n30214, n30217, n30218 );
nor U111275 ( n30217, n30222, n30223 );
nand U111276 ( n5191, n30233, n30234 );
nand U111277 ( n30234, n3072, n30235 );
nor U111278 ( n30233, n30236, n30237 );
nor U111279 ( n30236, n30241, n30242 );
nand U111280 ( n5181, n30252, n30253 );
nand U111281 ( n30253, n3072, n30254 );
nor U111282 ( n30252, n30255, n30256 );
nor U111283 ( n30255, n30260, n30261 );
nor U111284 ( n66614, n73296, n76717 );
nor U111285 ( n21253, n73060, n21259 );
nand U111286 ( n21259, n21208, n73527 );
nor U111287 ( n45713, n73304, n76669 );
nor U111288 ( n24804, n73291, n76765 );
nor U111289 ( n57938, n73290, n76698 );
nand U111290 ( n14785, n21251, n21252 );
nor U111291 ( n21251, n21294, n21295 );
nor U111292 ( n21252, n21253, n21254 );
nor U111293 ( n21295, n5147, n12837 );
nand U111294 ( n5246, n30127, n30128 );
or U111295 ( n30128, n30129, n30123 );
nor U111296 ( n30127, n30130, n30131 );
nor U111297 ( n30130, n30135, n30136 );
nand U111298 ( n5231, n30153, n30154 );
or U111299 ( n30154, n30155, n30123 );
nor U111300 ( n30153, n30156, n30157 );
nor U111301 ( n30156, n30161, n30162 );
nand U111302 ( n5221, n30172, n30173 );
or U111303 ( n30173, n30174, n30123 );
nor U111304 ( n30172, n30175, n30176 );
nor U111305 ( n30175, n30180, n30181 );
nand U111306 ( n16436, n43493, n43494 );
nand U111307 ( n43494, n7458, n43495 );
nor U111308 ( n43493, n43496, n43497 );
nor U111309 ( n43496, n43501, n43502 );
nand U111310 ( n16426, n43512, n43513 );
nand U111311 ( n43513, n7458, n43514 );
nor U111312 ( n43512, n43515, n43516 );
nor U111313 ( n43515, n43520, n43521 );
nand U111314 ( n16416, n43531, n43532 );
nand U111315 ( n43532, n7458, n43533 );
nor U111316 ( n43531, n43534, n43535 );
nor U111317 ( n43534, n43539, n43540 );
nand U111318 ( n16406, n43563, n43564 );
nand U111319 ( n43564, n7458, n43565 );
nor U111320 ( n43563, n43566, n43567 );
nor U111321 ( n43566, n43571, n43572 );
nand U111322 ( n11946, n64257, n64258 );
nand U111323 ( n64258, n5673, n64259 );
nor U111324 ( n64257, n64260, n64261 );
nor U111325 ( n64260, n64265, n64266 );
nand U111326 ( n11936, n64276, n64277 );
nand U111327 ( n64277, n5673, n64278 );
nor U111328 ( n64276, n64279, n64280 );
nor U111329 ( n64279, n64284, n64285 );
nand U111330 ( n11926, n64295, n64296 );
nand U111331 ( n64296, n5673, n64297 );
nor U111332 ( n64295, n64298, n64299 );
nor U111333 ( n64298, n64303, n64304 );
nand U111334 ( n11916, n64314, n64315 );
nand U111335 ( n64315, n5673, n64316 );
nor U111336 ( n64314, n64317, n64318 );
nor U111337 ( n64317, n64322, n64323 );
nor U111338 ( n31903, n73318, n76783 );
nand U111339 ( n9701, n9542, n9543 );
nand U111340 ( n9543, n4814, n9544 );
nor U111341 ( n9542, n9545, n9547 );
nor U111342 ( n9545, n9552, n9553 );
nand U111343 ( n9691, n9565, n9567 );
nand U111344 ( n9567, n4814, n9568 );
nor U111345 ( n9565, n9569, n9570 );
nor U111346 ( n9569, n9575, n9577 );
nand U111347 ( n9681, n9588, n9589 );
nand U111348 ( n9589, n4814, n9590 );
nor U111349 ( n9588, n9592, n9593 );
nor U111350 ( n9592, n9598, n9599 );
nand U111351 ( n9671, n9612, n9613 );
nand U111352 ( n9613, n4814, n9614 );
nor U111353 ( n9612, n9615, n9617 );
nor U111354 ( n9615, n9622, n9623 );
nor U111355 ( n24629, n75178, n76765 );
nor U111356 ( n57761, n75177, n76698 );
nor U111357 ( n66526, n73319, n76717 );
nor U111358 ( n45542, n75328, n76669 );
nor U111359 ( n31843, n75180, n76783 );
nand U111360 ( n16471, n43396, n43397 );
or U111361 ( n43397, n43398, n43392 );
nor U111362 ( n43396, n43399, n43400 );
nor U111363 ( n43399, n43404, n43405 );
nand U111364 ( n11981, n64140, n64141 );
or U111365 ( n64141, n64142, n64136 );
nor U111366 ( n64140, n64143, n64144 );
nor U111367 ( n64143, n64148, n64149 );
nand U111368 ( n7491, n22802, n22803 );
nand U111369 ( n22803, n22804, n76756 );
nor U111370 ( n22802, n22805, n22806 );
nor U111371 ( n22805, n22810, n22811 );
nand U111372 ( n14226, n55916, n55917 );
nand U111373 ( n55917, n55918, n76689 );
nor U111374 ( n55916, n55919, n55920 );
nor U111375 ( n55919, n55924, n55925 );
nand U111376 ( n7476, n22828, n22829 );
nand U111377 ( n22829, n22830, n76756 );
nor U111378 ( n22828, n22831, n22832 );
nor U111379 ( n22831, n22836, n22837 );
nand U111380 ( n14211, n55942, n55943 );
nand U111381 ( n55943, n55944, n76689 );
nor U111382 ( n55942, n55945, n55946 );
nor U111383 ( n55945, n55950, n55951 );
nand U111384 ( n16456, n43455, n43456 );
or U111385 ( n43456, n43457, n43392 );
nor U111386 ( n43455, n43458, n43459 );
nor U111387 ( n43458, n43463, n43464 );
nand U111388 ( n16446, n43474, n43475 );
or U111389 ( n43475, n43476, n43392 );
nor U111390 ( n43474, n43477, n43478 );
nor U111391 ( n43477, n43482, n43483 );
nand U111392 ( n11966, n64166, n64167 );
or U111393 ( n64167, n64168, n64136 );
nor U111394 ( n64166, n64169, n64170 );
nor U111395 ( n64169, n64174, n64175 );
nand U111396 ( n11956, n64238, n64239 );
or U111397 ( n64239, n64240, n64136 );
nor U111398 ( n64238, n64241, n64242 );
nor U111399 ( n64241, n64246, n64247 );
nand U111400 ( n9721, n9494, n9495 );
or U111401 ( n9495, n9497, n9457 );
nor U111402 ( n9494, n9498, n9499 );
nor U111403 ( n9498, n9504, n9505 );
nand U111404 ( n7466, n22847, n22848 );
or U111405 ( n22848, n22849, n22798 );
nor U111406 ( n22847, n22850, n22851 );
nor U111407 ( n22850, n22855, n22856 );
nand U111408 ( n14201, n55964, n55965 );
or U111409 ( n55965, n55966, n55912 );
nor U111410 ( n55964, n55967, n55968 );
nor U111411 ( n55967, n55972, n55973 );
nand U111412 ( n7456, n22868, n22869 );
nand U111413 ( n22869, n76756, n22870 );
nor U111414 ( n22868, n22871, n22872 );
nor U111415 ( n22871, n22876, n22877 );
nand U111416 ( n7446, n22887, n22888 );
nand U111417 ( n22888, n76756, n22889 );
nor U111418 ( n22887, n22890, n22891 );
nor U111419 ( n22890, n22895, n22896 );
nand U111420 ( n7436, n22906, n22907 );
nand U111421 ( n22907, n76756, n22908 );
nor U111422 ( n22906, n22909, n22910 );
nor U111423 ( n22909, n22914, n22915 );
nand U111424 ( n7426, n22925, n22926 );
nand U111425 ( n22926, n76756, n22927 );
nor U111426 ( n22925, n22928, n22929 );
nor U111427 ( n22928, n22933, n22934 );
nand U111428 ( n14191, n55983, n55984 );
nand U111429 ( n55984, n76689, n55985 );
nor U111430 ( n55983, n55986, n55987 );
nor U111431 ( n55986, n55991, n55992 );
nand U111432 ( n14181, n56002, n56003 );
nand U111433 ( n56003, n76689, n56004 );
nor U111434 ( n56002, n56005, n56006 );
nor U111435 ( n56005, n56010, n56011 );
nand U111436 ( n14171, n56021, n56022 );
nand U111437 ( n56022, n76689, n56023 );
nor U111438 ( n56021, n56024, n56025 );
nor U111439 ( n56024, n56029, n56030 );
nand U111440 ( n14161, n56040, n56041 );
nand U111441 ( n56041, n76689, n56042 );
nor U111442 ( n56040, n56043, n56044 );
nor U111443 ( n56043, n56048, n56049 );
nand U111444 ( n9736, n9462, n9463 );
or U111445 ( n9463, n9464, n9457 );
nor U111446 ( n9462, n9465, n9467 );
nor U111447 ( n9465, n9472, n9473 );
nand U111448 ( n9711, n9518, n9519 );
or U111449 ( n9519, n9520, n9457 );
nor U111450 ( n9518, n9522, n9523 );
nor U111451 ( n9522, n9528, n9529 );
nor U111452 ( n32036, n73293, n76783 );
nor U111453 ( n66466, n75179, n76717 );
nor U111454 ( n66639, n73292, n76717 );
nand U111455 ( n5151, n30313, n30314 );
nand U111456 ( n30314, n3072, n30315 );
nor U111457 ( n30313, n30316, n30317 );
nor U111458 ( n30316, n30321, n30322 );
nand U111459 ( n5171, n30271, n30272 );
nand U111460 ( n30272, n3072, n30273 );
nor U111461 ( n30271, n30274, n30275 );
nor U111462 ( n30274, n30279, n30280 );
nand U111463 ( n5161, n30290, n30291 );
nand U111464 ( n30291, n3072, n30292 );
nor U111465 ( n30290, n30293, n30294 );
nor U111466 ( n30293, n30298, n30299 );
nand U111467 ( n5141, n30332, n30333 );
nand U111468 ( n30333, n3072, n30334 );
nor U111469 ( n30332, n30335, n30336 );
nor U111470 ( n30335, n30340, n30341 );
nand U111471 ( n11886, n64432, n64433 );
nand U111472 ( n64433, n5673, n64434 );
nor U111473 ( n64432, n64435, n64436 );
nor U111474 ( n64435, n64440, n64441 );
nand U111475 ( n11906, n64394, n64395 );
nand U111476 ( n64395, n5673, n64396 );
nor U111477 ( n64394, n64397, n64398 );
nor U111478 ( n64397, n64402, n64403 );
nand U111479 ( n11896, n64413, n64414 );
nand U111480 ( n64414, n5673, n64415 );
nor U111481 ( n64413, n64416, n64417 );
nor U111482 ( n64416, n64421, n64422 );
nand U111483 ( n9631, n9710, n9712 );
nand U111484 ( n9712, n4814, n9713 );
nor U111485 ( n9710, n9714, n9715 );
nor U111486 ( n9714, n9720, n9722 );
nand U111487 ( n11876, n64451, n64452 );
nand U111488 ( n64452, n5673, n64453 );
nor U111489 ( n64451, n64454, n64455 );
nor U111490 ( n64454, n64459, n64460 );
nand U111491 ( n16396, n43582, n43583 );
nand U111492 ( n43583, n7458, n43584 );
nor U111493 ( n43582, n43585, n43586 );
nor U111494 ( n43585, n43590, n43591 );
nand U111495 ( n16386, n43601, n43602 );
nand U111496 ( n43602, n7458, n43603 );
nor U111497 ( n43601, n43604, n43605 );
nor U111498 ( n43604, n43609, n43610 );
nand U111499 ( n16376, n43620, n43621 );
nand U111500 ( n43621, n7458, n43622 );
nor U111501 ( n43620, n43623, n43624 );
nor U111502 ( n43623, n43628, n43629 );
nand U111503 ( n16366, n43639, n43640 );
nand U111504 ( n43640, n7458, n43641 );
nor U111505 ( n43639, n43642, n43643 );
nor U111506 ( n43642, n43647, n43648 );
nor U111507 ( n2221, n76401, n74742 );
nor U111508 ( n2296, n76401, n74741 );
nand U111509 ( n9661, n9635, n9637 );
nand U111510 ( n9637, n4814, n9638 );
nor U111511 ( n9635, n9639, n9640 );
nor U111512 ( n9639, n9645, n9647 );
nand U111513 ( n9651, n9663, n9664 );
nand U111514 ( n9664, n4814, n9665 );
nor U111515 ( n9663, n9667, n9668 );
nor U111516 ( n9667, n9673, n9674 );
nand U111517 ( n9641, n9687, n9688 );
nand U111518 ( n9688, n4814, n9689 );
nor U111519 ( n9687, n9690, n9692 );
nor U111520 ( n9690, n9697, n9698 );
nand U111521 ( n7396, n22984, n22985 );
nand U111522 ( n22985, n76757, n22986 );
nor U111523 ( n22984, n22987, n22988 );
nor U111524 ( n22987, n22992, n22993 );
nand U111525 ( n14131, n56100, n56101 );
nand U111526 ( n56101, n76690, n56102 );
nor U111527 ( n56100, n56103, n56104 );
nor U111528 ( n56103, n56108, n56109 );
nand U111529 ( n7416, n22944, n22945 );
nand U111530 ( n22945, n76757, n22946 );
nor U111531 ( n22944, n22947, n22948 );
nor U111532 ( n22947, n22952, n22953 );
nand U111533 ( n7406, n22965, n22966 );
nand U111534 ( n22966, n76757, n22967 );
nor U111535 ( n22965, n22968, n22969 );
nor U111536 ( n22968, n22973, n22974 );
nand U111537 ( n7386, n23003, n23004 );
nand U111538 ( n23004, n76757, n23005 );
nor U111539 ( n23003, n23006, n23007 );
nor U111540 ( n23006, n23011, n23012 );
nand U111541 ( n14151, n56062, n56063 );
nand U111542 ( n56063, n76690, n56064 );
nor U111543 ( n56062, n56065, n56066 );
nor U111544 ( n56065, n56070, n56071 );
nand U111545 ( n14141, n56081, n56082 );
nand U111546 ( n56082, n76690, n56083 );
nor U111547 ( n56081, n56084, n56085 );
nor U111548 ( n56084, n56089, n56090 );
nand U111549 ( n14121, n56119, n56120 );
nand U111550 ( n56120, n76690, n56121 );
nor U111551 ( n56119, n56122, n56123 );
nor U111552 ( n56122, n56127, n56128 );
xor U111553 ( n13848, n76035, n73176 );
xor U111554 ( n12472, n13817, n13848 );
and U111555 ( n11762, n12659, n4885 );
nor U111556 ( n12670, n75262, n76734 );
nand U111557 ( n45915, n45920, n76346 );
and U111558 ( n45920, n45921, n45922 );
nand U111559 ( n3596, n35635, n35636 );
nand U111560 ( n35635, P1_P3_STATE2_REG_3_, n35619 );
nand U111561 ( n35636, n185, n3078 );
nand U111562 ( n5841, n28456, n28457 );
nand U111563 ( n28456, P1_P2_STATE2_REG_3_, n28440 );
nand U111564 ( n28457, n148, n3922 );
nand U111565 ( n10331, n70361, n70362 );
nand U111566 ( n70361, P2_P3_STATE2_REG_3_, n70345 );
nand U111567 ( n70362, n457, n5679 );
nand U111568 ( n12576, n61761, n61762 );
nand U111569 ( n61761, P2_P2_STATE2_REG_3_, n61745 );
nand U111570 ( n61762, n420, n6554 );
nor U111571 ( n21133, n21134, n21135 );
nand U111572 ( n21135, n4770, n8297 );
nand U111573 ( n14821, n54133, n54134 );
nand U111574 ( n54133, n76176, n54117 );
nand U111575 ( n54134, n490, n7464 );
nand U111576 ( n8096, n21131, n21132 );
nor U111577 ( n21131, n21138, n21139 );
nor U111578 ( n21132, n9430, n21133 );
nor U111579 ( n21138, n21141, n74685 );
nand U111580 ( n66866, n66871, n76202 );
and U111581 ( n66871, n66872, n66873 );
nand U111582 ( n24990, n24995, n76526 );
and U111583 ( n24995, n24996, n24997 );
nand U111584 ( n58125, n58130, n76268 );
and U111585 ( n58130, n58131, n58132 );
not U111586 ( n2355, n16723 );
nor U111587 ( n17681, n73422, n17129 );
nor U111588 ( n12040, n74996, n76735 );
nor U111589 ( n12130, n74952, n76735 );
nor U111590 ( n12159, n73268, n76735 );
nor U111591 ( n12339, n73240, n76735 );
nor U111592 ( n12429, n74770, n76734 );
nor U111593 ( n12505, n73207, n76734 );
nor U111594 ( n12370, n74816, n76734 );
not U111595 ( n5165, n21608 );
not U111596 ( n5140, n21606 );
nand U111597 ( n14649, n21332, n21333 );
nand U111598 ( n21333, n5137, n21334 );
nand U111599 ( n21334, n21335, n21336 );
not U111600 ( n5137, n21339 );
nor U111601 ( n11947, n73309, n76736 );
nor U111602 ( n21139, n220, n8319 );
nor U111603 ( n11975, n73305, n76736 );
nor U111604 ( n11774, n75329, n76736 );
not U111605 ( n219, n21134 );
xnor U111606 ( n12498, n13853, n13905 );
xor U111607 ( n13905, n74658, n76034 );
nor U111608 ( n13897, n13899, n76594 );
nor U111609 ( n13899, n13900, n13902 );
nand U111610 ( n13900, n13923, n13924 );
nand U111611 ( n13902, n13903, n13904 );
nand U111612 ( n34261, n35720, n35721 );
nor U111613 ( n35720, n35749, n35750 );
nor U111614 ( n35721, n35722, n35723 );
nor U111615 ( n35750, n31497, n32707 );
nand U111616 ( n27018, n28541, n28542 );
nor U111617 ( n28541, n28570, n28571 );
nor U111618 ( n28542, n28543, n28544 );
nor U111619 ( n28571, n24203, n25467 );
nand U111620 ( n69015, n70446, n70447 );
nor U111621 ( n70446, n70475, n70476 );
nor U111622 ( n70447, n70448, n70449 );
nor U111623 ( n70476, n65747, n67472 );
nand U111624 ( n60159, n61846, n61847 );
nor U111625 ( n61846, n61875, n61876 );
nor U111626 ( n61847, n61848, n61849 );
nor U111627 ( n61876, n57325, n58604 );
nand U111628 ( n48007, n54218, n54219 );
nor U111629 ( n54218, n54247, n54248 );
nor U111630 ( n54219, n54220, n54221 );
nor U111631 ( n54248, n44882, n46408 );
nand U111632 ( n13800, n12463, n76727 );
nand U111633 ( n33467, n32415, n76774 );
nand U111634 ( n47187, n46114, n76660 );
nand U111635 ( n68218, n67078, n76708 );
nand U111636 ( n26217, n25180, n76754 );
nand U111637 ( n59356, n58316, n76687 );
and U111638 ( n21141, n21120, n21124 );
nor U111639 ( n21118, n21122, n21123 );
nor U111640 ( n21122, n8285, n14759 );
nand U111641 ( n21123, n21124, n74649 );
nand U111642 ( n45012, n45013, n45014 );
nand U111643 ( n45013, n45016, n45017 );
nand U111644 ( n45014, n45015, n857 );
nand U111645 ( n45016, n45018, n45019 );
not U111646 ( n7820, n54591 );
not U111647 ( n7795, n54589 );
nand U111648 ( n47880, n54315, n54316 );
nand U111649 ( n54316, n7792, n54317 );
nand U111650 ( n54317, n54318, n54319 );
not U111651 ( n7792, n54322 );
nand U111652 ( n63041, n64113, n64114 );
nor U111653 ( n64114, n5635, n64115 );
nor U111654 ( n64113, n62811, n64117 );
not U111655 ( n5635, n64116 );
nand U111656 ( n29274, n30096, n30097 );
nor U111657 ( n30097, n3034, n30098 );
nor U111658 ( n30096, n29144, n30100 );
not U111659 ( n3034, n30099 );
nand U111660 ( n21957, n22775, n22776 );
nor U111661 ( n22776, n3878, n22777 );
nor U111662 ( n22775, n21829, n22779 );
not U111663 ( n3878, n22778 );
nand U111664 ( n55069, n55889, n55890 );
nor U111665 ( n55890, n6510, n55891 );
nor U111666 ( n55889, n54905, n55893 );
not U111667 ( n6510, n55892 );
not U111668 ( n170, n21950 );
not U111669 ( n204, n29267 );
not U111670 ( n475, n63034 );
not U111671 ( n443, n55062 );
nor U111672 ( n22754, n74663, n3875 );
nor U111673 ( n30075, n74662, n3032 );
nor U111674 ( n64092, n74660, n5633 );
nor U111675 ( n55868, n74661, n6508 );
or U111676 ( n17648, n17077, n73422 );
nand U111677 ( n12121, n63180, n63181 );
nor U111678 ( n63181, n63182, n63183 );
nor U111679 ( n63180, n63195, n63196 );
nand U111680 ( n63183, n63184, n63185 );
nand U111681 ( n12101, n63349, n63350 );
nor U111682 ( n63350, n63351, n63352 );
nor U111683 ( n63349, n63362, n63363 );
nand U111684 ( n63352, n63353, n63354 );
nand U111685 ( n5386, n29417, n29418 );
nor U111686 ( n29418, n29419, n29420 );
nor U111687 ( n29417, n29432, n29433 );
nand U111688 ( n29420, n29421, n29422 );
nand U111689 ( n5366, n29520, n29521 );
nor U111690 ( n29521, n29522, n29523 );
nor U111691 ( n29520, n29533, n29534 );
nand U111692 ( n29523, n29524, n29525 );
nand U111693 ( n7611, n22201, n22202 );
nor U111694 ( n22202, n22203, n22204 );
nor U111695 ( n22201, n22214, n22215 );
nand U111696 ( n22204, n22205, n22206 );
nand U111697 ( n7631, n22098, n22099 );
nor U111698 ( n22099, n22100, n22101 );
nor U111699 ( n22098, n22113, n22114 );
nand U111700 ( n22101, n22102, n22103 );
nand U111701 ( n14346, n55315, n55316 );
nor U111702 ( n55316, n55317, n55318 );
nor U111703 ( n55315, n55328, n55329 );
nand U111704 ( n55318, n55319, n55320 );
nand U111705 ( n14366, n55208, n55209 );
nor U111706 ( n55209, n55210, n55211 );
nor U111707 ( n55208, n55223, n55224 );
nand U111708 ( n55211, n55212, n55213 );
nand U111709 ( n12081, n63526, n63527 );
nor U111710 ( n63526, n63537, n63538 );
nor U111711 ( n63527, n63528, n63529 );
nand U111712 ( n63538, n63539, n63540 );
nand U111713 ( n5346, n29627, n29628 );
nor U111714 ( n29627, n29638, n29639 );
nor U111715 ( n29628, n29629, n29630 );
nand U111716 ( n29639, n29640, n29641 );
nand U111717 ( n7591, n22306, n22307 );
nor U111718 ( n22306, n22317, n22318 );
nor U111719 ( n22307, n22308, n22309 );
nand U111720 ( n22318, n22319, n22320 );
nand U111721 ( n14326, n55418, n55419 );
nor U111722 ( n55418, n55429, n55430 );
nor U111723 ( n55419, n55420, n55421 );
nand U111724 ( n55430, n55431, n55432 );
nand U111725 ( n12111, n63231, n63232 );
nor U111726 ( n63231, n63245, n63246 );
nor U111727 ( n63232, n63233, n63234 );
nor U111728 ( n63245, n63070, n74751 );
nand U111729 ( n5376, n29468, n29469 );
nor U111730 ( n29468, n29482, n29483 );
nor U111731 ( n29469, n29470, n29471 );
nor U111732 ( n29482, n29303, n74752 );
nand U111733 ( n7621, n22149, n22150 );
nor U111734 ( n22149, n22163, n22164 );
nor U111735 ( n22150, n22151, n22152 );
nor U111736 ( n22163, n21988, n74753 );
nand U111737 ( n14356, n55263, n55264 );
nor U111738 ( n55263, n55277, n55278 );
nor U111739 ( n55264, n55265, n55266 );
nor U111740 ( n55277, n55098, n74754 );
nand U111741 ( n12041, n63795, n63796 );
nor U111742 ( n63796, n63797, n63798 );
nor U111743 ( n63795, n63806, n63807 );
nand U111744 ( n63798, n63799, n63800 );
nand U111745 ( n5306, n29839, n29840 );
nor U111746 ( n29840, n29841, n29842 );
nor U111747 ( n29839, n29850, n29851 );
nand U111748 ( n29842, n29843, n29844 );
nand U111749 ( n7551, n22516, n22517 );
nor U111750 ( n22517, n22518, n22519 );
nor U111751 ( n22516, n22527, n22528 );
nand U111752 ( n22519, n22520, n22521 );
nand U111753 ( n14286, n55629, n55630 );
nor U111754 ( n55630, n55631, n55632 );
nor U111755 ( n55629, n55640, n55641 );
nand U111756 ( n55632, n55633, n55634 );
nand U111757 ( n12131, n63130, n63131 );
nor U111758 ( n63131, n63132, n63133 );
nor U111759 ( n63130, n63143, n63144 );
nand U111760 ( n63133, n63134, n63135 );
nand U111761 ( n5396, n29367, n29368 );
nor U111762 ( n29368, n29369, n29370 );
nor U111763 ( n29367, n29380, n29381 );
nand U111764 ( n29370, n29371, n29372 );
nand U111765 ( n7641, n22048, n22049 );
nor U111766 ( n22049, n22050, n22051 );
nor U111767 ( n22048, n22061, n22062 );
nand U111768 ( n22051, n22052, n22053 );
nand U111769 ( n14376, n55158, n55159 );
nor U111770 ( n55159, n55160, n55161 );
nor U111771 ( n55158, n55171, n55172 );
nand U111772 ( n55161, n55162, n55163 );
nand U111773 ( n12091, n63472, n63473 );
nor U111774 ( n63473, n63474, n63475 );
nor U111775 ( n63472, n63485, n63486 );
nand U111776 ( n63474, n63480, n63481 );
nand U111777 ( n12061, n63629, n63630 );
nor U111778 ( n63630, n63631, n63632 );
nor U111779 ( n63629, n63640, n63641 );
nand U111780 ( n63631, n63637, n63481 );
nand U111781 ( n5356, n29573, n29574 );
nor U111782 ( n29574, n29575, n29576 );
nor U111783 ( n29573, n29586, n29587 );
nand U111784 ( n29575, n29581, n29582 );
nand U111785 ( n5326, n29730, n29731 );
nor U111786 ( n29731, n29732, n29733 );
nor U111787 ( n29730, n29741, n29742 );
nand U111788 ( n29732, n29738, n29582 );
nand U111789 ( n7571, n22409, n22410 );
nor U111790 ( n22410, n22411, n22412 );
nor U111791 ( n22409, n22420, n22421 );
nand U111792 ( n22411, n22417, n22261 );
nand U111793 ( n7601, n22252, n22253 );
nor U111794 ( n22253, n22254, n22255 );
nor U111795 ( n22252, n22265, n22266 );
nand U111796 ( n22254, n22260, n22261 );
nand U111797 ( n14306, n55524, n55525 );
nor U111798 ( n55525, n55526, n55527 );
nor U111799 ( n55524, n55535, n55536 );
nand U111800 ( n55526, n55532, n55373 );
nand U111801 ( n14336, n55364, n55365 );
nor U111802 ( n55365, n55366, n55367 );
nor U111803 ( n55364, n55377, n55378 );
nand U111804 ( n55366, n55372, n55373 );
nand U111805 ( n12071, n63578, n63579 );
nor U111806 ( n63579, n63580, n63581 );
nor U111807 ( n63578, n63588, n63589 );
nand U111808 ( n63580, n63586, n63481 );
nand U111809 ( n12051, n63742, n63743 );
nor U111810 ( n63743, n63744, n63745 );
nor U111811 ( n63742, n63751, n63752 );
nand U111812 ( n63744, n63750, n63481 );
nand U111813 ( n12031, n63846, n63847 );
nor U111814 ( n63847, n63848, n63849 );
nor U111815 ( n63846, n63857, n63858 );
nand U111816 ( n63848, n63854, n63481 );
nand U111817 ( n12021, n63898, n63899 );
nor U111818 ( n63899, n63900, n63901 );
nor U111819 ( n63898, n63907, n63908 );
nand U111820 ( n63900, n63906, n63481 );
nand U111821 ( n5336, n29679, n29680 );
nor U111822 ( n29680, n29681, n29682 );
nor U111823 ( n29679, n29689, n29690 );
nand U111824 ( n29681, n29687, n29582 );
nand U111825 ( n5316, n29782, n29783 );
nor U111826 ( n29783, n29784, n29785 );
nor U111827 ( n29782, n29791, n29792 );
nand U111828 ( n29784, n29790, n29582 );
nand U111829 ( n5296, n29890, n29891 );
nor U111830 ( n29891, n29892, n29893 );
nor U111831 ( n29890, n29901, n29902 );
nand U111832 ( n29892, n29898, n29582 );
nand U111833 ( n5286, n29942, n29943 );
nor U111834 ( n29943, n29944, n29945 );
nor U111835 ( n29942, n29951, n29952 );
nand U111836 ( n29944, n29950, n29582 );
nand U111837 ( n7541, n22567, n22568 );
nor U111838 ( n22568, n22569, n22570 );
nor U111839 ( n22567, n22578, n22579 );
nand U111840 ( n22569, n22575, n22261 );
nand U111841 ( n7581, n22358, n22359 );
nor U111842 ( n22359, n22360, n22361 );
nor U111843 ( n22358, n22368, n22369 );
nand U111844 ( n22360, n22366, n22261 );
nand U111845 ( n7561, n22461, n22462 );
nor U111846 ( n22462, n22463, n22464 );
nor U111847 ( n22461, n22470, n22471 );
nand U111848 ( n22463, n22469, n22261 );
nand U111849 ( n7531, n22619, n22620 );
nor U111850 ( n22620, n22621, n22622 );
nor U111851 ( n22619, n22628, n22629 );
nand U111852 ( n22621, n22627, n22261 );
nand U111853 ( n14276, n55680, n55681 );
nor U111854 ( n55681, n55682, n55683 );
nor U111855 ( n55680, n55691, n55692 );
nand U111856 ( n55682, n55688, n55373 );
nand U111857 ( n14316, n55470, n55471 );
nor U111858 ( n55471, n55472, n55473 );
nor U111859 ( n55470, n55480, n55481 );
nand U111860 ( n55472, n55478, n55373 );
nand U111861 ( n14296, n55576, n55577 );
nor U111862 ( n55577, n55578, n55579 );
nor U111863 ( n55576, n55585, n55586 );
nand U111864 ( n55578, n55584, n55373 );
nand U111865 ( n14266, n55732, n55733 );
nor U111866 ( n55733, n55734, n55735 );
nor U111867 ( n55732, n55741, n55742 );
nand U111868 ( n55734, n55740, n55373 );
nor U111869 ( n21323, n21339, n21335 );
and U111870 ( n11749, n75838, n21332 );
nand U111871 ( n75838, n21323, n21607 );
nand U111872 ( n8086, n21150, n21151 );
nand U111873 ( n21150, n76186, n21134 );
nand U111874 ( n21151, n219, n4820 );
and U111875 ( n25360, n26892, n26893 );
nand U111876 ( n26893, n21830, n74592 );
nand U111877 ( n26892, n3920, n26895 );
nand U111878 ( n26895, n26896, n26897 );
and U111879 ( n58497, n60032, n60033 );
nand U111880 ( n60033, n54906, n74594 );
nand U111881 ( n60032, n6553, n60035 );
nand U111882 ( n60035, n60036, n60037 );
not U111883 ( n450, n58496 );
nor U111884 ( n22748, n22757, n73120 );
nor U111885 ( n22757, n76909, n169 );
nor U111886 ( n30069, n30078, n73119 );
nor U111887 ( n30078, n76900, n203 );
nor U111888 ( n55862, n55871, n73122 );
nor U111889 ( n55871, n76883, n442 );
nor U111890 ( n64086, n64095, n73121 );
nor U111891 ( n64095, n76874, n474 );
not U111892 ( n179, n25359 );
and U111893 ( n32600, n34137, n34138 );
nand U111894 ( n34138, n29145, n74591 );
nand U111895 ( n34137, n3077, n34140 );
nand U111896 ( n34140, n34141, n34142 );
not U111897 ( n213, n32599 );
and U111898 ( n67365, n68891, n68892 );
nand U111899 ( n68892, n62812, n74593 );
nand U111900 ( n68891, n5678, n68894 );
nand U111901 ( n68894, n68895, n68896 );
not U111902 ( n484, n67364 );
nor U111903 ( n33930, n74622, n76897 );
nor U111904 ( n26685, n74620, n76906 );
nor U111905 ( n59827, n74619, n76880 );
nor U111906 ( n68686, n74621, n76871 );
nor U111907 ( n33853, n73169, n76897 );
nor U111908 ( n26608, n72961, n76906 );
nor U111909 ( n59750, n72960, n76880 );
nor U111910 ( n68609, n73168, n76871 );
nor U111911 ( n33768, n74643, n76897 );
nor U111912 ( n26523, n74641, n76906 );
nor U111913 ( n59665, n74640, n76880 );
nor U111914 ( n33689, n73194, n76897 );
nor U111915 ( n68524, n74642, n76871 );
nor U111916 ( n26444, n74694, n76906 );
nor U111917 ( n59583, n74693, n76880 );
nor U111918 ( n68445, n73193, n76871 );
nor U111919 ( n32592, n74662, n76468 );
nor U111920 ( n67357, n74660, n76195 );
nor U111921 ( n25352, n74663, n76519 );
nor U111922 ( n58489, n74661, n76261 );
nor U111923 ( n34005, n73164, n76897 );
nor U111924 ( n26762, n72958, n76906 );
nor U111925 ( n59902, n72959, n76880 );
nor U111926 ( n26809, n26810, n76903 );
nor U111927 ( n26810, n26811, n26812 );
nand U111928 ( n26811, n26819, n26820 );
nand U111929 ( n26812, n26813, n26814 );
nor U111930 ( n59949, n59950, n76877 );
nor U111931 ( n59950, n59951, n59952 );
nand U111932 ( n59951, n59959, n59960 );
nand U111933 ( n59952, n59953, n59954 );
nor U111934 ( n34054, n34055, n76894 );
nor U111935 ( n34055, n34056, n34057 );
nand U111936 ( n34056, n34064, n34065 );
nand U111937 ( n34057, n34058, n34059 );
nor U111938 ( n68761, n73163, n76871 );
nor U111939 ( n33595, n74712, n76897 );
nor U111940 ( n26350, n74710, n76906 );
nor U111941 ( n59489, n74709, n76880 );
nor U111942 ( n68808, n68809, n76868 );
nor U111943 ( n68809, n68810, n68811 );
nand U111944 ( n68810, n68818, n68819 );
nand U111945 ( n68811, n68812, n68813 );
nor U111946 ( n68351, n74711, n76871 );
nand U111947 ( n14658, n11749, n21322 );
nand U111948 ( n21322, n21323, n21324 );
not U111949 ( n7430, n45559 );
nand U111950 ( n64068, n63064, n64069 );
nand U111951 ( n64069, n76876, n73121 );
nand U111952 ( n30051, n29297, n30052 );
nand U111953 ( n30052, n76902, n73119 );
nand U111954 ( n22728, n21982, n22729 );
nand U111955 ( n22729, n76911, n73120 );
nand U111956 ( n55844, n55092, n55845 );
nand U111957 ( n55845, n76885, n73122 );
nand U111958 ( n12001, n64062, n64063 );
nor U111959 ( n64062, n64079, n64080 );
nor U111960 ( n64063, n64064, n64065 );
nor U111961 ( n64079, n73163, n63041 );
nand U111962 ( n5266, n30045, n30046 );
nor U111963 ( n30045, n30062, n30063 );
nor U111964 ( n30046, n30047, n30048 );
nor U111965 ( n30062, n73164, n29274 );
nand U111966 ( n7511, n22722, n22723 );
nor U111967 ( n22722, n22739, n22740 );
nor U111968 ( n22723, n22724, n22725 );
nor U111969 ( n22739, n72958, n21957 );
nand U111970 ( n14246, n55838, n55839 );
nor U111971 ( n55838, n55855, n55856 );
nor U111972 ( n55839, n55840, n55841 );
nor U111973 ( n55855, n72959, n55069 );
nand U111974 ( n10423, n10424, n10425 );
nand U111975 ( n10425, n76892, n74966 );
nand U111976 ( n44262, n44263, n44264 );
nand U111977 ( n44264, n76866, n74965 );
not U111978 ( n3055, n31861 );
nand U111979 ( n31838, n31866, n31867 );
or U111980 ( n31866, n31869, n31858 );
nand U111981 ( n31867, n31860, n3055 );
nand U111982 ( n12011, n63954, n63955 );
nor U111983 ( n63954, n63968, n63969 );
nor U111984 ( n63955, n63956, n63957 );
nand U111985 ( n63969, n63970, n63971 );
nand U111986 ( n5276, n29998, n29999 );
nor U111987 ( n29998, n30012, n30013 );
nor U111988 ( n29999, n30000, n30001 );
nand U111989 ( n30013, n30014, n30015 );
nand U111990 ( n7521, n22675, n22676 );
nor U111991 ( n22675, n22689, n22690 );
nor U111992 ( n22676, n22677, n22678 );
nand U111993 ( n22690, n22691, n22692 );
nand U111994 ( n14256, n55791, n55792 );
nor U111995 ( n55791, n55805, n55806 );
nor U111996 ( n55792, n55793, n55794 );
nand U111997 ( n55806, n55807, n55808 );
not U111998 ( n5657, n66484 );
not U111999 ( n3899, n24647 );
not U112000 ( n6532, n57783 );
nand U112001 ( n24624, n24652, n24653 );
or U112002 ( n24652, n24655, n24644 );
nand U112003 ( n24653, n24646, n3899 );
nand U112004 ( n57756, n57788, n57789 );
or U112005 ( n57788, n57791, n57780 );
nand U112006 ( n57789, n57782, n6532 );
nand U112007 ( n66461, n66489, n66490 );
or U112008 ( n66489, n66492, n66481 );
nand U112009 ( n66490, n66483, n5657 );
nand U112010 ( n10584, n10585, n10587 );
nand U112011 ( n10587, n76892, n74909 );
nand U112012 ( n10189, n10190, n10192 );
nand U112013 ( n10192, n76893, n75013 );
nand U112014 ( n44405, n44406, n44407 );
nand U112015 ( n44407, n76866, n74908 );
nand U112016 ( n44075, n44076, n44077 );
nand U112017 ( n44077, n76867, n75012 );
nand U112018 ( n10021, n10022, n10023 );
nand U112019 ( n10023, n76893, n75085 );
nand U112020 ( n43937, n43938, n43939 );
nand U112021 ( n43939, n76867, n75084 );
nand U112022 ( n9823, n9824, n9825 );
nand U112023 ( n9825, n76892, n75219 );
nand U112024 ( n43740, n43741, n43742 );
nand U112025 ( n43742, n76866, n75218 );
nand U112026 ( n7656, n21962, n21963 );
nor U112027 ( n21963, n21964, n21965 );
nor U112028 ( n21962, n21977, n21978 );
nand U112029 ( n21965, n21966, n21967 );
nand U112030 ( n5411, n29277, n29278 );
nor U112031 ( n29278, n29279, n29280 );
nor U112032 ( n29277, n29292, n29293 );
nand U112033 ( n29280, n29281, n29282 );
nand U112034 ( n23214, n23256, n23257 );
nand U112035 ( n23257, n76541, n23207 );
nand U112036 ( n12146, n63044, n63045 );
nor U112037 ( n63045, n63046, n63047 );
nor U112038 ( n63044, n63059, n63060 );
nand U112039 ( n63047, n63048, n63049 );
nand U112040 ( n14391, n55072, n55073 );
nor U112041 ( n55073, n55074, n55075 );
nor U112042 ( n55072, n55087, n55088 );
nand U112043 ( n55075, n55076, n55077 );
nand U112044 ( n56335, n56380, n56381 );
nand U112045 ( n56381, n76283, n56328 );
nand U112046 ( n34153, n31823, n35807 );
nand U112047 ( n35807, n35808, n35809 );
nand U112048 ( n33311, n3103, n32313 );
nand U112049 ( n30534, n30577, n30578 );
nand U112050 ( n30578, n76484, n30532 );
nand U112051 ( n64693, n64736, n64737 );
nand U112052 ( n64737, n76217, n64691 );
nand U112053 ( n13623, n4848, n12329 );
nand U112054 ( n26908, n24607, n28628 );
nand U112055 ( n28628, n28629, n28630 );
nand U112056 ( n68907, n66415, n70533 );
nand U112057 ( n70533, n70534, n70535 );
nand U112058 ( n60048, n57739, n61933 );
nand U112059 ( n61933, n61934, n61935 );
nand U112060 ( n47037, n7490, n46012 );
nand U112061 ( n10950, n10999, n11000 );
nand U112062 ( n11000, n76892, n74787 );
nand U112063 ( n44693, n44732, n44733 );
nand U112064 ( n44733, n76866, n74786 );
nand U112065 ( n10778, n10849, n10850 );
nand U112066 ( n10850, n76892, n74843 );
nand U112067 ( n44555, n44612, n44613 );
nand U112068 ( n44613, n76866, n74842 );
nand U112069 ( n68068, n5704, n66952 );
nand U112070 ( n26065, n3947, n25076 );
nand U112071 ( n59206, n6579, n58211 );
nand U112072 ( n11278, n11289, n11290 );
nand U112073 ( n11290, n76893, n74608 );
nand U112074 ( n44964, n44973, n44974 );
nand U112075 ( n44974, n76867, n74609 );
and U112076 ( n11289, n9965, n11299 );
nand U112077 ( n11299, n76893, n73162 );
and U112078 ( n44973, n43889, n44981 );
nand U112079 ( n44981, n76867, n73161 );
nand U112080 ( n11100, n11149, n11150 );
nand U112081 ( n11150, n76892, n74739 );
nand U112082 ( n11234, n11252, n11253 );
nand U112083 ( n11253, n76893, n74682 );
nand U112084 ( n44813, n44866, n44867 );
nand U112085 ( n44867, n76866, n74738 );
nand U112086 ( n44934, n44943, n44944 );
nand U112087 ( n44944, n76867, n74681 );
nand U112088 ( n10242, n10243, n10244 );
nand U112089 ( n10244, n10188, n75013 );
or U112090 ( n10243, n75013, n10190 );
nand U112091 ( n44117, n44118, n44119 );
nand U112092 ( n44119, n44074, n75012 );
or U112093 ( n44118, n75012, n44076 );
nand U112094 ( n44444, n44445, n44446 );
nand U112095 ( n44446, n44404, n74908 );
or U112096 ( n44445, n74908, n44406 );
nand U112097 ( n10633, n10634, n10635 );
nand U112098 ( n10635, n10583, n74909 );
or U112099 ( n10634, n74909, n10585 );
and U112100 ( n45522, n75839, n54315 );
nand U112101 ( n75839, n54306, n54590 );
nor U112102 ( n54306, n54322, n54318 );
not U112103 ( n1214, n49679 );
nand U112104 ( n10064, n10065, n10067 );
nand U112105 ( n10067, n10020, n75085 );
or U112106 ( n10065, n75085, n10022 );
nand U112107 ( n43979, n43980, n43981 );
nand U112108 ( n43981, n43936, n75084 );
or U112109 ( n43980, n75084, n43938 );
nand U112110 ( n32541, n32545, n32546 );
nand U112111 ( n32545, n30038, n32146 );
nand U112112 ( n32546, n32547, n76480 );
nand U112113 ( n67197, n67201, n67202 );
nand U112114 ( n67201, n64055, n66792 );
nand U112115 ( n67202, n67203, n76202 );
nand U112116 ( n46245, n46249, n46250 );
nand U112117 ( n46249, n43309, n45841 );
nand U112118 ( n46250, n46251, n76346 );
nand U112119 ( n25299, n25303, n25304 );
nand U112120 ( n25303, n22715, n24914 );
nand U112121 ( n25304, n25305, n76526 );
nand U112122 ( n58438, n58442, n58443 );
nand U112123 ( n58442, n55831, n58051 );
nand U112124 ( n58443, n58444, n76268 );
nand U112125 ( n32341, n32342, n76480 );
and U112126 ( n32342, n3173, n32343 );
nand U112127 ( n66980, n66981, n76202 );
and U112128 ( n66981, n5772, n66982 );
nand U112129 ( n46040, n46041, n76346 );
and U112130 ( n46041, n7559, n46042 );
nand U112131 ( n25104, n25105, n76526 );
and U112132 ( n25105, n4013, n25106 );
nand U112133 ( n58242, n58243, n76268 );
and U112134 ( n58243, n6645, n58244 );
not U112135 ( n4787, n11800 );
nor U112136 ( n16763, n17076, n73022 );
nand U112137 ( n47887, n45522, n54305 );
nand U112138 ( n54305, n54306, n54307 );
nand U112139 ( n30134, n30142, n30143 );
nand U112140 ( n30143, n76023, n75171 );
nand U112141 ( n43403, n43411, n43412 );
nand U112142 ( n43412, n76007, n75175 );
nand U112143 ( n64147, n64155, n64156 );
nand U112144 ( n64156, n75991, n75172 );
nand U112145 ( n22809, n22817, n22818 );
nand U112146 ( n22818, n76028, n75173 );
nand U112147 ( n55923, n55931, n55932 );
nand U112148 ( n55932, n75999, n75174 );
and U112149 ( n32385, n32386, n32387 );
nand U112150 ( n9470, n9480, n9482 );
nand U112151 ( n9482, n76036, n75176 );
and U112152 ( n46084, n46085, n46086 );
and U112153 ( n67048, n67049, n67050 );
and U112154 ( n25148, n25149, n25150 );
and U112155 ( n58286, n58287, n58288 );
nor U112156 ( n16513, n17129, n76788 );
nor U112157 ( n38303, n75428, n76432 );
nor U112158 ( n38468, n73432, n76432 );
nor U112159 ( n63435, n63436, n63437 );
nand U112160 ( n63436, n73034, n73455 );
nand U112161 ( n63437, n73032, n73445 );
nor U112162 ( n63417, n63432, n63433 );
nand U112163 ( n63432, n63439, n63440 );
nand U112164 ( n63433, n63434, n63435 );
nor U112165 ( n63440, n63441, n63442 );
nand U112166 ( n38306, n76436, n456 );
nand U112167 ( n38305, n456, n63374 );
nand U112168 ( n63374, n3794, n3797 );
nand U112169 ( n63419, n63426, n63427 );
nor U112170 ( n63427, n63428, n63429 );
nor U112171 ( n63426, n63430, n63431 );
nand U112172 ( n63428, n73039, n73463 );
nand U112173 ( n63431, n73490, n73044 );
nand U112174 ( n12612, n12617, n12618 );
nand U112175 ( n12617, n9354, n12118 );
nand U112176 ( n12618, n12619, n76607 );
nor U112177 ( n35784, n30103, n35786 );
nand U112178 ( n35786, n2978, n29171 );
nor U112179 ( n28605, n22782, n28607 );
nand U112180 ( n28607, n3822, n21858 );
nor U112181 ( n70510, n64120, n70512 );
nand U112182 ( n70512, n5579, n62893 );
nor U112183 ( n61910, n55896, n61912 );
nand U112184 ( n61912, n6454, n54949 );
nand U112185 ( n12364, n12365, n76607 );
and U112186 ( n12365, n4910, n12367 );
nand U112187 ( n45004, n45008, n45009 );
nand U112188 ( n45008, n45010, n45011 );
nand U112189 ( n14799, n21220, n21221 );
nor U112190 ( n21220, n21241, n21242 );
nor U112191 ( n21221, n21222, n21223 );
nor U112192 ( n21242, n11169, n12837 );
nor U112193 ( n54282, n43376, n54284 );
nand U112194 ( n54284, n7343, n42384 );
nand U112195 ( n63429, n73467, n73038 );
nor U112196 ( n17633, n17076, n73422 );
nand U112197 ( n45537, n45564, n45565 );
or U112198 ( n45564, n45567, n45556 );
nand U112199 ( n45565, n45558, n7430 );
nand U112200 ( n63745, n63746, n63747 );
nand U112201 ( n63746, n63749, n76226 );
nand U112202 ( n63747, n63748, n76875 );
nor U112203 ( n63749, n6148, n63731 );
nand U112204 ( n29785, n29786, n29787 );
nand U112205 ( n29786, n29789, n76493 );
nand U112206 ( n29787, n29788, n76901 );
nor U112207 ( n29789, n3533, n29771 );
nand U112208 ( n22464, n22465, n22466 );
nand U112209 ( n22465, n22468, n76546 );
nand U112210 ( n22466, n22467, n76910 );
nor U112211 ( n22468, n4370, n22450 );
nand U112212 ( n55579, n55580, n55581 );
nand U112213 ( n55580, n55583, n76292 );
nand U112214 ( n55581, n55582, n76884 );
nor U112215 ( n55583, n7003, n55565 );
nand U112216 ( n63717, n63718, n63719 );
nand U112217 ( n63718, n63639, n74800 );
nand U112218 ( n63719, n63720, n76875 );
nor U112219 ( n63720, n6332, n63721 );
nand U112220 ( n63873, n63874, n63875 );
nand U112221 ( n63874, n63856, n74711 );
nand U112222 ( n63875, n63876, n76875 );
nor U112223 ( n63876, n6335, n63877 );
nand U112224 ( n29757, n29758, n29759 );
nand U112225 ( n29758, n29740, n74801 );
nand U112226 ( n29759, n29760, n76901 );
nor U112227 ( n29760, n3698, n29761 );
nand U112228 ( n29917, n29918, n29919 );
nand U112229 ( n29918, n29900, n74712 );
nand U112230 ( n29919, n29920, n76901 );
nor U112231 ( n29920, n3702, n29921 );
nand U112232 ( n22436, n22437, n22438 );
nand U112233 ( n22437, n22419, n74799 );
nand U112234 ( n22438, n22439, n76910 );
nor U112235 ( n22439, n4592, n22440 );
nand U112236 ( n22594, n22595, n22596 );
nand U112237 ( n22595, n22577, n74710 );
nand U112238 ( n22596, n22597, n76910 );
nor U112239 ( n22597, n4595, n22598 );
nand U112240 ( n55551, n55552, n55553 );
nand U112241 ( n55552, n55534, n74798 );
nand U112242 ( n55553, n55554, n76884 );
nor U112243 ( n55554, n7224, n55555 );
nand U112244 ( n55707, n55708, n55709 );
nand U112245 ( n55708, n55690, n74709 );
nand U112246 ( n55709, n55710, n76884 );
nor U112247 ( n55710, n7228, n55711 );
nand U112248 ( n12056, n63714, n63715 );
nor U112249 ( n63714, n63734, n63735 );
nor U112250 ( n63715, n63716, n63717 );
nand U112251 ( n63735, n63736, n63737 );
nand U112252 ( n12026, n63870, n63871 );
nor U112253 ( n63870, n63890, n63891 );
nor U112254 ( n63871, n63872, n63873 );
nand U112255 ( n63891, n63892, n63893 );
nand U112256 ( n5321, n29754, n29755 );
nor U112257 ( n29754, n29774, n29775 );
nor U112258 ( n29755, n29756, n29757 );
nand U112259 ( n29775, n29776, n29777 );
nand U112260 ( n5291, n29914, n29915 );
nor U112261 ( n29914, n29934, n29935 );
nor U112262 ( n29915, n29916, n29917 );
nand U112263 ( n29935, n29936, n29937 );
nand U112264 ( n7566, n22433, n22434 );
nor U112265 ( n22433, n22453, n22454 );
nor U112266 ( n22434, n22435, n22436 );
nand U112267 ( n22454, n22455, n22456 );
nand U112268 ( n7536, n22591, n22592 );
nor U112269 ( n22591, n22611, n22612 );
nor U112270 ( n22592, n22593, n22594 );
nand U112271 ( n22612, n22613, n22614 );
nand U112272 ( n14301, n55548, n55549 );
nor U112273 ( n55548, n55568, n55569 );
nor U112274 ( n55549, n55550, n55551 );
nand U112275 ( n55569, n55570, n55571 );
nand U112276 ( n14271, n55704, n55705 );
nor U112277 ( n55704, n55724, n55725 );
nor U112278 ( n55705, n55706, n55707 );
nand U112279 ( n55725, n55726, n55727 );
nand U112280 ( n12016, n63920, n63921 );
nor U112281 ( n63920, n63946, n63947 );
nor U112282 ( n63921, n63922, n63923 );
nand U112283 ( n63946, n63950, n63951 );
nand U112284 ( n12006, n64039, n64040 );
nor U112285 ( n64039, n64056, n64057 );
nor U112286 ( n64040, n64041, n64042 );
nand U112287 ( n64056, n64060, n64061 );
nand U112288 ( n5281, n29964, n29965 );
nor U112289 ( n29964, n29990, n29991 );
nor U112290 ( n29965, n29966, n29967 );
nand U112291 ( n29990, n29994, n29995 );
nand U112292 ( n5271, n30022, n30023 );
nor U112293 ( n30022, n30039, n30040 );
nor U112294 ( n30023, n30024, n30025 );
nand U112295 ( n30039, n30043, n30044 );
nand U112296 ( n7526, n22641, n22642 );
nor U112297 ( n22641, n22667, n22668 );
nor U112298 ( n22642, n22643, n22644 );
nand U112299 ( n22667, n22671, n22672 );
nand U112300 ( n7516, n22699, n22700 );
nor U112301 ( n22699, n22716, n22717 );
nor U112302 ( n22700, n22701, n22702 );
nand U112303 ( n22716, n22720, n22721 );
nand U112304 ( n14261, n55754, n55755 );
nor U112305 ( n55754, n55780, n55781 );
nor U112306 ( n55755, n55756, n55757 );
nand U112307 ( n55780, n55784, n55785 );
nand U112308 ( n14251, n55815, n55816 );
nor U112309 ( n55815, n55832, n55833 );
nor U112310 ( n55816, n55817, n55818 );
nand U112311 ( n55832, n55836, n55837 );
nand U112312 ( n63956, n63964, n63965 );
nand U112313 ( n63964, n63967, n76226 );
nand U112314 ( n63965, n63966, n76875 );
nor U112315 ( n63967, n6153, n63940 );
nand U112316 ( n30000, n30008, n30009 );
nand U112317 ( n30008, n30011, n76493 );
nand U112318 ( n30009, n30010, n76901 );
nor U112319 ( n30011, n3538, n29984 );
nand U112320 ( n22677, n22685, n22686 );
nand U112321 ( n22685, n22688, n76546 );
nand U112322 ( n22686, n22687, n76910 );
nor U112323 ( n22688, n4375, n22661 );
nand U112324 ( n55793, n55801, n55802 );
nand U112325 ( n55801, n55804, n76292 );
nand U112326 ( n55802, n55803, n76884 );
nor U112327 ( n55804, n7008, n55774 );
nand U112328 ( n63475, n63476, n63477 );
nand U112329 ( n63476, n63479, n76227 );
nand U112330 ( n63477, n63478, n76874 );
nor U112331 ( n63479, n6143, n63460 );
nand U112332 ( n63581, n63582, n63583 );
nand U112333 ( n63582, n63585, n76226 );
nand U112334 ( n63583, n63584, n76874 );
nor U112335 ( n63585, n6145, n63557 );
nand U112336 ( n63632, n63633, n63634 );
nand U112337 ( n63633, n63636, n76226 );
nand U112338 ( n63634, n63635, n76874 );
nor U112339 ( n63636, n6147, n63616 );
nand U112340 ( n63849, n63850, n63851 );
nand U112341 ( n63850, n63853, n76226 );
nand U112342 ( n63851, n63852, n76874 );
nor U112343 ( n63853, n6150, n63827 );
nand U112344 ( n29576, n29577, n29578 );
nand U112345 ( n29577, n29580, n76494 );
nand U112346 ( n29578, n29579, n76900 );
nor U112347 ( n29580, n3528, n29557 );
nand U112348 ( n29682, n29683, n29684 );
nand U112349 ( n29683, n29686, n76493 );
nand U112350 ( n29684, n29685, n76900 );
nor U112351 ( n29686, n3530, n29658 );
nand U112352 ( n29733, n29734, n29735 );
nand U112353 ( n29734, n29737, n76493 );
nand U112354 ( n29735, n29736, n76900 );
nor U112355 ( n29737, n3532, n29717 );
nand U112356 ( n29893, n29894, n29895 );
nand U112357 ( n29894, n29897, n76493 );
nand U112358 ( n29895, n29896, n76900 );
nor U112359 ( n29897, n3535, n29871 );
nand U112360 ( n22412, n22413, n22414 );
nand U112361 ( n22413, n22416, n76546 );
nand U112362 ( n22414, n22415, n76909 );
nor U112363 ( n22416, n4369, n22396 );
nand U112364 ( n22570, n22571, n22572 );
nand U112365 ( n22571, n22574, n76546 );
nand U112366 ( n22572, n22573, n76909 );
nor U112367 ( n22574, n4373, n22548 );
nand U112368 ( n22255, n22256, n22257 );
nand U112369 ( n22256, n22259, n76547 );
nand U112370 ( n22257, n22258, n76909 );
nor U112371 ( n22259, n4365, n22240 );
nand U112372 ( n22361, n22362, n22363 );
nand U112373 ( n22362, n22365, n76546 );
nand U112374 ( n22363, n22364, n76909 );
nor U112375 ( n22365, n4368, n22337 );
nand U112376 ( n55527, n55528, n55529 );
nand U112377 ( n55528, n55531, n76292 );
nand U112378 ( n55529, n55530, n76883 );
nor U112379 ( n55531, n7002, n55508 );
nand U112380 ( n55683, n55684, n55685 );
nand U112381 ( n55684, n55687, n76292 );
nand U112382 ( n55685, n55686, n76883 );
nor U112383 ( n55687, n7005, n55661 );
nand U112384 ( n55367, n55368, n55369 );
nand U112385 ( n55368, n55371, n76293 );
nand U112386 ( n55369, n55370, n76883 );
nor U112387 ( n55371, n6998, n55352 );
nand U112388 ( n55473, n55474, n55475 );
nand U112389 ( n55474, n55477, n76292 );
nand U112390 ( n55475, n55476, n76883 );
nor U112391 ( n55477, n7000, n55449 );
nand U112392 ( n32309, n76481, n32313 );
nand U112393 ( n63603, n63604, n63605 );
nand U112394 ( n63604, n63568, n74830 );
nand U112395 ( n63605, n63606, n76874 );
nor U112396 ( n63606, n6330, n63607 );
nand U112397 ( n29704, n29705, n29706 );
nand U112398 ( n29705, n29669, n74829 );
nand U112399 ( n29706, n29707, n76900 );
nor U112400 ( n29707, n3697, n29708 );
nand U112401 ( n22383, n22384, n22385 );
nand U112402 ( n22384, n22348, n74828 );
nand U112403 ( n22385, n22386, n76909 );
nor U112404 ( n22386, n4590, n22387 );
nand U112405 ( n55495, n55496, n55497 );
nand U112406 ( n55496, n55460, n74827 );
nand U112407 ( n55497, n55498, n76883 );
nor U112408 ( n55498, n7223, n55499 );
nand U112409 ( n12086, n63498, n63499 );
nor U112410 ( n63498, n63518, n63519 );
nor U112411 ( n63499, n63500, n63501 );
nand U112412 ( n63519, n63520, n63521 );
nand U112413 ( n12066, n63600, n63601 );
nor U112414 ( n63600, n63619, n63620 );
nor U112415 ( n63601, n63602, n63603 );
nand U112416 ( n63619, n63623, n63624 );
nand U112417 ( n5351, n29599, n29600 );
nor U112418 ( n29599, n29619, n29620 );
nor U112419 ( n29600, n29601, n29602 );
nand U112420 ( n29620, n29621, n29622 );
nand U112421 ( n5331, n29701, n29702 );
nor U112422 ( n29701, n29720, n29721 );
nor U112423 ( n29702, n29703, n29704 );
nand U112424 ( n29720, n29724, n29725 );
nand U112425 ( n7576, n22380, n22381 );
nor U112426 ( n22380, n22399, n22400 );
nor U112427 ( n22381, n22382, n22383 );
nand U112428 ( n22399, n22403, n22404 );
nand U112429 ( n7596, n22278, n22279 );
nor U112430 ( n22278, n22298, n22299 );
nor U112431 ( n22279, n22280, n22281 );
nand U112432 ( n22299, n22300, n22301 );
nand U112433 ( n14311, n55492, n55493 );
nor U112434 ( n55492, n55511, n55512 );
nor U112435 ( n55493, n55494, n55495 );
nand U112436 ( n55511, n55515, n55516 );
nand U112437 ( n14331, n55390, n55391 );
nor U112438 ( n55390, n55410, n55411 );
nor U112439 ( n55391, n55392, n55393 );
nand U112440 ( n55411, n55412, n55413 );
nand U112441 ( n66948, n76203, n66952 );
nand U112442 ( n12324, n76607, n12329 );
nand U112443 ( n46008, n76347, n46012 );
nand U112444 ( n25072, n76527, n25076 );
nand U112445 ( n58207, n76269, n58211 );
nor U112446 ( n30208, n76489, n30212 );
nand U112447 ( n30212, n3677, n73283 );
nor U112448 ( n30246, n76489, n30250 );
nand U112449 ( n30250, n3679, n73256 );
nor U112450 ( n30265, n76489, n30269 );
nand U112451 ( n30269, n3680, n73242 );
nand U112452 ( n12106, n63319, n63320 );
nor U112453 ( n63319, n63345, n63346 );
nor U112454 ( n63320, n63321, n63322 );
nor U112455 ( n63345, n63070, n75240 );
nand U112456 ( n5371, n29490, n29491 );
nor U112457 ( n29490, n29516, n29517 );
nor U112458 ( n29491, n29492, n29493 );
nor U112459 ( n29516, n29303, n75239 );
nand U112460 ( n7616, n22171, n22172 );
nor U112461 ( n22171, n22197, n22198 );
nor U112462 ( n22172, n22173, n22174 );
nor U112463 ( n22197, n21988, n75241 );
nand U112464 ( n7646, n22018, n22019 );
nor U112465 ( n22018, n22044, n22045 );
nor U112466 ( n22019, n22020, n22021 );
nor U112467 ( n22044, n21988, n75243 );
nand U112468 ( n14351, n55285, n55286 );
nor U112469 ( n55285, n55311, n55312 );
nor U112470 ( n55286, n55287, n55288 );
nor U112471 ( n55311, n55098, n75242 );
nand U112472 ( n5401, n29337, n29338 );
nor U112473 ( n29337, n29363, n29364 );
nor U112474 ( n29338, n29339, n29340 );
nor U112475 ( n29363, n29303, n75246 );
nand U112476 ( n12136, n63100, n63101 );
nor U112477 ( n63100, n63126, n63127 );
nor U112478 ( n63101, n63102, n63103 );
nor U112479 ( n63126, n63070, n75244 );
nand U112480 ( n14381, n55128, n55129 );
nor U112481 ( n55128, n55154, n55155 );
nor U112482 ( n55129, n55130, n55131 );
nor U112483 ( n55154, n55098, n75245 );
nor U112484 ( n30227, n76490, n30231 );
nand U112485 ( n30231, n3678, n73270 );
nor U112486 ( n30284, n76490, n30288 );
nand U112487 ( n30288, n3682, n73227 );
nor U112488 ( n30307, n76490, n30311 );
nand U112489 ( n30311, n3683, n73208 );
nor U112490 ( n30326, n76490, n30330 );
nand U112491 ( n30330, n3684, n73200 );
nor U112492 ( n30344, n76490, n30348 );
nand U112493 ( n30348, n3685, n73170 );
nor U112494 ( n30361, n76490, n30365 );
nand U112495 ( n30365, n3687, n73152 );
nor U112496 ( n30378, n76489, n30382 );
nand U112497 ( n30382, n3688, n73144 );
nand U112498 ( n63233, n63241, n63242 );
nand U112499 ( n63241, n63244, n76227 );
nand U112500 ( n63242, n63243, n76874 );
nor U112501 ( n63244, n6140, n63219 );
nand U112502 ( n29470, n29478, n29479 );
nand U112503 ( n29478, n29481, n76494 );
nand U112504 ( n29479, n29480, n76900 );
nor U112505 ( n29481, n3525, n29456 );
nand U112506 ( n22151, n22159, n22160 );
nand U112507 ( n22159, n22162, n76547 );
nand U112508 ( n22160, n22161, n76909 );
nor U112509 ( n22162, n4363, n22137 );
nand U112510 ( n55265, n55273, n55274 );
nand U112511 ( n55273, n55276, n76293 );
nand U112512 ( n55274, n55275, n76883 );
nor U112513 ( n55276, n6995, n55247 );
nand U112514 ( n63901, n63902, n63903 );
nand U112515 ( n63903, n63904, n76226 );
nand U112516 ( n63902, n63905, n76875 );
nor U112517 ( n63904, n6152, n63887 );
nand U112518 ( n29945, n29946, n29947 );
nand U112519 ( n29947, n29948, n76493 );
nand U112520 ( n29946, n29949, n76901 );
nor U112521 ( n29948, n3537, n29931 );
nand U112522 ( n22622, n22623, n22624 );
nand U112523 ( n22624, n22625, n76546 );
nand U112524 ( n22623, n22626, n76910 );
nor U112525 ( n22625, n4374, n22608 );
nand U112526 ( n55735, n55736, n55737 );
nand U112527 ( n55737, n55738, n76292 );
nand U112528 ( n55736, n55739, n76884 );
nor U112529 ( n55738, n7007, n55721 );
nor U112530 ( n43544, n76363, n43548 );
nand U112531 ( n43548, n8094, n73255 );
nor U112532 ( n43576, n76363, n43580 );
nand U112533 ( n43580, n8095, n73241 );
nor U112534 ( n64270, n76222, n64274 );
nand U112535 ( n64274, n6310, n73284 );
nor U112536 ( n64308, n76222, n64312 );
nand U112537 ( n64312, n6313, n73257 );
nor U112538 ( n64327, n76222, n64331 );
nand U112539 ( n64331, n6314, n73243 );
nand U112540 ( n5236, n30145, n30146 );
or U112541 ( n30146, n30147, n30123 );
nor U112542 ( n30145, n30148, n30149 );
nor U112543 ( n30149, n30142, n75171 );
nor U112544 ( n43506, n76363, n43510 );
nand U112545 ( n43510, n8092, n73282 );
nor U112546 ( n30166, n76490, n30170 );
nand U112547 ( n30170, n3674, n73311 );
nor U112548 ( n30185, n76489, n30189 );
nand U112549 ( n30189, n3675, n73299 );
nor U112550 ( n9558, n76633, n9563 );
nand U112551 ( n9563, n5437, n73287 );
nor U112552 ( n9604, n76633, n9609 );
nand U112553 ( n9609, n5439, n73260 );
nor U112554 ( n9628, n76633, n9633 );
nand U112555 ( n9633, n5440, n73246 );
nand U112556 ( n63820, n63821, n63822 );
nand U112557 ( n63822, n63823, n76226 );
nand U112558 ( n63821, n63830, n76875 );
nor U112559 ( n63823, n6149, n63824 );
nand U112560 ( n29864, n29865, n29866 );
nand U112561 ( n29866, n29867, n76493 );
nand U112562 ( n29865, n29874, n76901 );
nor U112563 ( n29867, n3534, n29868 );
nand U112564 ( n22541, n22542, n22543 );
nand U112565 ( n22543, n22544, n76546 );
nand U112566 ( n22542, n22551, n76910 );
nor U112567 ( n22544, n4372, n22545 );
nand U112568 ( n55654, n55655, n55656 );
nand U112569 ( n55656, n55657, n76292 );
nand U112570 ( n55655, n55664, n76884 );
nor U112571 ( n55657, n7004, n55658 );
nand U112572 ( n12036, n63817, n63818 );
nor U112573 ( n63817, n63836, n63837 );
nor U112574 ( n63818, n63819, n63820 );
nand U112575 ( n63836, n63840, n63841 );
nand U112576 ( n5301, n29861, n29862 );
nor U112577 ( n29861, n29880, n29881 );
nor U112578 ( n29862, n29863, n29864 );
nand U112579 ( n29880, n29884, n29885 );
nand U112580 ( n7546, n22538, n22539 );
nor U112581 ( n22538, n22557, n22558 );
nor U112582 ( n22539, n22540, n22541 );
nand U112583 ( n22557, n22561, n22562 );
nand U112584 ( n14281, n55651, n55652 );
nor U112585 ( n55651, n55670, n55671 );
nor U112586 ( n55652, n55653, n55654 );
nand U112587 ( n55670, n55674, n55675 );
nand U112588 ( n7651, n21989, n21990 );
nor U112589 ( n21989, n22014, n22015 );
nor U112590 ( n21990, n21991, n21992 );
nor U112591 ( n22014, n21988, n74910 );
nand U112592 ( n14386, n55099, n55100 );
nor U112593 ( n55099, n55124, n55125 );
nor U112594 ( n55100, n55101, n55102 );
nor U112595 ( n55124, n55098, n74911 );
nand U112596 ( n5406, n29308, n29309 );
nor U112597 ( n29308, n29333, n29334 );
nor U112598 ( n29309, n29310, n29311 );
nor U112599 ( n29333, n29303, n74912 );
nand U112600 ( n12141, n63071, n63072 );
nor U112601 ( n63071, n63096, n63097 );
nor U112602 ( n63072, n63073, n63074 );
nor U112603 ( n63096, n63070, n74913 );
nor U112604 ( n43525, n76364, n43529 );
nand U112605 ( n43529, n8093, n73269 );
nor U112606 ( n64289, n76223, n64293 );
nand U112607 ( n64293, n6312, n73271 );
nor U112608 ( n64407, n76223, n64411 );
nand U112609 ( n64411, n6315, n73228 );
nor U112610 ( n64426, n76223, n64430 );
nand U112611 ( n64430, n6317, n73209 );
nor U112612 ( n22881, n76542, n22885 );
nand U112613 ( n22885, n4570, n73285 );
nor U112614 ( n22919, n76542, n22923 );
nand U112615 ( n22923, n4573, n73258 );
nor U112616 ( n22938, n76542, n22942 );
nand U112617 ( n22942, n4574, n73244 );
nor U112618 ( n9582, n76634, n9586 );
nand U112619 ( n9586, n5438, n73274 );
nor U112620 ( n9655, n76634, n9660 );
nand U112621 ( n9660, n5442, n73231 );
nor U112622 ( n9679, n76634, n9684 );
nand U112623 ( n9684, n5443, n73213 );
nor U112624 ( n9703, n76634, n9708 );
nand U112625 ( n9708, n5444, n73205 );
nor U112626 ( n9725, n76634, n9730 );
nand U112627 ( n9730, n5445, n73175 );
nor U112628 ( n9747, n76634, n9752 );
nand U112629 ( n9752, n5447, n73157 );
nor U112630 ( n9772, n76633, n9777 );
nand U112631 ( n9777, n5448, n73143 );
nor U112632 ( n64445, n76223, n64449 );
nand U112633 ( n64449, n6318, n73201 );
nor U112634 ( n64463, n76223, n64467 );
nand U112635 ( n64467, n6319, n73172 );
nor U112636 ( n64480, n76223, n64484 );
nand U112637 ( n64484, n6320, n73154 );
nor U112638 ( n64541, n76222, n64545 );
nand U112639 ( n64545, n6322, n73146 );
nor U112640 ( n43595, n76364, n43599 );
nand U112641 ( n43599, n8097, n73226 );
nor U112642 ( n43614, n76364, n43618 );
nand U112643 ( n43618, n8098, n73212 );
nor U112644 ( n43633, n76364, n43637 );
nand U112645 ( n43637, n8099, n73204 );
nor U112646 ( n43651, n76364, n43655 );
nand U112647 ( n43655, n8100, n73174 );
nor U112648 ( n43682, n76364, n43686 );
nand U112649 ( n43686, n8102, n73156 );
nor U112650 ( n43699, n76363, n43703 );
nand U112651 ( n43703, n8103, n73142 );
nor U112652 ( n55996, n76284, n56000 );
nand U112653 ( n56000, n7203, n73286 );
nor U112654 ( n56034, n76284, n56038 );
nand U112655 ( n56038, n7205, n73259 );
nor U112656 ( n56056, n76284, n56060 );
nand U112657 ( n56060, n7207, n73245 );
nand U112658 ( n16461, n43414, n43415 );
or U112659 ( n43415, n43416, n43392 );
nor U112660 ( n43414, n43417, n43418 );
nor U112661 ( n43418, n43411, n75175 );
nand U112662 ( n11971, n64158, n64159 );
or U112663 ( n64159, n64160, n64136 );
nor U112664 ( n64158, n64161, n64162 );
nor U112665 ( n64162, n64155, n75172 );
nand U112666 ( n9726, n9484, n9485 );
or U112667 ( n9485, n9487, n9457 );
nor U112668 ( n9484, n9488, n9489 );
nor U112669 ( n9489, n9480, n75176 );
nand U112670 ( n7481, n22820, n22821 );
or U112671 ( n22821, n22822, n22798 );
nor U112672 ( n22820, n22823, n22824 );
nor U112673 ( n22824, n22817, n75173 );
nand U112674 ( n14216, n55934, n55935 );
or U112675 ( n55935, n55936, n55912 );
nor U112676 ( n55934, n55937, n55938 );
nor U112677 ( n55938, n55931, n75174 );
nor U112678 ( n43468, n76364, n43472 );
nand U112679 ( n43472, n8089, n73310 );
nor U112680 ( n43487, n76363, n43491 );
nand U112681 ( n43491, n8090, n73298 );
nor U112682 ( n64179, n76223, n64183 );
nand U112683 ( n64183, n6308, n73312 );
nor U112684 ( n64251, n76222, n64255 );
nand U112685 ( n64255, n6309, n73300 );
nor U112686 ( n22841, n76543, n22845 );
nand U112687 ( n22845, n4568, n73313 );
nor U112688 ( n22860, n76543, n22864 );
nand U112689 ( n22864, n4569, n73301 );
nor U112690 ( n55958, n76285, n55962 );
nand U112691 ( n55962, n7200, n73314 );
nor U112692 ( n22900, n76543, n22904 );
nand U112693 ( n22904, n4572, n73272 );
nor U112694 ( n22957, n76543, n22961 );
nand U112695 ( n22961, n4575, n73229 );
nor U112696 ( n22978, n76543, n22982 );
nand U112697 ( n22982, n4577, n73210 );
nor U112698 ( n22997, n76543, n23001 );
nand U112699 ( n23001, n4578, n73202 );
nor U112700 ( n23015, n76542, n23019 );
nand U112701 ( n23019, n4579, n73171 );
nor U112702 ( n23032, n76543, n23036 );
nand U112703 ( n23036, n4580, n73153 );
nor U112704 ( n23049, n76542, n23053 );
nand U112705 ( n23053, n4582, n73145 );
nor U112706 ( n55977, n76285, n55981 );
nand U112707 ( n55981, n7202, n73302 );
nor U112708 ( n9510, n76634, n9515 );
nand U112709 ( n9515, n5434, n73315 );
nor U112710 ( n9534, n76633, n9539 );
nand U112711 ( n9539, n5435, n73303 );
nor U112712 ( n56015, n76285, n56019 );
nand U112713 ( n56019, n7204, n73273 );
nor U112714 ( n56075, n76285, n56079 );
nand U112715 ( n56079, n7208, n73230 );
nor U112716 ( n56094, n76285, n56098 );
nand U112717 ( n56098, n7209, n73211 );
nor U112718 ( n56131, n76285, n56135 );
nand U112719 ( n56135, n7212, n73173 );
nor U112720 ( n56151, n76284, n56155 );
nand U112721 ( n56155, n7213, n73155 );
nor U112722 ( n56172, n76285, n56176 );
nand U112723 ( n56176, n7214, n73147 );
nor U112724 ( n56113, n76284, n56117 );
nand U112725 ( n56117, n7210, n73203 );
nand U112726 ( n63550, n63551, n63552 );
nand U112727 ( n63552, n63553, n76226 );
nand U112728 ( n63551, n63560, n76874 );
nor U112729 ( n63553, n6144, n63554 );
nand U112730 ( n63768, n63769, n63770 );
nand U112731 ( n63770, n63771, n76226 );
nand U112732 ( n63769, n63778, n76874 );
nor U112733 ( n63771, n6148, n63772 );
nand U112734 ( n29651, n29652, n29653 );
nand U112735 ( n29653, n29654, n76493 );
nand U112736 ( n29652, n29661, n76900 );
nor U112737 ( n29654, n3529, n29655 );
nand U112738 ( n29808, n29809, n29810 );
nand U112739 ( n29810, n29811, n76493 );
nand U112740 ( n29809, n29818, n76900 );
nor U112741 ( n29811, n3533, n29812 );
nand U112742 ( n22489, n22490, n22491 );
nand U112743 ( n22491, n22492, n76546 );
nand U112744 ( n22490, n22499, n76909 );
nor U112745 ( n22492, n4370, n22493 );
nand U112746 ( n22330, n22331, n22332 );
nand U112747 ( n22332, n22333, n76546 );
nand U112748 ( n22331, n22340, n76909 );
nor U112749 ( n22333, n4367, n22334 );
nand U112750 ( n55602, n55603, n55604 );
nand U112751 ( n55604, n55605, n76292 );
nand U112752 ( n55603, n55612, n76883 );
nor U112753 ( n55605, n7003, n55606 );
nand U112754 ( n55442, n55443, n55444 );
nand U112755 ( n55444, n55445, n76292 );
nand U112756 ( n55443, n55452, n76883 );
nor U112757 ( n55445, n6999, n55446 );
nand U112758 ( n12076, n63547, n63548 );
nor U112759 ( n63547, n63569, n63570 );
nor U112760 ( n63548, n63549, n63550 );
nand U112761 ( n63570, n63571, n63572 );
nand U112762 ( n12046, n63765, n63766 );
nor U112763 ( n63765, n63786, n63787 );
nor U112764 ( n63766, n63767, n63768 );
nand U112765 ( n63787, n63788, n63789 );
nand U112766 ( n5341, n29648, n29649 );
nor U112767 ( n29648, n29670, n29671 );
nor U112768 ( n29649, n29650, n29651 );
nand U112769 ( n29671, n29672, n29673 );
nand U112770 ( n5311, n29805, n29806 );
nor U112771 ( n29805, n29826, n29827 );
nor U112772 ( n29806, n29807, n29808 );
nand U112773 ( n29827, n29828, n29829 );
nand U112774 ( n7556, n22486, n22487 );
nor U112775 ( n22486, n22507, n22508 );
nor U112776 ( n22487, n22488, n22489 );
nand U112777 ( n22508, n22509, n22510 );
nand U112778 ( n7586, n22327, n22328 );
nor U112779 ( n22327, n22349, n22350 );
nor U112780 ( n22328, n22329, n22330 );
nand U112781 ( n22350, n22351, n22352 );
nand U112782 ( n14291, n55599, n55600 );
nor U112783 ( n55599, n55620, n55621 );
nor U112784 ( n55600, n55601, n55602 );
nand U112785 ( n55621, n55622, n55623 );
nand U112786 ( n14321, n55439, n55440 );
nor U112787 ( n55439, n55461, n55462 );
nor U112788 ( n55440, n55441, n55442 );
nand U112789 ( n55462, n55463, n55464 );
nand U112790 ( n63153, n63162, n63163 );
nand U112791 ( n63163, n63164, n76227 );
nand U112792 ( n63162, n63171, n76874 );
nor U112793 ( n63164, n6138, n63165 );
nand U112794 ( n29390, n29399, n29400 );
nand U112795 ( n29400, n29401, n76494 );
nand U112796 ( n29399, n29408, n76900 );
nor U112797 ( n29401, n3523, n29402 );
nand U112798 ( n22071, n22080, n22081 );
nand U112799 ( n22081, n22082, n76547 );
nand U112800 ( n22080, n22089, n76909 );
nor U112801 ( n22082, n4360, n22083 );
nand U112802 ( n55181, n55190, n55191 );
nand U112803 ( n55191, n55192, n76293 );
nand U112804 ( n55190, n55199, n76883 );
nor U112805 ( n55192, n6993, n55193 );
nand U112806 ( n12116, n63204, n63205 );
nor U112807 ( n63204, n63227, n63228 );
nor U112808 ( n63205, n63206, n63207 );
nor U112809 ( n63227, n63070, n75210 );
nand U112810 ( n5381, n29441, n29442 );
nor U112811 ( n29441, n29464, n29465 );
nor U112812 ( n29442, n29443, n29444 );
nor U112813 ( n29464, n29303, n75209 );
nand U112814 ( n7626, n22122, n22123 );
nor U112815 ( n22122, n22145, n22146 );
nor U112816 ( n22123, n22124, n22125 );
nor U112817 ( n22145, n21988, n75211 );
nand U112818 ( n14361, n55232, n55233 );
nor U112819 ( n55232, n55255, n55256 );
nor U112820 ( n55233, n55234, n55235 );
nor U112821 ( n55255, n55098, n75212 );
nand U112822 ( n63206, n63213, n63214 );
nand U112823 ( n63214, n63215, n76227 );
nand U112824 ( n63213, n63222, n76874 );
nor U112825 ( n63215, n6139, n63216 );
nand U112826 ( n63446, n63454, n63455 );
nand U112827 ( n63455, n63456, n76227 );
nand U112828 ( n63454, n63463, n76874 );
nor U112829 ( n63456, n6142, n63457 );
nand U112830 ( n29443, n29450, n29451 );
nand U112831 ( n29451, n29452, n76494 );
nand U112832 ( n29450, n29459, n76900 );
nor U112833 ( n29452, n3524, n29453 );
nand U112834 ( n29543, n29551, n29552 );
nand U112835 ( n29552, n29553, n76494 );
nand U112836 ( n29551, n29560, n76900 );
nor U112837 ( n29553, n3527, n29554 );
nand U112838 ( n22226, n22234, n22235 );
nand U112839 ( n22235, n22236, n76547 );
nand U112840 ( n22234, n22243, n76909 );
nor U112841 ( n22236, n4364, n22237 );
nand U112842 ( n22124, n22131, n22132 );
nand U112843 ( n22132, n22133, n76547 );
nand U112844 ( n22131, n22140, n76909 );
nor U112845 ( n22133, n4362, n22134 );
nand U112846 ( n55338, n55346, n55347 );
nand U112847 ( n55347, n55348, n76293 );
nand U112848 ( n55346, n55355, n76883 );
nor U112849 ( n55348, n6997, n55349 );
nand U112850 ( n55234, n55241, n55242 );
nand U112851 ( n55242, n55243, n76293 );
nand U112852 ( n55241, n55250, n76883 );
nor U112853 ( n55243, n6994, n55244 );
nand U112854 ( n12126, n63151, n63152 );
nor U112855 ( n63151, n63176, n63177 );
nor U112856 ( n63152, n63153, n63154 );
nor U112857 ( n63176, n63070, n75045 );
nand U112858 ( n12096, n63444, n63445 );
nor U112859 ( n63444, n63468, n63469 );
nor U112860 ( n63445, n63446, n63447 );
nor U112861 ( n63468, n63070, n74940 );
nand U112862 ( n5391, n29388, n29389 );
nor U112863 ( n29388, n29413, n29414 );
nor U112864 ( n29389, n29390, n29391 );
nor U112865 ( n29413, n29303, n75044 );
nand U112866 ( n5361, n29541, n29542 );
nor U112867 ( n29541, n29565, n29566 );
nor U112868 ( n29542, n29543, n29544 );
nor U112869 ( n29565, n29303, n74941 );
nand U112870 ( n7636, n22069, n22070 );
nor U112871 ( n22069, n22094, n22095 );
nor U112872 ( n22070, n22071, n22072 );
nor U112873 ( n22094, n21988, n75043 );
nand U112874 ( n7606, n22224, n22225 );
nor U112875 ( n22224, n22248, n22249 );
nor U112876 ( n22225, n22226, n22227 );
nor U112877 ( n22248, n21988, n74942 );
nand U112878 ( n14371, n55179, n55180 );
nor U112879 ( n55179, n55204, n55205 );
nor U112880 ( n55180, n55181, n55182 );
nor U112881 ( n55204, n55098, n75046 );
nand U112882 ( n14341, n55336, n55337 );
nor U112883 ( n55336, n55360, n55361 );
nor U112884 ( n55337, n55338, n55339 );
nor U112885 ( n55360, n55098, n74943 );
nor U112886 ( n10470, n10424, n74966 );
nor U112887 ( n44300, n44263, n74965 );
nor U112888 ( n37094, n38601, n37303 );
nand U112889 ( n63430, n73477, n73041 );
nor U112890 ( n66951, n66989, n74463 );
nor U112891 ( n32312, n32350, n74465 );
nor U112892 ( n25075, n25113, n74466 );
nor U112893 ( n58210, n58251, n74464 );
nor U112894 ( n66831, n74563, n66845 );
nor U112895 ( n32185, n74564, n32199 );
nor U112896 ( n24955, n74565, n24969 );
nor U112897 ( n58090, n74566, n58104 );
nor U112898 ( n66914, n66916, n6177 );
nor U112899 ( n32275, n32277, n3562 );
nor U112900 ( n25038, n25040, n4399 );
nor U112901 ( n58173, n58175, n7032 );
nor U112902 ( n66785, n66784, n6175 );
nor U112903 ( n32139, n32138, n3560 );
nor U112904 ( n24907, n24906, n4398 );
nor U112905 ( n58044, n58043, n7030 );
nor U112906 ( n24860, n24849, n74689 );
nor U112907 ( n32092, n32081, n74688 );
nor U112908 ( n66695, n66684, n74687 );
nor U112909 ( n57994, n57983, n74690 );
nor U112910 ( n67022, n67057, n73110 );
nor U112911 ( n32359, n32394, n73112 );
nor U112912 ( n25122, n25157, n73113 );
nor U112913 ( n58260, n58295, n73111 );
nor U112914 ( n67064, n67099, n73100 );
nor U112915 ( n32401, n32443, n73102 );
nor U112916 ( n25166, n25201, n73103 );
nor U112917 ( n58302, n58337, n73101 );
nor U112918 ( n67158, n67166, n73080 );
nor U112919 ( n32502, n32510, n73082 );
nor U112920 ( n25260, n25268, n73083 );
nor U112921 ( n58396, n58404, n73081 );
nor U112922 ( n24739, n24783, n74806 );
nor U112923 ( n31971, n32015, n74804 );
nor U112924 ( n66574, n66618, n74805 );
nor U112925 ( n57873, n57917, n74807 );
nor U112926 ( n24696, n24729, n74850 );
nor U112927 ( n31908, n31961, n74849 );
nor U112928 ( n66531, n66564, n74848 );
nor U112929 ( n57830, n57863, n74851 );
nor U112930 ( n67118, n67138, n73091 );
nor U112931 ( n32462, n32482, n73093 );
nor U112932 ( n25220, n25240, n73094 );
nor U112933 ( n58356, n58376, n73092 );
nor U112934 ( n24808, n24818, n74753 );
nor U112935 ( n32040, n32050, n74752 );
nor U112936 ( n66643, n66653, n74751 );
nor U112937 ( n57942, n57952, n74754 );
nor U112938 ( n24618, n24648, n74910 );
nor U112939 ( n31832, n31862, n74912 );
nor U112940 ( n66455, n66485, n74913 );
nor U112941 ( n57750, n57784, n74911 );
or U112942 ( n66845, n66847, n66878 );
or U112943 ( n32199, n32201, n32240 );
or U112944 ( n24969, n24971, n25002 );
or U112945 ( n58104, n58106, n58137 );
nand U112946 ( n11768, n11807, n11808 );
or U112947 ( n11807, n11810, n11797 );
nand U112948 ( n11808, n11799, n4787 );
nand U112949 ( n48033, n76326, n45392 );
nand U112950 ( n42495, n43357, n43358 );
nor U112951 ( n43358, n503, n43350 );
nor U112952 ( n43357, n43347, n74992 );
nor U112953 ( n21299, n9437, n21301 );
nand U112954 ( n21301, n4711, n8297 );
nor U112955 ( n45190, n905, n42344 );
not U112956 ( n905, n42302 );
nand U112957 ( n30390, n3075, n30401 );
nand U112958 ( n30401, n76023, n73119 );
nand U112959 ( n23063, n3919, n23070 );
nand U112960 ( n23070, n76028, n73120 );
nand U112961 ( n9787, n4818, n9795 );
nand U112962 ( n9795, n76036, n73126 );
nand U112963 ( n64553, n5677, n64560 );
nand U112964 ( n64560, n75991, n73121 );
nand U112965 ( n56184, n6552, n56191 );
nand U112966 ( n56191, n75999, n73122 );
nand U112967 ( n43711, n7462, n43718 );
nand U112968 ( n43718, n76007, n73123 );
nand U112969 ( n11747, n11749, n8297 );
nand U112970 ( n30373, n3075, n30380 );
nand U112971 ( n30380, n76024, n30381 );
nand U112972 ( n64536, n5677, n64543 );
nand U112973 ( n64543, n75992, n64544 );
nand U112974 ( n23044, n3919, n23051 );
nand U112975 ( n23051, n76029, n23052 );
nand U112976 ( n9762, n4818, n9774 );
nand U112977 ( n9774, n76037, n9775 );
nand U112978 ( n56163, n6552, n56174 );
nand U112979 ( n56174, n76000, n56175 );
nand U112980 ( n43694, n7462, n43701 );
nand U112981 ( n43701, n76008, n43702 );
nor U112982 ( n45255, n904, n42344 );
not U112983 ( n904, n42309 );
nand U112984 ( n71097, n71329, n71330 );
nor U112985 ( n71329, n71333, n71334 );
nor U112986 ( n71330, n71331, n71332 );
nor U112987 ( n71334, n74489, n73026 );
nand U112988 ( n71095, n71096, n71097 );
nor U112989 ( n71331, n73124, n71105 );
nand U112990 ( n24605, n24607, n21858 );
nand U112991 ( n57737, n57739, n54949 );
nor U112992 ( n24600, n74780, n76529 );
nor U112993 ( n57732, n74779, n76271 );
nand U112994 ( n66413, n66415, n62893 );
nor U112995 ( n66407, n74776, n76205 );
nand U112996 ( n8408, n9413, n9414 );
nor U112997 ( n9414, n232, n9404 );
nor U112998 ( n9413, n9400, n74985 );
nand U112999 ( n9372, n76890, n73126 );
nor U113000 ( n22765, n22770, n75222 );
nor U113001 ( n22770, n76546, n22771 );
nand U113002 ( n22771, n21970, n21988 );
nor U113003 ( n55879, n55884, n75224 );
nor U113004 ( n55884, n76292, n55885 );
nand U113005 ( n55885, n55080, n55098 );
nor U113006 ( n30086, n30091, n75221 );
nor U113007 ( n30091, n76493, n30092 );
nand U113008 ( n30092, n29285, n29303 );
nor U113009 ( n64103, n64108, n75223 );
nor U113010 ( n64108, n76226, n64109 );
nand U113011 ( n64109, n63052, n63070 );
nand U113012 ( n8429, n76890, n8410 );
buf U113013 ( n76548, n21935 );
buf U113014 ( n76495, n29252 );
buf U113015 ( n76228, n63019 );
buf U113016 ( n76294, n55047 );
nor U113017 ( n43341, n43351, n73123 );
nor U113018 ( n43351, n76862, n500 );
xnor U113019 ( n46134, n47193, n47238 );
xor U113020 ( n47238, n73178, n47194 );
xnor U113021 ( n12488, n13805, n13854 );
xor U113022 ( n13854, n73176, n13807 );
xnor U113023 ( n67098, n68224, n68269 );
xor U113024 ( n68269, n73187, n68225 );
xnor U113025 ( n25200, n26223, n26268 );
xor U113026 ( n26268, n73188, n26224 );
xnor U113027 ( n58336, n59362, n59407 );
xor U113028 ( n59407, n73189, n59363 );
nand U113029 ( n71099, n71100, n71101 );
nor U113030 ( n71100, n71106, n71107 );
nor U113031 ( n71101, n71102, n71103 );
nor U113032 ( n71107, n74496, n73026 );
xnor U113033 ( n32442, n33473, n33514 );
xor U113034 ( n33514, n73197, n33474 );
nand U113035 ( n45520, n45522, n42384 );
nor U113036 ( n71102, n74493, n71105 );
nand U113037 ( n42303, n903, n74217 );
not U113038 ( n903, n42299 );
nor U113039 ( n63645, n63740, n63741 );
nor U113040 ( n63862, n63896, n63897 );
nor U113041 ( n29746, n29780, n29781 );
nor U113042 ( n29906, n29940, n29941 );
nor U113043 ( n22425, n22459, n22460 );
nor U113044 ( n22583, n22617, n22618 );
nor U113045 ( n55540, n55574, n55575 );
nor U113046 ( n55696, n55730, n55731 );
nor U113047 ( n63932, n63976, n63977 );
nor U113048 ( n29976, n30020, n30021 );
nor U113049 ( n55766, n55813, n55814 );
nor U113050 ( n22653, n22697, n22698 );
nand U113051 ( n42308, n903, n74219 );
nand U113052 ( n43323, n76864, n73123 );
nand U113053 ( n64071, n76228, n75223 );
nand U113054 ( n30054, n76495, n75221 );
nand U113055 ( n22731, n76548, n75222 );
nand U113056 ( n55847, n76294, n75224 );
nand U113057 ( n8438, n9427, n9425 );
nor U113058 ( n9427, n4762, n74685 );
nor U113059 ( n9415, n9422, n75226 );
nor U113060 ( n9422, n4759, n9423 );
nand U113061 ( n9423, n8480, n8414 );
nand U113062 ( n32384, n73115, n33459 );
or U113063 ( n33459, n33458, n73114 );
nand U113064 ( n9751, n9390, n9392 );
nor U113065 ( n9392, n9393, n9394 );
nor U113066 ( n9390, n9415, n9417 );
nor U113067 ( n9394, n9395, n75262 );
nand U113068 ( n42512, n43368, n43367 );
nor U113069 ( n43368, n7407, n74686 );
nor U113070 ( n43359, n43364, n75225 );
nor U113071 ( n43364, n7404, n43365 );
nand U113072 ( n43365, n43338, n42500 );
nor U113073 ( n9393, n9405, n73126 );
nor U113074 ( n9405, n76889, n229 );
nor U113075 ( n10897, n10849, n74843 );
nor U113076 ( n11047, n10999, n74787 );
nor U113077 ( n44650, n44612, n74842 );
nor U113078 ( n44770, n44732, n74786 );
nand U113079 ( n12424, n74735, n13789 );
or U113080 ( n13789, n13788, n73109 );
nand U113081 ( n46083, n74734, n47179 );
or U113082 ( n47179, n47178, n73078 );
nor U113083 ( n11298, n11289, n74608 );
nor U113084 ( n44980, n44973, n74609 );
nand U113085 ( n23640, n23256, n23682 );
nand U113086 ( n23682, n76541, n23595 );
nand U113087 ( n23551, n23256, n23593 );
nand U113088 ( n23593, n76541, n23451 );
nand U113089 ( n23729, n23256, n23771 );
nand U113090 ( n23771, n76541, n23684 );
nand U113091 ( n56673, n56380, n56715 );
nand U113092 ( n56715, n76283, n56573 );
nand U113093 ( n56762, n56380, n56804 );
nand U113094 ( n56804, n76283, n56717 );
nand U113095 ( n56851, n56380, n56896 );
nand U113096 ( n56896, n76283, n56806 );
nand U113097 ( n67047, n74758, n68210 );
or U113098 ( n68210, n68209, n73084 );
nand U113099 ( n25147, n74759, n26209 );
or U113100 ( n26209, n26208, n73085 );
nand U113101 ( n58285, n74760, n59348 );
or U113102 ( n59348, n59347, n73086 );
nor U113103 ( n11218, n11149, n74739 );
nor U113104 ( n44921, n44866, n74738 );
nor U113105 ( n44951, n44943, n74681 );
nor U113106 ( n11262, n11252, n74682 );
nand U113107 ( n31030, n30577, n31070 );
nand U113108 ( n31070, n76484, n30987 );
nand U113109 ( n65062, n64736, n65102 );
nand U113110 ( n65102, n76217, n64964 );
nand U113111 ( n65147, n64736, n65187 );
nand U113112 ( n65187, n76217, n65104 );
nand U113113 ( n65232, n64736, n65272 );
nand U113114 ( n65272, n76217, n65189 );
nand U113115 ( n31841, n31861, n31869 );
nand U113116 ( n30945, n30577, n30985 );
nand U113117 ( n30985, n76484, n30902 );
nand U113118 ( n30860, n30577, n30900 );
nand U113119 ( n30900, n76484, n30762 );
nand U113120 ( n24627, n24647, n24655 );
nand U113121 ( n66464, n66484, n66492 );
nand U113122 ( n57759, n57783, n57791 );
nand U113123 ( n23404, n23256, n23449 );
nand U113124 ( n23449, n76540, n23354 );
nand U113125 ( n23307, n23256, n23352 );
nand U113126 ( n23352, n76540, n23259 );
nand U113127 ( n56431, n56380, n56476 );
nand U113128 ( n56476, n76282, n56383 );
nand U113129 ( n56526, n56380, n56571 );
nand U113130 ( n56571, n76282, n56478 );
nand U113131 ( n45540, n45559, n45567 );
nand U113132 ( n24727, n24627, n74850 );
nand U113133 ( n31959, n31841, n74849 );
nand U113134 ( n66562, n66464, n74848 );
nand U113135 ( n57861, n57759, n74851 );
nand U113136 ( n63922, n63934, n63935 );
nand U113137 ( n63935, n63936, n76226 );
nor U113138 ( n63934, n5634, n63943 );
nor U113139 ( n63936, n6152, n63937 );
nand U113140 ( n29966, n29978, n29979 );
nand U113141 ( n29979, n29980, n76493 );
nor U113142 ( n29978, n3033, n29987 );
nor U113143 ( n29980, n3537, n29981 );
nand U113144 ( n22643, n22655, n22656 );
nand U113145 ( n22656, n22657, n76546 );
nor U113146 ( n22655, n3877, n22664 );
nor U113147 ( n22657, n4374, n22658 );
nand U113148 ( n55756, n55768, n55769 );
nand U113149 ( n55769, n55770, n76292 );
nor U113150 ( n55768, n6509, n55777 );
nor U113151 ( n55770, n7007, n55771 );
nand U113152 ( n32027, n31841, n75209 );
nand U113153 ( n45705, n45540, n74740 );
nand U113154 ( n64831, n64736, n64873 );
nand U113155 ( n64873, n76216, n64739 );
nand U113156 ( n64920, n64736, n64962 );
nand U113157 ( n64962, n76216, n64875 );
nand U113158 ( n66630, n66464, n75210 );
nand U113159 ( n24795, n24627, n75211 );
nand U113160 ( n57929, n57759, n75212 );
nand U113161 ( n45638, n45540, n75208 );
nor U113162 ( n63793, n63810, n63811 );
nor U113163 ( n29833, n29854, n29855 );
nor U113164 ( n22514, n22531, n22532 );
nor U113165 ( n55627, n55644, n55645 );
nand U113166 ( n30625, n30577, n30667 );
nand U113167 ( n30667, n76483, n30580 );
nand U113168 ( n30714, n30577, n30760 );
nand U113169 ( n30760, n76483, n30669 );
nor U113170 ( n71333, n73125, n71108 );
nand U113171 ( n43874, n43666, n43668 );
nand U113172 ( n43871, n43872, n43873 );
nand U113173 ( n43873, n43874, n74397 );
nor U113174 ( n43867, n43868, n43869 );
nor U113175 ( n43868, n867, n43875 );
nor U113176 ( n43869, n43870, n43871 );
not U113177 ( n867, n43870 );
nand U113178 ( n43872, n870, n864 );
not U113179 ( n870, n43668 );
nand U113180 ( n65650, n64736, n65689 );
nand U113181 ( n65689, n76217, n65611 );
nand U113182 ( n57228, n56380, n57267 );
nand U113183 ( n57267, n76283, n57189 );
nand U113184 ( n24106, n23256, n24145 );
nand U113185 ( n24145, n76541, n24067 );
nand U113186 ( n31400, n30577, n31439 );
nand U113187 ( n31439, n76484, n31361 );
nand U113188 ( n65569, n64736, n65608 );
nand U113189 ( n65608, n76217, n65530 );
nand U113190 ( n31319, n30577, n31358 );
nand U113191 ( n31358, n76484, n31280 );
nand U113192 ( n24025, n23256, n24064 );
nand U113193 ( n24064, n76541, n23986 );
nand U113194 ( n57147, n56380, n57186 );
nand U113195 ( n57186, n76283, n57108 );
nand U113196 ( n31570, n30577, n31583 );
nand U113197 ( n31583, n76484, n31561 );
nand U113198 ( n65488, n64736, n65527 );
nand U113199 ( n65527, n76217, n65432 );
nand U113200 ( n65731, n64736, n65787 );
nand U113201 ( n65787, n76217, n65692 );
nand U113202 ( n65839, n64736, n65848 );
nand U113203 ( n65848, n76217, n65790 );
nand U113204 ( n65860, n64736, n65869 );
nand U113205 ( n65869, n76217, n65851 );
nand U113206 ( n31234, n30577, n31277 );
nand U113207 ( n31277, n76484, n31178 );
nand U113208 ( n57066, n56380, n57105 );
nand U113209 ( n57105, n76283, n57059 );
nand U113210 ( n57309, n56380, n57368 );
nand U113211 ( n57368, n76283, n57270 );
nand U113212 ( n57380, n56380, n57389 );
nand U113213 ( n57389, n76283, n57371 );
nand U113214 ( n57401, n56380, n57410 );
nand U113215 ( n57410, n76283, n57392 );
nand U113216 ( n24187, n23256, n24243 );
nand U113217 ( n24243, n76541, n24148 );
nand U113218 ( n24255, n23256, n24264 );
nand U113219 ( n24264, n76541, n24246 );
nand U113220 ( n24278, n23256, n24287 );
nand U113221 ( n24287, n76541, n24267 );
nand U113222 ( n31481, n30577, n31537 );
nand U113223 ( n31537, n76484, n31442 );
nand U113224 ( n31549, n30577, n31558 );
nand U113225 ( n31558, n76484, n31540 );
nand U113226 ( n23944, n23256, n23983 );
nand U113227 ( n23983, n76541, n23935 );
and U113228 ( n23817, n23256, n23933 );
nand U113229 ( n23933, n76541, n23773 );
and U113230 ( n56942, n56380, n57057 );
nand U113231 ( n57057, n76283, n56898 );
nor U113232 ( n71106, n74494, n71108 );
and U113233 ( n31114, n30577, n31175 );
nand U113234 ( n31175, n76484, n31072 );
and U113235 ( n65368, n64736, n65429 );
nand U113236 ( n65429, n76217, n65274 );
nand U113237 ( n57421, n56380, n57430 );
nand U113238 ( n57430, n76282, n74490 );
nand U113239 ( n24298, n23256, n24307 );
nand U113240 ( n24307, n76540, n74491 );
nand U113241 ( n31594, n30577, n31603 );
nand U113242 ( n31603, n76483, n74488 );
nand U113243 ( n65880, n64736, n65889 );
nand U113244 ( n65889, n76216, n74487 );
nand U113245 ( n11772, n11800, n11810 );
nand U113246 ( n11863, n11772, n75207 );
nand U113247 ( n43860, n43666, n43664 );
nor U113248 ( n43855, n43856, n43857 );
nand U113249 ( n43857, n43858, n43859 );
nand U113250 ( n43859, n43860, n74396 );
nand U113251 ( n54200, n54166, n54169 );
nand U113252 ( n35702, n35668, n35671 );
nand U113253 ( n28523, n28489, n28492 );
nand U113254 ( n70428, n70394, n70397 );
nand U113255 ( n61828, n61794, n61797 );
nand U113256 ( n12149, n11772, n74785 );
nand U113257 ( n71091, n71326, n71096 );
or U113258 ( n17098, n17076, n73423 );
xnor U113259 ( n67107, n68317, n68276 );
xor U113260 ( n68317, n68275, n74695 );
xnor U113261 ( n25209, n26316, n26275 );
xor U113262 ( n26316, n26274, n74697 );
xnor U113263 ( n58345, n59455, n59414 );
xor U113264 ( n59455, n59413, n74698 );
xnor U113265 ( n46143, n47286, n47245 );
xor U113266 ( n47286, n47244, n74659 );
xnor U113267 ( n32451, n33561, n33521 );
xor U113268 ( n33561, n33520, n74696 );
xnor U113269 ( n12499, n13913, n13863 );
xor U113270 ( n13913, n13862, n74658 );
nand U113271 ( n13712, n4848, n12402 );
nand U113272 ( n33396, n3103, n32371 );
nand U113273 ( n43858, n874, n864 );
not U113274 ( n874, n43664 );
nand U113275 ( n47117, n7490, n46070 );
nand U113276 ( n68148, n5704, n67034 );
nand U113277 ( n26147, n3947, n25134 );
nand U113278 ( n59286, n6579, n58272 );
nor U113279 ( n32569, n32575, n75221 );
nor U113280 ( n32575, n31841, n32576 );
nand U113281 ( n32576, n31969, n31830 );
nor U113282 ( n25327, n25333, n75222 );
nor U113283 ( n25333, n24627, n25334 );
nand U113284 ( n25334, n24737, n24616 );
nor U113285 ( n67334, n67340, n75223 );
nor U113286 ( n67340, n66464, n67341 );
nand U113287 ( n67341, n66572, n66453 );
nor U113288 ( n58466, n58472, n75224 );
nor U113289 ( n58472, n57759, n58473 );
nand U113290 ( n58473, n57871, n57748 );
nor U113291 ( n46273, n46279, n75225 );
nor U113292 ( n46279, n45540, n46280 );
nand U113293 ( n46280, n45648, n45529 );
nand U113294 ( n21217, n21188, n21183 );
nand U113295 ( n43018, n43019, n43020 );
nand U113296 ( n43019, n43001, n74815 );
nand U113297 ( n43020, n43021, n76863 );
nor U113298 ( n43021, n8113, n43022 );
nand U113299 ( n43174, n43175, n43176 );
nand U113300 ( n43175, n43157, n74728 );
nand U113301 ( n43176, n43177, n76863 );
nor U113302 ( n43177, n8117, n43178 );
nand U113303 ( n42965, n42966, n42967 );
nand U113304 ( n42966, n42916, n74860 );
nand U113305 ( n42967, n42968, n76862 );
nor U113306 ( n42968, n8112, n42969 );
nand U113307 ( n28642, n28630, n4249 );
not U113308 ( n4249, n28643 );
nand U113309 ( n61947, n61935, n6882 );
not U113310 ( n6882, n61948 );
nand U113311 ( n70547, n70535, n6027 );
not U113312 ( n6027, n70548 );
nand U113313 ( n35821, n35809, n3412 );
not U113314 ( n3412, n35822 );
nand U113315 ( n32146, n31861, n31830 );
nand U113316 ( n66792, n66484, n66453 );
nand U113317 ( n24914, n24647, n24616 );
nand U113318 ( n58051, n57783, n57748 );
nand U113319 ( n32145, n29556, n32146 );
nand U113320 ( n66791, n63459, n66792 );
nand U113321 ( n24913, n22239, n24914 );
nand U113322 ( n58050, n55351, n58051 );
nand U113323 ( n8859, n8865, n8867 );
nand U113324 ( n8865, n8793, n74905 );
nand U113325 ( n8867, n4759, n8832 );
nand U113326 ( n42885, n42890, n42891 );
nand U113327 ( n42890, n42832, n74904 );
nand U113328 ( n42891, n7404, n42863 );
nand U113329 ( n45841, n45559, n45529 );
nand U113330 ( n45840, n42807, n45841 );
nand U113331 ( n9896, n8450, n8452 );
nor U113332 ( n8452, n8453, n8454 );
nor U113333 ( n8450, n8482, n8483 );
nand U113334 ( n8454, n8455, n8457 );
nor U113335 ( n16549, n17077, n76788 );
and U113336 ( n71337, n71326, n71098 );
xnor U113337 ( n44858, n44859, n44860 );
xor U113338 ( n44860, n74413, n44857 );
nand U113339 ( n8942, n8943, n8944 );
nand U113340 ( n8943, n8898, n74861 );
nand U113341 ( n8944, n8945, n76889 );
nor U113342 ( n8945, n5458, n8947 );
nand U113343 ( n9008, n9009, n9010 );
nand U113344 ( n9009, n8987, n74816 );
nand U113345 ( n9010, n9012, n76889 );
nor U113346 ( n9012, n5459, n9013 );
nand U113347 ( n9203, n9204, n9205 );
nand U113348 ( n9204, n9182, n74729 );
nand U113349 ( n9205, n9207, n76889 );
nor U113350 ( n9207, n5463, n9208 );
nand U113351 ( n7321, n23249, n23250 );
nor U113352 ( n23249, n23292, n23293 );
nor U113353 ( n23250, n23251, n23252 );
nor U113354 ( n23292, n23296, n23152 );
nand U113355 ( n14056, n56373, n56374 );
nor U113356 ( n56373, n56416, n56417 );
nor U113357 ( n56374, n56375, n56376 );
nor U113358 ( n56416, n56420, n56273 );
nand U113359 ( n11811, n64729, n64730 );
nor U113360 ( n64729, n64772, n64773 );
nor U113361 ( n64730, n64731, n64732 );
nor U113362 ( n64772, n75307, n64640 );
nand U113363 ( n5076, n30570, n30571 );
nor U113364 ( n30570, n30613, n30614 );
nor U113365 ( n30571, n30572, n30573 );
nor U113366 ( n30613, n75318, n30481 );
nor U113367 ( n12655, n12663, n75226 );
nor U113368 ( n12663, n11772, n12664 );
nand U113369 ( n12664, n11899, n11758 );
nand U113370 ( n7281, n23675, n23676 );
nor U113371 ( n23675, n23685, n23686 );
nor U113372 ( n23676, n23677, n23678 );
nor U113373 ( n23685, n19, n23152 );
nand U113374 ( n7291, n23586, n23587 );
nor U113375 ( n23586, n23596, n23597 );
nor U113376 ( n23587, n23588, n23589 );
nor U113377 ( n23596, n29, n23152 );
nand U113378 ( n14026, n56708, n56709 );
nor U113379 ( n56708, n56718, n56719 );
nor U113380 ( n56709, n56710, n56711 );
nor U113381 ( n56718, n280, n56273 );
nand U113382 ( n14016, n56797, n56798 );
nor U113383 ( n56797, n56807, n56808 );
nor U113384 ( n56798, n56799, n56800 );
nor U113385 ( n56807, n268, n56273 );
nand U113386 ( n7271, n23764, n23765 );
nor U113387 ( n23764, n23774, n23775 );
nor U113388 ( n23765, n23766, n23767 );
nor U113389 ( n23774, n9, n23152 );
nand U113390 ( n14006, n56889, n56890 );
nor U113391 ( n56889, n56899, n56900 );
nor U113392 ( n56890, n56891, n56892 );
nor U113393 ( n56899, n255, n56273 );
nand U113394 ( n5026, n31063, n31064 );
nor U113395 ( n31063, n31103, n31104 );
nor U113396 ( n31064, n31065, n31066 );
nor U113397 ( n31103, n75297, n30481 );
nand U113398 ( n5046, n30893, n30894 );
nor U113399 ( n30893, n30933, n30934 );
nor U113400 ( n30894, n30895, n30896 );
nor U113401 ( n30933, n75312, n30481 );
nand U113402 ( n11781, n65095, n65096 );
nor U113403 ( n65095, n65135, n65136 );
nor U113404 ( n65096, n65097, n65098 );
nor U113405 ( n65135, n75291, n64640 );
nand U113406 ( n11771, n65180, n65181 );
nor U113407 ( n65180, n65220, n65221 );
nor U113408 ( n65181, n65182, n65183 );
nor U113409 ( n65220, n75289, n64640 );
nand U113410 ( n5036, n30978, n30979 );
nor U113411 ( n30978, n31018, n31019 );
nor U113412 ( n30979, n30980, n30981 );
nor U113413 ( n31018, n75298, n30481 );
nand U113414 ( n11761, n65265, n65266 );
nor U113415 ( n65265, n65305, n65306 );
nor U113416 ( n65266, n65267, n65268 );
nor U113417 ( n65305, n75295, n64640 );
nand U113418 ( n7301, n23442, n23443 );
nor U113419 ( n23442, n23452, n23453 );
nor U113420 ( n23443, n23444, n23445 );
nor U113421 ( n23452, n38, n23152 );
nand U113422 ( n14046, n56469, n56470 );
nor U113423 ( n56469, n56479, n56480 );
nor U113424 ( n56470, n56471, n56472 );
nor U113425 ( n56479, n56515, n56273 );
nand U113426 ( n14036, n56564, n56565 );
nor U113427 ( n56564, n56574, n56575 );
nor U113428 ( n56565, n56566, n56567 );
nor U113429 ( n56574, n292, n56273 );
nand U113430 ( n7311, n23345, n23346 );
nor U113431 ( n23345, n23355, n23356 );
nor U113432 ( n23346, n23347, n23348 );
nor U113433 ( n23355, n23391, n23152 );
nand U113434 ( n5066, n30660, n30661 );
nor U113435 ( n30660, n30702, n30703 );
nor U113436 ( n30661, n30662, n30663 );
nor U113437 ( n30702, n75319, n30481 );
nand U113438 ( n5056, n30753, n30754 );
nor U113439 ( n30753, n30848, n30849 );
nor U113440 ( n30754, n30755, n30756 );
nor U113441 ( n30848, n75315, n30481 );
nand U113442 ( n11801, n64866, n64867 );
nor U113443 ( n64866, n64908, n64909 );
nor U113444 ( n64867, n64868, n64869 );
nor U113445 ( n64908, n75308, n64640 );
nand U113446 ( n11791, n64955, n64956 );
nor U113447 ( n64955, n65050, n65051 );
nor U113448 ( n64956, n64957, n64958 );
nor U113449 ( n65050, n75294, n64640 );
nand U113450 ( n42539, n43344, n43345 );
nor U113451 ( n43345, n42390, n43346 );
nor U113452 ( n43344, n43347, n43348 );
nor U113453 ( n43007, n43041, n43042 );
nor U113454 ( n43163, n43197, n43198 );
nor U113455 ( n43247, n43291, n43292 );
nand U113456 ( n23818, n76541, n74780 );
nand U113457 ( n56943, n76283, n74779 );
nand U113458 ( n31115, n76484, n74778 );
not U113459 ( n7409, n43347 );
nand U113460 ( n23639, n76541, n74878 );
nand U113461 ( n23728, n76541, n74820 );
nand U113462 ( n23550, n76541, n74923 );
nand U113463 ( n65369, n76217, n74776 );
nand U113464 ( n56761, n76283, n74877 );
nand U113465 ( n56672, n76283, n74922 );
nand U113466 ( n56850, n76283, n74819 );
nand U113467 ( n12118, n11800, n11758 );
nand U113468 ( n12117, n8762, n12118 );
nand U113469 ( n65061, n76217, n74921 );
nand U113470 ( n65146, n76217, n74875 );
nand U113471 ( n65231, n76217, n74814 );
nand U113472 ( n31029, n76484, n74817 );
nor U113473 ( n31174, n31114, n74778 );
nor U113474 ( n65428, n65368, n74776 );
nand U113475 ( n30944, n76484, n74876 );
nand U113476 ( n23306, n76540, n75037 );
nand U113477 ( n56430, n76282, n75036 );
nand U113478 ( n56525, n76282, n74971 );
nand U113479 ( n23403, n76540, n74972 );
nand U113480 ( n64830, n76216, n75028 );
nand U113481 ( n64919, n76216, n74968 );
nand U113482 ( n30859, n76484, n74927 );
nand U113483 ( n31821, n31823, n29171 );
nand U113484 ( n30624, n76483, n75041 );
nand U113485 ( n30713, n76483, n74984 );
nor U113486 ( n43094, n43111, n43112 );
nor U113487 ( n57009, n56942, n74779 );
nor U113488 ( n23885, n23817, n74780 );
nor U113489 ( n8994, n9037, n9038 );
nor U113490 ( n9189, n9232, n9233 );
nand U113491 ( n8463, n9397, n9398 );
nor U113492 ( n9398, n8304, n9399 );
nor U113493 ( n9397, n9400, n9402 );
and U113494 ( n32556, n74470, n32146 );
nor U113495 ( n9277, n9332, n9333 );
and U113496 ( n67321, n74469, n66792 );
and U113497 ( n25314, n74471, n24914 );
and U113498 ( n58453, n74472, n58051 );
and U113499 ( n46260, n74467, n45841 );
not U113500 ( n4764, n9400 );
nor U113501 ( n9103, n9124, n9125 );
or U113502 ( n43110, n73221, n43094 );
and U113503 ( n12630, n74477, n12118 );
nor U113504 ( n11397, n11398, n933 );
nor U113505 ( n11398, n11399, n76626 );
nand U113506 ( n936, n11392, n11393 );
nand U113507 ( n11393, n11394, n76628 );
nor U113508 ( n11392, n1834, n11395 );
nor U113509 ( n11395, n11397, n73506 );
or U113510 ( n43040, n74815, n43007 );
or U113511 ( n43196, n74728, n43163 );
or U113512 ( n9123, n73222, n9103 );
xor U113513 ( n32402, n33458, n73114 );
xor U113514 ( n46101, n47178, n73078 );
nand U113515 ( n30115, n76024, n75213 );
xor U113516 ( n67065, n68209, n73084 );
xor U113517 ( n25167, n26208, n73085 );
xor U113518 ( n58303, n59347, n73086 );
nand U113519 ( n64128, n75992, n75214 );
nand U113520 ( n22790, n76029, n75215 );
nand U113521 ( n55904, n76000, n75216 );
nand U113522 ( n43384, n76008, n75220 );
nand U113523 ( n9447, n76037, n75217 );
nand U113524 ( n63819, n63835, n63481 );
nand U113525 ( n63835, n63811, n6379 );
not U113526 ( n6379, n63758 );
nand U113527 ( n29863, n29879, n29582 );
nand U113528 ( n29879, n29855, n3745 );
not U113529 ( n3745, n29798 );
nand U113530 ( n22540, n22556, n22261 );
nand U113531 ( n22556, n22532, n4639 );
not U113532 ( n4639, n22477 );
nand U113533 ( n55653, n55669, n55373 );
nand U113534 ( n55669, n55645, n7272 );
not U113535 ( n7272, n55592 );
nand U113536 ( n63750, n63741, n6380 );
not U113537 ( n6380, n63628 );
nand U113538 ( n63906, n63897, n6378 );
not U113539 ( n6378, n63845 );
nand U113540 ( n29790, n29781, n3747 );
not U113541 ( n3747, n29729 );
nand U113542 ( n29950, n29941, n3744 );
not U113543 ( n3744, n29889 );
nand U113544 ( n22469, n22460, n4640 );
not U113545 ( n4640, n22408 );
nand U113546 ( n22627, n22618, n4638 );
not U113547 ( n4638, n22566 );
nand U113548 ( n55584, n55575, n7273 );
not U113549 ( n7273, n55520 );
nand U113550 ( n55740, n55731, n7270 );
not U113551 ( n7270, n55679 );
not U113552 ( n3059, n31830 );
nand U113553 ( n32310, n3059, n29717 );
not U113554 ( n3903, n24616 );
not U113555 ( n5660, n66453 );
not U113556 ( n6535, n57748 );
not U113557 ( n7434, n45529 );
nand U113558 ( n66949, n5660, n63616 );
nand U113559 ( n46009, n7434, n42978 );
nand U113560 ( n25073, n3903, n22396 );
nand U113561 ( n58208, n6535, n55508 );
not U113562 ( n247, n45392 );
or U113563 ( n9035, n74816, n8994 );
or U113564 ( n9230, n74729, n9189 );
nor U113565 ( n32150, n32152, n31869 );
nor U113566 ( n32293, n32295, n31869 );
xor U113567 ( n12447, n13788, n73109 );
nand U113568 ( n63537, n63542, n63543 );
nand U113569 ( n63543, n5630, n63515 );
nand U113570 ( n63542, n63484, n74884 );
nand U113571 ( n29638, n29643, n29644 );
nand U113572 ( n29644, n3029, n29616 );
nand U113573 ( n29643, n29585, n74885 );
nand U113574 ( n22317, n22322, n22323 );
nand U113575 ( n22323, n3873, n22295 );
nand U113576 ( n22322, n22264, n74883 );
nand U113577 ( n55429, n55434, n55435 );
nand U113578 ( n55435, n6505, n55407 );
nand U113579 ( n55434, n55376, n74882 );
nor U113580 ( n66796, n66798, n66492 );
nor U113581 ( n66932, n66934, n66492 );
nor U113582 ( n45845, n45847, n45567 );
nor U113583 ( n45981, n45983, n45567 );
nor U113584 ( n24918, n24920, n24655 );
nor U113585 ( n25056, n25058, n24655 );
nor U113586 ( n58055, n58057, n57791 );
nor U113587 ( n58191, n58193, n57791 );
or U113588 ( n42871, n74914, n42838 );
nor U113589 ( n32230, n32232, n31869 );
nor U113590 ( n8445, n8480, n8400 );
or U113591 ( n8842, n74915, n8800 );
nand U113592 ( n16166, n44986, n44987 );
nor U113593 ( n44986, n44991, n44992 );
nor U113594 ( n44987, n44988, n44989 );
nor U113595 ( n44992, n43889, n73161 );
nor U113596 ( n16583, n17076, n76788 );
not U113597 ( n4790, n11758 );
nand U113598 ( n12325, n4790, n8958 );
nor U113599 ( n12123, n12125, n11810 );
nor U113600 ( n12304, n12307, n11810 );
buf U113601 ( n76926, n72968 );
nor U113602 ( n12225, n12228, n11810 );
nand U113603 ( MUL_1411_U15, n71498, n71499 );
nand U113604 ( n71499, n71500, n71096 );
nand U113605 ( n71498, n71502, n71098 );
nand U113606 ( n71500, n71272, n71501 );
nand U113607 ( n21982, n22754, n22758 );
nand U113608 ( n22758, n22759, n22760 );
nand U113609 ( n22760, n22761, n4060 );
nand U113610 ( n22759, n4058, n22762 );
nand U113611 ( n29297, n30075, n30079 );
nand U113612 ( n30079, n30080, n30081 );
nand U113613 ( n30081, n30082, n3233 );
nand U113614 ( n30080, n3230, n30083 );
nand U113615 ( n63064, n64092, n64096 );
nand U113616 ( n64096, n64097, n64098 );
nand U113617 ( n64098, n64099, n5832 );
nand U113618 ( n64097, n5829, n64100 );
nand U113619 ( n55092, n55868, n55872 );
nand U113620 ( n55872, n55873, n55874 );
nand U113621 ( n55874, n55875, n6693 );
nand U113622 ( n55873, n6690, n55876 );
nand U113623 ( n63020, n63022, n63023 );
nor U113624 ( n63023, n63024, n63025 );
nor U113625 ( n63022, n63037, n63038 );
nor U113626 ( n63024, n63034, n63035 );
nand U113627 ( n29253, n29255, n29256 );
nor U113628 ( n29256, n29257, n29258 );
nor U113629 ( n29255, n29270, n29271 );
nor U113630 ( n29257, n29267, n29268 );
nand U113631 ( n21936, n21938, n21939 );
nor U113632 ( n21939, n21940, n21941 );
nor U113633 ( n21938, n21953, n21954 );
nor U113634 ( n21940, n21950, n21951 );
nand U113635 ( n55048, n55050, n55051 );
nor U113636 ( n55051, n55052, n55053 );
nor U113637 ( n55050, n55065, n55066 );
nor U113638 ( n55052, n55062, n55063 );
xnor U113639 ( n12523, n13962, n13922 );
xor U113640 ( n13962, n13920, n73090 );
nor U113641 ( n13953, n13955, n76594 );
nor U113642 ( n13955, n13957, n13958 );
nand U113643 ( n13957, n13985, n13987 );
nand U113644 ( n13958, n13959, n13960 );
xnor U113645 ( n67137, n68363, n68324 );
xor U113646 ( n68363, n68323, n73066 );
xnor U113647 ( n46173, n47331, n47293 );
xor U113648 ( n47331, n47292, n73065 );
xnor U113649 ( n25239, n26362, n26323 );
xor U113650 ( n26362, n26322, n73067 );
xnor U113651 ( n58375, n59501, n59462 );
xor U113652 ( n59501, n59461, n73068 );
nor U113653 ( n68352, n68353, n68354 );
nand U113654 ( n68353, n68376, n68377 );
nand U113655 ( n68354, n68355, n68356 );
nand U113656 ( n68377, n5704, n67125 );
nor U113657 ( n26351, n26352, n26353 );
nand U113658 ( n26352, n26375, n26376 );
nand U113659 ( n26353, n26354, n26355 );
nand U113660 ( n26376, n3947, n25227 );
nor U113661 ( n59490, n59491, n59492 );
nand U113662 ( n59491, n59514, n59515 );
nand U113663 ( n59492, n59493, n59494 );
nand U113664 ( n59515, n6579, n58363 );
nor U113665 ( n47318, n47320, n76328 );
nor U113666 ( n47320, n47321, n47322 );
nand U113667 ( n47321, n47344, n47345 );
nand U113668 ( n47322, n47323, n47324 );
xnor U113669 ( n32481, n33607, n33568 );
xor U113670 ( n33607, n33567, n73088 );
nor U113671 ( n33596, n33597, n33598 );
nand U113672 ( n33597, n33620, n33621 );
nand U113673 ( n33598, n33599, n33600 );
nand U113674 ( n33621, n3103, n32469 );
not U113675 ( n7959, n42581 );
and U113676 ( n42553, n42584, n7925 );
nor U113677 ( n42584, n7959, n42582 );
nand U113678 ( n71055, n71098, n71097 );
xor U113679 ( n17073, n17074, n17075 );
nor U113680 ( n17075, n75919, n17076 );
nor U113681 ( n17074, n73020, n17077 );
nand U113682 ( n12772, n12773, n12774 );
nand U113683 ( n12774, n12775, n74946 );
nand U113684 ( n12773, n12733, n73279 );
nor U113685 ( n12720, n12724, n12725 );
nor U113686 ( n12724, n74989, n12734 );
nor U113687 ( n12725, n12727, n75051 );
nand U113688 ( n12734, n12735, n75051 );
xor U113689 ( n44392, n44393, n44394 );
xor U113690 ( n44394, n74430, n859 );
nand U113691 ( n64049, n76082, n73163 );
nand U113692 ( n30032, n76154, n73164 );
nand U113693 ( n55825, n76085, n72959 );
nand U113694 ( n22709, n76157, n72958 );
nor U113695 ( n17404, n17080, n73422 );
nand U113696 ( n46362, n46363, n46364 );
nand U113697 ( n46364, n46365, n74974 );
nand U113698 ( n46363, n46332, n74986 );
nor U113699 ( n46322, n46325, n46326 );
nor U113700 ( n46325, n75016, n46333 );
nor U113701 ( n46326, n46327, n75052 );
nand U113702 ( n46333, n46334, n75052 );
nand U113703 ( n43448, n43230, n43232 );
nand U113704 ( n43445, n43446, n43447 );
nand U113705 ( n43447, n43448, n74386 );
nor U113706 ( n43441, n43442, n43443 );
nor U113707 ( n43442, n878, n43449 );
nor U113708 ( n43443, n43444, n43445 );
not U113709 ( n878, n43444 );
nand U113710 ( n30099, n35604, P1_P3_STATE2_REG_3_ );
nor U113711 ( n35604, n74591, n29162 );
nand U113712 ( n22778, n28427, P1_P2_STATE2_REG_3_ );
nor U113713 ( n28427, n74592, n21849 );
nand U113714 ( n64116, n70332, P2_P3_STATE2_REG_3_ );
nor U113715 ( n70332, n74593, n62884 );
nand U113716 ( n55892, n61732, P2_P2_STATE2_REG_3_ );
nor U113717 ( n61732, n74594, n54940 );
nand U113718 ( n43120, n43136, n42829 );
nand U113719 ( n43136, n43112, n8162 );
not U113720 ( n8162, n43059 );
nand U113721 ( n43051, n43042, n8163 );
not U113722 ( n8163, n42990 );
nand U113723 ( n43207, n43198, n8160 );
not U113724 ( n8160, n43146 );
nand U113725 ( n43446, n884, n888 );
not U113726 ( n884, n43232 );
nor U113727 ( n54224, n54230, n54231 );
nor U113728 ( n54230, n73497, n44894 );
nor U113729 ( n35726, n35732, n35733 );
nor U113730 ( n35732, n73524, n31509 );
nor U113731 ( n28547, n28553, n28554 );
nor U113732 ( n28553, n73503, n24215 );
nor U113733 ( n70452, n70458, n70459 );
nor U113734 ( n70458, n73502, n65759 );
nor U113735 ( n61852, n61858, n61859 );
nor U113736 ( n61858, n73504, n57337 );
not U113737 ( n893, n45184 );
nand U113738 ( n42425, n893, n74281 );
not U113739 ( n7958, n42627 );
nand U113740 ( n42583, n42630, n7927 );
nor U113741 ( n42630, n7958, n42628 );
nand U113742 ( n42433, n893, n74282 );
nand U113743 ( n9135, n9155, n8789 );
nand U113744 ( n9155, n9125, n5508 );
not U113745 ( n5508, n9059 );
nand U113746 ( n9049, n9038, n5509 );
not U113747 ( n5509, n8973 );
nand U113748 ( n9244, n9233, n5507 );
not U113749 ( n5507, n9168 );
nor U113750 ( n45183, n895, n42678 );
not U113751 ( n895, n42424 );
nand U113752 ( n8479, n8518, n5270 );
nor U113753 ( n8518, n5304, n8515 );
not U113754 ( n5304, n8514 );
nor U113755 ( n45249, n894, n42678 );
not U113756 ( n894, n42432 );
nand U113757 ( n71501, n1218, n71274 );
nor U113758 ( n43430, n43431, n43432 );
nand U113759 ( n43432, n43433, n43434 );
nand U113760 ( n43434, n43435, n74384 );
nand U113761 ( n43435, n43230, n43228 );
not U113762 ( n7957, n42702 );
nand U113763 ( n42629, n42705, n7928 );
nor U113764 ( n42705, n7957, n42703 );
nand U113765 ( n43433, n885, n888 );
not U113766 ( n885, n43228 );
nor U113767 ( n66319, n75304, n66323 );
nor U113768 ( n66315, n75305, n66323 );
nor U113769 ( n66311, n75306, n66323 );
nor U113770 ( n66307, n75307, n66323 );
nor U113771 ( n66237, n75289, n66323 );
nor U113772 ( n66249, n75290, n66323 );
nor U113773 ( n66261, n75308, n66323 );
nor U113774 ( n66245, n75291, n66323 );
nor U113775 ( n66257, n75309, n66323 );
nor U113776 ( n66233, n75292, n66323 );
nor U113777 ( n66241, n75293, n66323 );
nor U113778 ( n66253, n75294, n66323 );
nor U113779 ( n66229, n75295, n66323 );
nor U113780 ( n66167, n75287, n66323 );
nor U113781 ( n66265, n75310, n66323 );
nor U113782 ( n24515, n23248, n24530 );
nor U113783 ( n24511, n23296, n24530 );
nor U113784 ( n24499, n23441, n24530 );
nor U113785 ( n24525, n23151, n24530 );
nor U113786 ( n24521, n23199, n24530 );
nor U113787 ( n57645, n56369, n57658 );
nor U113788 ( n57641, n56420, n57658 );
nor U113789 ( n57626, n56563, n57658 );
nor U113790 ( n57649, n56320, n57658 );
nor U113791 ( n57630, n56515, n57658 );
nor U113792 ( n57653, n56272, n57658 );
nor U113793 ( n24503, n23391, n24530 );
nor U113794 ( n57637, n56468, n57658 );
nor U113795 ( n24507, n23344, n24530 );
nand U113796 ( n21970, n22772, n22773 );
nor U113797 ( n22772, n3875, n73181 );
nand U113798 ( n29285, n30093, n30094 );
nor U113799 ( n30093, n3032, n73182 );
nand U113800 ( n63052, n64110, n64111 );
nor U113801 ( n64110, n5633, n73183 );
nand U113802 ( n55080, n55886, n55887 );
nor U113803 ( n55886, n6508, n73180 );
nand U113804 ( n63521, n5630, n63514 );
nand U113805 ( n29622, n3029, n29615 );
nand U113806 ( n22301, n3873, n22294 );
nand U113807 ( n55413, n6505, n55406 );
nor U113808 ( n40475, n40362, n76399 );
nor U113809 ( n40655, n2212, n76399 );
not U113810 ( n2212, n40315 );
nor U113811 ( n40545, n40415, n76398 );
nor U113812 ( n40537, n40418, n76398 );
not U113813 ( n7955, n42763 );
nand U113814 ( n42704, n42766, n7929 );
nor U113815 ( n42766, n7955, n42764 );
nor U113816 ( n40567, n76397, n40569 );
nand U113817 ( n40569, n39627, n39626 );
and U113818 ( n8399, n8400, n8402 );
nor U113819 ( n40648, n76398, n40650 );
nand U113820 ( n40650, n40290, n40289 );
nor U113821 ( n13169, n76626, n13172 );
nand U113822 ( n13172, n13173, n13174 );
nor U113823 ( n14370, n76626, n14373 );
nand U113824 ( n14373, n14374, n14375 );
nor U113825 ( n14918, n76625, n14920 );
nand U113826 ( n14920, n14922, n14923 );
nor U113827 ( n15209, n76625, n15212 );
nand U113828 ( n15212, n15213, n15214 );
nor U113829 ( n15477, n76625, n15479 );
nand U113830 ( n15479, n15480, n15482 );
nor U113831 ( n15740, n76625, n15743 );
nand U113832 ( n15743, n15744, n15745 );
nor U113833 ( n15997, n76625, n15999 );
nand U113834 ( n15999, n16000, n16002 );
nor U113835 ( n16265, n76625, n16268 );
nand U113836 ( n16268, n16269, n16270 );
nor U113837 ( n40637, n76397, n40639 );
nand U113838 ( n40639, n40206, n40205 );
nor U113839 ( n40626, n76397, n40628 );
nand U113840 ( n40628, n40129, n40128 );
nor U113841 ( n40611, n76397, n40613 );
nand U113842 ( n40613, n40036, n40035 );
nor U113843 ( n40589, n76397, n40591 );
nand U113844 ( n40591, n39857, n39856 );
nor U113845 ( n40578, n76397, n40580 );
nand U113846 ( n40580, n39756, n39755 );
nor U113847 ( n40507, n76397, n40509 );
nand U113848 ( n40509, n40458, n40457 );
nor U113849 ( n12647, n76625, n12649 );
or U113850 ( n12649, n12650, n12652 );
nor U113851 ( n40600, n76397, n40602 );
nand U113852 ( n40602, n39956, n39955 );
not U113853 ( n5303, n8572 );
nand U113854 ( n8517, n8575, n5272 );
nor U113855 ( n8575, n5303, n8573 );
nand U113856 ( n42864, n42907, n7933 );
nor U113857 ( n42907, n7950, n42905 );
not U113858 ( n7950, n42904 );
not U113859 ( n7952, n45928 );
nand U113860 ( n42765, n42810, n7930 );
nor U113861 ( n42810, n42807, n42808 );
nor U113862 ( n16698, n76626, n16700 );
nand U113863 ( n16700, n16702, n16703 );
xor U113864 ( n42554, n75077, n45560 );
nor U113865 ( n26916, n26917, n26905 );
nor U113866 ( n26917, n26918, n24460 );
nor U113867 ( n60056, n60057, n60045 );
nor U113868 ( n60057, n60058, n57586 );
nor U113869 ( n34161, n34162, n34150 );
nor U113870 ( n34162, n34163, n31722 );
nor U113871 ( n68915, n68916, n68904 );
nor U113872 ( n68916, n68917, n66162 );
nand U113873 ( n25421, n25422, n25423 );
nand U113874 ( n25423, n25424, n74975 );
nand U113875 ( n25422, n25391, n75007 );
nand U113876 ( n58558, n58559, n58560 );
nand U113877 ( n58560, n58561, n74977 );
nand U113878 ( n58559, n58528, n75008 );
nand U113879 ( n32661, n32662, n32663 );
nand U113880 ( n32663, n32664, n74973 );
nand U113881 ( n32662, n32631, n75010 );
nand U113882 ( n67426, n67427, n67428 );
nand U113883 ( n67428, n67429, n74976 );
nand U113884 ( n67427, n67396, n75009 );
nand U113885 ( n46298, n47786, n73190 );
nand U113886 ( n12687, n14532, n73191 );
nand U113887 ( n47786, n47871, n47872 );
nand U113888 ( n47872, n42324, n74648 );
nand U113889 ( n47871, n7463, n47874 );
nand U113890 ( n47874, n47875, n47876 );
nand U113891 ( n14532, n14638, n14639 );
nand U113892 ( n14639, n8264, n74649 );
nand U113893 ( n14638, n4819, n14642 );
nand U113894 ( n14642, n14643, n14644 );
nor U113895 ( n47788, n47789, n76328 );
nor U113896 ( n47789, n47790, n47791 );
nand U113897 ( n47790, n47798, n47799 );
nand U113898 ( n47791, n47792, n47793 );
nor U113899 ( n14534, n14535, n76594 );
nor U113900 ( n14535, n14537, n14538 );
nand U113901 ( n14537, n14547, n14548 );
nand U113902 ( n14538, n14539, n14540 );
nor U113903 ( n14380, n74656, n76598 );
nor U113904 ( n47665, n74655, n76332 );
nor U113905 ( n47588, n72964, n76332 );
nor U113906 ( n14275, n72965, n76598 );
nor U113907 ( n14169, n74673, n76598 );
nor U113908 ( n47503, n74672, n76332 );
nor U113909 ( n14072, n74727, n76598 );
nor U113910 ( n47424, n74726, n76332 );
nor U113911 ( n47740, n72962, n76332 );
nor U113912 ( n14474, n72963, n76598 );
nor U113913 ( n32621, n32624, n32625 );
nor U113914 ( n32624, n75042, n32632 );
nor U113915 ( n32625, n32626, n75065 );
nand U113916 ( n32632, n32633, n75065 );
nor U113917 ( n25381, n25384, n25385 );
nor U113918 ( n25384, n75038, n25392 );
nor U113919 ( n25385, n25386, n75066 );
nand U113920 ( n25392, n25393, n75066 );
nor U113921 ( n67386, n67389, n67390 );
nor U113922 ( n67389, n75039, n67397 );
nor U113923 ( n67390, n67391, n75068 );
nand U113924 ( n67397, n67398, n75068 );
nor U113925 ( n58518, n58521, n58522 );
nor U113926 ( n58521, n75040, n58529 );
nor U113927 ( n58522, n58523, n75067 );
nand U113928 ( n58529, n58530, n75067 );
nor U113929 ( n22034, n74999, n22036 );
nor U113930 ( n55144, n75000, n55146 );
nor U113931 ( n29353, n75004, n29355 );
nor U113932 ( n63116, n75003, n63118 );
buf U113933 ( n76330, n76327 );
buf U113934 ( n76596, n76593 );
not U113935 ( n5302, n8635 );
nand U113936 ( n8574, n8639, n5273 );
nor U113937 ( n8639, n5302, n8637 );
nor U113938 ( n32907, n32908, n32909 );
nand U113939 ( n32908, n32912, n32852 );
nand U113940 ( n32909, n3095, n32910 );
nand U113941 ( n32912, n32664, n74652 );
nor U113942 ( n67668, n67669, n67670 );
nand U113943 ( n67669, n67673, n67617 );
nand U113944 ( n67670, n5697, n67671 );
nand U113945 ( n67673, n67429, n74595 );
nor U113946 ( n25663, n25664, n25665 );
nand U113947 ( n25664, n25668, n25612 );
nand U113948 ( n25665, n3939, n25666 );
nand U113949 ( n25668, n25424, n74596 );
nor U113950 ( n58803, n58804, n58805 );
nand U113951 ( n58804, n58808, n58749 );
nand U113952 ( n58805, n6572, n58806 );
nand U113953 ( n58808, n58561, n74597 );
nor U113954 ( n33254, n33255, n33181 );
nor U113955 ( n33255, n33257, n73160 );
nor U113956 ( n68013, n68014, n67932 );
nor U113957 ( n68014, n68016, n74431 );
nor U113958 ( n26010, n26011, n25929 );
nor U113959 ( n26011, n26013, n74432 );
nor U113960 ( n59148, n59149, n59067 );
nor U113961 ( n59149, n59151, n74433 );
nor U113962 ( n13298, n13299, n13300 );
nand U113963 ( n13299, n13304, n4863 );
nand U113964 ( n13300, n4828, n13302 );
nand U113965 ( n13304, n12732, n74599 );
xor U113966 ( n43075, n74554, n46058 );
nand U113967 ( n42906, n42980, n7934 );
nor U113968 ( n42980, n42977, n42978 );
nor U113969 ( n25552, n25553, n25506 );
nor U113970 ( n25553, n25558, n74949 );
nor U113971 ( n32792, n32793, n32746 );
nor U113972 ( n32793, n32798, n74948 );
nor U113973 ( n67557, n67558, n67511 );
nor U113974 ( n67558, n67563, n74947 );
nor U113975 ( n58689, n58690, n58643 );
nor U113976 ( n58690, n58695, n74950 );
nor U113977 ( n13484, n13485, n13428 );
nor U113978 ( n13485, n13489, n74823 );
nor U113979 ( n13489, n13490, n13440 );
nor U113980 ( n13490, n73117, n13492 );
not U113981 ( n200, n29171 );
nor U113982 ( n46494, n46495, n46447 );
nor U113983 ( n46495, n46500, n74919 );
nor U113984 ( n46500, n46501, n7483 );
not U113985 ( n7483, n46457 );
nor U113986 ( n46501, n73220, n46502 );
not U113987 ( n5300, n8707 );
nand U113988 ( n8638, n8710, n5274 );
nor U113989 ( n8710, n5300, n8708 );
nor U113990 ( n12953, n12893, n12997 );
nor U113991 ( n12997, n12998, n74774 );
and U113992 ( n12994, n75840, n12953 );
or U113993 ( n75840, n12952, n13003 );
nor U113994 ( n21226, n21232, n21233 );
nor U113995 ( n21232, n73525, n11184 );
nor U113996 ( n13090, n13092, n13093 );
nand U113997 ( n13092, n13097, n12993 );
nand U113998 ( n13093, n4839, n13094 );
nand U113999 ( n13097, n12775, n74625 );
nor U114000 ( n46621, n46622, n46623 );
nand U114001 ( n46622, n46626, n46570 );
nand U114002 ( n46623, n7482, n46624 );
nand U114003 ( n46626, n46365, n74585 );
nand U114004 ( n68245, n67396, n73187 );
nand U114005 ( n26244, n25391, n73188 );
nand U114006 ( n59383, n58528, n73189 );
nor U114007 ( n68242, n68243, n68244 );
nand U114008 ( n68243, n68248, n68249 );
nand U114009 ( n68244, n5692, n68245 );
nand U114010 ( n68248, n67429, n74695 );
nor U114011 ( n26241, n26242, n26243 );
nand U114012 ( n26242, n26247, n26248 );
nand U114013 ( n26243, n3934, n26244 );
nand U114014 ( n26247, n25424, n74697 );
nor U114015 ( n59380, n59381, n59382 );
nand U114016 ( n59381, n59386, n59387 );
nand U114017 ( n59382, n6567, n59383 );
nand U114018 ( n59386, n58561, n74698 );
nor U114019 ( n13537, n13538, n13440 );
nor U114020 ( n13538, n13540, n73117 );
nand U114021 ( n33490, n32631, n73197 );
nand U114022 ( n33136, n32631, n74879 );
nor U114023 ( n33487, n33488, n33489 );
nand U114024 ( n33488, n33493, n33494 );
nand U114025 ( n33489, n3090, n33490 );
nand U114026 ( n33493, n32664, n74696 );
nor U114027 ( n33133, n33134, n33135 );
nand U114028 ( n33134, n33138, n3122 );
nand U114029 ( n33135, n3094, n33136 );
nand U114030 ( n33138, n32664, n74845 );
nand U114031 ( n8833, n8887, n5278 );
nor U114032 ( n8887, n5295, n8884 );
not U114033 ( n5295, n8883 );
nand U114034 ( n32910, n32631, n75050 );
nand U114035 ( n67892, n67396, n74872 );
nand U114036 ( n25889, n25391, n74873 );
nand U114037 ( n59027, n58528, n74874 );
not U114038 ( n5297, n12238 );
nand U114039 ( n8709, n8765, n5275 );
nor U114040 ( n8765, n8762, n8763 );
nor U114041 ( n67889, n67890, n67891 );
nand U114042 ( n67890, n67894, n5722 );
nand U114043 ( n67891, n5695, n67892 );
nand U114044 ( n67894, n67429, n73130 );
nor U114045 ( n25886, n25887, n25888 );
nand U114046 ( n25887, n25891, n3964 );
nand U114047 ( n25888, n3938, n25889 );
nand U114048 ( n25891, n25424, n73131 );
nor U114049 ( n59024, n59025, n59026 );
nand U114050 ( n59025, n59029, n6597 );
nand U114051 ( n59026, n6570, n59027 );
nand U114052 ( n59029, n58561, n73132 );
nand U114053 ( n67671, n67396, n74637 );
nand U114054 ( n25666, n25391, n74638 );
nand U114055 ( n58806, n58528, n74639 );
or U114056 ( n68009, n68011, n75841 );
and U114057 ( n75841, n67396, n74431 );
or U114058 ( n26006, n26008, n75842 );
and U114059 ( n75842, n25391, n74432 );
or U114060 ( n59144, n59146, n75843 );
and U114061 ( n75843, n58528, n74433 );
xor U114062 ( n43127, n74522, n46100 );
or U114063 ( n33250, n33252, n75844 );
and U114064 ( n75844, n32631, n73160 );
nor U114065 ( n46978, n46979, n46885 );
nor U114066 ( n46979, n46981, n74417 );
not U114067 ( n888, n43230 );
nand U114068 ( n45174, n45177, n45168 );
nand U114069 ( n45177, n888, n74384 );
nor U114070 ( n68674, n68675, n68676 );
nand U114071 ( n68676, n68677, n68600 );
nand U114072 ( n68677, n67396, n74587 );
nor U114073 ( n33918, n33919, n33920 );
nand U114074 ( n33920, n33921, n33844 );
nand U114075 ( n33921, n32631, n74588 );
nor U114076 ( n26673, n26674, n26675 );
nand U114077 ( n26675, n26676, n26599 );
nand U114078 ( n26676, n25391, n74589 );
nor U114079 ( n59815, n59816, n59817 );
nand U114080 ( n59817, n59818, n59741 );
nand U114081 ( n59818, n58528, n74590 );
nor U114082 ( n68610, n68611, n68612 );
nand U114083 ( n68612, n68613, n68614 );
nand U114084 ( n68611, n68633, n68634 );
nand U114085 ( n68613, n67194, n76708 );
nor U114086 ( n33854, n33855, n33856 );
nand U114087 ( n33856, n33857, n33858 );
nand U114088 ( n33855, n33877, n33878 );
nand U114089 ( n33857, n32538, n76774 );
nor U114090 ( n26609, n26610, n26611 );
nand U114091 ( n26611, n26612, n26613 );
nand U114092 ( n26610, n26632, n26633 );
nand U114093 ( n26612, n25296, n76754 );
nor U114094 ( n59751, n59752, n59753 );
nand U114095 ( n59753, n59754, n59755 );
nand U114096 ( n59752, n59774, n59775 );
nand U114097 ( n59754, n58432, n76687 );
not U114098 ( n472, n62893 );
nand U114099 ( n68675, n68713, n68714 );
nand U114100 ( n68714, n67429, n73076 );
nand U114101 ( n68713, n67396, n75054 );
nand U114102 ( n33919, n33957, n33958 );
nand U114103 ( n33958, n32664, n73077 );
nand U114104 ( n33957, n32631, n75055 );
nand U114105 ( n26674, n26712, n26713 );
nand U114106 ( n26713, n25424, n73075 );
nand U114107 ( n26712, n25391, n75056 );
nand U114108 ( n59816, n59854, n59855 );
nand U114109 ( n59855, n58561, n73074 );
nand U114110 ( n59854, n58528, n75057 );
nand U114111 ( n43303, n76102, n72962 );
nand U114112 ( n45239, n45242, n45233 );
nand U114113 ( n45242, n888, n74386 );
nor U114114 ( n68431, n68338, n68432 );
nand U114115 ( n68432, n68433, n68434 );
or U114116 ( n68434, n5714, n68343 );
nand U114117 ( n68433, n67396, n74452 );
nor U114118 ( n33675, n33582, n33676 );
nand U114119 ( n33676, n33677, n33678 );
or U114120 ( n33678, n3113, n33587 );
nand U114121 ( n33677, n32631, n74455 );
nor U114122 ( n26430, n26337, n26431 );
nand U114123 ( n26431, n26432, n26433 );
or U114124 ( n26433, n3957, n26342 );
nand U114125 ( n26432, n25391, n74453 );
nor U114126 ( n59569, n59476, n59570 );
nand U114127 ( n59570, n59571, n59572 );
or U114128 ( n59572, n6589, n59481 );
nand U114129 ( n59571, n58528, n74454 );
or U114130 ( n42503, n42528, n75845 );
and U114131 ( n75845, n42527, n73391 );
xnor U114132 ( n8478, n75170, n11802 );
nor U114133 ( n8510, n5269, n8512 );
nor U114134 ( n8512, n8513, n8514 );
not U114135 ( n5269, n8479 );
nor U114136 ( n8513, n8515, n8517 );
nand U114137 ( n63516, n63559, n6145 );
nor U114138 ( n63559, n6163, n63557 );
nand U114139 ( n29617, n29660, n3530 );
nor U114140 ( n29660, n3548, n29658 );
nand U114141 ( n22296, n22339, n4368 );
nor U114142 ( n22339, n4385, n22337 );
nand U114143 ( n55408, n55451, n7000 );
nor U114144 ( n55451, n7018, n55449 );
not U114145 ( n6163, n63556 );
not U114146 ( n3548, n29657 );
not U114147 ( n4385, n22336 );
not U114148 ( n7018, n55448 );
nand U114149 ( n63043, n63094, n63095 );
nand U114150 ( n29276, n29331, n29332 );
nand U114151 ( n21959, n22012, n22013 );
nand U114152 ( n55071, n55122, n55123 );
nand U114153 ( n63169, n63221, n6140 );
nor U114154 ( n63221, n63218, n63219 );
nand U114155 ( n63220, n63344, n6142 );
nor U114156 ( n63344, n63341, n63342 );
nand U114157 ( n63343, n63462, n6143 );
nor U114158 ( n63462, n63459, n63460 );
nand U114159 ( n29406, n29458, n3525 );
nor U114160 ( n29458, n29455, n29456 );
nand U114161 ( n29457, n29515, n3527 );
nor U114162 ( n29515, n29512, n29513 );
nand U114163 ( n29514, n29559, n3528 );
nor U114164 ( n29559, n29556, n29557 );
nand U114165 ( n22087, n22139, n4363 );
nor U114166 ( n22139, n22136, n22137 );
nand U114167 ( n22138, n22196, n4364 );
nor U114168 ( n22196, n22193, n22194 );
nand U114169 ( n55197, n55249, n6995 );
nor U114170 ( n55249, n55246, n55247 );
nand U114171 ( n55248, n55310, n6997 );
nor U114172 ( n55310, n55307, n55308 );
nand U114173 ( n63124, n63170, n6139 );
nor U114174 ( n63170, n63167, n63168 );
nand U114175 ( n29361, n29407, n3524 );
nor U114176 ( n29407, n29404, n29405 );
nand U114177 ( n22042, n22088, n4362 );
nor U114178 ( n22088, n22085, n22086 );
nand U114179 ( n22195, n22242, n4365 );
nor U114180 ( n22242, n22239, n22240 );
nand U114181 ( n55152, n55198, n6994 );
nor U114182 ( n55198, n55195, n55196 );
nand U114183 ( n55309, n55354, n6998 );
nor U114184 ( n55354, n55351, n55352 );
nand U114185 ( n63461, n63517, n6144 );
nor U114186 ( n63517, n63515, n63514 );
nand U114187 ( n29558, n29618, n3529 );
nor U114188 ( n29618, n29616, n29615 );
nand U114189 ( n22241, n22297, n4367 );
nor U114190 ( n22297, n22295, n22294 );
nand U114191 ( n55353, n55409, n6999 );
nor U114192 ( n55409, n55407, n55406 );
not U114193 ( n6164, n66878 );
not U114194 ( n3549, n32240 );
not U114195 ( n4387, n25002 );
not U114196 ( n7019, n58137 );
and U114197 ( n22012, n22043, n4360 );
nor U114198 ( n22043, n22040, n22041 );
and U114199 ( n29331, n29362, n3523 );
nor U114200 ( n29362, n29359, n29360 );
and U114201 ( n63094, n63125, n6138 );
nor U114202 ( n63125, n63122, n63123 );
and U114203 ( n55122, n55153, n6993 );
nor U114204 ( n55153, n55150, n55151 );
nand U114205 ( n9347, n76172, n72963 );
or U114206 ( n8418, n8449, n75846 );
and U114207 ( n75846, n8448, n73392 );
nand U114208 ( n13824, n12733, n73176 );
nor U114209 ( n13820, n13822, n13823 );
nand U114210 ( n13822, n13828, n13829 );
nand U114211 ( n13823, n4834, n13824 );
nand U114212 ( n13828, n12775, n74658 );
nand U114213 ( n13094, n12733, n74920 );
nand U114214 ( n63025, n63026, n63027 );
nand U114215 ( n63027, n482, n63028 );
nand U114216 ( n63026, n483, n63032 );
xor U114217 ( n63028, n75179, n63029 );
nand U114218 ( n29258, n29259, n29260 );
nand U114219 ( n29260, n210, n29261 );
nand U114220 ( n29259, n212, n29265 );
xor U114221 ( n29261, n75180, n29262 );
nand U114222 ( n21941, n21942, n21943 );
nand U114223 ( n21943, n177, n21944 );
nand U114224 ( n21942, n178, n21948 );
xor U114225 ( n21944, n75178, n21945 );
nand U114226 ( n55053, n55054, n55055 );
nand U114227 ( n55055, n448, n55056 );
nand U114228 ( n55054, n449, n55060 );
xor U114229 ( n55056, n75177, n55057 );
nand U114230 ( n13384, n12733, n74847 );
nor U114231 ( n13380, n13382, n13383 );
nand U114232 ( n13382, n13387, n4863 );
nand U114233 ( n13383, n4838, n13384 );
nand U114234 ( n13387, n12775, n74818 );
or U114235 ( n13532, n13534, n75847 );
and U114236 ( n75847, n12733, n73117 );
nand U114237 ( n25544, n25550, n25551 );
nand U114238 ( n25551, n25424, n73224 );
nand U114239 ( n25550, n25391, n74949 );
nand U114240 ( n32784, n32790, n32791 );
nand U114241 ( n32791, n32664, n73232 );
nand U114242 ( n32790, n32631, n74948 );
nand U114243 ( n67549, n67555, n67556 );
nand U114244 ( n67556, n67429, n73223 );
nand U114245 ( n67555, n67396, n74947 );
nand U114246 ( n58681, n58687, n58688 );
nand U114247 ( n58688, n58561, n73225 );
nand U114248 ( n58687, n58528, n74950 );
nand U114249 ( n68510, n67826, n75937 );
nand U114250 ( n33754, n33070, n75940 );
nand U114251 ( n26509, n25823, n75938 );
nand U114252 ( n59648, n58961, n75939 );
nor U114253 ( n68446, n68447, n68448 );
nand U114254 ( n68448, n68449, n68450 );
nand U114255 ( n68447, n68467, n68468 );
nand U114256 ( n68450, n76705, n67146 );
nor U114257 ( n33690, n33691, n33692 );
nand U114258 ( n33692, n33693, n33694 );
nand U114259 ( n33691, n33711, n33712 );
nand U114260 ( n33694, n76772, n32490 );
nor U114261 ( n26445, n26446, n26447 );
nand U114262 ( n26447, n26448, n26449 );
nand U114263 ( n26446, n26466, n26467 );
nand U114264 ( n26449, n76751, n25248 );
nor U114265 ( n59584, n59585, n59586 );
nand U114266 ( n59586, n59587, n59588 );
nand U114267 ( n59585, n59605, n59606 );
nand U114268 ( n59588, n76684, n58384 );
nor U114269 ( n41966, n41967, n41968 );
nor U114270 ( n41967, n41969, n41460 );
nor U114271 ( n41969, n41970, n41971 );
nand U114272 ( n41971, n839, n41471 );
nor U114273 ( n68507, n68508, n68509 );
nand U114274 ( n68508, n68435, n68512 );
nand U114275 ( n68509, n5715, n68510 );
nand U114276 ( n68512, n67395, n74408 );
nor U114277 ( n33751, n33752, n33753 );
nand U114278 ( n33752, n33679, n33756 );
nand U114279 ( n33753, n3114, n33754 );
nand U114280 ( n33756, n32630, n74412 );
nor U114281 ( n26506, n26507, n26508 );
nand U114282 ( n26507, n26434, n26511 );
nand U114283 ( n26508, n3958, n26509 );
nand U114284 ( n26511, n25390, n74409 );
nor U114285 ( n59645, n59646, n59647 );
nand U114286 ( n59646, n59573, n59650 );
nand U114287 ( n59647, n6590, n59648 );
nand U114288 ( n59650, n58527, n74410 );
nor U114289 ( n14357, n14358, n14359 );
nand U114290 ( n14359, n14360, n14264 );
nand U114291 ( n14360, n12733, n74579 );
nor U114292 ( n14277, n14278, n14279 );
nand U114293 ( n14279, n14280, n14282 );
nand U114294 ( n14278, n14305, n14307 );
nand U114295 ( n14280, n12608, n76727 );
nand U114296 ( n14358, n14414, n14415 );
nand U114297 ( n14415, n12775, n73079 );
nand U114298 ( n14414, n12733, n75059 );
nand U114299 ( n67825, n67826, n74574 );
nand U114300 ( n25822, n25823, n74575 );
nand U114301 ( n58960, n58961, n74576 );
nor U114302 ( n67822, n67823, n67824 );
nand U114303 ( n67823, n67828, n5722 );
nand U114304 ( n67824, n5687, n67825 );
nand U114305 ( n67828, n67395, n74546 );
nor U114306 ( n25819, n25820, n25821 );
nand U114307 ( n25820, n25825, n3964 );
nand U114308 ( n25821, n3929, n25822 );
nand U114309 ( n25825, n25390, n74547 );
nor U114310 ( n58957, n58958, n58959 );
nand U114311 ( n58958, n58963, n6597 );
nand U114312 ( n58959, n6562, n58960 );
nand U114313 ( n58963, n58527, n74548 );
nand U114314 ( n68289, n67826, n74695 );
nand U114315 ( n26288, n25823, n74697 );
nand U114316 ( n59427, n58961, n74698 );
nand U114317 ( n33069, n33070, n74610 );
nor U114318 ( n33066, n33067, n33068 );
nand U114319 ( n33067, n33072, n3122 );
nand U114320 ( n33068, n3085, n33069 );
nand U114321 ( n33072, n32630, n74635 );
nor U114322 ( n14054, n13939, n14055 );
nand U114323 ( n14055, n14057, n14058 );
or U114324 ( n14058, n4855, n13944 );
nand U114325 ( n14057, n12733, n74461 );
nand U114326 ( n68161, n67826, n74758 );
nand U114327 ( n26160, n25823, n74759 );
nand U114328 ( n59299, n58961, n74760 );
xor U114329 ( n43187, n74500, n46154 );
nand U114330 ( n33533, n33070, n74696 );
nand U114331 ( n47214, n46332, n73178 );
nand U114332 ( n33411, n33070, n73115 );
nor U114333 ( n47211, n47212, n47213 );
nand U114334 ( n47212, n47217, n47218 );
nand U114335 ( n47213, n7477, n47214 );
nand U114336 ( n47217, n46365, n74659 );
nand U114337 ( n46845, n46332, n74841 );
nor U114338 ( n46842, n46843, n46844 );
nand U114339 ( n46843, n46847, n7508 );
nand U114340 ( n46844, n7480, n46845 );
nand U114341 ( n46847, n46365, n73118 );
nand U114342 ( n46624, n46332, n73159 );
or U114343 ( n46974, n46976, n75848 );
and U114344 ( n75848, n46332, n74417 );
nor U114345 ( n13389, n13393, n74847 );
nand U114346 ( n22031, n76157, n74999 );
nand U114347 ( n29350, n76154, n75004 );
nand U114348 ( n63113, n76082, n75003 );
nand U114349 ( n55141, n76085, n75000 );
nor U114350 ( n13103, n13048, n13153 );
nor U114351 ( n13153, n13154, n74625 );
nor U114352 ( n13100, n13103, n74920 );
nor U114353 ( n47653, n47654, n47655 );
nand U114354 ( n47655, n47656, n47579 );
nand U114355 ( n47656, n46332, n74580 );
nand U114356 ( n63491, n76082, n74900 );
nand U114357 ( n63646, n76082, n74800 );
nand U114358 ( n63863, n76082, n74711 );
nand U114359 ( n29592, n76154, n74901 );
nand U114360 ( n29747, n76154, n74801 );
nand U114361 ( n29907, n76154, n74712 );
nor U114362 ( n47589, n47590, n47591 );
nand U114363 ( n47591, n47592, n47593 );
nand U114364 ( n47590, n47612, n47613 );
nand U114365 ( n47592, n46242, n76660 );
nand U114366 ( n22426, n76157, n74799 );
nand U114367 ( n22584, n76157, n74710 );
nand U114368 ( n22271, n76157, n74899 );
nand U114369 ( n55541, n76085, n74798 );
nand U114370 ( n55697, n76085, n74709 );
nand U114371 ( n55383, n76085, n74898 );
nand U114372 ( n21985, n21986, n73317 );
nand U114373 ( n29300, n29301, n73318 );
nand U114374 ( n63067, n63068, n73319 );
nand U114375 ( n55095, n55096, n73316 );
nand U114376 ( n63332, n76082, n74944 );
nand U114377 ( n29503, n76154, n74945 );
nand U114378 ( n22184, n76157, n74939 );
nand U114379 ( n55298, n76085, n74938 );
xor U114380 ( n63939, n74479, n67158 );
xor U114381 ( n29983, n74478, n32502 );
xor U114382 ( n22660, n74480, n25260 );
xor U114383 ( n55773, n74481, n58396 );
nand U114384 ( n47654, n47692, n47693 );
nand U114385 ( n47693, n46365, n73071 );
nand U114386 ( n47692, n46332, n75058 );
nand U114387 ( n63558, n63618, n6147 );
nor U114388 ( n63618, n63615, n63616 );
nand U114389 ( n29659, n29719, n3532 );
nor U114390 ( n29719, n29716, n29717 );
nand U114391 ( n22338, n22398, n4369 );
nor U114392 ( n22398, n22395, n22396 );
nand U114393 ( n55450, n55510, n7002 );
nor U114394 ( n55510, n55507, n55508 );
nand U114395 ( n63794, n76082, n73216 );
nand U114396 ( n29678, n76154, n74839 );
nand U114397 ( n29834, n76154, n73217 );
nand U114398 ( n63577, n76082, n74840 );
nand U114399 ( n22515, n76157, n73215 );
nand U114400 ( n22357, n76157, n74838 );
nand U114401 ( n55628, n76085, n73214 );
nand U114402 ( n55469, n76085, n74837 );
xnor U114403 ( n43031, n74607, n46011 );
nor U114404 ( n47399, n47307, n47400 );
nand U114405 ( n47400, n47401, n47402 );
or U114406 ( n47402, n7500, n47311 );
nand U114407 ( n47401, n46332, n74443 );
nor U114408 ( n17091, n17080, n73423 );
nand U114409 ( n63933, n76082, n73168 );
nand U114410 ( n29977, n76154, n73169 );
nand U114411 ( n22654, n76157, n72961 );
nand U114412 ( n55767, n76085, n72960 );
xor U114413 ( n63826, n74526, n67064 );
xor U114414 ( n29870, n74527, n32401 );
xor U114415 ( n22547, n74528, n25166 );
xor U114416 ( n55660, n74529, n58302 );
xor U114417 ( n63886, n74502, n67118 );
xor U114418 ( n29930, n74503, n32462 );
xor U114419 ( n22607, n74504, n25220 );
xor U114420 ( n55720, n74505, n58356 );
nand U114421 ( n63203, n76082, n74993 );
nand U114422 ( n29440, n76154, n74994 );
nand U114423 ( n22121, n76157, n74991 );
nand U114424 ( n55231, n76085, n74990 );
xor U114425 ( n63774, n74558, n67022 );
xor U114426 ( n29814, n74557, n32359 );
xor U114427 ( n22495, n74559, n25122 );
xor U114428 ( n55608, n74560, n58260 );
nor U114429 ( n33540, n3113, n74696 );
xor U114430 ( n9079, n74577, n12387 );
nand U114431 ( n8885, n8960, n5279 );
nor U114432 ( n8960, n8957, n8958 );
nand U114433 ( n14152, n12828, n75941 );
nor U114434 ( n14073, n14074, n14075 );
nand U114435 ( n14075, n14076, n14077 );
nand U114436 ( n14074, n14098, n14099 );
nand U114437 ( n14077, n76724, n12548 );
nor U114438 ( n14148, n14149, n14150 );
nand U114439 ( n14149, n14059, n14154 );
nand U114440 ( n14150, n4857, n14152 );
nand U114441 ( n14154, n12732, n74429 );
or U114442 ( n12988, n12938, n75849 );
and U114443 ( n75849, n12828, n74774 );
not U114444 ( n880, n45243 );
nor U114445 ( n68296, n5714, n74695 );
nor U114446 ( n26295, n3957, n74697 );
nor U114447 ( n59434, n6589, n74698 );
nand U114448 ( n45168, n880, n74381 );
nand U114449 ( n13302, n12828, n74586 );
nand U114450 ( n14832, n76592, n11595 );
nand U114451 ( n13878, n12828, n74658 );
xor U114452 ( n42490, n45531, n74931 );
xor U114453 ( n43560, n872, n43561 );
xor U114454 ( n43561, n74379, n43559 );
nand U114455 ( n45233, n880, n74380 );
nand U114456 ( n13728, n12828, n74735 );
nand U114457 ( n781, n21768, n6429 );
nor U114458 ( n21768, n76682, n21769 );
not U114459 ( n7319, n796 );
xnor U114460 ( n42862, n74772, n45880 );
xor U114461 ( n43254, n74473, n46194 );
nand U114462 ( n9431, n11305, n11307 );
nor U114463 ( n11305, n11312, n11313 );
nor U114464 ( n11307, n11308, n11309 );
nor U114465 ( n11313, n9965, n73162 );
nand U114466 ( n47489, n46779, n75934 );
nor U114467 ( n47486, n47487, n47488 );
nand U114468 ( n47487, n47403, n47491 );
nand U114469 ( n47488, n7502, n47489 );
nand U114470 ( n47491, n46331, n74400 );
nor U114471 ( n47425, n47426, n47427 );
nand U114472 ( n47427, n47428, n47429 );
nand U114473 ( n47426, n47446, n47447 );
nand U114474 ( n47429, n76657, n46182 );
nand U114475 ( n46486, n46492, n46493 );
nand U114476 ( n46493, n46365, n73220 );
nand U114477 ( n46492, n46332, n74919 );
nand U114478 ( n46778, n46779, n74550 );
nor U114479 ( n46775, n46776, n46777 );
nand U114480 ( n46776, n46781, n7508 );
nand U114481 ( n46777, n7472, n46778 );
nand U114482 ( n46781, n46331, n74524 );
nand U114483 ( n47258, n46779, n74659 );
nand U114484 ( n42524, n7409, n43352 );
nand U114485 ( n43352, n43353, n43354 );
nand U114486 ( n43354, n43355, n7619 );
nand U114487 ( n43353, n7617, n43356 );
nor U114488 ( n42484, n42493, n74992 );
nor U114489 ( n42493, n42494, n500 );
nor U114490 ( n42494, n42495, n42496 );
nand U114491 ( n42496, n42497, n75220 );
nor U114492 ( n42578, n42553, n42579 );
nor U114493 ( n42579, n42580, n42581 );
nor U114494 ( n42580, n42582, n42583 );
nand U114495 ( n47130, n46779, n74734 );
nor U114496 ( n16623, n17080, n76788 );
nand U114497 ( n8428, n4764, n9407 );
nand U114498 ( n9407, n9408, n9409 );
nand U114499 ( n9409, n9410, n4965 );
nand U114500 ( n9408, n4963, n9412 );
nand U114501 ( n12764, n12880, n12775 );
nor U114502 ( n12757, n12760, n73279 );
nor U114503 ( n12760, n12762, n12763 );
nor U114504 ( n12762, n74946, n12764 );
nor U114505 ( n8394, n8405, n74985 );
nor U114506 ( n8405, n8407, n229 );
nor U114507 ( n8407, n8408, n8409 );
nand U114508 ( n8409, n8410, n75217 );
nor U114509 ( n46350, n46353, n74986 );
nor U114510 ( n46353, n46354, n46355 );
nor U114511 ( n46354, n74974, n46356 );
nand U114512 ( n12825, n12828, n74946 );
xor U114513 ( n9144, n74541, n12445 );
nor U114514 ( n13627, n13628, n13629 );
nand U114515 ( n13628, n13633, n13575 );
nand U114516 ( n13629, n4835, n13630 );
nand U114517 ( n13633, n12999, n73116 );
nand U114518 ( n13630, n13214, n74476 );
xor U114519 ( n12504, n13870, n13925 );
xor U114520 ( n13925, n74658, n13907 );
xor U114521 ( n67111, n68283, n68327 );
xor U114522 ( n68327, n74695, n68312 );
nand U114523 ( n13938, n13214, n73090 );
nor U114524 ( n13934, n13935, n13937 );
nand U114525 ( n13935, n13940, n13829 );
nand U114526 ( n13937, n4833, n13938 );
nand U114527 ( n13940, n12999, n74461 );
xor U114528 ( n25213, n26282, n26326 );
xor U114529 ( n26326, n74697, n26311 );
xor U114530 ( n58349, n59421, n59465 );
xor U114531 ( n59465, n74698, n59450 );
xor U114532 ( n46147, n47252, n47296 );
xor U114533 ( n47296, n74659, n47281 );
xor U114534 ( n32455, n33527, n33571 );
xor U114535 ( n33571, n74696, n33556 );
nor U114536 ( n14257, n14153, n14258 );
nand U114537 ( n14258, n14259, n14260 );
nand U114538 ( n14260, n12999, n14262 );
nand U114539 ( n14259, n13214, n74429 );
nor U114540 ( n14170, n14172, n14173 );
nand U114541 ( n14173, n14174, n14175 );
nand U114542 ( n14172, n14208, n14209 );
nand U114543 ( n14175, n76724, n12585 );
nand U114544 ( n13478, n13479, n13480 );
nand U114545 ( n13480, n12999, n73117 );
nand U114546 ( n13479, n13214, n74823 );
nor U114547 ( n33216, n33217, n33171 );
nor U114548 ( n33217, n33220, n74855 );
nor U114549 ( n33220, n33221, n33181 );
nor U114550 ( n33221, n73160, n33222 );
nor U114551 ( n22749, n22750, n75260 );
nor U114552 ( n22750, n3875, n21986 );
nor U114553 ( n55863, n55864, n75261 );
nor U114554 ( n55864, n6508, n55096 );
nor U114555 ( n30070, n30071, n75258 );
nor U114556 ( n30071, n3032, n29301 );
nor U114557 ( n64087, n64088, n75257 );
nor U114558 ( n64088, n5633, n63068 );
xor U114559 ( MUL_1421_A1_U5, n71002, n71003 );
nor U114560 ( n71002, n2360, n71023 );
xor U114561 ( n71003, n71004, n71005 );
nand U114562 ( n71023, n71000, n70997 );
not U114563 ( n2359, n71001 );
nor U114564 ( n67971, n67972, n67934 );
nor U114565 ( n67972, n67975, n74852 );
nor U114566 ( n67975, n67976, n67932 );
nor U114567 ( n67976, n74431, n67977 );
nor U114568 ( n46924, n46925, n46887 );
nor U114569 ( n46925, n46928, n74822 );
nor U114570 ( n46928, n46929, n46885 );
nor U114571 ( n46929, n74417, n46930 );
nor U114572 ( n25968, n25969, n25931 );
nor U114573 ( n25969, n25972, n74853 );
nor U114574 ( n25972, n25973, n25929 );
nor U114575 ( n25973, n74432, n25974 );
nor U114576 ( n59106, n59107, n59069 );
nor U114577 ( n59107, n59110, n74854 );
nor U114578 ( n59110, n59111, n59067 );
nor U114579 ( n59111, n74433, n59112 );
nor U114580 ( n13208, n13209, n13210 );
nand U114581 ( n13210, n13212, n13213 );
nand U114582 ( n13209, n13215, n13217 );
nand U114583 ( n13213, n12999, n75053 );
not U114584 ( n3077, n29193 );
xnor U114585 ( n37838, n37839, n37840 );
xor U114586 ( n37840, n74371, n37841 );
nor U114587 ( n32994, n32995, n32996 );
nand U114588 ( n32996, n32997, n32998 );
nand U114589 ( n32995, n32999, n33000 );
nand U114590 ( n32998, n76128, n75060 );
nor U114591 ( n67750, n67751, n67752 );
nand U114592 ( n67752, n67753, n67754 );
nand U114593 ( n67751, n67755, n67756 );
nand U114594 ( n67754, n76058, n75017 );
nor U114595 ( n25745, n25746, n25747 );
nand U114596 ( n25747, n25748, n25749 );
nand U114597 ( n25746, n25750, n25751 );
nand U114598 ( n25749, n76156, n75018 );
nor U114599 ( n58885, n58886, n58887 );
nand U114600 ( n58887, n58888, n58889 );
nand U114601 ( n58886, n58890, n58891 );
nand U114602 ( n58889, n76084, n75019 );
not U114603 ( n1220, n71018 );
nand U114604 ( n13212, n13214, n73158 );
not U114605 ( n3920, n21876 );
not U114606 ( n6553, n54967 );
xor U114607 ( n9219, n74506, n12513 );
not U114608 ( n5678, n62911 );
nor U114609 ( n33335, n33336, n33278 );
nor U114610 ( n33336, n33339, n74458 );
nor U114611 ( n33339, n33340, n33341 );
nor U114612 ( n33340, n33342, n33343 );
nor U114613 ( n68092, n68093, n68037 );
nor U114614 ( n68093, n68096, n74438 );
nor U114615 ( n68096, n68097, n68098 );
nor U114616 ( n68097, n68099, n68100 );
nor U114617 ( n47061, n47062, n47002 );
nor U114618 ( n47062, n47065, n74427 );
nor U114619 ( n47065, n47066, n47067 );
nor U114620 ( n47066, n47068, n47069 );
nor U114621 ( n26089, n26090, n26034 );
nor U114622 ( n26090, n26093, n74439 );
nor U114623 ( n26093, n26094, n26095 );
nor U114624 ( n26094, n26096, n26097 );
nor U114625 ( n59230, n59231, n59175 );
nor U114626 ( n59231, n59234, n74440 );
nor U114627 ( n59234, n59235, n59236 );
nor U114628 ( n59235, n59237, n59238 );
nor U114629 ( n47309, n47310, n47268 );
nor U114630 ( n47310, n47312, n73065 );
nor U114631 ( n47312, n47313, n47314 );
nor U114632 ( n47313, n47267, n47315 );
xnor U114633 ( n9024, n74644, n12328 );
nor U114634 ( n68340, n68341, n68342 );
nor U114635 ( n68342, n5714, n68202 );
nor U114636 ( n68341, n68344, n73066 );
nor U114637 ( n68344, n68345, n68346 );
nor U114638 ( n33584, n33585, n33586 );
nor U114639 ( n33586, n3113, n33451 );
nor U114640 ( n33585, n33588, n73088 );
nor U114641 ( n33588, n33589, n33590 );
nor U114642 ( n26339, n26340, n26341 );
nor U114643 ( n26341, n3957, n26201 );
nor U114644 ( n26340, n26343, n73067 );
nor U114645 ( n26343, n26344, n26345 );
nor U114646 ( n59478, n59479, n59480 );
nor U114647 ( n59480, n6589, n59340 );
nor U114648 ( n59479, n59482, n73068 );
nor U114649 ( n59482, n59483, n59484 );
nor U114650 ( n46703, n46704, n46705 );
nand U114651 ( n46705, n46706, n46707 );
nand U114652 ( n46704, n46708, n46709 );
nand U114653 ( n46707, n76101, n75020 );
xnor U114654 ( n8830, n74785, n12167 );
xor U114655 ( n9285, n74484, n12563 );
or U114656 ( n33331, n33333, n75850 );
and U114657 ( n75850, n32738, n74458 );
or U114658 ( n47057, n47059, n75851 );
and U114659 ( n75851, n46439, n74427 );
or U114660 ( n68088, n68090, n75852 );
and U114661 ( n75852, n67503, n74438 );
or U114662 ( n26085, n26087, n75853 );
and U114663 ( n75853, n25498, n74439 );
or U114664 ( n59226, n59228, n75854 );
and U114665 ( n75854, n58635, n74440 );
or U114666 ( n68336, n68338, n75855 );
and U114667 ( n75855, n67503, n73066 );
or U114668 ( n33580, n33582, n75856 );
and U114669 ( n75856, n32738, n73088 );
or U114670 ( n26335, n26337, n75857 );
and U114671 ( n75857, n25498, n73067 );
or U114672 ( n59474, n59476, n75858 );
and U114673 ( n75858, n58635, n73068 );
or U114674 ( n47305, n47307, n75859 );
and U114675 ( n75859, n46439, n73065 );
nor U114676 ( n68687, n68688, n68689 );
nand U114677 ( n68688, n68715, n68716 );
nand U114678 ( n68689, n68690, n68691 );
nand U114679 ( n68716, n5704, n67203 );
nor U114680 ( n33931, n33932, n33933 );
nand U114681 ( n33932, n33959, n33960 );
nand U114682 ( n33933, n33934, n33935 );
nand U114683 ( n33960, n3103, n32547 );
nor U114684 ( n26686, n26687, n26688 );
nand U114685 ( n26687, n26714, n26715 );
nand U114686 ( n26688, n26689, n26690 );
nand U114687 ( n26715, n3947, n25305 );
nor U114688 ( n59828, n59829, n59830 );
nand U114689 ( n59829, n59856, n59857 );
nand U114690 ( n59830, n59831, n59832 );
nand U114691 ( n59857, n6579, n58444 );
xor U114692 ( n22041, n24729, n74850 );
xor U114693 ( n29360, n31961, n74849 );
xor U114694 ( n63123, n66564, n74848 );
xor U114695 ( n55151, n57863, n74851 );
nor U114696 ( n42575, n75014, n42577 );
nor U114697 ( n68594, n68511, n68595 );
nand U114698 ( n68595, n68596, n68597 );
nand U114699 ( n68597, n76057, n68598 );
nand U114700 ( n68596, n67503, n74408 );
nor U114701 ( n33838, n33755, n33839 );
nand U114702 ( n33839, n33840, n33841 );
nand U114703 ( n33841, n76127, n33842 );
nand U114704 ( n33840, n32738, n74412 );
nor U114705 ( n47573, n47490, n47574 );
nand U114706 ( n47574, n47575, n47576 );
nand U114707 ( n47576, n76100, n47577 );
nand U114708 ( n47575, n46439, n74400 );
nor U114709 ( n26593, n26510, n26594 );
nand U114710 ( n26594, n26595, n26596 );
nand U114711 ( n26596, n76155, n26597 );
nand U114712 ( n26595, n25498, n74409 );
nor U114713 ( n59735, n59649, n59736 );
nand U114714 ( n59736, n59737, n59738 );
nand U114715 ( n59738, n76083, n59739 );
nand U114716 ( n59737, n58635, n74410 );
nor U114717 ( n47504, n47505, n47506 );
nand U114718 ( n47506, n47507, n47508 );
nand U114719 ( n47505, n47534, n47535 );
nand U114720 ( n47508, n76657, n46212 );
nor U114721 ( n68525, n68526, n68527 );
nand U114722 ( n68527, n68528, n68529 );
nand U114723 ( n68526, n68555, n68556 );
nand U114724 ( n68529, n76705, n67176 );
nor U114725 ( n33769, n33770, n33771 );
nand U114726 ( n33771, n33772, n33773 );
nand U114727 ( n33770, n33799, n33800 );
nand U114728 ( n33773, n76772, n32520 );
nor U114729 ( n26524, n26525, n26526 );
nand U114730 ( n26526, n26527, n26528 );
nand U114731 ( n26525, n26554, n26555 );
nand U114732 ( n26528, n76751, n25278 );
nor U114733 ( n59666, n59667, n59668 );
nand U114734 ( n59668, n59669, n59670 );
nand U114735 ( n59667, n59696, n59697 );
nand U114736 ( n59670, n76684, n58414 );
nand U114737 ( n67966, n67967, n67968 );
nand U114738 ( n67968, n67502, n74431 );
nand U114739 ( n67967, n67503, n74852 );
nand U114740 ( n46919, n46920, n46921 );
nand U114741 ( n46921, n46438, n74417 );
nand U114742 ( n46920, n46439, n74822 );
nand U114743 ( n25963, n25964, n25965 );
nand U114744 ( n25965, n25497, n74432 );
nand U114745 ( n25964, n25498, n74853 );
nand U114746 ( n59101, n59102, n59103 );
nand U114747 ( n59103, n58634, n74433 );
nand U114748 ( n59102, n58635, n74854 );
xnor U114749 ( n63730, n74616, n66951 );
xnor U114750 ( n29770, n74615, n32312 );
xnor U114751 ( n22449, n74617, n25075 );
xnor U114752 ( n55564, n74618, n58210 );
nor U114753 ( n22011, n22012, n22013 );
nor U114754 ( n29330, n29331, n29332 );
nor U114755 ( n63093, n63094, n63095 );
nor U114756 ( n55121, n55122, n55123 );
nand U114757 ( n33211, n33212, n33213 );
nand U114758 ( n33213, n32737, n73160 );
nand U114759 ( n33212, n32738, n74855 );
not U114760 ( n5305, n8402 );
xor U114761 ( n63219, n66653, n74751 );
xor U114762 ( n29456, n32050, n74752 );
xor U114763 ( n22137, n24818, n74753 );
xor U114764 ( n55247, n57952, n74754 );
xor U114765 ( n63342, n66684, n74687 );
xor U114766 ( n29513, n32081, n74688 );
xor U114767 ( n22194, n24849, n74689 );
xor U114768 ( n55308, n57983, n74690 );
xor U114769 ( n63168, n66618, n74805 );
xor U114770 ( n29405, n32015, n74804 );
xor U114771 ( n22086, n24783, n74806 );
xor U114772 ( n55196, n57917, n74807 );
nor U114773 ( n54987, n842, n41466 );
nand U114774 ( n41970, n41449, n41972 );
nor U114775 ( n68460, n68368, n68462 );
nor U114776 ( n68462, n68375, n5807 );
nor U114777 ( n47439, n47336, n47441 );
nor U114778 ( n47441, n47343, n7594 );
nor U114779 ( n26459, n26367, n26461 );
nor U114780 ( n26461, n26374, n4040 );
nor U114781 ( n59598, n59506, n59600 );
nor U114782 ( n59600, n59513, n6673 );
nor U114783 ( n33704, n33612, n33706 );
nor U114784 ( n33706, n33619, n3208 );
nor U114785 ( n14089, n13968, n14092 );
nor U114786 ( n14092, n13977, n4940 );
nor U114787 ( n8507, n75015, n8509 );
nor U114788 ( n33415, n33419, n3118 );
nor U114789 ( n68165, n68169, n5719 );
nor U114790 ( n47134, n47138, n7505 );
nor U114791 ( n26164, n26168, n3962 );
nor U114792 ( n59303, n59307, n6594 );
nand U114793 ( n32997, n32738, n73167 );
nor U114794 ( n14382, n14383, n14384 );
nand U114795 ( n14383, n14417, n14418 );
nand U114796 ( n14384, n14385, n14387 );
nand U114797 ( n14418, n4848, n12619 );
nand U114798 ( n67753, n67503, n73149 );
nand U114799 ( n46706, n46439, n73148 );
nand U114800 ( n25748, n25498, n73150 );
nand U114801 ( n58888, n58635, n73151 );
nor U114802 ( n46631, n46587, n46664 );
nor U114803 ( n46664, n46665, n74585 );
nor U114804 ( n46629, n46631, n73159 );
nor U114805 ( n67678, n67636, n67711 );
nor U114806 ( n67711, n67712, n74595 );
nor U114807 ( n25673, n25631, n25706 );
nor U114808 ( n25706, n25707, n74596 );
nor U114809 ( n58813, n58768, n58846 );
nor U114810 ( n58846, n58847, n74597 );
nor U114811 ( n67676, n67678, n74637 );
nor U114812 ( n25671, n25673, n74638 );
nor U114813 ( n58811, n58813, n74639 );
nor U114814 ( n32917, n32875, n32957 );
nor U114815 ( n32957, n32958, n74652 );
nor U114816 ( n32915, n32917, n75050 );
nor U114817 ( n33140, n33143, n74879 );
nor U114818 ( n67896, n67899, n74872 );
nor U114819 ( n46849, n46852, n74841 );
nor U114820 ( n25893, n25896, n74873 );
nor U114821 ( n59031, n59034, n74874 );
nand U114822 ( n43256, n43308, n7967 );
not U114823 ( n7967, n43309 );
nor U114824 ( n68762, n68763, n68764 );
nand U114825 ( n68764, n68765, n68766 );
nand U114826 ( n68763, n68800, n68801 );
nand U114827 ( n68766, n67326, n68767 );
nor U114828 ( n34006, n34007, n34008 );
nand U114829 ( n34008, n34009, n34010 );
nand U114830 ( n34007, n34044, n34045 );
nand U114831 ( n34010, n32561, n34011 );
nor U114832 ( n26763, n26764, n26765 );
nand U114833 ( n26765, n26766, n26767 );
nand U114834 ( n26764, n26801, n26802 );
nand U114835 ( n26767, n25319, n26768 );
nor U114836 ( n59903, n59904, n59905 );
nand U114837 ( n59905, n59906, n59907 );
nand U114838 ( n59904, n59941, n59942 );
nand U114839 ( n59907, n58458, n59908 );
nand U114840 ( n21336, n21324, n5159 );
not U114841 ( n5159, n21337 );
nor U114842 ( n47666, n47667, n47668 );
nand U114843 ( n47667, n47694, n47695 );
nand U114844 ( n47668, n47669, n47670 );
nand U114845 ( n47695, n7490, n46251 );
nand U114846 ( n63941, n64054, n6178 );
nand U114847 ( n29985, n30037, n3563 );
nand U114848 ( n22662, n22714, n4400 );
nand U114849 ( n55775, n55830, n7033 );
not U114850 ( n6178, n64055 );
not U114851 ( n3563, n30038 );
not U114852 ( n4400, n22715 );
not U114853 ( n7033, n55831 );
nor U114854 ( n33093, n33033, n3123 );
nor U114855 ( n67849, n67788, n5723 );
nor U114856 ( n46802, n46741, n7509 );
nor U114857 ( n25846, n25785, n3965 );
nor U114858 ( n58984, n58923, n6598 );
nand U114859 ( n37607, n37080, n37609 );
nor U114860 ( n37602, n37604, n37605 );
nor U114861 ( n37605, n2198, n2083 );
nor U114862 ( n37604, n37606, n37091 );
nor U114863 ( n37606, n37607, n37608 );
nor U114864 ( n12932, n12945, n12947 );
and U114865 ( n12947, n72970, n12895 );
nor U114866 ( n12945, n12953, n12915 );
nor U114867 ( n13733, n13738, n4859 );
nand U114868 ( n54319, n54307, n7814 );
not U114869 ( n7814, n54320 );
nor U114870 ( n47741, n47742, n47743 );
nand U114871 ( n47743, n47744, n47745 );
nand U114872 ( n47742, n47779, n47780 );
nand U114873 ( n47745, n46265, n47746 );
or U114874 ( n67495, n5689, n67474 );
or U114875 ( n32730, n3088, n32709 );
or U114876 ( n25490, n3932, n25469 );
or U114877 ( n58627, n6564, n58606 );
nor U114878 ( n13330, n13258, n4864 );
nand U114879 ( n67499, n67500, n67501 );
nand U114880 ( n67501, n76057, n74947 );
nand U114881 ( n67500, n67503, n74962 );
nand U114882 ( n32734, n32735, n32736 );
nand U114883 ( n32736, n76127, n74948 );
nand U114884 ( n32735, n32738, n74961 );
nand U114885 ( n25494, n25495, n25496 );
nand U114886 ( n25496, n76155, n74949 );
nand U114887 ( n25495, n25498, n74960 );
nand U114888 ( n58631, n58632, n58633 );
nand U114889 ( n58633, n76083, n74950 );
nand U114890 ( n58632, n58635, n74963 );
nand U114891 ( n46435, n46436, n46437 );
nand U114892 ( n46437, n76100, n74919 );
nand U114893 ( n46436, n46439, n74930 );
nor U114894 ( n42624, n7925, n42625 );
nor U114895 ( n42625, n42626, n42627 );
nor U114896 ( n42626, n42628, n42629 );
nor U114897 ( n8568, n5270, n8569 );
nor U114898 ( n8569, n8570, n8572 );
nor U114899 ( n8570, n8573, n8574 );
nor U114900 ( n11809, n11813, n11845 );
nor U114901 ( n45566, n45569, n45592 );
nor U114902 ( n45656, n45658, n45681 );
nor U114903 ( n11909, n11912, n11945 );
nor U114904 ( n12000, n12003, n12032 );
nor U114905 ( n45733, n45735, n45776 );
nor U114906 ( n45558, n75077, n7963 );
not U114907 ( n7963, n45566 );
nor U114908 ( n11799, n75170, n5308 );
not U114909 ( n5308, n11809 );
nand U114910 ( n42572, n76102, n75014 );
nand U114911 ( n43008, n76102, n74815 );
nand U114912 ( n43164, n76102, n74728 );
nand U114913 ( n42839, n76102, n74914 );
nand U114914 ( n42754, n76102, n74958 );
not U114915 ( n6323, n63109 );
not U114916 ( n3689, n29346 );
not U114917 ( n4583, n22027 );
not U114918 ( n7215, n55137 );
not U114919 ( n6324, n63174 );
not U114920 ( n6325, n63225 );
not U114921 ( n6327, n63328 );
not U114922 ( n6328, n63466 );
not U114923 ( n6329, n63507 );
not U114924 ( n6330, n63563 );
not U114925 ( n6332, n63609 );
not U114926 ( n6333, n63723 );
not U114927 ( n6334, n63781 );
not U114928 ( n6335, n63833 );
not U114929 ( n6337, n63879 );
not U114930 ( n6338, n63929 );
not U114931 ( n3690, n29411 );
not U114932 ( n3692, n29462 );
not U114933 ( n3693, n29499 );
not U114934 ( n3694, n29563 );
not U114935 ( n3695, n29608 );
not U114936 ( n3697, n29664 );
not U114937 ( n3698, n29710 );
not U114938 ( n3699, n29763 );
not U114939 ( n3700, n29821 );
not U114940 ( n3702, n29877 );
not U114941 ( n3703, n29923 );
not U114942 ( n3704, n29973 );
not U114943 ( n4587, n22180 );
not U114944 ( n4594, n22502 );
not U114945 ( n4584, n22092 );
not U114946 ( n4585, n22143 );
not U114947 ( n4588, n22246 );
not U114948 ( n4589, n22287 );
not U114949 ( n4590, n22343 );
not U114950 ( n4592, n22389 );
not U114951 ( n4593, n22442 );
not U114952 ( n4595, n22554 );
not U114953 ( n4597, n22600 );
not U114954 ( n4598, n22650 );
not U114955 ( n7219, n55294 );
not U114956 ( n7227, n55615 );
not U114957 ( n7230, n55763 );
not U114958 ( n7217, n55202 );
not U114959 ( n7218, n55253 );
not U114960 ( n7220, n55358 );
not U114961 ( n7222, n55399 );
not U114962 ( n7223, n55455 );
not U114963 ( n7224, n55501 );
not U114964 ( n7225, n55557 );
not U114965 ( n7228, n55667 );
not U114966 ( n7229, n55713 );
and U114967 ( n21952, n22009, n75183 );
and U114968 ( n29269, n29328, n75181 );
and U114969 ( n63036, n63091, n75182 );
and U114970 ( n55064, n55119, n75184 );
nand U114971 ( n43248, n76102, n72964 );
nand U114972 ( n63035, n63036, n75214 );
nand U114973 ( n29268, n29269, n75213 );
nand U114974 ( n21951, n21952, n75215 );
nand U114975 ( n55063, n55064, n75216 );
nand U114976 ( n42663, n76102, n75005 );
nor U114977 ( n12933, n12934, n12935 );
and U114978 ( n12935, n12733, n12913 );
nor U114979 ( n12934, n12937, n72970 );
nor U114980 ( n12937, n12938, n12939 );
nand U114981 ( n8503, n76172, n75015 );
nor U114982 ( n68463, n68375, n68465 );
nor U114983 ( n68465, n68368, n68466 );
nor U114984 ( n47442, n47343, n47444 );
nor U114985 ( n47444, n47336, n47445 );
nor U114986 ( n26462, n26374, n26464 );
nor U114987 ( n26464, n26367, n26465 );
nor U114988 ( n59601, n59513, n59603 );
nor U114989 ( n59603, n59506, n59604 );
nand U114990 ( n8995, n76172, n74816 );
nand U114991 ( n9190, n76172, n74729 );
nand U114992 ( n8802, n76172, n74915 );
nor U114993 ( n33707, n33619, n33709 );
nor U114994 ( n33709, n33612, n33710 );
nor U114995 ( n14093, n13977, n14095 );
nor U114996 ( n14095, n13968, n14097 );
nand U114997 ( n8695, n76172, n74959 );
nor U114998 ( n40336, n2042, n37300 );
nand U114999 ( n9278, n76172, n72965 );
nand U115000 ( n8617, n76172, n75006 );
nor U115001 ( n14475, n14477, n14478 );
nand U115002 ( n14478, n14479, n14480 );
nand U115003 ( n14477, n14523, n14524 );
nand U115004 ( n14480, n12637, n14482 );
nor U115005 ( n66491, n66494, n66517 );
nor U115006 ( n31868, n31871, n31894 );
nor U115007 ( n24654, n24657, n24682 );
nor U115008 ( n57790, n57793, n57816 );
nor U115009 ( n66659, n66661, n66684 );
nor U115010 ( n32056, n32058, n32081 );
nor U115011 ( n24824, n24826, n24849 );
nor U115012 ( n57958, n57960, n57983 );
nor U115013 ( n66580, n66582, n66605 );
nor U115014 ( n31977, n31979, n32002 );
nor U115015 ( n24745, n24747, n24770 );
nor U115016 ( n57879, n57881, n57904 );
nor U115017 ( n32649, n32652, n75010 );
nor U115018 ( n32652, n32653, n32654 );
nor U115019 ( n32653, n74973, n32655 );
nor U115020 ( n25409, n25412, n75007 );
nor U115021 ( n25412, n25413, n25414 );
nor U115022 ( n25413, n74975, n25415 );
nor U115023 ( n67414, n67417, n75009 );
nor U115024 ( n67417, n67418, n67419 );
nor U115025 ( n67418, n74976, n67420 );
nor U115026 ( n58546, n58549, n75008 );
nor U115027 ( n58549, n58550, n58551 );
nor U115028 ( n58550, n74977, n58552 );
nor U115029 ( n24646, n74910, n4397 );
not U115030 ( n4397, n24654 );
nor U115031 ( n57782, n74911, n7029 );
not U115032 ( n7029, n57790 );
nor U115033 ( n31860, n74912, n3559 );
not U115034 ( n3559, n31868 );
nor U115035 ( n66483, n74913, n6174 );
not U115036 ( n6174, n66491 );
nand U115037 ( n65905, n66159, n66160 );
nand U115038 ( n66159, n5679, n74593 );
nand U115039 ( n66160, n66161, n5700 );
nor U115040 ( n66161, n62911, n66162 );
nand U115041 ( n57446, n57583, n57584 );
nand U115042 ( n57583, n6554, n74594 );
nand U115043 ( n57584, n57585, n6575 );
nor U115044 ( n57585, n54967, n57586 );
nand U115045 ( n65910, n65905, n74593 );
nand U115046 ( n57451, n57446, n74594 );
nand U115047 ( n41490, n41460, n76925 );
nand U115048 ( n9288, n9353, n5312 );
not U115049 ( n5312, n9354 );
nand U115050 ( n24323, n24457, n24458 );
nand U115051 ( n24457, n3922, n74592 );
nand U115052 ( n24458, n24459, n3943 );
nor U115053 ( n24459, n21876, n24460 );
nand U115054 ( n70997, n71001, n71018 );
nand U115055 ( n24328, n24323, n74592 );
nor U115056 ( n22037, n22012, n22038 );
nor U115057 ( n22038, n22039, n4394 );
not U115058 ( n4394, n22040 );
nor U115059 ( n22039, n22041, n22042 );
nor U115060 ( n29356, n29331, n29357 );
nor U115061 ( n29357, n29358, n3557 );
not U115062 ( n3557, n29359 );
nor U115063 ( n29358, n29360, n29361 );
nor U115064 ( n63119, n63094, n63120 );
nor U115065 ( n63120, n63121, n6172 );
not U115066 ( n6172, n63122 );
nor U115067 ( n63121, n63123, n63124 );
nor U115068 ( n55147, n55122, n55148 );
nor U115069 ( n55148, n55149, n7027 );
not U115070 ( n7027, n55150 );
nor U115071 ( n55149, n55151, n55152 );
xnor U115072 ( n67126, n68316, n68357 );
xnor U115073 ( n46162, n47285, n47325 );
xnor U115074 ( n25228, n26315, n26356 );
xnor U115075 ( n58364, n59454, n59495 );
xnor U115076 ( n32470, n33560, n33601 );
not U115077 ( n8104, n42568 );
not U115078 ( n5453, n8644 );
not U115079 ( n5454, n8690 );
not U115080 ( n5458, n8892 );
not U115081 ( n5459, n8949 );
not U115082 ( n5460, n9015 );
not U115083 ( n5462, n9088 );
not U115084 ( n5465, n9273 );
not U115085 ( n8108, n42750 );
not U115086 ( n8112, n42911 );
not U115087 ( n8113, n42971 );
not U115088 ( n8114, n43024 );
not U115089 ( n8115, n43082 );
not U115090 ( n8119, n43244 );
not U115091 ( n8105, n42634 );
not U115092 ( n8107, n42709 );
not U115093 ( n8109, n42814 );
not U115094 ( n8110, n42855 );
not U115095 ( n5450, n8498 );
not U115096 ( n5452, n8580 );
not U115097 ( n5455, n8770 );
not U115098 ( n5457, n8822 );
not U115099 ( n8117, n43134 );
not U115100 ( n8118, n43180 );
not U115101 ( n5463, n9153 );
not U115102 ( n5464, n9210 );
and U115103 ( n42497, n42550, n75190 );
not U115104 ( n865, n43866 );
nand U115105 ( n45317, n45320, n45321 );
nand U115106 ( n45320, n7464, n74648 );
nand U115107 ( n45321, n45322, n7487 );
nor U115108 ( n45322, n42402, n43348 );
nand U115109 ( n45161, n45164, n45155 );
nand U115110 ( n45164, n864, n74396 );
nand U115111 ( n45155, n865, n74401 );
nand U115112 ( n45025, n45317, n74648 );
xor U115113 ( n63515, n66845, n74563 );
xor U115114 ( n29616, n32199, n74564 );
xor U115115 ( n22295, n24969, n74565 );
xor U115116 ( n55407, n58104, n74566 );
xnor U115117 ( n12538, n13912, n13978 );
xor U115118 ( n8832, n12184, n74512 );
nor U115119 ( n43342, n43343, n75259 );
nor U115120 ( n43343, n7407, n42527 );
nand U115121 ( n45226, n45229, n45220 );
nand U115122 ( n45229, n864, n74397 );
nand U115123 ( n45220, n865, n74406 );
xnor U115124 ( n12522, n13978, n13929 );
xnor U115125 ( n67125, n68357, n68330 );
xnor U115126 ( n46161, n47325, n47299 );
xnor U115127 ( n25227, n26356, n26329 );
xnor U115128 ( n58363, n59495, n59468 );
xnor U115129 ( n32469, n33601, n33574 );
nand U115130 ( n67592, n67593, n74947 );
nand U115131 ( n67593, n67563, n67594 );
nand U115132 ( n67594, n5729, n6124 );
nand U115133 ( n32827, n32828, n74948 );
nand U115134 ( n32828, n32798, n32829 );
nand U115135 ( n32829, n3128, n3509 );
nand U115136 ( n25587, n25588, n74949 );
nand U115137 ( n25588, n25558, n25589 );
nand U115138 ( n25589, n3972, n4347 );
nand U115139 ( n58724, n58725, n74950 );
nand U115140 ( n58725, n58695, n58726 );
nand U115141 ( n58726, n6604, n6979 );
nand U115142 ( n13773, n13774, n5224 );
nor U115143 ( n13774, n4832, n73176 );
nand U115144 ( n11494, n11498, n11499 );
nand U115145 ( n11498, n4820, n74649 );
nand U115146 ( n11499, n11500, n4844 );
nor U115147 ( n11500, n8319, n9402 );
nand U115148 ( n11324, n11494, n74649 );
nand U115149 ( n12818, n12775, n5220 );
not U115150 ( n5220, n12880 );
xnor U115151 ( n63042, n66455, n75188 );
xnor U115152 ( n29275, n31832, n75185 );
xnor U115153 ( n21958, n24618, n75186 );
xnor U115154 ( n55070, n57750, n75187 );
nand U115155 ( n12752, n12735, n74989 );
and U115156 ( n16463, n18706, n76591 );
nor U115157 ( n18706, n18707, n18708 );
nor U115158 ( n18708, n5195, n4813 );
nor U115159 ( n18707, n18710, n18711 );
not U115160 ( n5204, n14705 );
nand U115161 ( n15390, n5193, n15273 );
nand U115162 ( n15272, n14735, n14739 );
nor U115163 ( n18703, n18704, n18705 );
nor U115164 ( n18704, n14934, n18709 );
nor U115165 ( n18705, n16463, n74361 );
nand U115166 ( n46345, n46334, n75016 );
nand U115167 ( n25404, n25393, n75038 );
nand U115168 ( n58541, n58530, n75040 );
nand U115169 ( n32644, n32633, n75042 );
nand U115170 ( n67409, n67398, n75039 );
nand U115171 ( n53885, n74442, n7863 );
nor U115172 ( n48130, n47908, n48711 );
nand U115173 ( n48718, n48780, n76325 );
nor U115174 ( n48780, n48781, n48782 );
nor U115175 ( n48782, n7849, n7457 );
nor U115176 ( n48781, n48783, n48779 );
nor U115177 ( n42209, n73633, n73024 );
xor U115178 ( U154, n70998, n70999 );
and U115179 ( n70998, n71000, n71001 );
nor U115180 ( n70999, n2360, n1220 );
nand U115181 ( n13147, n13148, n74920 );
nand U115182 ( n13148, n13103, n13149 );
nand U115183 ( n13149, n13150, n4867 );
nor U115184 ( n13150, n74625, n73158 );
not U115185 ( n864, n43666 );
nand U115186 ( n8457, n8435, n73392 );
nor U115187 ( n33280, n33281, n33282 );
nor U115188 ( n33281, n3119, n33289 );
nor U115189 ( n33282, n33283, n73160 );
or U115190 ( n33289, n33271, n74458 );
nor U115191 ( n47004, n47005, n47006 );
nor U115192 ( n47005, n7507, n47013 );
nor U115193 ( n47006, n47007, n74417 );
or U115194 ( n47013, n46995, n74427 );
nor U115195 ( n68039, n68040, n68041 );
nor U115196 ( n68040, n5720, n68048 );
nor U115197 ( n68041, n68042, n74431 );
or U115198 ( n68048, n68030, n74438 );
nor U115199 ( n26036, n26037, n26038 );
nor U115200 ( n26037, n3963, n26045 );
nor U115201 ( n26038, n26039, n74432 );
or U115202 ( n26045, n26027, n74439 );
nor U115203 ( n59177, n59178, n59179 );
nor U115204 ( n59178, n6595, n59186 );
nor U115205 ( n59179, n59180, n74433 );
or U115206 ( n59186, n59168, n74440 );
nand U115207 ( n63951, n5632, n63952 );
nand U115208 ( n63952, n63953, n74613 );
nand U115209 ( n29995, n3030, n29996 );
nand U115210 ( n29996, n29997, n74611 );
nand U115211 ( n22672, n3874, n22673 );
nand U115212 ( n22673, n22674, n74612 );
nand U115213 ( n55785, n6507, n55786 );
nand U115214 ( n55786, n55787, n74614 );
not U115215 ( n167, n21858 );
and U115216 ( n8320, n8270, n21166 );
nand U115217 ( n21166, n21167, n8297 );
nand U115218 ( n21167, n21168, n21169 );
nand U115219 ( n21169, n4964, n14654 );
not U115220 ( n2360, n71024 );
not U115221 ( n2, n11595 );
xnor U115222 ( n67145, n68469, n68382 );
xor U115223 ( n68469, n68381, n74452 );
xnor U115224 ( n12547, n14100, n13993 );
xor U115225 ( n14100, n13992, n74461 );
xnor U115226 ( n46181, n47448, n47350 );
xor U115227 ( n47448, n47349, n74443 );
xnor U115228 ( n25247, n26468, n26381 );
xor U115229 ( n26468, n26380, n74453 );
xnor U115230 ( n58383, n59607, n59520 );
xor U115231 ( n59607, n59519, n74454 );
xnor U115232 ( n32489, n33713, n33626 );
xor U115233 ( n33713, n33625, n74455 );
nand U115234 ( n49280, n49346, n47920 );
nor U115235 ( n49346, n7833, n7855 );
nand U115236 ( n15827, n15917, n14690 );
nand U115237 ( n16039, n15917, n14717 );
nand U115238 ( n67177, n68539, n68540 );
nand U115239 ( n68539, n68543, n68466 );
nand U115240 ( n68540, n68541, n5807 );
or U115241 ( n68543, n68368, n68375 );
nand U115242 ( n46213, n47518, n47519 );
nand U115243 ( n47518, n47522, n47445 );
nand U115244 ( n47519, n47520, n7594 );
or U115245 ( n47522, n47336, n47343 );
nand U115246 ( n25279, n26538, n26539 );
nand U115247 ( n26538, n26542, n26465 );
nand U115248 ( n26539, n26540, n4040 );
or U115249 ( n26542, n26367, n26374 );
nand U115250 ( n58415, n59680, n59681 );
nand U115251 ( n59680, n59684, n59604 );
nand U115252 ( n59681, n59682, n6673 );
or U115253 ( n59684, n59506, n59513 );
nand U115254 ( n32521, n33783, n33784 );
nand U115255 ( n33783, n33787, n33710 );
nand U115256 ( n33784, n33785, n3208 );
or U115257 ( n33787, n33612, n33619 );
nand U115258 ( n12587, n14188, n14189 );
nand U115259 ( n14188, n14193, n14097 );
nand U115260 ( n14189, n14190, n4940 );
or U115261 ( n14193, n13968, n13977 );
nand U115262 ( n16242, n16332, n14690 );
nor U115263 ( n16332, n5178, n5200 );
and U115264 ( n29194, n29150, n35651 );
nand U115265 ( n35651, n35652, n29171 );
nand U115266 ( n35652, n35653, n35654 );
nand U115267 ( n35654, n3232, n34150 );
and U115268 ( n21877, n21835, n28472 );
nand U115269 ( n28472, n28473, n21858 );
nand U115270 ( n28473, n28474, n28475 );
nand U115271 ( n28475, n4059, n26905 );
and U115272 ( n62912, n62817, n70377 );
nand U115273 ( n70377, n70378, n62893 );
nand U115274 ( n70378, n70379, n70380 );
nand U115275 ( n70380, n5830, n68904 );
and U115276 ( n54968, n54928, n61777 );
nand U115277 ( n61777, n61778, n54949 );
nand U115278 ( n61778, n61779, n61780 );
nand U115279 ( n61780, n6692, n60045 );
nand U115280 ( n46583, n46584, n73220 );
nand U115281 ( n46584, n7499, n46585 );
nand U115282 ( n46585, n46586, n46587 );
not U115283 ( n7499, n46534 );
not U115284 ( n439, n54949 );
nand U115285 ( n13689, n13734, n13735 );
nand U115286 ( n13735, n5223, n12999 );
or U115287 ( n13734, n13739, n74735 );
nand U115288 ( n68130, n68166, n68167 );
nand U115289 ( n68167, n6088, n67502 );
or U115290 ( n68166, n68170, n74758 );
nand U115291 ( n33378, n33416, n33417 );
nand U115292 ( n33417, n3473, n32737 );
or U115293 ( n33416, n33420, n73115 );
nand U115294 ( n47099, n47135, n47136 );
nand U115295 ( n47136, n7877, n46438 );
or U115296 ( n47135, n47139, n74734 );
nand U115297 ( n26127, n26165, n26166 );
nand U115298 ( n26166, n4310, n25497 );
or U115299 ( n26165, n26169, n74759 );
nand U115300 ( n59268, n59304, n59305 );
nand U115301 ( n59305, n6943, n58634 );
or U115302 ( n59304, n59308, n74760 );
nand U115303 ( n15710, n15797, n76591 );
nor U115304 ( n15797, n15798, n15799 );
nor U115305 ( n15799, n5198, n4813 );
nor U115306 ( n15798, n15802, n15803 );
nand U115307 ( n16129, n16213, n76591 );
nor U115308 ( n16213, n16214, n16215 );
nor U115309 ( n16215, n5197, n4813 );
nor U115310 ( n16214, n16218, n16219 );
nand U115311 ( n49179, n49241, n76325 );
nor U115312 ( n49241, n49242, n49243 );
nor U115313 ( n49243, n7852, n7457 );
nor U115314 ( n49242, n49245, n49246 );
nand U115315 ( n48810, n48872, n76325 );
nor U115316 ( n48872, n48873, n48874 );
nor U115317 ( n48874, n7853, n7457 );
nor U115318 ( n48873, n48876, n48877 );
nand U115319 ( n26989, P1_P2_STATE2_REG_3_, n74612 );
and U115320 ( n28286, n28395, n23824 );
and U115321 ( n26979, n74592, n28402 );
nand U115322 ( n28402, n28403, n26989 );
nand U115323 ( n28403, n27028, n21849 );
nor U115324 ( n13569, n13570, n13572 );
nor U115325 ( n13570, n4860, n13580 );
nor U115326 ( n13572, n13573, n73117 );
or U115327 ( n13580, n13558, n74476 );
nand U115328 ( n6181, n27693, n27694 );
nor U115329 ( n27693, n27707, n27708 );
nor U115330 ( n27694, n27695, n27696 );
nor U115331 ( n27707, n26970, n27128 );
nand U115332 ( n5901, n28262, n28263 );
nor U115333 ( n28263, n28264, n28265 );
nor U115334 ( n28262, n28275, n28276 );
nor U115335 ( n28264, n27133, n28205 );
nand U115336 ( n5941, n28181, n28182 );
nor U115337 ( n28182, n28183, n28184 );
nor U115338 ( n28181, n28194, n28195 );
nor U115339 ( n28183, n27133, n28124 );
nand U115340 ( n5981, n28099, n28100 );
nor U115341 ( n28100, n28101, n28102 );
nor U115342 ( n28099, n28113, n28114 );
nor U115343 ( n28101, n27128, n28042 );
nand U115344 ( n6021, n28019, n28020 );
nor U115345 ( n28020, n28021, n28022 );
nor U115346 ( n28019, n28032, n28033 );
nor U115347 ( n28021, n27133, n27966 );
nand U115348 ( n6061, n27937, n27938 );
nor U115349 ( n27938, n27939, n27940 );
nor U115350 ( n27937, n27950, n27951 );
nor U115351 ( n27939, n27133, n27884 );
nand U115352 ( n6101, n27859, n27860 );
nor U115353 ( n27860, n27861, n27862 );
nor U115354 ( n27859, n27872, n27873 );
nor U115355 ( n27861, n27133, n27802 );
nand U115356 ( n6141, n27776, n27777 );
nor U115357 ( n27777, n27778, n27779 );
nor U115358 ( n27776, n27790, n27791 );
nor U115359 ( n27778, n27128, n27717 );
nand U115360 ( n6221, n27616, n27617 );
nor U115361 ( n27617, n27618, n27619 );
nor U115362 ( n27616, n27629, n27630 );
nor U115363 ( n27618, n27133, n27563 );
nand U115364 ( n6261, n27536, n27537 );
nor U115365 ( n27537, n27538, n27539 );
nor U115366 ( n27536, n27550, n27551 );
nor U115367 ( n27538, n27133, n27477 );
nor U115368 ( n15804, n15273, n5193 );
nand U115369 ( n48896, n48983, n47920 );
nor U115370 ( n48983, n7833, n47935 );
nand U115371 ( n14468, n14469, n74579 );
nand U115372 ( n14469, n4832, n14367 );
nor U115373 ( n14417, n14462, n14463 );
nor U115374 ( n14463, n4864, n14464 );
nor U115375 ( n14462, n75059, n14468 );
nor U115376 ( n14464, n14465, n5219 );
and U115377 ( n42403, n42363, n54149 );
nand U115378 ( n54149, n54150, n42384 );
nand U115379 ( n54150, n54151, n54152 );
nand U115380 ( n54152, n7618, n47884 );
nand U115381 ( n6211, n27643, n27644 );
nor U115382 ( n27643, n27649, n27650 );
nor U115383 ( n27644, n27645, n27646 );
nor U115384 ( n27649, n26970, n27052 );
nand U115385 ( n6186, n27685, n27686 );
nor U115386 ( n27685, n27691, n27692 );
nor U115387 ( n27686, n27687, n27688 );
nor U115388 ( n27691, n26970, n27107 );
nand U115389 ( n6216, n27632, n27633 );
nor U115390 ( n27632, n27640, n27641 );
nor U115391 ( n27633, n27634, n27635 );
nor U115392 ( n27640, n26970, n27039 );
nand U115393 ( n6191, n27677, n27678 );
nor U115394 ( n27677, n27683, n27684 );
nor U115395 ( n27678, n27679, n27680 );
nor U115396 ( n27683, n26970, n27096 );
nand U115397 ( n6201, n27661, n27662 );
nor U115398 ( n27661, n27667, n27668 );
nor U115399 ( n27662, n27663, n27664 );
nor U115400 ( n27667, n26970, n27074 );
nand U115401 ( n6196, n27669, n27670 );
nor U115402 ( n27669, n27675, n27676 );
nor U115403 ( n27670, n27671, n27672 );
nor U115404 ( n27675, n26970, n27085 );
nand U115405 ( n6206, n27653, n27654 );
nor U115406 ( n27653, n27659, n27660 );
nor U115407 ( n27654, n27655, n27656 );
nor U115408 ( n27659, n26970, n27063 );
nand U115409 ( n60132, P2_P2_STATE2_REG_3_, n74614 );
and U115410 ( n61508, n61676, n31914 );
and U115411 ( n60119, n74594, n61711 );
nand U115412 ( n61711, n61712, n60132 );
nand U115413 ( n61712, n60169, n54940 );
nand U115414 ( n12926, n60828, n60829 );
nor U115415 ( n60828, n60834, n60835 );
nor U115416 ( n60829, n60830, n60831 );
nor U115417 ( n60834, n60110, n60240 );
nand U115418 ( n12936, n60812, n60813 );
nor U115419 ( n60812, n60818, n60819 );
nor U115420 ( n60813, n60814, n60815 );
nor U115421 ( n60818, n60110, n60215 );
nand U115422 ( n12921, n60836, n60837 );
nor U115423 ( n60836, n60842, n60843 );
nor U115424 ( n60837, n60838, n60839 );
nor U115425 ( n60842, n60110, n60251 );
nand U115426 ( n12946, n60796, n60797 );
nor U115427 ( n60796, n60802, n60803 );
nor U115428 ( n60797, n60798, n60799 );
nor U115429 ( n60802, n60110, n60193 );
nand U115430 ( n12951, n60785, n60786 );
nor U115431 ( n60785, n60793, n60794 );
nor U115432 ( n60786, n60787, n60788 );
nor U115433 ( n60793, n60110, n60180 );
nand U115434 ( n12941, n60804, n60805 );
nor U115435 ( n60804, n60810, n60811 );
nor U115436 ( n60805, n60806, n60807 );
nor U115437 ( n60810, n60110, n60204 );
nand U115438 ( n12931, n60820, n60821 );
nor U115439 ( n60820, n60826, n60827 );
nor U115440 ( n60821, n60822, n60823 );
nor U115441 ( n60826, n60110, n60226 );
nand U115442 ( n12916, n60844, n60845 );
nor U115443 ( n60844, n60858, n60859 );
nor U115444 ( n60845, n60846, n60847 );
nor U115445 ( n60858, n60110, n60272 );
nand U115446 ( n5986, n28091, n28092 );
nor U115447 ( n28092, n28093, n28094 );
nor U115448 ( n28091, n28097, n28098 );
nor U115449 ( n28093, n27107, n28042 );
nand U115450 ( n6146, n27768, n27769 );
nor U115451 ( n27769, n27770, n27771 );
nor U115452 ( n27768, n27774, n27775 );
nor U115453 ( n27770, n27107, n27717 );
nand U115454 ( n6016, n28034, n28035 );
nor U115455 ( n28035, n28036, n28037 );
nor U115456 ( n28034, n28043, n28044 );
nor U115457 ( n28036, n27039, n28042 );
nand U115458 ( n6176, n27709, n27710 );
nor U115459 ( n27710, n27711, n27712 );
nor U115460 ( n27709, n27718, n27719 );
nor U115461 ( n27711, n27039, n27717 );
nand U115462 ( n5991, n28083, n28084 );
nor U115463 ( n28084, n28085, n28086 );
nor U115464 ( n28083, n28089, n28090 );
nor U115465 ( n28085, n27096, n28042 );
nand U115466 ( n6151, n27760, n27761 );
nor U115467 ( n27761, n27762, n27763 );
nor U115468 ( n27760, n27766, n27767 );
nor U115469 ( n27762, n27096, n27717 );
nand U115470 ( n5921, n28226, n28227 );
nor U115471 ( n28227, n28228, n28229 );
nor U115472 ( n28226, n28232, n28233 );
nor U115473 ( n28228, n27077, n28205 );
nand U115474 ( n5961, n28145, n28146 );
nor U115475 ( n28146, n28147, n28148 );
nor U115476 ( n28145, n28151, n28152 );
nor U115477 ( n28147, n27077, n28124 );
nand U115478 ( n6041, n27987, n27988 );
nor U115479 ( n27988, n27989, n27990 );
nor U115480 ( n27987, n27993, n27994 );
nor U115481 ( n27989, n27077, n27966 );
nand U115482 ( n6081, n27905, n27906 );
nor U115483 ( n27906, n27907, n27908 );
nor U115484 ( n27905, n27911, n27912 );
nor U115485 ( n27907, n27077, n27884 );
nand U115486 ( n6121, n27823, n27824 );
nor U115487 ( n27824, n27825, n27826 );
nor U115488 ( n27823, n27829, n27830 );
nor U115489 ( n27825, n27077, n27802 );
nand U115490 ( n6241, n27584, n27585 );
nor U115491 ( n27585, n27586, n27587 );
nor U115492 ( n27584, n27590, n27591 );
nor U115493 ( n27586, n27077, n27563 );
nand U115494 ( n6281, n27500, n27501 );
nor U115495 ( n27501, n27502, n27503 );
nor U115496 ( n27500, n27507, n27508 );
nor U115497 ( n27502, n27077, n27477 );
nand U115498 ( n5926, n28218, n28219 );
nor U115499 ( n28219, n28220, n28221 );
nor U115500 ( n28218, n28224, n28225 );
nor U115501 ( n28220, n27066, n28205 );
nand U115502 ( n5966, n28137, n28138 );
nor U115503 ( n28138, n28139, n28140 );
nor U115504 ( n28137, n28143, n28144 );
nor U115505 ( n28139, n27066, n28124 );
nand U115506 ( n6046, n27979, n27980 );
nor U115507 ( n27980, n27981, n27982 );
nor U115508 ( n27979, n27985, n27986 );
nor U115509 ( n27981, n27066, n27966 );
nand U115510 ( n6086, n27897, n27898 );
nor U115511 ( n27898, n27899, n27900 );
nor U115512 ( n27897, n27903, n27904 );
nor U115513 ( n27899, n27066, n27884 );
nand U115514 ( n6126, n27815, n27816 );
nor U115515 ( n27816, n27817, n27818 );
nor U115516 ( n27815, n27821, n27822 );
nor U115517 ( n27817, n27066, n27802 );
nand U115518 ( n6246, n27576, n27577 );
nor U115519 ( n27577, n27578, n27579 );
nor U115520 ( n27576, n27582, n27583 );
nor U115521 ( n27578, n27066, n27563 );
nand U115522 ( n6286, n27491, n27492 );
nor U115523 ( n27492, n27493, n27494 );
nor U115524 ( n27491, n27498, n27499 );
nor U115525 ( n27493, n27066, n27477 );
nand U115526 ( n5951, n28165, n28166 );
nor U115527 ( n28166, n28167, n28168 );
nor U115528 ( n28165, n28171, n28172 );
nor U115529 ( n28167, n27099, n28124 );
nand U115530 ( n6031, n28003, n28004 );
nor U115531 ( n28004, n28005, n28006 );
nor U115532 ( n28003, n28009, n28010 );
nor U115533 ( n28005, n27099, n27966 );
nand U115534 ( n6071, n27921, n27922 );
nor U115535 ( n27922, n27923, n27924 );
nor U115536 ( n27921, n27927, n27928 );
nor U115537 ( n27923, n27099, n27884 );
nand U115538 ( n6111, n27839, n27840 );
nor U115539 ( n27840, n27841, n27842 );
nor U115540 ( n27839, n27845, n27846 );
nor U115541 ( n27841, n27099, n27802 );
nand U115542 ( n6231, n27600, n27601 );
nor U115543 ( n27601, n27602, n27603 );
nor U115544 ( n27600, n27606, n27607 );
nor U115545 ( n27602, n27099, n27563 );
nand U115546 ( n6271, n27518, n27519 );
nor U115547 ( n27519, n27520, n27521 );
nor U115548 ( n27518, n27525, n27526 );
nor U115549 ( n27520, n27099, n27477 );
nand U115550 ( n5911, n28242, n28243 );
nor U115551 ( n28243, n28244, n28245 );
nor U115552 ( n28242, n28248, n28249 );
nor U115553 ( n28244, n27099, n28205 );
nand U115554 ( n5971, n28129, n28130 );
nor U115555 ( n28130, n28131, n28132 );
nor U115556 ( n28129, n28135, n28136 );
nor U115557 ( n28131, n27055, n28124 );
nand U115558 ( n6051, n27971, n27972 );
nor U115559 ( n27972, n27973, n27974 );
nor U115560 ( n27971, n27977, n27978 );
nor U115561 ( n27973, n27055, n27966 );
nand U115562 ( n6091, n27889, n27890 );
nor U115563 ( n27890, n27891, n27892 );
nor U115564 ( n27889, n27895, n27896 );
nor U115565 ( n27891, n27055, n27884 );
nand U115566 ( n6131, n27807, n27808 );
nor U115567 ( n27808, n27809, n27810 );
nor U115568 ( n27807, n27813, n27814 );
nor U115569 ( n27809, n27055, n27802 );
nand U115570 ( n6251, n27568, n27569 );
nor U115571 ( n27569, n27570, n27571 );
nor U115572 ( n27568, n27574, n27575 );
nor U115573 ( n27570, n27055, n27563 );
nand U115574 ( n6291, n27482, n27483 );
nor U115575 ( n27483, n27484, n27485 );
nor U115576 ( n27482, n27489, n27490 );
nor U115577 ( n27484, n27055, n27477 );
nand U115578 ( n5916, n28234, n28235 );
nor U115579 ( n28235, n28236, n28237 );
nor U115580 ( n28234, n28240, n28241 );
nor U115581 ( n28236, n27088, n28205 );
nand U115582 ( n5956, n28157, n28158 );
nor U115583 ( n28158, n28159, n28160 );
nor U115584 ( n28157, n28163, n28164 );
nor U115585 ( n28159, n27088, n28124 );
nand U115586 ( n6036, n27995, n27996 );
nor U115587 ( n27996, n27997, n27998 );
nor U115588 ( n27995, n28001, n28002 );
nor U115589 ( n27997, n27088, n27966 );
nand U115590 ( n6076, n27913, n27914 );
nor U115591 ( n27914, n27915, n27916 );
nor U115592 ( n27913, n27919, n27920 );
nor U115593 ( n27915, n27088, n27884 );
nand U115594 ( n6116, n27831, n27832 );
nor U115595 ( n27832, n27833, n27834 );
nor U115596 ( n27831, n27837, n27838 );
nor U115597 ( n27833, n27088, n27802 );
nand U115598 ( n6236, n27592, n27593 );
nor U115599 ( n27593, n27594, n27595 );
nor U115600 ( n27592, n27598, n27599 );
nor U115601 ( n27594, n27088, n27563 );
nand U115602 ( n6276, n27509, n27510 );
nor U115603 ( n27510, n27511, n27512 );
nor U115604 ( n27509, n27516, n27517 );
nor U115605 ( n27511, n27088, n27477 );
nand U115606 ( n5931, n28210, n28211 );
nor U115607 ( n28211, n28212, n28213 );
nor U115608 ( n28210, n28216, n28217 );
nor U115609 ( n28212, n27055, n28205 );
nand U115610 ( n12726, n61238, n61239 );
nor U115611 ( n61239, n61240, n61241 );
nor U115612 ( n61238, n61244, n61245 );
nor U115613 ( n61240, n60240, n61201 );
nand U115614 ( n12886, n60908, n60909 );
nor U115615 ( n60909, n60910, n60911 );
nor U115616 ( n60908, n60914, n60915 );
nor U115617 ( n60910, n60240, n60868 );
nand U115618 ( n12696, n61313, n61314 );
nor U115619 ( n61314, n61315, n61316 );
nor U115620 ( n61313, n61319, n61320 );
nor U115621 ( n61315, n60218, n61279 );
nand U115622 ( n12776, n61136, n61137 );
nor U115623 ( n61137, n61138, n61139 );
nor U115624 ( n61136, n61142, n61143 );
nor U115625 ( n61138, n60218, n61115 );
nand U115626 ( n12816, n61052, n61053 );
nor U115627 ( n61053, n61054, n61055 );
nor U115628 ( n61052, n61058, n61059 );
nor U115629 ( n61054, n60218, n61031 );
nand U115630 ( n12856, n60974, n60975 );
nor U115631 ( n60975, n60976, n60977 );
nor U115632 ( n60974, n60980, n60981 );
nor U115633 ( n60976, n60218, n60950 );
nand U115634 ( n12976, n60734, n60735 );
nor U115635 ( n60735, n60736, n60737 );
nor U115636 ( n60734, n60740, n60741 );
nor U115637 ( n60736, n60218, n60713 );
nand U115638 ( n13016, n60649, n60650 );
nor U115639 ( n60650, n60651, n60652 );
nor U115640 ( n60649, n60656, n60657 );
nor U115641 ( n60651, n60218, n60626 );
nand U115642 ( n12721, n61246, n61247 );
nor U115643 ( n61247, n61248, n61249 );
nor U115644 ( n61246, n61252, n61253 );
nor U115645 ( n61248, n60251, n61201 );
nand U115646 ( n12881, n60916, n60917 );
nor U115647 ( n60917, n60918, n60919 );
nor U115648 ( n60916, n60922, n60923 );
nor U115649 ( n60918, n60251, n60868 );
nand U115650 ( n12751, n61193, n61194 );
nor U115651 ( n61194, n61195, n61196 );
nor U115652 ( n61193, n61202, n61203 );
nor U115653 ( n61195, n60180, n61201 );
nand U115654 ( n12911, n60860, n60861 );
nor U115655 ( n60861, n60862, n60863 );
nor U115656 ( n60860, n60869, n60870 );
nor U115657 ( n60862, n60180, n60868 );
nand U115658 ( n12661, n61382, n61383 );
nor U115659 ( n61383, n61384, n61385 );
nor U115660 ( n61382, n61388, n61389 );
nor U115661 ( n61384, n60207, n61369 );
nand U115662 ( n12701, n61305, n61306 );
nor U115663 ( n61306, n61307, n61308 );
nor U115664 ( n61305, n61311, n61312 );
nor U115665 ( n61307, n60207, n61279 );
nand U115666 ( n12781, n61128, n61129 );
nor U115667 ( n61129, n61130, n61131 );
nor U115668 ( n61128, n61134, n61135 );
nor U115669 ( n61130, n60207, n61115 );
nand U115670 ( n12821, n61044, n61045 );
nor U115671 ( n61045, n61046, n61047 );
nor U115672 ( n61044, n61050, n61051 );
nor U115673 ( n61046, n60207, n61031 );
nand U115674 ( n12861, n60963, n60964 );
nor U115675 ( n60964, n60965, n60966 );
nor U115676 ( n60963, n60969, n60970 );
nor U115677 ( n60965, n60207, n60950 );
nand U115678 ( n12981, n60726, n60727 );
nor U115679 ( n60727, n60728, n60729 );
nor U115680 ( n60726, n60732, n60733 );
nor U115681 ( n60728, n60207, n60713 );
nand U115682 ( n13021, n60640, n60641 );
nor U115683 ( n60641, n60642, n60643 );
nor U115684 ( n60640, n60647, n60648 );
nor U115685 ( n60642, n60207, n60626 );
nand U115686 ( n12651, n61460, n61461 );
nor U115687 ( n61461, n61462, n61463 );
nor U115688 ( n61460, n61466, n61467 );
nor U115689 ( n61462, n60229, n61369 );
nand U115690 ( n12691, n61321, n61322 );
nor U115691 ( n61322, n61323, n61324 );
nor U115692 ( n61321, n61327, n61328 );
nor U115693 ( n61323, n60229, n61279 );
nand U115694 ( n12771, n61144, n61145 );
nor U115695 ( n61145, n61146, n61147 );
nor U115696 ( n61144, n61150, n61151 );
nor U115697 ( n61146, n60229, n61115 );
nand U115698 ( n12811, n61060, n61061 );
nor U115699 ( n61061, n61062, n61063 );
nor U115700 ( n61060, n61066, n61067 );
nor U115701 ( n61062, n60229, n61031 );
nand U115702 ( n12851, n60982, n60983 );
nor U115703 ( n60983, n60984, n60985 );
nor U115704 ( n60982, n60988, n60989 );
nor U115705 ( n60984, n60229, n60950 );
nand U115706 ( n12971, n60742, n60743 );
nor U115707 ( n60743, n60744, n60745 );
nor U115708 ( n60742, n60748, n60749 );
nor U115709 ( n60744, n60229, n60713 );
nand U115710 ( n13011, n60658, n60659 );
nor U115711 ( n60659, n60660, n60661 );
nor U115712 ( n60658, n60665, n60666 );
nor U115713 ( n60660, n60229, n60626 );
nand U115714 ( n12656, n61452, n61453 );
nor U115715 ( n61453, n61454, n61455 );
nor U115716 ( n61452, n61458, n61459 );
nor U115717 ( n61454, n60218, n61369 );
nand U115718 ( n12676, n61345, n61346 );
nor U115719 ( n61346, n61347, n61348 );
nor U115720 ( n61345, n61358, n61359 );
nor U115721 ( n61347, n60277, n61279 );
nand U115722 ( n12716, n61254, n61255 );
nor U115723 ( n61255, n61256, n61257 );
nor U115724 ( n61254, n61268, n61269 );
nor U115725 ( n61256, n60272, n61201 );
nand U115726 ( n12756, n61178, n61179 );
nor U115727 ( n61179, n61180, n61181 );
nor U115728 ( n61178, n61191, n61192 );
nor U115729 ( n61180, n60277, n61115 );
nand U115730 ( n12796, n61090, n61091 );
nor U115731 ( n61091, n61092, n61093 );
nor U115732 ( n61090, n61103, n61104 );
nor U115733 ( n61092, n60277, n61031 );
nand U115734 ( n12836, n61006, n61007 );
nor U115735 ( n61007, n61008, n61009 );
nor U115736 ( n61006, n61019, n61020 );
nor U115737 ( n61008, n60277, n60950 );
nand U115738 ( n12876, n60924, n60925 );
nor U115739 ( n60925, n60926, n60927 );
nor U115740 ( n60924, n60938, n60939 );
nor U115741 ( n60926, n60272, n60868 );
nand U115742 ( n12956, n60769, n60770 );
nor U115743 ( n60770, n60771, n60772 );
nor U115744 ( n60769, n60782, n60783 );
nor U115745 ( n60771, n60277, n60713 );
nand U115746 ( n12996, n60688, n60689 );
nor U115747 ( n60689, n60690, n60691 );
nor U115748 ( n60688, n60702, n60703 );
nor U115749 ( n60690, n60277, n60626 );
nand U115750 ( n12636, n61484, n61485 );
nor U115751 ( n61485, n61486, n61487 );
nor U115752 ( n61484, n61497, n61498 );
nor U115753 ( n61486, n60277, n61369 );
nand U115754 ( n5946, n28173, n28174 );
nor U115755 ( n28174, n28175, n28176 );
nor U115756 ( n28173, n28179, n28180 );
nor U115757 ( n28175, n27110, n28124 );
nand U115758 ( n5976, n28116, n28117 );
nor U115759 ( n28117, n28118, n28119 );
nor U115760 ( n28116, n28125, n28126 );
nor U115761 ( n28118, n27043, n28124 );
nand U115762 ( n6026, n28011, n28012 );
nor U115763 ( n28012, n28013, n28014 );
nor U115764 ( n28011, n28017, n28018 );
nor U115765 ( n28013, n27110, n27966 );
nand U115766 ( n6066, n27929, n27930 );
nor U115767 ( n27930, n27931, n27932 );
nor U115768 ( n27929, n27935, n27936 );
nor U115769 ( n27931, n27110, n27884 );
nand U115770 ( n6106, n27851, n27852 );
nor U115771 ( n27852, n27853, n27854 );
nor U115772 ( n27851, n27857, n27858 );
nor U115773 ( n27853, n27110, n27802 );
nand U115774 ( n6226, n27608, n27609 );
nor U115775 ( n27609, n27610, n27611 );
nor U115776 ( n27608, n27614, n27615 );
nor U115777 ( n27610, n27110, n27563 );
nand U115778 ( n6266, n27527, n27528 );
nor U115779 ( n27528, n27529, n27530 );
nor U115780 ( n27527, n27534, n27535 );
nor U115781 ( n27529, n27110, n27477 );
nand U115782 ( n5936, n28197, n28198 );
nor U115783 ( n28198, n28199, n28200 );
nor U115784 ( n28197, n28206, n28207 );
nor U115785 ( n28199, n27043, n28205 );
nand U115786 ( n6056, n27958, n27959 );
nor U115787 ( n27959, n27960, n27961 );
nor U115788 ( n27958, n27967, n27968 );
nor U115789 ( n27960, n27043, n27966 );
nand U115790 ( n6096, n27876, n27877 );
nor U115791 ( n27877, n27878, n27879 );
nor U115792 ( n27876, n27885, n27886 );
nor U115793 ( n27878, n27043, n27884 );
nand U115794 ( n6136, n27794, n27795 );
nor U115795 ( n27795, n27796, n27797 );
nor U115796 ( n27794, n27803, n27804 );
nor U115797 ( n27796, n27043, n27802 );
nand U115798 ( n6296, n27468, n27469 );
nor U115799 ( n27469, n27470, n27471 );
nor U115800 ( n27468, n27478, n27479 );
nor U115801 ( n27470, n27043, n27477 );
nand U115802 ( n6001, n28067, n28068 );
nor U115803 ( n28068, n28069, n28070 );
nor U115804 ( n28067, n28073, n28074 );
nor U115805 ( n28069, n27074, n28042 );
nand U115806 ( n6161, n27738, n27739 );
nor U115807 ( n27739, n27740, n27741 );
nor U115808 ( n27738, n27744, n27745 );
nor U115809 ( n27740, n27074, n27717 );
nand U115810 ( n5996, n28075, n28076 );
nor U115811 ( n28076, n28077, n28078 );
nor U115812 ( n28075, n28081, n28082 );
nor U115813 ( n28077, n27085, n28042 );
nand U115814 ( n6156, n27752, n27753 );
nor U115815 ( n27753, n27754, n27755 );
nor U115816 ( n27752, n27758, n27759 );
nor U115817 ( n27754, n27085, n27717 );
nand U115818 ( n6006, n28059, n28060 );
nor U115819 ( n28060, n28061, n28062 );
nor U115820 ( n28059, n28065, n28066 );
nor U115821 ( n28061, n27063, n28042 );
nand U115822 ( n12646, n61468, n61469 );
nor U115823 ( n61469, n61470, n61471 );
nor U115824 ( n61468, n61474, n61475 );
nor U115825 ( n61470, n60243, n61369 );
nand U115826 ( n12686, n61329, n61330 );
nor U115827 ( n61330, n61331, n61332 );
nor U115828 ( n61329, n61335, n61336 );
nor U115829 ( n61331, n60243, n61279 );
nand U115830 ( n12766, n61152, n61153 );
nor U115831 ( n61153, n61154, n61155 );
nor U115832 ( n61152, n61158, n61159 );
nor U115833 ( n61154, n60243, n61115 );
nand U115834 ( n12806, n61074, n61075 );
nor U115835 ( n61075, n61076, n61077 );
nor U115836 ( n61074, n61080, n61081 );
nor U115837 ( n61076, n60243, n61031 );
nand U115838 ( n12846, n60990, n60991 );
nor U115839 ( n60991, n60992, n60993 );
nor U115840 ( n60990, n60996, n60997 );
nor U115841 ( n60992, n60243, n60950 );
nand U115842 ( n12966, n60750, n60751 );
nor U115843 ( n60751, n60752, n60753 );
nor U115844 ( n60750, n60756, n60757 );
nor U115845 ( n60752, n60243, n60713 );
nand U115846 ( n13006, n60670, n60671 );
nor U115847 ( n60671, n60672, n60673 );
nor U115848 ( n60670, n60677, n60678 );
nor U115849 ( n60672, n60243, n60626 );
nand U115850 ( n12666, n61374, n61375 );
nor U115851 ( n61375, n61376, n61377 );
nor U115852 ( n61374, n61380, n61381 );
nor U115853 ( n61376, n60196, n61369 );
nand U115854 ( n12706, n61297, n61298 );
nor U115855 ( n61298, n61299, n61300 );
nor U115856 ( n61297, n61303, n61304 );
nor U115857 ( n61299, n60196, n61279 );
nand U115858 ( n12786, n61120, n61121 );
nor U115859 ( n61121, n61122, n61123 );
nor U115860 ( n61120, n61126, n61127 );
nor U115861 ( n61122, n60196, n61115 );
nand U115862 ( n12826, n61036, n61037 );
nor U115863 ( n61037, n61038, n61039 );
nor U115864 ( n61036, n61042, n61043 );
nor U115865 ( n61038, n60196, n61031 );
nand U115866 ( n12866, n60955, n60956 );
nor U115867 ( n60956, n60957, n60958 );
nor U115868 ( n60955, n60961, n60962 );
nor U115869 ( n60957, n60196, n60950 );
nand U115870 ( n12986, n60718, n60719 );
nor U115871 ( n60719, n60720, n60721 );
nor U115872 ( n60718, n60724, n60725 );
nor U115873 ( n60720, n60196, n60713 );
nand U115874 ( n13026, n60631, n60632 );
nor U115875 ( n60632, n60633, n60634 );
nor U115876 ( n60631, n60638, n60639 );
nor U115877 ( n60633, n60196, n60626 );
nand U115878 ( n41602, n829, n41466 );
nand U115879 ( n6011, n28047, n28048 );
nor U115880 ( n28048, n28049, n28050 );
nor U115881 ( n28047, n28053, n28054 );
nor U115882 ( n28049, n27052, n28042 );
nand U115883 ( n6171, n27722, n27723 );
nor U115884 ( n27723, n27724, n27725 );
nor U115885 ( n27722, n27728, n27729 );
nor U115886 ( n27724, n27052, n27717 );
nand U115887 ( n6256, n27555, n27556 );
nor U115888 ( n27556, n27557, n27558 );
nor U115889 ( n27555, n27564, n27565 );
nor U115890 ( n27557, n27043, n27563 );
nand U115891 ( n6166, n27730, n27731 );
nor U115892 ( n27731, n27732, n27733 );
nor U115893 ( n27730, n27736, n27737 );
nor U115894 ( n27732, n27063, n27717 );
nand U115895 ( n12681, n61337, n61338 );
nor U115896 ( n61338, n61339, n61340 );
nor U115897 ( n61337, n61343, n61344 );
nor U115898 ( n61339, n60254, n61279 );
nand U115899 ( n12711, n61271, n61272 );
nor U115900 ( n61272, n61273, n61274 );
nor U115901 ( n61271, n61280, n61281 );
nor U115902 ( n61273, n60184, n61279 );
nand U115903 ( n5906, n28254, n28255 );
nor U115904 ( n28255, n28256, n28257 );
nor U115905 ( n28254, n28260, n28261 );
nor U115906 ( n28256, n27110, n28205 );
nand U115907 ( n12736, n61222, n61223 );
nor U115908 ( n61223, n61224, n61225 );
nor U115909 ( n61222, n61228, n61229 );
nor U115910 ( n61224, n60215, n61201 );
nand U115911 ( n12896, n60892, n60893 );
nor U115912 ( n60893, n60894, n60895 );
nor U115913 ( n60892, n60898, n60899 );
nor U115914 ( n60894, n60215, n60868 );
nand U115915 ( n12746, n61206, n61207 );
nor U115916 ( n61207, n61208, n61209 );
nor U115917 ( n61206, n61212, n61213 );
nor U115918 ( n61208, n60193, n61201 );
nand U115919 ( n12906, n60876, n60877 );
nor U115920 ( n60877, n60878, n60879 );
nor U115921 ( n60876, n60882, n60883 );
nor U115922 ( n60878, n60193, n60868 );
nand U115923 ( n12741, n61214, n61215 );
nor U115924 ( n61215, n61216, n61217 );
nor U115925 ( n61214, n61220, n61221 );
nor U115926 ( n61216, n60204, n61201 );
nand U115927 ( n12901, n60884, n60885 );
nor U115928 ( n60885, n60886, n60887 );
nor U115929 ( n60884, n60890, n60891 );
nor U115930 ( n60886, n60204, n60868 );
nand U115931 ( n12731, n61230, n61231 );
nor U115932 ( n61231, n61232, n61233 );
nor U115933 ( n61230, n61236, n61237 );
nor U115934 ( n61232, n60226, n61201 );
nand U115935 ( n12891, n60900, n60901 );
nor U115936 ( n60901, n60902, n60903 );
nor U115937 ( n60900, n60906, n60907 );
nor U115938 ( n60902, n60226, n60868 );
nand U115939 ( n12641, n61476, n61477 );
nor U115940 ( n61477, n61478, n61479 );
nor U115941 ( n61476, n61482, n61483 );
nor U115942 ( n61478, n60254, n61369 );
nand U115943 ( n12761, n61160, n61161 );
nor U115944 ( n61161, n61162, n61163 );
nor U115945 ( n61160, n61166, n61167 );
nor U115946 ( n61162, n60254, n61115 );
nand U115947 ( n12801, n61082, n61083 );
nor U115948 ( n61083, n61084, n61085 );
nor U115949 ( n61082, n61088, n61089 );
nor U115950 ( n61084, n60254, n61031 );
nand U115951 ( n12841, n60998, n60999 );
nor U115952 ( n60999, n61000, n61001 );
nor U115953 ( n60998, n61004, n61005 );
nor U115954 ( n61000, n60254, n60950 );
nand U115955 ( n12961, n60758, n60759 );
nor U115956 ( n60759, n60760, n60761 );
nor U115957 ( n60758, n60764, n60765 );
nor U115958 ( n60760, n60254, n60713 );
nand U115959 ( n13001, n60679, n60680 );
nor U115960 ( n60680, n60681, n60682 );
nor U115961 ( n60679, n60686, n60687 );
nor U115962 ( n60681, n60254, n60626 );
nand U115963 ( n12671, n61361, n61362 );
nor U115964 ( n61362, n61363, n61364 );
nor U115965 ( n61361, n61370, n61371 );
nor U115966 ( n61363, n60184, n61369 );
nand U115967 ( n12791, n61107, n61108 );
nor U115968 ( n61108, n61109, n61110 );
nor U115969 ( n61107, n61116, n61117 );
nor U115970 ( n61109, n60184, n61115 );
nand U115971 ( n12831, n61023, n61024 );
nor U115972 ( n61024, n61025, n61026 );
nor U115973 ( n61023, n61032, n61033 );
nor U115974 ( n61025, n60184, n61031 );
nand U115975 ( n12871, n60942, n60943 );
nor U115976 ( n60943, n60944, n60945 );
nor U115977 ( n60942, n60951, n60952 );
nor U115978 ( n60944, n60184, n60950 );
nand U115979 ( n12991, n60705, n60706 );
nor U115980 ( n60706, n60707, n60708 );
nor U115981 ( n60705, n60714, n60715 );
nor U115982 ( n60707, n60184, n60713 );
nand U115983 ( n13031, n60617, n60618 );
nor U115984 ( n60618, n60619, n60620 );
nor U115985 ( n60617, n60627, n60628 );
nor U115986 ( n60619, n60184, n60626 );
nand U115987 ( n68197, n68198, n6089 );
nor U115988 ( n68198, n5689, n73187 );
nand U115989 ( n33446, n33447, n3474 );
nor U115990 ( n33447, n3088, n73197 );
nand U115991 ( n47166, n47167, n7878 );
nor U115992 ( n47167, n7474, n73178 );
nand U115993 ( n26196, n26197, n4312 );
nor U115994 ( n26197, n3932, n73188 );
nand U115995 ( n59335, n59336, n6944 );
nor U115996 ( n59336, n6564, n73189 );
nor U115997 ( n8430, n8408, n8410 );
not U115998 ( n7865, n47926 );
nand U115999 ( n48518, n7848, n48413 );
nand U116000 ( n48412, n47941, n47951 );
not U116001 ( n52, n27497 );
not U116002 ( n58, n27524 );
not U116003 ( n54, n27506 );
not U116004 ( n50, n27488 );
not U116005 ( n56, n27515 );
not U116006 ( n48, n27475 );
not U116007 ( n60, n27533 );
not U116008 ( n62, n27542 );
not U116009 ( n312, n60655 );
not U116010 ( n317, n60676 );
not U116011 ( n309, n60646 );
not U116012 ( n307, n60637 );
not U116013 ( n314, n60664 );
not U116014 ( n319, n60685 );
not U116015 ( n322, n60694 );
not U116016 ( n304, n60624 );
nand U116017 ( n6371, n27316, n27317 );
nor U116018 ( n27316, n27322, n27323 );
nor U116019 ( n27317, n27318, n27319 );
nor U116020 ( n27322, n27055, n27315 );
nand U116021 ( n6411, n27234, n27235 );
nor U116022 ( n27234, n27240, n27241 );
nor U116023 ( n27235, n27236, n27237 );
nor U116024 ( n27240, n27055, n27233 );
nand U116025 ( n6451, n27152, n27153 );
nor U116026 ( n27152, n27158, n27159 );
nor U116027 ( n27153, n27154, n27155 );
nor U116028 ( n27158, n27055, n27151 );
nand U116029 ( n6341, n27366, n27367 );
nor U116030 ( n27366, n27380, n27381 );
nor U116031 ( n27367, n27368, n27369 );
nor U116032 ( n27380, n27133, n27315 );
nand U116033 ( n6381, n27284, n27285 );
nor U116034 ( n27284, n27298, n27299 );
nor U116035 ( n27285, n27286, n27287 );
nor U116036 ( n27298, n27133, n27233 );
nand U116037 ( n6421, n27200, n27201 );
nor U116038 ( n27200, n27215, n27216 );
nor U116039 ( n27201, n27202, n27203 );
nor U116040 ( n27215, n27133, n27151 );
nand U116041 ( n6346, n27358, n27359 );
nor U116042 ( n27358, n27364, n27365 );
nor U116043 ( n27359, n27360, n27361 );
nor U116044 ( n27364, n27110, n27315 );
nand U116045 ( n6386, n27276, n27277 );
nor U116046 ( n27276, n27282, n27283 );
nor U116047 ( n27277, n27278, n27279 );
nor U116048 ( n27282, n27110, n27233 );
nand U116049 ( n6426, n27192, n27193 );
nor U116050 ( n27192, n27198, n27199 );
nor U116051 ( n27193, n27194, n27195 );
nor U116052 ( n27198, n27110, n27151 );
nand U116053 ( n6376, n27303, n27304 );
nor U116054 ( n27303, n27312, n27313 );
nor U116055 ( n27304, n27305, n27306 );
nor U116056 ( n27312, n27043, n27315 );
nand U116057 ( n6416, n27221, n27222 );
nor U116058 ( n27221, n27230, n27231 );
nor U116059 ( n27222, n27223, n27224 );
nor U116060 ( n27230, n27043, n27233 );
nand U116061 ( n6456, n27139, n27140 );
nor U116062 ( n27139, n27148, n27149 );
nor U116063 ( n27140, n27141, n27142 );
nor U116064 ( n27148, n27043, n27151 );
nand U116065 ( n6351, n27350, n27351 );
nor U116066 ( n27350, n27356, n27357 );
nor U116067 ( n27351, n27352, n27353 );
nor U116068 ( n27356, n27099, n27315 );
nand U116069 ( n6391, n27268, n27269 );
nor U116070 ( n27268, n27274, n27275 );
nor U116071 ( n27269, n27270, n27271 );
nor U116072 ( n27274, n27099, n27233 );
nand U116073 ( n6431, n27184, n27185 );
nor U116074 ( n27184, n27190, n27191 );
nor U116075 ( n27185, n27186, n27187 );
nor U116076 ( n27190, n27099, n27151 );
nand U116077 ( n6361, n27332, n27333 );
nor U116078 ( n27332, n27338, n27339 );
nor U116079 ( n27333, n27334, n27335 );
nor U116080 ( n27338, n27077, n27315 );
nand U116081 ( n6401, n27252, n27253 );
nor U116082 ( n27252, n27258, n27259 );
nor U116083 ( n27253, n27254, n27255 );
nor U116084 ( n27258, n27077, n27233 );
nand U116085 ( n6441, n27168, n27169 );
nor U116086 ( n27168, n27174, n27175 );
nor U116087 ( n27169, n27170, n27171 );
nor U116088 ( n27174, n27077, n27151 );
nand U116089 ( n6356, n27342, n27343 );
nor U116090 ( n27342, n27348, n27349 );
nor U116091 ( n27343, n27344, n27345 );
nor U116092 ( n27348, n27088, n27315 );
nand U116093 ( n6396, n27260, n27261 );
nor U116094 ( n27260, n27266, n27267 );
nor U116095 ( n27261, n27262, n27263 );
nor U116096 ( n27266, n27088, n27233 );
nand U116097 ( n6436, n27176, n27177 );
nor U116098 ( n27176, n27182, n27183 );
nor U116099 ( n27177, n27178, n27179 );
nor U116100 ( n27182, n27088, n27151 );
nand U116101 ( n6366, n27324, n27325 );
nor U116102 ( n27324, n27330, n27331 );
nor U116103 ( n27325, n27326, n27327 );
nor U116104 ( n27330, n27066, n27315 );
nand U116105 ( n6406, n27244, n27245 );
nor U116106 ( n27244, n27250, n27251 );
nor U116107 ( n27245, n27246, n27247 );
nor U116108 ( n27250, n27066, n27233 );
nand U116109 ( n6446, n27160, n27161 );
nor U116110 ( n27160, n27166, n27167 );
nor U116111 ( n27161, n27162, n27163 );
nor U116112 ( n27166, n27066, n27151 );
nand U116113 ( n13086, n60498, n60499 );
nor U116114 ( n60498, n60504, n60505 );
nor U116115 ( n60499, n60500, n60501 );
nor U116116 ( n60504, n60243, n60458 );
nand U116117 ( n13126, n60411, n60412 );
nor U116118 ( n60411, n60417, n60418 );
nor U116119 ( n60412, n60413, n60414 );
nor U116120 ( n60417, n60243, n60378 );
nand U116121 ( n13166, n60326, n60327 );
nor U116122 ( n60326, n60332, n60333 );
nor U116123 ( n60327, n60328, n60329 );
nor U116124 ( n60332, n60243, n60293 );
nand U116125 ( n13096, n60482, n60483 );
nor U116126 ( n60482, n60488, n60489 );
nor U116127 ( n60483, n60484, n60485 );
nor U116128 ( n60488, n60218, n60458 );
nand U116129 ( n13136, n60395, n60396 );
nor U116130 ( n60395, n60401, n60402 );
nor U116131 ( n60396, n60397, n60398 );
nor U116132 ( n60401, n60218, n60378 );
nand U116133 ( n13176, n60310, n60311 );
nor U116134 ( n60310, n60316, n60317 );
nor U116135 ( n60311, n60312, n60313 );
nor U116136 ( n60316, n60218, n60293 );
nand U116137 ( n13081, n60506, n60507 );
nor U116138 ( n60506, n60512, n60513 );
nor U116139 ( n60507, n60508, n60509 );
nor U116140 ( n60512, n60254, n60458 );
nand U116141 ( n13121, n60419, n60420 );
nor U116142 ( n60419, n60425, n60426 );
nor U116143 ( n60420, n60421, n60422 );
nor U116144 ( n60425, n60254, n60378 );
nand U116145 ( n13161, n60334, n60335 );
nor U116146 ( n60334, n60340, n60341 );
nor U116147 ( n60335, n60336, n60337 );
nor U116148 ( n60340, n60254, n60293 );
nand U116149 ( n13106, n60462, n60463 );
nor U116150 ( n60462, n60468, n60469 );
nor U116151 ( n60463, n60464, n60465 );
nor U116152 ( n60468, n60196, n60458 );
nand U116153 ( n13146, n60379, n60380 );
nor U116154 ( n60379, n60385, n60386 );
nor U116155 ( n60380, n60381, n60382 );
nor U116156 ( n60385, n60196, n60378 );
nand U116157 ( n13186, n60294, n60295 );
nor U116158 ( n60294, n60300, n60301 );
nor U116159 ( n60295, n60296, n60297 );
nor U116160 ( n60300, n60196, n60293 );
nand U116161 ( n13111, n60446, n60447 );
nor U116162 ( n60446, n60455, n60456 );
nor U116163 ( n60447, n60448, n60449 );
nor U116164 ( n60455, n60184, n60458 );
nand U116165 ( n13151, n60366, n60367 );
nor U116166 ( n60366, n60375, n60376 );
nor U116167 ( n60367, n60368, n60369 );
nor U116168 ( n60375, n60184, n60378 );
nand U116169 ( n13191, n60281, n60282 );
nor U116170 ( n60281, n60290, n60291 );
nor U116171 ( n60282, n60283, n60284 );
nor U116172 ( n60290, n60184, n60293 );
nand U116173 ( n13101, n60470, n60471 );
nor U116174 ( n60470, n60476, n60477 );
nor U116175 ( n60471, n60472, n60473 );
nor U116176 ( n60476, n60207, n60458 );
nand U116177 ( n13141, n60387, n60388 );
nor U116178 ( n60387, n60393, n60394 );
nor U116179 ( n60388, n60389, n60390 );
nor U116180 ( n60393, n60207, n60378 );
nand U116181 ( n13181, n60302, n60303 );
nor U116182 ( n60302, n60308, n60309 );
nor U116183 ( n60303, n60304, n60305 );
nor U116184 ( n60308, n60207, n60293 );
nand U116185 ( n13091, n60490, n60491 );
nor U116186 ( n60490, n60496, n60497 );
nor U116187 ( n60491, n60492, n60493 );
nor U116188 ( n60496, n60229, n60458 );
nand U116189 ( n13131, n60403, n60404 );
nor U116190 ( n60403, n60409, n60410 );
nor U116191 ( n60404, n60405, n60406 );
nor U116192 ( n60409, n60229, n60378 );
nand U116193 ( n13171, n60318, n60319 );
nor U116194 ( n60318, n60324, n60325 );
nor U116195 ( n60319, n60320, n60321 );
nor U116196 ( n60324, n60229, n60293 );
nand U116197 ( n13076, n60514, n60515 );
nor U116198 ( n60514, n60528, n60529 );
nor U116199 ( n60515, n60516, n60517 );
nor U116200 ( n60528, n60277, n60458 );
nand U116201 ( n13116, n60427, n60428 );
nor U116202 ( n60427, n60441, n60442 );
nor U116203 ( n60428, n60429, n60430 );
nor U116204 ( n60441, n60277, n60378 );
nand U116205 ( n13156, n60345, n60346 );
nor U116206 ( n60345, n60360, n60361 );
nor U116207 ( n60346, n60347, n60348 );
nor U116208 ( n60360, n60277, n60293 );
nand U116209 ( n26814, n25823, n73075 );
nand U116210 ( n59954, n58961, n73074 );
nand U116211 ( n34059, n33070, n73077 );
nand U116212 ( n68813, n67826, n73076 );
nand U116213 ( n6301, n27448, n27449 );
nor U116214 ( n27449, n27450, n27451 );
nor U116215 ( n27448, n27465, n27466 );
nor U116216 ( n27450, n27128, n27393 );
nand U116217 ( n6336, n27385, n27386 );
nor U116218 ( n27386, n27387, n27388 );
nor U116219 ( n27385, n27394, n27395 );
nor U116220 ( n27387, n27039, n27393 );
nand U116221 ( n6311, n27430, n27431 );
nor U116222 ( n27431, n27432, n27433 );
nor U116223 ( n27430, n27436, n27437 );
nor U116224 ( n27432, n27096, n27393 );
nand U116225 ( n6306, n27440, n27441 );
nor U116226 ( n27441, n27442, n27443 );
nor U116227 ( n27440, n27446, n27447 );
nor U116228 ( n27442, n27107, n27393 );
nand U116229 ( n6461, n27111, n27112 );
nor U116230 ( n27112, n27113, n27114 );
nor U116231 ( n27111, n27131, n27132 );
nor U116232 ( n27113, n27038, n27128 );
nand U116233 ( n6466, n27100, n27101 );
nor U116234 ( n27101, n27102, n27103 );
nor U116235 ( n27100, n27108, n27109 );
nor U116236 ( n27102, n27038, n27107 );
nand U116237 ( n6496, n27029, n27030 );
nor U116238 ( n27030, n27031, n27032 );
nor U116239 ( n27029, n27040, n27041 );
nor U116240 ( n27031, n27038, n27039 );
nand U116241 ( n6471, n27089, n27090 );
nor U116242 ( n27090, n27091, n27092 );
nor U116243 ( n27089, n27097, n27098 );
nor U116244 ( n27091, n27038, n27096 );
nand U116245 ( n13046, n60581, n60582 );
nor U116246 ( n60582, n60583, n60584 );
nor U116247 ( n60581, n60587, n60588 );
nor U116248 ( n60583, n60240, n60541 );
nand U116249 ( n13071, n60533, n60534 );
nor U116250 ( n60534, n60535, n60536 );
nor U116251 ( n60533, n60542, n60543 );
nor U116252 ( n60535, n60180, n60541 );
nand U116253 ( n13041, n60589, n60590 );
nor U116254 ( n60590, n60591, n60592 );
nor U116255 ( n60589, n60595, n60596 );
nor U116256 ( n60591, n60251, n60541 );
nand U116257 ( n13036, n60597, n60598 );
nor U116258 ( n60598, n60599, n60600 );
nor U116259 ( n60597, n60614, n60615 );
nor U116260 ( n60599, n60272, n60541 );
nand U116261 ( n13206, n60233, n60234 );
nor U116262 ( n60234, n60235, n60236 );
nor U116263 ( n60233, n60241, n60242 );
nor U116264 ( n60235, n60179, n60240 );
nand U116265 ( n13201, n60244, n60245 );
nor U116266 ( n60245, n60246, n60247 );
nor U116267 ( n60244, n60252, n60253 );
nor U116268 ( n60246, n60179, n60251 );
nand U116269 ( n13231, n60170, n60171 );
nor U116270 ( n60171, n60172, n60173 );
nor U116271 ( n60170, n60181, n60182 );
nor U116272 ( n60172, n60179, n60180 );
nand U116273 ( n13196, n60255, n60256 );
nor U116274 ( n60256, n60257, n60258 );
nor U116275 ( n60255, n60275, n60276 );
nor U116276 ( n60257, n60179, n60272 );
nand U116277 ( n6331, n27398, n27399 );
nor U116278 ( n27399, n27400, n27401 );
nor U116279 ( n27398, n27404, n27405 );
nor U116280 ( n27400, n27052, n27393 );
nand U116281 ( n6321, n27414, n27415 );
nor U116282 ( n27415, n27416, n27417 );
nor U116283 ( n27414, n27420, n27421 );
nor U116284 ( n27416, n27074, n27393 );
nand U116285 ( n6316, n27422, n27423 );
nor U116286 ( n27423, n27424, n27425 );
nor U116287 ( n27422, n27428, n27429 );
nor U116288 ( n27424, n27085, n27393 );
nand U116289 ( n6326, n27406, n27407 );
nor U116290 ( n27407, n27408, n27409 );
nor U116291 ( n27406, n27412, n27413 );
nor U116292 ( n27408, n27063, n27393 );
nand U116293 ( n6491, n27045, n27046 );
nor U116294 ( n27046, n27047, n27048 );
nor U116295 ( n27045, n27053, n27054 );
nor U116296 ( n27047, n27038, n27052 );
nand U116297 ( n6481, n27067, n27068 );
nor U116298 ( n27068, n27069, n27070 );
nor U116299 ( n27067, n27075, n27076 );
nor U116300 ( n27069, n27038, n27074 );
nand U116301 ( n6476, n27078, n27079 );
nor U116302 ( n27079, n27080, n27081 );
nor U116303 ( n27078, n27086, n27087 );
nor U116304 ( n27080, n27038, n27085 );
nand U116305 ( n6486, n27056, n27057 );
nor U116306 ( n27057, n27058, n27059 );
nor U116307 ( n27056, n27064, n27065 );
nor U116308 ( n27058, n27038, n27063 );
nor U116309 ( n48878, n48413, n7848 );
nand U116310 ( n13056, n60565, n60566 );
nor U116311 ( n60566, n60567, n60568 );
nor U116312 ( n60565, n60571, n60572 );
nor U116313 ( n60567, n60215, n60541 );
nand U116314 ( n13061, n60554, n60555 );
nor U116315 ( n60555, n60556, n60557 );
nor U116316 ( n60554, n60560, n60561 );
nor U116317 ( n60556, n60204, n60541 );
nand U116318 ( n13051, n60573, n60574 );
nor U116319 ( n60574, n60575, n60576 );
nor U116320 ( n60573, n60579, n60580 );
nor U116321 ( n60575, n60226, n60541 );
nand U116322 ( n13066, n60546, n60547 );
nor U116323 ( n60547, n60548, n60549 );
nor U116324 ( n60546, n60552, n60553 );
nor U116325 ( n60548, n60193, n60541 );
nand U116326 ( n13216, n60208, n60209 );
nor U116327 ( n60209, n60210, n60211 );
nor U116328 ( n60208, n60216, n60217 );
nor U116329 ( n60210, n60179, n60215 );
nand U116330 ( n13226, n60186, n60187 );
nor U116331 ( n60187, n60188, n60189 );
nor U116332 ( n60186, n60194, n60195 );
nor U116333 ( n60188, n60179, n60193 );
nand U116334 ( n13221, n60197, n60198 );
nor U116335 ( n60198, n60199, n60200 );
nor U116336 ( n60197, n60205, n60206 );
nor U116337 ( n60199, n60179, n60204 );
nand U116338 ( n13211, n60219, n60220 );
nor U116339 ( n60220, n60221, n60222 );
nor U116340 ( n60219, n60227, n60228 );
nor U116341 ( n60221, n60179, n60226 );
nor U116342 ( n22007, n21952, n22008 );
nor U116343 ( n22008, n22009, n75183 );
nor U116344 ( n29326, n29269, n29327 );
nor U116345 ( n29327, n29328, n75181 );
nor U116346 ( n63089, n63036, n63090 );
nor U116347 ( n63090, n63091, n75182 );
nor U116348 ( n55117, n55064, n55118 );
nor U116349 ( n55118, n55119, n75184 );
nand U116350 ( n23209, n23819, n23824 );
nand U116351 ( n441, n33042, n3794 );
nor U116352 ( n33042, n76749, n23824 );
not U116353 ( n4687, n456 );
nor U116354 ( n68679, n68598, n68682 );
nor U116355 ( n33923, n33842, n33926 );
nor U116356 ( n26678, n26597, n26681 );
nor U116357 ( n59820, n59739, n59823 );
nor U116358 ( n47658, n47577, n47661 );
nor U116359 ( n14363, n14262, n14367 );
nor U116360 ( n23299, n75391, n23162 );
nor U116361 ( n23444, n75394, n23162 );
nor U116362 ( n23632, n75395, n23162 );
nor U116363 ( n23677, n75397, n23162 );
nor U116364 ( n23721, n75396, n23162 );
nor U116365 ( n23588, n75398, n23162 );
nor U116366 ( n23543, n75400, n23162 );
nor U116367 ( n23155, n75392, n23162 );
nor U116368 ( n23347, n75393, n23162 );
nor U116369 ( n23766, n75401, n23162 );
nor U116370 ( n23810, n75399, n23162 );
nand U116371 ( n14540, n12828, n73079 );
not U116372 ( n7907, n46668 );
nor U116373 ( n47916, n48315, n48233 );
nand U116374 ( n56330, n56944, n31914 );
nand U116375 ( n67928, n67929, n74872 );
nand U116376 ( n67929, n67899, n67930 );
nand U116377 ( n67930, n67931, n67932 );
nor U116378 ( n67931, n73130, n74852 );
nand U116379 ( n46881, n46882, n74841 );
nand U116380 ( n46882, n46852, n46883 );
nand U116381 ( n46883, n46884, n46885 );
nor U116382 ( n46884, n73118, n74822 );
nand U116383 ( n25925, n25926, n74873 );
nand U116384 ( n25926, n25896, n25927 );
nand U116385 ( n25927, n25928, n25929 );
nor U116386 ( n25928, n73131, n74853 );
nand U116387 ( n59063, n59064, n74874 );
nand U116388 ( n59064, n59034, n59065 );
nand U116389 ( n59065, n59066, n59067 );
nor U116390 ( n59066, n73132, n74854 );
nor U116391 ( n56710, n75375, n56283 );
nor U116392 ( n56754, n75370, n56283 );
nor U116393 ( n56276, n75367, n56283 );
nor U116394 ( n56423, n75366, n56283 );
nor U116395 ( n56471, n75368, n56283 );
nor U116396 ( n56566, n75376, n56283 );
nor U116397 ( n56665, n75374, n56283 );
nor U116398 ( n56799, n75369, n56283 );
nor U116399 ( n56843, n75371, n56283 );
nor U116400 ( n56891, n75373, n56283 );
nor U116401 ( n56935, n75372, n56283 );
nand U116402 ( n13204, n13205, n13154 );
or U116403 ( n13205, n13207, n13158 );
nand U116404 ( n47793, n46779, n73071 );
nor U116405 ( n42549, n42550, n75190 );
nand U116406 ( n25515, n25469, n25497 );
nand U116407 ( n32755, n32709, n32737 );
nand U116408 ( n67520, n67474, n67502 );
nand U116409 ( n58652, n58606, n58634 );
nand U116410 ( n21161, n21209, n8322 );
nand U116411 ( n21209, n4842, n14805 );
nand U116412 ( n46659, n46660, n73159 );
nand U116413 ( n46660, n46631, n46661 );
nand U116414 ( n46661, n46662, n7513 );
nor U116415 ( n46662, n74585, n73148 );
nand U116416 ( n67706, n67707, n74637 );
nand U116417 ( n67707, n67678, n67708 );
nand U116418 ( n67708, n67709, n5727 );
nor U116419 ( n67709, n74595, n73149 );
nand U116420 ( n25701, n25702, n74638 );
nand U116421 ( n25702, n25673, n25703 );
nand U116422 ( n25703, n25704, n3969 );
nor U116423 ( n25704, n74596, n73150 );
nand U116424 ( n58841, n58842, n74639 );
nand U116425 ( n58842, n58813, n58843 );
nand U116426 ( n58843, n58844, n6602 );
nor U116427 ( n58844, n74597, n73151 );
nand U116428 ( n32952, n32953, n75050 );
nand U116429 ( n32953, n32917, n32954 );
nand U116430 ( n32954, n32955, n3125 );
nor U116431 ( n32955, n74652, n73167 );
nand U116432 ( n37608, n2007, n37102 );
nor U116433 ( n42699, n7927, n42700 );
nor U116434 ( n42700, n42701, n42702 );
nor U116435 ( n42701, n42703, n42704 );
nor U116436 ( n8632, n5272, n8633 );
nor U116437 ( n8633, n8634, n8635 );
nor U116438 ( n8634, n8637, n8638 );
not U116439 ( n4395, n22013 );
not U116440 ( n3558, n29332 );
not U116441 ( n6173, n63095 );
not U116442 ( n7028, n55123 );
xor U116443 ( n51671, n53885, n48413 );
not U116444 ( n4298, n26946 );
not U116445 ( n6930, n60086 );
nand U116446 ( n27460, n4283, n27384 );
nand U116447 ( n60609, n6915, n60532 );
nand U116448 ( n27383, n26970, n26973 );
nand U116449 ( n60531, n60110, n60113 );
not U116450 ( n6118, n67715 );
not U116451 ( n4340, n25710 );
not U116452 ( n6973, n58850 );
not U116453 ( n3460, n34191 );
not U116454 ( n6075, n68945 );
nand U116455 ( n34705, n3445, n34629 );
nand U116456 ( n69449, n6060, n69375 );
nand U116457 ( n34628, n34215, n34218 );
nand U116458 ( n69374, n68969, n68972 );
nand U116459 ( n3691, n35430, n35431 );
nor U116460 ( n35430, n35439, n35440 );
nor U116461 ( n35431, n35432, n35433 );
nor U116462 ( n35439, n34283, n35442 );
nand U116463 ( n3851, n35115, n35116 );
nor U116464 ( n35115, n35124, n35125 );
nor U116465 ( n35116, n35117, n35118 );
nor U116466 ( n35124, n34283, n35127 );
nand U116467 ( n10426, n70160, n70161 );
nor U116468 ( n70160, n70169, n70170 );
nor U116469 ( n70161, n70162, n70163 );
nor U116470 ( n70169, n69035, n70172 );
nand U116471 ( n10586, n69851, n69852 );
nor U116472 ( n69851, n69860, n69861 );
nor U116473 ( n69852, n69853, n69854 );
nor U116474 ( n69860, n69035, n69863 );
nand U116475 ( n3686, n35443, n35444 );
nor U116476 ( n35443, n35449, n35450 );
nor U116477 ( n35444, n35445, n35446 );
nor U116478 ( n35450, n34735, n35441 );
nand U116479 ( n3846, n35128, n35129 );
nor U116480 ( n35128, n35134, n35135 );
nor U116481 ( n35129, n35130, n35131 );
nor U116482 ( n35135, n34735, n35126 );
nand U116483 ( n3826, n35160, n35161 );
nor U116484 ( n35160, n35166, n35167 );
nor U116485 ( n35161, n35162, n35163 );
nor U116486 ( n35167, n34771, n35126 );
nand U116487 ( n3666, n35475, n35476 );
nor U116488 ( n35475, n35481, n35482 );
nor U116489 ( n35476, n35477, n35478 );
nor U116490 ( n35482, n34771, n35441 );
nand U116491 ( n3821, n35168, n35169 );
nor U116492 ( n35168, n35174, n35175 );
nor U116493 ( n35169, n35170, n35171 );
nor U116494 ( n35175, n34780, n35126 );
nand U116495 ( n3661, n35483, n35484 );
nor U116496 ( n35483, n35489, n35490 );
nor U116497 ( n35484, n35485, n35486 );
nor U116498 ( n35490, n34780, n35441 );
nand U116499 ( n3656, n35493, n35494 );
nor U116500 ( n35493, n35506, n35507 );
nor U116501 ( n35494, n35495, n35496 );
nor U116502 ( n35507, n34796, n35441 );
nand U116503 ( n3816, n35176, n35177 );
nor U116504 ( n35176, n35189, n35190 );
nor U116505 ( n35177, n35178, n35179 );
nor U116506 ( n35190, n34796, n35126 );
nand U116507 ( n3676, n35459, n35460 );
nor U116508 ( n35459, n35465, n35466 );
nor U116509 ( n35460, n35461, n35462 );
nor U116510 ( n35466, n34753, n35441 );
nand U116511 ( n3836, n35144, n35145 );
nor U116512 ( n35144, n35150, n35151 );
nor U116513 ( n35145, n35146, n35147 );
nor U116514 ( n35151, n34753, n35126 );
nand U116515 ( n3671, n35467, n35468 );
nor U116516 ( n35467, n35473, n35474 );
nor U116517 ( n35468, n35469, n35470 );
nor U116518 ( n35474, n34762, n35441 );
nand U116519 ( n3831, n35152, n35153 );
nor U116520 ( n35152, n35158, n35159 );
nor U116521 ( n35153, n35154, n35155 );
nor U116522 ( n35159, n34762, n35126 );
nand U116523 ( n3841, n35136, n35137 );
nor U116524 ( n35136, n35142, n35143 );
nor U116525 ( n35137, n35138, n35139 );
nor U116526 ( n35143, n34744, n35126 );
nand U116527 ( n10421, n70173, n70174 );
nor U116528 ( n70173, n70179, n70180 );
nor U116529 ( n70174, n70175, n70176 );
nor U116530 ( n70180, n69479, n70171 );
nand U116531 ( n10581, n69864, n69865 );
nor U116532 ( n69864, n69870, n69871 );
nor U116533 ( n69865, n69866, n69867 );
nor U116534 ( n69871, n69479, n69862 );
nand U116535 ( n10576, n69872, n69873 );
nor U116536 ( n69872, n69878, n69879 );
nor U116537 ( n69873, n69874, n69875 );
nor U116538 ( n69879, n69488, n69862 );
nand U116539 ( n10411, n70189, n70190 );
nor U116540 ( n70189, n70195, n70196 );
nor U116541 ( n70190, n70191, n70192 );
nor U116542 ( n70196, n69497, n70171 );
nand U116543 ( n10571, n69880, n69881 );
nor U116544 ( n69880, n69886, n69887 );
nor U116545 ( n69881, n69882, n69883 );
nor U116546 ( n69887, n69497, n69862 );
nand U116547 ( n10556, n69904, n69905 );
nor U116548 ( n69904, n69910, n69911 );
nor U116549 ( n69905, n69906, n69907 );
nor U116550 ( n69911, n69524, n69862 );
nand U116551 ( n10396, n70213, n70214 );
nor U116552 ( n70213, n70219, n70220 );
nor U116553 ( n70214, n70215, n70216 );
nor U116554 ( n70220, n69524, n70171 );
nand U116555 ( n10391, n70221, n70222 );
nor U116556 ( n70221, n70234, n70235 );
nor U116557 ( n70222, n70223, n70224 );
nor U116558 ( n70235, n69540, n70171 );
nand U116559 ( n10551, n69912, n69913 );
nor U116560 ( n69912, n69925, n69926 );
nor U116561 ( n69913, n69914, n69915 );
nor U116562 ( n69926, n69540, n69862 );
nand U116563 ( n10561, n69896, n69897 );
nor U116564 ( n69896, n69902, n69903 );
nor U116565 ( n69897, n69898, n69899 );
nor U116566 ( n69903, n69515, n69862 );
nand U116567 ( n10401, n70205, n70206 );
nor U116568 ( n70205, n70211, n70212 );
nor U116569 ( n70206, n70207, n70208 );
nor U116570 ( n70212, n69515, n70171 );
nand U116571 ( n10406, n70197, n70198 );
nor U116572 ( n70197, n70203, n70204 );
nor U116573 ( n70198, n70199, n70200 );
nor U116574 ( n70204, n69506, n70171 );
nand U116575 ( n10566, n69888, n69889 );
nor U116576 ( n69888, n69894, n69895 );
nor U116577 ( n69889, n69890, n69891 );
nor U116578 ( n69895, n69506, n69862 );
nand U116579 ( n10416, n70181, n70182 );
nor U116580 ( n70181, n70187, n70188 );
nor U116581 ( n70182, n70183, n70184 );
nor U116582 ( n70188, n69488, n70171 );
nand U116583 ( n3681, n35451, n35452 );
nor U116584 ( n35451, n35457, n35458 );
nor U116585 ( n35452, n35453, n35454 );
nor U116586 ( n35458, n34744, n35441 );
nand U116587 ( n35646, n35694, n29195 );
nand U116588 ( n35694, n3097, n34268 );
nand U116589 ( n28467, n28515, n21878 );
nand U116590 ( n28515, n3940, n27023 );
nand U116591 ( n70372, n70420, n62913 );
nand U116592 ( n70420, n5698, n69020 );
nand U116593 ( n61772, n61820, n54969 );
nand U116594 ( n61820, n6573, n60164 );
nand U116595 ( n34234, P1_P3_STATE2_REG_3_, n74611 );
nand U116596 ( n68988, P2_P3_STATE2_REG_3_, n74613 );
not U116597 ( n385, n69052 );
not U116598 ( n390, n69074 );
not U116599 ( n398, n69107 );
not U116600 ( n400, n69131 );
not U116601 ( n395, n69096 );
not U116602 ( n393, n69085 );
not U116603 ( n383, n69041 );
not U116604 ( n388, n69063 );
not U116605 ( n114, n34300 );
not U116606 ( n123, n34344 );
not U116607 ( n125, n34355 );
not U116608 ( n128, n34379 );
not U116609 ( n118, n34322 );
not U116610 ( n120, n34333 );
not U116611 ( n112, n34289 );
not U116612 ( n116, n34311 );
and U116613 ( n68978, n74593, n70311 );
nand U116614 ( n70311, n70312, n68988 );
nand U116615 ( n70312, n69025, n62884 );
and U116616 ( n34224, n74591, n35583 );
nand U116617 ( n35583, n35584, n34234 );
nand U116618 ( n35584, n34273, n29162 );
nand U116619 ( n3766, n35284, n35285 );
nor U116620 ( n35284, n35290, n35291 );
nor U116621 ( n35285, n35286, n35287 );
nor U116622 ( n35290, n34299, n35283 );
nand U116623 ( n3926, n34967, n34968 );
nor U116624 ( n34967, n34973, n34974 );
nor U116625 ( n34968, n34969, n34970 );
nor U116626 ( n34973, n34299, n34966 );
nand U116627 ( n3746, n35318, n35319 );
nor U116628 ( n35318, n35324, n35325 );
nor U116629 ( n35319, n35320, n35321 );
nor U116630 ( n35324, n34343, n35283 );
nand U116631 ( n3906, n35001, n35002 );
nor U116632 ( n35001, n35007, n35008 );
nor U116633 ( n35002, n35003, n35004 );
nor U116634 ( n35007, n34343, n34966 );
nand U116635 ( n3741, n35326, n35327 );
nor U116636 ( n35326, n35332, n35333 );
nor U116637 ( n35327, n35328, n35329 );
nor U116638 ( n35332, n34354, n35283 );
nand U116639 ( n3901, n35009, n35010 );
nor U116640 ( n35009, n35015, n35016 );
nor U116641 ( n35010, n35011, n35012 );
nor U116642 ( n35015, n34354, n34966 );
nand U116643 ( n3736, n35334, n35335 );
nor U116644 ( n35334, n35348, n35349 );
nor U116645 ( n35335, n35336, n35337 );
nor U116646 ( n35348, n34377, n35283 );
nand U116647 ( n3896, n35017, n35018 );
nor U116648 ( n35017, n35031, n35032 );
nor U116649 ( n35018, n35019, n35020 );
nor U116650 ( n35031, n34377, n34966 );
nand U116651 ( n3756, n35302, n35303 );
nor U116652 ( n35302, n35308, n35309 );
nor U116653 ( n35303, n35304, n35305 );
nor U116654 ( n35308, n34321, n35283 );
nand U116655 ( n3916, n34983, n34984 );
nor U116656 ( n34983, n34989, n34990 );
nor U116657 ( n34984, n34985, n34986 );
nor U116658 ( n34989, n34321, n34966 );
nand U116659 ( n3751, n35310, n35311 );
nor U116660 ( n35310, n35316, n35317 );
nor U116661 ( n35311, n35312, n35313 );
nor U116662 ( n35316, n34332, n35283 );
nand U116663 ( n3911, n34991, n34992 );
nor U116664 ( n34991, n34997, n34998 );
nor U116665 ( n34992, n34993, n34994 );
nor U116666 ( n34997, n34332, n34966 );
nand U116667 ( n3731, n35351, n35352 );
nor U116668 ( n35351, n35360, n35361 );
nor U116669 ( n35352, n35353, n35354 );
nor U116670 ( n35360, n34283, n35363 );
nand U116671 ( n3811, n35193, n35194 );
nor U116672 ( n35193, n35202, n35203 );
nor U116673 ( n35194, n35195, n35196 );
nor U116674 ( n35202, n34283, n35205 );
nand U116675 ( n3891, n35035, n35036 );
nor U116676 ( n35035, n35044, n35045 );
nor U116677 ( n35036, n35037, n35038 );
nor U116678 ( n35044, n34283, n35047 );
nand U116679 ( n4011, n34798, n34799 );
nor U116680 ( n34798, n34807, n34808 );
nor U116681 ( n34799, n34800, n34801 );
nor U116682 ( n34807, n34283, n34810 );
nand U116683 ( n4051, n34713, n34714 );
nor U116684 ( n34713, n34722, n34723 );
nor U116685 ( n34714, n34715, n34716 );
nor U116686 ( n34722, n34283, n34726 );
nand U116687 ( n3761, n35292, n35293 );
nor U116688 ( n35292, n35298, n35299 );
nor U116689 ( n35293, n35294, n35295 );
nor U116690 ( n35298, n34310, n35283 );
nand U116691 ( n3921, n34975, n34976 );
nor U116692 ( n34975, n34981, n34982 );
nor U116693 ( n34976, n34977, n34978 );
nor U116694 ( n34981, n34310, n34966 );
nand U116695 ( n10501, n70018, n70019 );
nor U116696 ( n70018, n70024, n70025 );
nor U116697 ( n70019, n70020, n70021 );
nor U116698 ( n70024, n69051, n70017 );
nand U116699 ( n10661, n69707, n69708 );
nor U116700 ( n69707, n69713, n69714 );
nor U116701 ( n69708, n69709, n69710 );
nor U116702 ( n69713, n69051, n69706 );
nand U116703 ( n10496, n70026, n70027 );
nor U116704 ( n70026, n70032, n70033 );
nor U116705 ( n70027, n70028, n70029 );
nor U116706 ( n70032, n69062, n70017 );
nand U116707 ( n10656, n69715, n69716 );
nor U116708 ( n69715, n69721, n69722 );
nor U116709 ( n69716, n69717, n69718 );
nor U116710 ( n69721, n69062, n69706 );
nand U116711 ( n10491, n70034, n70035 );
nor U116712 ( n70034, n70040, n70041 );
nor U116713 ( n70035, n70036, n70037 );
nor U116714 ( n70040, n69073, n70017 );
nand U116715 ( n10651, n69723, n69724 );
nor U116716 ( n69723, n69729, n69730 );
nor U116717 ( n69724, n69725, n69726 );
nor U116718 ( n69729, n69073, n69706 );
nand U116719 ( n10476, n70058, n70059 );
nor U116720 ( n70058, n70064, n70065 );
nor U116721 ( n70059, n70060, n70061 );
nor U116722 ( n70064, n69106, n70017 );
nand U116723 ( n10636, n69747, n69748 );
nor U116724 ( n69747, n69753, n69754 );
nor U116725 ( n69748, n69749, n69750 );
nor U116726 ( n69753, n69106, n69706 );
nand U116727 ( n10471, n70066, n70067 );
nor U116728 ( n70066, n70080, n70081 );
nor U116729 ( n70067, n70068, n70069 );
nor U116730 ( n70080, n69129, n70017 );
nand U116731 ( n10631, n69755, n69756 );
nor U116732 ( n69755, n69769, n69770 );
nor U116733 ( n69756, n69757, n69758 );
nor U116734 ( n69769, n69129, n69706 );
nand U116735 ( n10481, n70050, n70051 );
nor U116736 ( n70050, n70056, n70057 );
nor U116737 ( n70051, n70052, n70053 );
nor U116738 ( n70056, n69095, n70017 );
nand U116739 ( n10641, n69739, n69740 );
nor U116740 ( n69739, n69745, n69746 );
nor U116741 ( n69740, n69741, n69742 );
nor U116742 ( n69745, n69095, n69706 );
nand U116743 ( n10486, n70042, n70043 );
nor U116744 ( n70042, n70048, n70049 );
nor U116745 ( n70043, n70044, n70045 );
nor U116746 ( n70048, n69084, n70017 );
nand U116747 ( n10646, n69731, n69732 );
nor U116748 ( n69731, n69737, n69738 );
nor U116749 ( n69732, n69733, n69734 );
nor U116750 ( n69737, n69084, n69706 );
nand U116751 ( n10466, n70083, n70084 );
nor U116752 ( n70083, n70092, n70093 );
nor U116753 ( n70084, n70085, n70086 );
nor U116754 ( n70092, n69035, n70095 );
nand U116755 ( n10546, n69929, n69930 );
nor U116756 ( n69929, n69938, n69939 );
nor U116757 ( n69930, n69931, n69932 );
nor U116758 ( n69938, n69035, n69941 );
nand U116759 ( n10626, n69773, n69774 );
nor U116760 ( n69773, n69782, n69783 );
nor U116761 ( n69774, n69775, n69776 );
nor U116762 ( n69782, n69035, n69785 );
nand U116763 ( n10746, n69542, n69543 );
nor U116764 ( n69542, n69551, n69552 );
nor U116765 ( n69543, n69544, n69545 );
nor U116766 ( n69551, n69035, n69554 );
nand U116767 ( n10786, n69457, n69458 );
nor U116768 ( n69457, n69466, n69467 );
nor U116769 ( n69458, n69459, n69460 );
nor U116770 ( n69466, n69035, n69470 );
nand U116771 ( n3726, n35364, n35365 );
nor U116772 ( n35364, n35370, n35371 );
nor U116773 ( n35365, n35366, n35367 );
nor U116774 ( n35371, n34735, n35362 );
nand U116775 ( n3806, n35208, n35209 );
nor U116776 ( n35208, n35214, n35215 );
nor U116777 ( n35209, n35210, n35211 );
nor U116778 ( n35215, n34735, n35204 );
nand U116779 ( n3886, n35048, n35049 );
nor U116780 ( n35048, n35054, n35055 );
nor U116781 ( n35049, n35050, n35051 );
nor U116782 ( n35055, n34735, n35046 );
nand U116783 ( n4006, n34813, n34814 );
nor U116784 ( n34813, n34819, n34820 );
nor U116785 ( n34814, n34815, n34816 );
nor U116786 ( n34820, n34735, n34809 );
nand U116787 ( n4046, n34727, n34728 );
nor U116788 ( n34727, n34733, n34734 );
nor U116789 ( n34728, n34729, n34730 );
nor U116790 ( n34734, n34735, n34725 );
nand U116791 ( n3706, n35398, n35399 );
nor U116792 ( n35398, n35404, n35405 );
nor U116793 ( n35399, n35400, n35401 );
nor U116794 ( n35405, n34771, n35362 );
nand U116795 ( n3786, n35240, n35241 );
nor U116796 ( n35240, n35246, n35247 );
nor U116797 ( n35241, n35242, n35243 );
nor U116798 ( n35247, n34771, n35204 );
nand U116799 ( n3866, n35080, n35081 );
nor U116800 ( n35080, n35086, n35087 );
nor U116801 ( n35081, n35082, n35083 );
nor U116802 ( n35087, n34771, n35046 );
nand U116803 ( n3986, n34845, n34846 );
nor U116804 ( n34845, n34851, n34852 );
nor U116805 ( n34846, n34847, n34848 );
nor U116806 ( n34852, n34771, n34809 );
nand U116807 ( n4026, n34763, n34764 );
nor U116808 ( n34763, n34769, n34770 );
nor U116809 ( n34764, n34765, n34766 );
nor U116810 ( n34770, n34771, n34725 );
nand U116811 ( n3701, n35406, n35407 );
nor U116812 ( n35406, n35412, n35413 );
nor U116813 ( n35407, n35408, n35409 );
nor U116814 ( n35413, n34780, n35362 );
nand U116815 ( n3781, n35248, n35249 );
nor U116816 ( n35248, n35254, n35255 );
nor U116817 ( n35249, n35250, n35251 );
nor U116818 ( n35255, n34780, n35204 );
nand U116819 ( n3861, n35088, n35089 );
nor U116820 ( n35088, n35094, n35095 );
nor U116821 ( n35089, n35090, n35091 );
nor U116822 ( n35095, n34780, n35046 );
nand U116823 ( n3981, n34853, n34854 );
nor U116824 ( n34853, n34859, n34860 );
nor U116825 ( n34854, n34855, n34856 );
nor U116826 ( n34860, n34780, n34809 );
nand U116827 ( n4021, n34772, n34773 );
nor U116828 ( n34772, n34778, n34779 );
nor U116829 ( n34773, n34774, n34775 );
nor U116830 ( n34779, n34780, n34725 );
nand U116831 ( n3696, n35414, n35415 );
nor U116832 ( n35414, n35427, n35428 );
nor U116833 ( n35415, n35416, n35417 );
nor U116834 ( n35428, n34796, n35362 );
nand U116835 ( n3776, n35256, n35257 );
nor U116836 ( n35256, n35269, n35270 );
nor U116837 ( n35257, n35258, n35259 );
nor U116838 ( n35270, n34796, n35204 );
nand U116839 ( n3856, n35098, n35099 );
nor U116840 ( n35098, n35111, n35112 );
nor U116841 ( n35099, n35100, n35101 );
nor U116842 ( n35112, n34796, n35046 );
nand U116843 ( n3976, n34861, n34862 );
nor U116844 ( n34861, n34874, n34875 );
nor U116845 ( n34862, n34863, n34864 );
nor U116846 ( n34875, n34796, n34809 );
nand U116847 ( n4016, n34781, n34782 );
nor U116848 ( n34781, n34794, n34795 );
nor U116849 ( n34782, n34783, n34784 );
nor U116850 ( n34795, n34796, n34725 );
nand U116851 ( n3716, n35380, n35381 );
nor U116852 ( n35380, n35386, n35387 );
nor U116853 ( n35381, n35382, n35383 );
nor U116854 ( n35387, n34753, n35362 );
nand U116855 ( n3796, n35224, n35225 );
nor U116856 ( n35224, n35230, n35231 );
nor U116857 ( n35225, n35226, n35227 );
nor U116858 ( n35231, n34753, n35204 );
nand U116859 ( n3876, n35064, n35065 );
nor U116860 ( n35064, n35070, n35071 );
nor U116861 ( n35065, n35066, n35067 );
nor U116862 ( n35071, n34753, n35046 );
nand U116863 ( n3996, n34829, n34830 );
nor U116864 ( n34829, n34835, n34836 );
nor U116865 ( n34830, n34831, n34832 );
nor U116866 ( n34836, n34753, n34809 );
nand U116867 ( n4036, n34745, n34746 );
nor U116868 ( n34745, n34751, n34752 );
nor U116869 ( n34746, n34747, n34748 );
nor U116870 ( n34752, n34753, n34725 );
nand U116871 ( n3711, n35388, n35389 );
nor U116872 ( n35388, n35394, n35395 );
nor U116873 ( n35389, n35390, n35391 );
nor U116874 ( n35395, n34762, n35362 );
nand U116875 ( n3791, n35232, n35233 );
nor U116876 ( n35232, n35238, n35239 );
nor U116877 ( n35233, n35234, n35235 );
nor U116878 ( n35239, n34762, n35204 );
nand U116879 ( n3871, n35072, n35073 );
nor U116880 ( n35072, n35078, n35079 );
nor U116881 ( n35073, n35074, n35075 );
nor U116882 ( n35079, n34762, n35046 );
nand U116883 ( n3991, n34837, n34838 );
nor U116884 ( n34837, n34843, n34844 );
nor U116885 ( n34838, n34839, n34840 );
nor U116886 ( n34844, n34762, n34809 );
nand U116887 ( n4031, n34754, n34755 );
nor U116888 ( n34754, n34760, n34761 );
nor U116889 ( n34755, n34756, n34757 );
nor U116890 ( n34761, n34762, n34725 );
nand U116891 ( n3771, n35271, n35272 );
nor U116892 ( n35271, n35280, n35281 );
nor U116893 ( n35272, n35273, n35274 );
nor U116894 ( n35280, n34287, n35283 );
nand U116895 ( n3931, n34954, n34955 );
nor U116896 ( n34954, n34963, n34964 );
nor U116897 ( n34955, n34956, n34957 );
nor U116898 ( n34963, n34287, n34966 );
nand U116899 ( n3721, n35372, n35373 );
nor U116900 ( n35372, n35378, n35379 );
nor U116901 ( n35373, n35374, n35375 );
nor U116902 ( n35379, n34744, n35362 );
nand U116903 ( n3801, n35216, n35217 );
nor U116904 ( n35216, n35222, n35223 );
nor U116905 ( n35217, n35218, n35219 );
nor U116906 ( n35223, n34744, n35204 );
nand U116907 ( n3881, n35056, n35057 );
nor U116908 ( n35056, n35062, n35063 );
nor U116909 ( n35057, n35058, n35059 );
nor U116910 ( n35063, n34744, n35046 );
nand U116911 ( n4001, n34821, n34822 );
nor U116912 ( n34821, n34827, n34828 );
nor U116913 ( n34822, n34823, n34824 );
nor U116914 ( n34828, n34744, n34809 );
nand U116915 ( n4041, n34736, n34737 );
nor U116916 ( n34736, n34742, n34743 );
nor U116917 ( n34737, n34738, n34739 );
nor U116918 ( n34743, n34744, n34725 );
nand U116919 ( n10461, n70096, n70097 );
nor U116920 ( n70096, n70102, n70103 );
nor U116921 ( n70097, n70098, n70099 );
nor U116922 ( n70103, n69479, n70094 );
nand U116923 ( n10541, n69942, n69943 );
nor U116924 ( n69942, n69948, n69949 );
nor U116925 ( n69943, n69944, n69945 );
nor U116926 ( n69949, n69479, n69940 );
nand U116927 ( n10621, n69786, n69787 );
nor U116928 ( n69786, n69792, n69793 );
nor U116929 ( n69787, n69788, n69789 );
nor U116930 ( n69793, n69479, n69784 );
nand U116931 ( n10741, n69555, n69556 );
nor U116932 ( n69555, n69561, n69562 );
nor U116933 ( n69556, n69557, n69558 );
nor U116934 ( n69562, n69479, n69553 );
nand U116935 ( n10781, n69471, n69472 );
nor U116936 ( n69471, n69477, n69478 );
nor U116937 ( n69472, n69473, n69474 );
nor U116938 ( n69478, n69479, n69469 );
nand U116939 ( n10456, n70104, n70105 );
nor U116940 ( n70104, n70110, n70111 );
nor U116941 ( n70105, n70106, n70107 );
nor U116942 ( n70111, n69488, n70094 );
nand U116943 ( n10536, n69950, n69951 );
nor U116944 ( n69950, n69956, n69957 );
nor U116945 ( n69951, n69952, n69953 );
nor U116946 ( n69957, n69488, n69940 );
nand U116947 ( n10616, n69794, n69795 );
nor U116948 ( n69794, n69800, n69801 );
nor U116949 ( n69795, n69796, n69797 );
nor U116950 ( n69801, n69488, n69784 );
nand U116951 ( n10736, n69563, n69564 );
nor U116952 ( n69563, n69569, n69570 );
nor U116953 ( n69564, n69565, n69566 );
nor U116954 ( n69570, n69488, n69553 );
nand U116955 ( n10776, n69480, n69481 );
nor U116956 ( n69480, n69486, n69487 );
nor U116957 ( n69481, n69482, n69483 );
nor U116958 ( n69487, n69488, n69469 );
nand U116959 ( n10451, n70112, n70113 );
nor U116960 ( n70112, n70118, n70119 );
nor U116961 ( n70113, n70114, n70115 );
nor U116962 ( n70119, n69497, n70094 );
nand U116963 ( n10531, n69958, n69959 );
nor U116964 ( n69958, n69964, n69965 );
nor U116965 ( n69959, n69960, n69961 );
nor U116966 ( n69965, n69497, n69940 );
nand U116967 ( n10611, n69802, n69803 );
nor U116968 ( n69802, n69808, n69809 );
nor U116969 ( n69803, n69804, n69805 );
nor U116970 ( n69809, n69497, n69784 );
nand U116971 ( n10731, n69571, n69572 );
nor U116972 ( n69571, n69577, n69578 );
nor U116973 ( n69572, n69573, n69574 );
nor U116974 ( n69578, n69497, n69553 );
nand U116975 ( n10771, n69489, n69490 );
nor U116976 ( n69489, n69495, n69496 );
nor U116977 ( n69490, n69491, n69492 );
nor U116978 ( n69496, n69497, n69469 );
nand U116979 ( n10436, n70136, n70137 );
nor U116980 ( n70136, n70142, n70143 );
nor U116981 ( n70137, n70138, n70139 );
nor U116982 ( n70143, n69524, n70094 );
nand U116983 ( n10516, n69982, n69983 );
nor U116984 ( n69982, n69988, n69989 );
nor U116985 ( n69983, n69984, n69985 );
nor U116986 ( n69989, n69524, n69940 );
nand U116987 ( n10596, n69826, n69827 );
nor U116988 ( n69826, n69832, n69833 );
nor U116989 ( n69827, n69828, n69829 );
nor U116990 ( n69833, n69524, n69784 );
nand U116991 ( n10716, n69595, n69596 );
nor U116992 ( n69595, n69601, n69602 );
nor U116993 ( n69596, n69597, n69598 );
nor U116994 ( n69602, n69524, n69553 );
nand U116995 ( n10756, n69516, n69517 );
nor U116996 ( n69516, n69522, n69523 );
nor U116997 ( n69517, n69518, n69519 );
nor U116998 ( n69523, n69524, n69469 );
nand U116999 ( n10431, n70144, n70145 );
nor U117000 ( n70144, n70157, n70158 );
nor U117001 ( n70145, n70146, n70147 );
nor U117002 ( n70158, n69540, n70094 );
nand U117003 ( n10511, n69990, n69991 );
nor U117004 ( n69990, n70003, n70004 );
nor U117005 ( n69991, n69992, n69993 );
nor U117006 ( n70004, n69540, n69940 );
nand U117007 ( n10591, n69834, n69835 );
nor U117008 ( n69834, n69847, n69848 );
nor U117009 ( n69835, n69836, n69837 );
nor U117010 ( n69848, n69540, n69784 );
nand U117011 ( n10711, n69603, n69604 );
nor U117012 ( n69603, n69616, n69617 );
nor U117013 ( n69604, n69605, n69606 );
nor U117014 ( n69617, n69540, n69553 );
nand U117015 ( n10751, n69525, n69526 );
nor U117016 ( n69525, n69538, n69539 );
nor U117017 ( n69526, n69527, n69528 );
nor U117018 ( n69539, n69540, n69469 );
nand U117019 ( n10441, n70128, n70129 );
nor U117020 ( n70128, n70134, n70135 );
nor U117021 ( n70129, n70130, n70131 );
nor U117022 ( n70135, n69515, n70094 );
nand U117023 ( n10521, n69974, n69975 );
nor U117024 ( n69974, n69980, n69981 );
nor U117025 ( n69975, n69976, n69977 );
nor U117026 ( n69981, n69515, n69940 );
nand U117027 ( n10601, n69818, n69819 );
nor U117028 ( n69818, n69824, n69825 );
nor U117029 ( n69819, n69820, n69821 );
nor U117030 ( n69825, n69515, n69784 );
nand U117031 ( n10721, n69587, n69588 );
nor U117032 ( n69587, n69593, n69594 );
nor U117033 ( n69588, n69589, n69590 );
nor U117034 ( n69594, n69515, n69553 );
nand U117035 ( n10761, n69507, n69508 );
nor U117036 ( n69507, n69513, n69514 );
nor U117037 ( n69508, n69509, n69510 );
nor U117038 ( n69514, n69515, n69469 );
nand U117039 ( n10446, n70120, n70121 );
nor U117040 ( n70120, n70126, n70127 );
nor U117041 ( n70121, n70122, n70123 );
nor U117042 ( n70127, n69506, n70094 );
nand U117043 ( n10526, n69966, n69967 );
nor U117044 ( n69966, n69972, n69973 );
nor U117045 ( n69967, n69968, n69969 );
nor U117046 ( n69973, n69506, n69940 );
nand U117047 ( n10606, n69810, n69811 );
nor U117048 ( n69810, n69816, n69817 );
nor U117049 ( n69811, n69812, n69813 );
nor U117050 ( n69817, n69506, n69784 );
nand U117051 ( n10726, n69579, n69580 );
nor U117052 ( n69579, n69585, n69586 );
nor U117053 ( n69580, n69581, n69582 );
nor U117054 ( n69586, n69506, n69553 );
nand U117055 ( n10766, n69498, n69499 );
nor U117056 ( n69498, n69504, n69505 );
nor U117057 ( n69499, n69500, n69501 );
nor U117058 ( n69505, n69506, n69469 );
nand U117059 ( n10506, n70005, n70006 );
nor U117060 ( n70005, n70014, n70015 );
nor U117061 ( n70006, n70007, n70008 );
nor U117062 ( n70014, n69039, n70017 );
nand U117063 ( n10666, n69694, n69695 );
nor U117064 ( n69694, n69703, n69704 );
nor U117065 ( n69695, n69696, n69697 );
nor U117066 ( n69703, n69039, n69706 );
nand U117067 ( n43266, n7408, n43267 );
nand U117068 ( n43267, n43268, n74626 );
nand U117069 ( n43326, n7408, n43329 );
nand U117070 ( n43329, n43330, n43331 );
not U117071 ( n408, n69488 );
not U117072 ( n410, n69497 );
not U117073 ( n418, n69524 );
not U117074 ( n415, n69515 );
not U117075 ( n403, n69468 );
not U117076 ( n405, n69479 );
not U117077 ( n143, n34771 );
not U117078 ( n145, n34780 );
not U117079 ( n138, n34753 );
not U117080 ( n135, n34744 );
not U117081 ( n130, n34724 );
not U117082 ( n133, n34735 );
not U117083 ( n140, n34762 );
not U117084 ( n413, n69506 );
not U117085 ( n147, n34796 );
not U117086 ( n419, n69540 );
nand U117087 ( n3626, n35557, n35558 );
nor U117088 ( n35557, n35563, n35564 );
nor U117089 ( n35558, n35559, n35560 );
nor U117090 ( n35563, n34343, n35523 );
nand U117091 ( n3621, n35565, n35566 );
nor U117092 ( n35565, n35571, n35572 );
nor U117093 ( n35566, n35567, n35568 );
nor U117094 ( n35571, n34354, n35523 );
nand U117095 ( n3636, n35540, n35541 );
nor U117096 ( n35540, n35547, n35548 );
nor U117097 ( n35541, n35542, n35543 );
nor U117098 ( n35547, n34321, n35523 );
nand U117099 ( n3631, n35549, n35550 );
nor U117100 ( n35549, n35555, n35556 );
nor U117101 ( n35550, n35551, n35552 );
nor U117102 ( n35555, n34332, n35523 );
nand U117103 ( n3641, n35532, n35533 );
nor U117104 ( n35532, n35538, n35539 );
nor U117105 ( n35533, n35534, n35535 );
nor U117106 ( n35538, n34310, n35523 );
nand U117107 ( n10376, n70260, n70261 );
nor U117108 ( n70260, n70266, n70267 );
nor U117109 ( n70261, n70262, n70263 );
nor U117110 ( n70266, n69062, n70251 );
nand U117111 ( n10371, n70268, n70269 );
nor U117112 ( n70268, n70275, n70276 );
nor U117113 ( n70269, n70270, n70271 );
nor U117114 ( n70275, n69073, n70251 );
nand U117115 ( n10356, n70293, n70294 );
nor U117116 ( n70293, n70299, n70300 );
nor U117117 ( n70294, n70295, n70296 );
nor U117118 ( n70299, n69106, n70251 );
nand U117119 ( n10361, n70285, n70286 );
nor U117120 ( n70285, n70291, n70292 );
nor U117121 ( n70286, n70287, n70288 );
nor U117122 ( n70291, n69095, n70251 );
nand U117123 ( n10366, n70277, n70278 );
nor U117124 ( n70277, n70283, n70284 );
nor U117125 ( n70278, n70279, n70280 );
nor U117126 ( n70283, n69084, n70251 );
nand U117127 ( n3651, n35508, n35509 );
nor U117128 ( n35508, n35520, n35521 );
nor U117129 ( n35509, n35510, n35511 );
nor U117130 ( n35520, n34287, n35523 );
nand U117131 ( n10386, n70236, n70237 );
nor U117132 ( n70236, n70248, n70249 );
nor U117133 ( n70237, n70238, n70239 );
nor U117134 ( n70248, n69039, n70251 );
nand U117135 ( n3616, n35573, n35574 );
nor U117136 ( n35573, n35579, n35580 );
nor U117137 ( n35574, n35575, n35576 );
nor U117138 ( n35580, n34377, n35523 );
nand U117139 ( n3646, n35524, n35525 );
nor U117140 ( n35524, n35530, n35531 );
nor U117141 ( n35525, n35526, n35527 );
nor U117142 ( n35530, n34299, n35523 );
nand U117143 ( n10351, n70301, n70302 );
nor U117144 ( n70301, n70307, n70308 );
nor U117145 ( n70302, n70303, n70304 );
nor U117146 ( n70308, n69129, n70251 );
nand U117147 ( n10381, n70252, n70253 );
nor U117148 ( n70252, n70258, n70259 );
nor U117149 ( n70253, n70254, n70255 );
nor U117150 ( n70258, n69051, n70251 );
or U117151 ( n24329, n24390, n4067 );
or U117152 ( n65911, n66054, n5842 );
or U117153 ( n57452, n57515, n6699 );
xnor U117154 ( n67146, n68361, n68451 );
xor U117155 ( n68451, n74452, n68362 );
xnor U117156 ( n46182, n47329, n47430 );
xor U117157 ( n47430, n74443, n47330 );
xnor U117158 ( n25248, n26360, n26450 );
xor U117159 ( n26450, n74453, n26361 );
xnor U117160 ( n58384, n59499, n59589 );
xor U117161 ( n59589, n74454, n59500 );
nand U117162 ( n27716, n27782, n76517 );
nor U117163 ( n27782, n27783, n27784 );
and U117164 ( n27784, n27717, P1_P2_STATE2_REG_3_ );
nor U117165 ( n27783, n27785, n27786 );
nand U117166 ( n60867, n60930, n76259 );
nor U117167 ( n60930, n60931, n60932 );
and U117168 ( n60932, n60868, P2_P2_STATE2_REG_3_ );
nor U117169 ( n60931, n60933, n60934 );
nand U117170 ( n29169, n76918, n73182 );
nand U117171 ( n21856, n76916, n73181 );
nand U117172 ( n62891, n76914, n73183 );
nand U117173 ( n54947, n76912, n73180 );
nand U117174 ( n34961, n35023, n76461 );
nor U117175 ( n35023, n35024, n35025 );
and U117176 ( n35025, n34962, P1_P3_STATE2_REG_3_ );
nor U117177 ( n35024, n35026, n35027 );
nand U117178 ( n69701, n69761, n76193 );
nor U117179 ( n69761, n69762, n69763 );
and U117180 ( n69763, n69702, P2_P3_STATE2_REG_3_ );
nor U117181 ( n69762, n69764, n69765 );
xnor U117182 ( n32490, n33605, n33695 );
xor U117183 ( n33695, n74455, n33606 );
xnor U117184 ( n12548, n13983, n14078 );
xor U117185 ( n14078, n74461, n13984 );
nand U117186 ( n46700, n46701, n46665 );
or U117187 ( n46701, n46702, n46668 );
nand U117188 ( n58882, n58883, n58847 );
or U117189 ( n58883, n58884, n58850 );
nand U117190 ( n67747, n67748, n67712 );
or U117191 ( n67748, n67749, n67715 );
nand U117192 ( n25742, n25743, n25707 );
or U117193 ( n25743, n25744, n25710 );
nand U117194 ( n32991, n32992, n32958 );
or U117195 ( n32992, n32993, n32961 );
nand U117196 ( n9300, n4763, n9302 );
nand U117197 ( n9302, n9303, n74646 );
nand U117198 ( n9375, n4763, n9379 );
nand U117199 ( n9379, n9380, n9382 );
nand U117200 ( n69784, n69849, n68933 );
and U117201 ( n29402, n75860, n29404 );
or U117202 ( n75860, n29405, n29406 );
and U117203 ( n22083, n75861, n22085 );
or U117204 ( n75861, n22086, n22087 );
and U117205 ( n55193, n75862, n55195 );
or U117206 ( n75862, n55196, n55197 );
nand U117207 ( n4076, n34659, n34660 );
nor U117208 ( n34659, n34665, n34666 );
nor U117209 ( n34660, n34661, n34662 );
nor U117210 ( n34666, n34321, n34641 );
nand U117211 ( n4081, n34651, n34652 );
nor U117212 ( n34651, n34657, n34658 );
nor U117213 ( n34652, n34653, n34654 );
nor U117214 ( n34658, n34310, n34641 );
nand U117215 ( n10816, n69397, n69398 );
nor U117216 ( n69397, n69403, n69404 );
nor U117217 ( n69398, n69399, n69400 );
nor U117218 ( n69404, n69062, n69387 );
nand U117219 ( n10811, n69405, n69406 );
nor U117220 ( n69405, n69411, n69412 );
nor U117221 ( n69406, n69407, n69408 );
nor U117222 ( n69412, n69073, n69387 );
nand U117223 ( n35046, n35113, n34179 );
nand U117224 ( n4086, n34643, n34644 );
nor U117225 ( n34643, n34649, n34650 );
nor U117226 ( n34644, n34645, n34646 );
nor U117227 ( n34650, n34299, n34641 );
nand U117228 ( n4066, n34675, n34676 );
nor U117229 ( n34675, n34681, n34682 );
nor U117230 ( n34676, n34677, n34678 );
nor U117231 ( n34682, n34343, n34641 );
nand U117232 ( n4061, n34683, n34684 );
nor U117233 ( n34683, n34689, n34690 );
nor U117234 ( n34684, n34685, n34686 );
nor U117235 ( n34690, n34354, n34641 );
nor U117236 ( n28196, n4268, n4287 );
nand U117237 ( n35204, n35113, n34200 );
and U117238 ( n63165, n75863, n63167 );
or U117239 ( n75863, n63168, n63169 );
nor U117240 ( n61360, n6900, n6919 );
nand U117241 ( n69940, n69849, n68954 );
nand U117242 ( n4071, n34667, n34668 );
nor U117243 ( n34667, n34673, n34674 );
nor U117244 ( n34668, n34669, n34670 );
nor U117245 ( n34674, n34332, n34641 );
nand U117246 ( n10821, n69389, n69390 );
nor U117247 ( n69389, n69395, n69396 );
nor U117248 ( n69390, n69391, n69392 );
nor U117249 ( n69396, n69051, n69387 );
nand U117250 ( n10801, n69421, n69422 );
nor U117251 ( n69421, n69427, n69428 );
nor U117252 ( n69422, n69423, n69424 );
nor U117253 ( n69428, n69095, n69387 );
nand U117254 ( n4056, n34693, n34694 );
nor U117255 ( n34693, n34710, n34711 );
nor U117256 ( n34694, n34695, n34696 );
nor U117257 ( n34711, n34377, n34641 );
nand U117258 ( n10796, n69429, n69430 );
nor U117259 ( n69429, n69435, n69436 );
nor U117260 ( n69430, n69431, n69432 );
nor U117261 ( n69436, n69106, n69387 );
nand U117262 ( n10806, n69413, n69414 );
nor U117263 ( n69413, n69419, n69420 );
nor U117264 ( n69414, n69415, n69416 );
nor U117265 ( n69420, n69084, n69387 );
nand U117266 ( n10791, n69437, n69438 );
nor U117267 ( n69437, n69454, n69455 );
nor U117268 ( n69438, n69439, n69440 );
nor U117269 ( n69455, n69129, n69387 );
nand U117270 ( n35362, n35429, n34179 );
nor U117271 ( n35429, n3430, n3449 );
nand U117272 ( n70094, n70159, n68933 );
nor U117273 ( n70159, n6045, n6064 );
nand U117274 ( n4091, n34630, n34631 );
nor U117275 ( n34630, n34639, n34640 );
nor U117276 ( n34631, n34632, n34633 );
nor U117277 ( n34640, n34287, n34641 );
nand U117278 ( n10826, n69376, n69377 );
nor U117279 ( n69376, n69385, n69386 );
nor U117280 ( n69377, n69378, n69379 );
nor U117281 ( n69386, n69039, n69387 );
nand U117282 ( n4126, n34561, n34562 );
nor U117283 ( n34561, n34567, n34568 );
nor U117284 ( n34562, n34563, n34564 );
nor U117285 ( n34567, n34299, n34560 );
nand U117286 ( n4166, n34479, n34480 );
nor U117287 ( n34479, n34485, n34486 );
nor U117288 ( n34480, n34481, n34482 );
nor U117289 ( n34485, n34299, n34478 );
nand U117290 ( n4206, n34397, n34398 );
nor U117291 ( n34397, n34403, n34404 );
nor U117292 ( n34398, n34399, n34400 );
nor U117293 ( n34403, n34299, n34394 );
nand U117294 ( n4106, n34595, n34596 );
nor U117295 ( n34595, n34601, n34602 );
nor U117296 ( n34596, n34597, n34598 );
nor U117297 ( n34601, n34343, n34560 );
nand U117298 ( n4146, n34513, n34514 );
nor U117299 ( n34513, n34519, n34520 );
nor U117300 ( n34514, n34515, n34516 );
nor U117301 ( n34519, n34343, n34478 );
nand U117302 ( n4186, n34429, n34430 );
nor U117303 ( n34429, n34435, n34436 );
nor U117304 ( n34430, n34431, n34432 );
nor U117305 ( n34435, n34343, n34394 );
nand U117306 ( n4101, n34603, n34604 );
nor U117307 ( n34603, n34609, n34610 );
nor U117308 ( n34604, n34605, n34606 );
nor U117309 ( n34609, n34354, n34560 );
nand U117310 ( n4141, n34521, n34522 );
nor U117311 ( n34521, n34527, n34528 );
nor U117312 ( n34522, n34523, n34524 );
nor U117313 ( n34527, n34354, n34478 );
nand U117314 ( n4181, n34437, n34438 );
nor U117315 ( n34437, n34443, n34444 );
nor U117316 ( n34438, n34439, n34440 );
nor U117317 ( n34443, n34354, n34394 );
nand U117318 ( n4096, n34611, n34612 );
nor U117319 ( n34611, n34625, n34626 );
nor U117320 ( n34612, n34613, n34614 );
nor U117321 ( n34625, n34377, n34560 );
nand U117322 ( n4136, n34529, n34530 );
nor U117323 ( n34529, n34543, n34544 );
nor U117324 ( n34530, n34531, n34532 );
nor U117325 ( n34543, n34377, n34478 );
nand U117326 ( n4176, n34445, n34446 );
nor U117327 ( n34445, n34460, n34461 );
nor U117328 ( n34446, n34447, n34448 );
nor U117329 ( n34460, n34377, n34394 );
nand U117330 ( n4116, n34577, n34578 );
nor U117331 ( n34577, n34583, n34584 );
nor U117332 ( n34578, n34579, n34580 );
nor U117333 ( n34583, n34321, n34560 );
nand U117334 ( n4156, n34497, n34498 );
nor U117335 ( n34497, n34503, n34504 );
nor U117336 ( n34498, n34499, n34500 );
nor U117337 ( n34503, n34321, n34478 );
nand U117338 ( n4196, n34413, n34414 );
nor U117339 ( n34413, n34419, n34420 );
nor U117340 ( n34414, n34415, n34416 );
nor U117341 ( n34419, n34321, n34394 );
nand U117342 ( n4111, n34585, n34586 );
nor U117343 ( n34585, n34591, n34592 );
nor U117344 ( n34586, n34587, n34588 );
nor U117345 ( n34591, n34332, n34560 );
nand U117346 ( n4151, n34505, n34506 );
nor U117347 ( n34505, n34511, n34512 );
nor U117348 ( n34506, n34507, n34508 );
nor U117349 ( n34511, n34332, n34478 );
nand U117350 ( n4191, n34421, n34422 );
nor U117351 ( n34421, n34427, n34428 );
nor U117352 ( n34422, n34423, n34424 );
nor U117353 ( n34427, n34332, n34394 );
nand U117354 ( n4131, n34548, n34549 );
nor U117355 ( n34548, n34557, n34558 );
nor U117356 ( n34549, n34550, n34551 );
nor U117357 ( n34557, n34287, n34560 );
nand U117358 ( n4171, n34466, n34467 );
nor U117359 ( n34466, n34475, n34476 );
nor U117360 ( n34467, n34468, n34469 );
nor U117361 ( n34475, n34287, n34478 );
nand U117362 ( n4211, n34382, n34383 );
nor U117363 ( n34382, n34391, n34392 );
nor U117364 ( n34383, n34384, n34385 );
nor U117365 ( n34391, n34287, n34394 );
nand U117366 ( n4121, n34569, n34570 );
nor U117367 ( n34569, n34575, n34576 );
nor U117368 ( n34570, n34571, n34572 );
nor U117369 ( n34575, n34310, n34560 );
nand U117370 ( n4161, n34487, n34488 );
nor U117371 ( n34487, n34493, n34494 );
nor U117372 ( n34488, n34489, n34490 );
nor U117373 ( n34493, n34310, n34478 );
nand U117374 ( n4201, n34405, n34406 );
nor U117375 ( n34405, n34411, n34412 );
nor U117376 ( n34406, n34407, n34408 );
nor U117377 ( n34411, n34310, n34394 );
nand U117378 ( n10861, n69309, n69310 );
nor U117379 ( n69309, n69315, n69316 );
nor U117380 ( n69310, n69311, n69312 );
nor U117381 ( n69315, n69051, n69308 );
nand U117382 ( n10901, n69229, n69230 );
nor U117383 ( n69229, n69235, n69236 );
nor U117384 ( n69230, n69231, n69232 );
nor U117385 ( n69235, n69051, n69228 );
nand U117386 ( n10941, n69147, n69148 );
nor U117387 ( n69147, n69153, n69154 );
nor U117388 ( n69148, n69149, n69150 );
nor U117389 ( n69153, n69051, n69146 );
nand U117390 ( n10856, n69317, n69318 );
nor U117391 ( n69317, n69323, n69324 );
nor U117392 ( n69318, n69319, n69320 );
nor U117393 ( n69323, n69062, n69308 );
nand U117394 ( n10896, n69237, n69238 );
nor U117395 ( n69237, n69243, n69244 );
nor U117396 ( n69238, n69239, n69240 );
nor U117397 ( n69243, n69062, n69228 );
nand U117398 ( n10936, n69155, n69156 );
nor U117399 ( n69155, n69161, n69162 );
nor U117400 ( n69156, n69157, n69158 );
nor U117401 ( n69161, n69062, n69146 );
nand U117402 ( n10851, n69325, n69326 );
nor U117403 ( n69325, n69331, n69332 );
nor U117404 ( n69326, n69327, n69328 );
nor U117405 ( n69331, n69073, n69308 );
nand U117406 ( n10891, n69245, n69246 );
nor U117407 ( n69245, n69251, n69252 );
nor U117408 ( n69246, n69247, n69248 );
nor U117409 ( n69251, n69073, n69228 );
nand U117410 ( n10931, n69163, n69164 );
nor U117411 ( n69163, n69169, n69170 );
nor U117412 ( n69164, n69165, n69166 );
nor U117413 ( n69169, n69073, n69146 );
nand U117414 ( n10836, n69349, n69350 );
nor U117415 ( n69349, n69355, n69356 );
nor U117416 ( n69350, n69351, n69352 );
nor U117417 ( n69355, n69106, n69308 );
nand U117418 ( n10876, n69269, n69270 );
nor U117419 ( n69269, n69275, n69276 );
nor U117420 ( n69270, n69271, n69272 );
nor U117421 ( n69275, n69106, n69228 );
nand U117422 ( n10916, n69187, n69188 );
nor U117423 ( n69187, n69193, n69194 );
nor U117424 ( n69188, n69189, n69190 );
nor U117425 ( n69193, n69106, n69146 );
nand U117426 ( n10831, n69357, n69358 );
nor U117427 ( n69357, n69371, n69372 );
nor U117428 ( n69358, n69359, n69360 );
nor U117429 ( n69371, n69129, n69308 );
nand U117430 ( n10871, n69277, n69278 );
nor U117431 ( n69277, n69291, n69292 );
nor U117432 ( n69278, n69279, n69280 );
nor U117433 ( n69291, n69129, n69228 );
nand U117434 ( n10911, n69195, n69196 );
nor U117435 ( n69195, n69210, n69211 );
nor U117436 ( n69196, n69197, n69198 );
nor U117437 ( n69210, n69129, n69146 );
nand U117438 ( n10841, n69341, n69342 );
nor U117439 ( n69341, n69347, n69348 );
nor U117440 ( n69342, n69343, n69344 );
nor U117441 ( n69347, n69095, n69308 );
nand U117442 ( n10881, n69261, n69262 );
nor U117443 ( n69261, n69267, n69268 );
nor U117444 ( n69262, n69263, n69264 );
nor U117445 ( n69267, n69095, n69228 );
nand U117446 ( n10921, n69179, n69180 );
nor U117447 ( n69179, n69185, n69186 );
nor U117448 ( n69180, n69181, n69182 );
nor U117449 ( n69185, n69095, n69146 );
nand U117450 ( n10846, n69333, n69334 );
nor U117451 ( n69333, n69339, n69340 );
nor U117452 ( n69334, n69335, n69336 );
nor U117453 ( n69339, n69084, n69308 );
nand U117454 ( n10886, n69253, n69254 );
nor U117455 ( n69253, n69259, n69260 );
nor U117456 ( n69254, n69255, n69256 );
nor U117457 ( n69259, n69084, n69228 );
nand U117458 ( n10926, n69171, n69172 );
nor U117459 ( n69171, n69177, n69178 );
nor U117460 ( n69172, n69173, n69174 );
nor U117461 ( n69177, n69084, n69146 );
nand U117462 ( n10866, n69296, n69297 );
nor U117463 ( n69296, n69305, n69306 );
nor U117464 ( n69297, n69298, n69299 );
nor U117465 ( n69305, n69039, n69308 );
nand U117466 ( n10906, n69216, n69217 );
nor U117467 ( n69216, n69225, n69226 );
nor U117468 ( n69217, n69218, n69219 );
nor U117469 ( n69225, n69039, n69228 );
nand U117470 ( n10946, n69134, n69135 );
nor U117471 ( n69134, n69143, n69144 );
nor U117472 ( n69135, n69136, n69137 );
nor U117473 ( n69143, n69039, n69146 );
nand U117474 ( n4236, n34312, n34313 );
nor U117475 ( n34312, n34319, n34320 );
nor U117476 ( n34313, n34314, n34315 );
nor U117477 ( n34320, n34286, n34321 );
nand U117478 ( n4241, n34301, n34302 );
nor U117479 ( n34301, n34308, n34309 );
nor U117480 ( n34302, n34303, n34304 );
nor U117481 ( n34309, n34286, n34310 );
nand U117482 ( n10981, n69042, n69043 );
nor U117483 ( n69042, n69049, n69050 );
nor U117484 ( n69043, n69044, n69045 );
nor U117485 ( n69050, n69038, n69051 );
nand U117486 ( n10976, n69053, n69054 );
nor U117487 ( n69053, n69060, n69061 );
nor U117488 ( n69054, n69055, n69056 );
nor U117489 ( n69061, n69038, n69062 );
nand U117490 ( n10971, n69064, n69065 );
nor U117491 ( n69064, n69071, n69072 );
nor U117492 ( n69065, n69066, n69067 );
nor U117493 ( n69072, n69038, n69073 );
nand U117494 ( n4246, n34290, n34291 );
nor U117495 ( n34290, n34297, n34298 );
nor U117496 ( n34291, n34292, n34293 );
nor U117497 ( n34298, n34286, n34299 );
nand U117498 ( n4226, n34334, n34335 );
nor U117499 ( n34334, n34341, n34342 );
nor U117500 ( n34335, n34336, n34337 );
nor U117501 ( n34342, n34286, n34343 );
nand U117502 ( n4221, n34345, n34346 );
nor U117503 ( n34345, n34352, n34353 );
nor U117504 ( n34346, n34347, n34348 );
nor U117505 ( n34353, n34286, n34354 );
nand U117506 ( n4216, n34356, n34357 );
nor U117507 ( n34356, n34375, n34376 );
nor U117508 ( n34357, n34358, n34359 );
nor U117509 ( n34376, n34286, n34377 );
nand U117510 ( n4231, n34323, n34324 );
nor U117511 ( n34323, n34330, n34331 );
nor U117512 ( n34324, n34325, n34326 );
nor U117513 ( n34331, n34286, n34332 );
nand U117514 ( n10956, n69097, n69098 );
nor U117515 ( n69097, n69104, n69105 );
nor U117516 ( n69098, n69099, n69100 );
nor U117517 ( n69105, n69038, n69106 );
nand U117518 ( n10951, n69108, n69109 );
nor U117519 ( n69108, n69127, n69128 );
nor U117520 ( n69109, n69110, n69111 );
nor U117521 ( n69128, n69038, n69129 );
nand U117522 ( n10961, n69086, n69087 );
nor U117523 ( n69086, n69093, n69094 );
nor U117524 ( n69087, n69088, n69089 );
nor U117525 ( n69094, n69038, n69095 );
nand U117526 ( n10966, n69075, n69076 );
nor U117527 ( n69075, n69082, n69083 );
nor U117528 ( n69076, n69077, n69078 );
nor U117529 ( n69083, n69038, n69084 );
nand U117530 ( n4251, n34274, n34275 );
nor U117531 ( n34274, n34284, n34285 );
nor U117532 ( n34275, n34276, n34277 );
nor U117533 ( n34285, n34286, n34287 );
nand U117534 ( n10986, n69026, n69027 );
nor U117535 ( n69026, n69036, n69037 );
nor U117536 ( n69027, n69028, n69029 );
nor U117537 ( n69037, n69038, n69039 );
nand U117538 ( n68335, n68339, n68249 );
nand U117539 ( n68339, n76057, n74452 );
nand U117540 ( n33579, n33583, n33494 );
nand U117541 ( n33583, n76127, n74455 );
nand U117542 ( n47304, n47308, n47218 );
nand U117543 ( n47308, n76100, n74443 );
nand U117544 ( n26334, n26338, n26248 );
nand U117545 ( n26338, n76155, n74453 );
nand U117546 ( n59473, n59477, n59387 );
nand U117547 ( n59477, n76083, n74454 );
nand U117548 ( n54144, n54192, n42404 );
nand U117549 ( n54192, n7484, n48012 );
nand U117550 ( n68893, n76914, n74660 );
nand U117551 ( n34139, n76918, n74662 );
nand U117552 ( n60034, n76912, n74661 );
nand U117553 ( n26894, n76916, n74663 );
xor U117554 ( n68357, n5774, n73066 );
xor U117555 ( n47325, n7562, n73065 );
xor U117556 ( n26356, n4015, n73067 );
xor U117557 ( n59495, n6648, n73068 );
nor U117558 ( n68619, n68620, n74408 );
xor U117559 ( n68620, n68617, n68538 );
nand U117560 ( n48247, n48310, n76325 );
nor U117561 ( n48310, n48311, n48312 );
and U117562 ( n48312, n48253, n76182 );
nor U117563 ( n48311, n48313, n48309 );
nor U117564 ( n26618, n26619, n74409 );
xor U117565 ( n26619, n26616, n26537 );
nor U117566 ( n59760, n59761, n74410 );
xor U117567 ( n59761, n59758, n59679 );
nor U117568 ( n47598, n47599, n74400 );
xor U117569 ( n47599, n47596, n47517 );
nand U117570 ( n67193, n68615, n68616 );
nand U117571 ( n68616, n68537, n68617 );
nor U117572 ( n68615, n68618, n68619 );
nor U117573 ( n68618, n68617, n68621 );
xor U117574 ( n33601, n3175, n73088 );
nand U117575 ( n25295, n26614, n26615 );
nand U117576 ( n26615, n26536, n26616 );
nor U117577 ( n26614, n26617, n26618 );
nor U117578 ( n26617, n26616, n26620 );
nand U117579 ( n58431, n59756, n59757 );
nand U117580 ( n59757, n59678, n59758 );
nor U117581 ( n59756, n59759, n59760 );
nor U117582 ( n59759, n59758, n59762 );
nand U117583 ( n46241, n47594, n47595 );
nand U117584 ( n47595, n47516, n47596 );
nor U117585 ( n47594, n47597, n47598 );
nor U117586 ( n47597, n47596, n47600 );
nor U117587 ( n33863, n33864, n74412 );
xor U117588 ( n33864, n33861, n33782 );
nor U117589 ( n14288, n14289, n74429 );
xor U117590 ( n14289, n14285, n14187 );
nand U117591 ( n32537, n33859, n33860 );
nand U117592 ( n33860, n33781, n33861 );
nor U117593 ( n33859, n33862, n33863 );
nor U117594 ( n33862, n33861, n33865 );
nand U117595 ( n12607, n14283, n14284 );
nand U117596 ( n14284, n14185, n14285 );
nor U117597 ( n14283, n14287, n14288 );
nor U117598 ( n14287, n14285, n14290 );
xor U117599 ( n13978, n4912, n73090 );
or U117600 ( n45026, n45111, n7629 );
nand U117601 ( n48024, n48123, n76325 );
nor U117602 ( n48123, n48124, n48125 );
and U117603 ( n48125, n48026, n76176 );
nor U117604 ( n48124, n48128, n48129 );
nand U117605 ( n20929, n74435, n15389 );
nor U117606 ( n27793, n27384, n4283 );
nor U117607 ( n35034, n34629, n3445 );
nor U117608 ( n69772, n69375, n6060 );
nor U117609 ( n60941, n60532, n6915 );
nor U117610 ( n68715, n68751, n68752 );
nor U117611 ( n68752, n5723, n68753 );
nor U117612 ( n68751, n75054, n68756 );
nor U117613 ( n68753, n68754, n6083 );
nor U117614 ( n33959, n33995, n33996 );
nor U117615 ( n33996, n3123, n33997 );
nor U117616 ( n33995, n75055, n34000 );
nor U117617 ( n33997, n33998, n3468 );
nor U117618 ( n47694, n47730, n47731 );
nor U117619 ( n47731, n7509, n47732 );
nor U117620 ( n47730, n75058, n47735 );
nor U117621 ( n47732, n47733, n7873 );
nor U117622 ( n26714, n26750, n26751 );
nor U117623 ( n26751, n3965, n26752 );
nor U117624 ( n26750, n75056, n26755 );
nor U117625 ( n26752, n26753, n4305 );
nor U117626 ( n59856, n59892, n59893 );
nor U117627 ( n59893, n6598, n59894 );
nor U117628 ( n59892, n75057, n59897 );
nor U117629 ( n59894, n59895, n6938 );
nand U117630 ( n68756, n68757, n74587 );
nand U117631 ( n68757, n5689, n68682 );
nand U117632 ( n34000, n34001, n74588 );
nand U117633 ( n34001, n3088, n33926 );
nand U117634 ( n47735, n47736, n74580 );
nand U117635 ( n47736, n7474, n47661 );
nand U117636 ( n26755, n26756, n74589 );
nand U117637 ( n26756, n3932, n26681 );
nand U117638 ( n59897, n59898, n74590 );
nand U117639 ( n59898, n6564, n59823 );
nand U117640 ( n68087, n68091, n68044 );
nand U117641 ( n68091, n76057, n72950 );
nand U117642 ( n33330, n33334, n33285 );
nand U117643 ( n33334, n76127, n74755 );
nand U117644 ( n26084, n26088, n26041 );
nand U117645 ( n26088, n76155, n72951 );
nand U117646 ( n59225, n59229, n59182 );
nand U117647 ( n59229, n76083, n72952 );
nand U117648 ( n63481, n62812, n63041 );
nand U117649 ( n29582, n29145, n29274 );
nand U117650 ( n47056, n47060, n47009 );
nand U117651 ( n47060, n76100, n72948 );
nand U117652 ( n22261, n21830, n21957 );
nand U117653 ( n55373, n54906, n55069 );
or U117654 ( n11325, n11410, n4975 );
nor U117655 ( n57005, n57006, n57007 );
nor U117656 ( n23881, n23882, n23883 );
and U117657 ( n15179, n15279, n5178 );
and U117658 ( n15279, n14717, n5200 );
nand U117659 ( n28317, n28318, n28319 );
nand U117660 ( n28319, n28283, n27062 );
or U117661 ( n28318, n28288, n27063 );
nand U117662 ( n28360, n28361, n28362 );
nand U117663 ( n28362, n28283, n27095 );
or U117664 ( n28361, n28288, n27096 );
nand U117665 ( n28331, n28332, n28333 );
nand U117666 ( n28333, n28283, n27073 );
or U117667 ( n28332, n28288, n27074 );
nand U117668 ( n61553, n61554, n61555 );
nand U117669 ( n61555, n61505, n60214 );
or U117670 ( n61554, n61510, n60215 );
nand U117671 ( n61637, n61638, n61639 );
nand U117672 ( n61639, n61505, n60239 );
or U117673 ( n61638, n61510, n60240 );
nand U117674 ( n61539, n61540, n61541 );
nand U117675 ( n61541, n61505, n60203 );
or U117676 ( n61540, n61510, n60204 );
nand U117677 ( n61568, n61569, n61570 );
nand U117678 ( n61570, n61505, n60225 );
or U117679 ( n61569, n61510, n60226 );
nand U117680 ( n28346, n28347, n28348 );
nand U117681 ( n28348, n28283, n27084 );
or U117682 ( n28347, n28288, n27085 );
nand U117683 ( n28388, n28389, n28390 );
nand U117684 ( n28390, n28283, n27125 );
or U117685 ( n28389, n28288, n27128 );
nand U117686 ( n61669, n61670, n61671 );
nand U117687 ( n61671, n61505, n60269 );
or U117688 ( n61670, n61510, n60272 );
nand U117689 ( n61525, n61526, n61527 );
nand U117690 ( n61527, n61505, n60192 );
or U117691 ( n61526, n61510, n60193 );
nand U117692 ( n28303, n28304, n28305 );
nand U117693 ( n28305, n28283, n27051 );
or U117694 ( n28304, n28288, n27052 );
nand U117695 ( n14163, n14365, n12732 );
and U117696 ( n64117, n74593, n62812 );
and U117697 ( n30100, n74591, n29145 );
and U117698 ( n22779, n74592, n21830 );
and U117699 ( n55893, n74594, n54906 );
nand U117700 ( n68691, n76708, n67208 );
nand U117701 ( n33935, n76774, n32552 );
nand U117702 ( n47670, n76660, n46256 );
nand U117703 ( n26690, n76754, n25310 );
nand U117704 ( n59832, n76687, n58449 );
nand U117705 ( n42829, n42324, n42617 );
nand U117706 ( n48535, n48617, n47920 );
nor U117707 ( n48617, n7855, n48240 );
nand U117708 ( n12939, n12817, n12940 );
nand U117709 ( n12940, n12775, n74774 );
nor U117710 ( n31107, n75288, n30481 );
nor U117711 ( n65361, n75287, n64640 );
nor U117712 ( n30569, n75327, n30480 );
nor U117713 ( n64728, n75326, n64639 );
nand U117714 ( n28280, n28281, n28282 );
or U117715 ( n28281, n28288, n27039 );
nand U117716 ( n28282, n28283, n27037 );
nand U117717 ( n28374, n28375, n28376 );
or U117718 ( n28375, n28288, n27107 );
nand U117719 ( n28376, n28283, n27106 );
nand U117720 ( n61651, n61652, n61653 );
or U117721 ( n61652, n61510, n60251 );
nand U117722 ( n61653, n61505, n60250 );
nand U117723 ( n61502, n61503, n61504 );
or U117724 ( n61503, n61510, n60180 );
nand U117725 ( n61504, n61505, n60178 );
nand U117726 ( n47498, n47660, n46331 );
nand U117727 ( n68519, n68681, n67395 );
nand U117728 ( n33763, n33925, n32630 );
nand U117729 ( n26518, n26680, n25390 );
nand U117730 ( n59657, n59822, n58527 );
nand U117731 ( n8789, n8264, n8559 );
nand U117732 ( n15070, n15155, n76591 );
nor U117733 ( n15155, n15157, n15158 );
and U117734 ( n15158, n15078, n76192 );
nor U117735 ( n15157, n15159, n15154 );
nand U117736 ( n13530, n13535, n13413 );
nand U117737 ( n13535, n12775, n74468 );
nand U117738 ( n68008, n68012, n67913 );
nand U117739 ( n68012, n67429, n73104 );
nand U117740 ( n33249, n33253, n33159 );
nand U117741 ( n33253, n32664, n74460 );
nand U117742 ( n46973, n46977, n46866 );
nand U117743 ( n46977, n46365, n73099 );
nand U117744 ( n26005, n26009, n25910 );
nand U117745 ( n26009, n25424, n73105 );
nand U117746 ( n59143, n59147, n59048 );
nand U117747 ( n59147, n58561, n73106 );
and U117748 ( n48150, n48239, n47920 );
nor U117749 ( n48239, n48240, n47935 );
nor U117750 ( n8482, n75170, n8414 );
nand U117751 ( n14820, n14935, n76591 );
nor U117752 ( n14935, n14937, n14938 );
and U117753 ( n14938, n14823, n76186 );
nor U117754 ( n14937, n14942, n14943 );
nand U117755 ( n31619, n31719, n31720 );
nand U117756 ( n31719, n3078, n74591 );
nand U117757 ( n31720, n31721, n3099 );
nor U117758 ( n31721, n29193, n31722 );
or U117759 ( n31625, n31646, n3242 );
nor U117760 ( n31640, n74817, n31625 );
nor U117761 ( n31632, n74876, n31625 );
nor U117762 ( n31644, n75421, n31625 );
nor U117763 ( n31636, n75422, n31625 );
nor U117764 ( n31622, n75447, n31625 );
nor U117765 ( n16614, n16463, n74243 );
nor U117766 ( n16540, n16463, n74111 );
nor U117767 ( n16578, n16463, n74143 );
nor U117768 ( n16650, n16463, n74297 );
nor U117769 ( n16462, n16463, n74019 );
nor U117770 ( n16504, n16463, n73998 );
nor U117771 ( n16688, n16463, n74333 );
not U117772 ( n6513, n60062 );
not U117773 ( n3880, n26922 );
not U117774 ( n3037, n34167 );
not U117775 ( n5638, n68921 );
nand U117776 ( n13276, n60067, n60068 );
nor U117777 ( n60068, n60069, n60070 );
nor U117778 ( n60067, n60077, n60078 );
nor U117779 ( n60069, n6515, n60076 );
nand U117780 ( n6541, n26927, n26928 );
nor U117781 ( n26928, n26929, n26930 );
nor U117782 ( n26927, n26937, n26938 );
nor U117783 ( n26929, n3883, n26936 );
nand U117784 ( n4296, n34172, n34173 );
nor U117785 ( n34173, n34174, n34175 );
nor U117786 ( n34172, n34182, n34183 );
nor U117787 ( n34174, n3039, n34181 );
nand U117788 ( n11031, n68926, n68927 );
nor U117789 ( n68927, n68928, n68929 );
nor U117790 ( n68926, n68936, n68937 );
nor U117791 ( n68928, n5640, n68935 );
nand U117792 ( n13266, n60097, n60098 );
nor U117793 ( n60097, n60111, n60112 );
nor U117794 ( n60098, n60099, n60100 );
nor U117795 ( n60111, n76912, n60113 );
nand U117796 ( n6531, n26957, n26958 );
nor U117797 ( n26957, n26971, n26972 );
nor U117798 ( n26958, n26959, n26960 );
nor U117799 ( n26971, n76916, n26973 );
nand U117800 ( n4286, n34202, n34203 );
nor U117801 ( n34202, n34216, n34217 );
nor U117802 ( n34203, n34204, n34205 );
nor U117803 ( n34216, n76918, n34218 );
nand U117804 ( n11021, n68956, n68957 );
nor U117805 ( n68956, n68970, n68971 );
nor U117806 ( n68957, n68958, n68959 );
nor U117807 ( n68970, n76914, n68972 );
nor U117808 ( n13203, n73158, n13152 );
nand U117809 ( n15412, n15503, n14690 );
nor U117810 ( n15503, n5200, n14734 );
nor U117811 ( n34292, n34282, n34296 );
nor U117812 ( n34336, n34282, n34340 );
nor U117813 ( n34347, n34282, n34351 );
nor U117814 ( n34358, n34282, n34372 );
nor U117815 ( n34314, n34282, n34318 );
nor U117816 ( n34325, n34282, n34329 );
nor U117817 ( n34303, n34282, n34307 );
nor U117818 ( n69044, n69034, n69048 );
nor U117819 ( n69055, n69034, n69059 );
nor U117820 ( n69066, n69034, n69070 );
nor U117821 ( n69099, n69034, n69103 );
nor U117822 ( n69110, n69034, n69124 );
nor U117823 ( n69088, n69034, n69092 );
nor U117824 ( n69077, n69034, n69081 );
nor U117825 ( n48237, n7860, n74442 );
nand U117826 ( n47934, n74442, n7859 );
nor U117827 ( n47921, n48319, n48237 );
nor U117828 ( n60063, n60066, n74424 );
nor U117829 ( n60066, n6513, n58486 );
nor U117830 ( n26923, n26926, n74423 );
nor U117831 ( n26926, n3880, n25347 );
nor U117832 ( n34168, n34171, n74426 );
nor U117833 ( n34171, n3037, n32589 );
nor U117834 ( n68922, n68925, n74425 );
nor U117835 ( n68925, n5638, n67354 );
nand U117836 ( n3936, n34938, n34939 );
nor U117837 ( n34939, n34940, n34941 );
nor U117838 ( n34938, n34952, n34953 );
nand U117839 ( n34941, n34942, n34943 );
nand U117840 ( n3956, n34906, n34907 );
nor U117841 ( n34907, n34908, n34909 );
nor U117842 ( n34906, n34912, n34913 );
nand U117843 ( n34909, n34910, n34911 );
nand U117844 ( n3961, n34896, n34897 );
nor U117845 ( n34897, n34898, n34899 );
nor U117846 ( n34896, n34902, n34903 );
nand U117847 ( n34899, n34900, n34901 );
nand U117848 ( n10696, n69638, n69639 );
nor U117849 ( n69639, n69640, n69641 );
nor U117850 ( n69638, n69644, n69645 );
nand U117851 ( n69641, n69642, n69643 );
nand U117852 ( n10691, n69646, n69647 );
nor U117853 ( n69647, n69648, n69649 );
nor U117854 ( n69646, n69652, n69653 );
nand U117855 ( n69649, n69650, n69651 );
nand U117856 ( n10671, n69678, n69679 );
nor U117857 ( n69679, n69680, n69681 );
nor U117858 ( n69678, n69692, n69693 );
nand U117859 ( n69681, n69682, n69683 );
nand U117860 ( n3966, n34888, n34889 );
nor U117861 ( n34889, n34890, n34891 );
nor U117862 ( n34888, n34894, n34895 );
nand U117863 ( n34891, n34892, n34893 );
nand U117864 ( n3946, n34922, n34923 );
nor U117865 ( n34923, n34924, n34925 );
nor U117866 ( n34922, n34928, n34929 );
nand U117867 ( n34925, n34926, n34927 );
nand U117868 ( n3941, n34930, n34931 );
nor U117869 ( n34931, n34932, n34933 );
nor U117870 ( n34930, n34936, n34937 );
nand U117871 ( n34933, n34934, n34935 );
nand U117872 ( n10701, n69630, n69631 );
nor U117873 ( n69631, n69632, n69633 );
nor U117874 ( n69630, n69636, n69637 );
nand U117875 ( n69633, n69634, n69635 );
nand U117876 ( n10676, n69670, n69671 );
nor U117877 ( n69671, n69672, n69673 );
nor U117878 ( n69670, n69676, n69677 );
nand U117879 ( n69673, n69674, n69675 );
nand U117880 ( n10681, n69662, n69663 );
nor U117881 ( n69663, n69664, n69665 );
nor U117882 ( n69662, n69668, n69669 );
nand U117883 ( n69665, n69666, n69667 );
nand U117884 ( n3951, n34914, n34915 );
nor U117885 ( n34915, n34916, n34917 );
nor U117886 ( n34914, n34920, n34921 );
nand U117887 ( n34917, n34918, n34919 );
nand U117888 ( n10686, n69654, n69655 );
nor U117889 ( n69655, n69656, n69657 );
nor U117890 ( n69654, n69660, n69661 );
nand U117891 ( n69657, n69658, n69659 );
and U117892 ( n14968, n15060, n14690 );
nor U117893 ( n15060, n14734, n15062 );
nor U117894 ( n67746, n73149, n67710 );
nor U117895 ( n46699, n73148, n46663 );
nor U117896 ( n25741, n73150, n25705 );
nor U117897 ( n58881, n73151, n58845 );
not U117898 ( n4819, n8319 );
not U117899 ( n7463, n42402 );
nor U117900 ( n32990, n73167, n32956 );
nand U117901 ( n13314, n13258, n12732 );
nor U117902 ( n13307, n13313, n13314 );
nor U117903 ( n27267, n27085, n27232 );
nor U117904 ( n60410, n60226, n60377 );
nor U117905 ( n27241, n27052, n27232 );
nor U117906 ( n27299, n27128, n27232 );
nor U117907 ( n27275, n27096, n27232 );
nor U117908 ( n60418, n60240, n60377 );
nor U117909 ( n60386, n60193, n60377 );
nor U117910 ( n60442, n60272, n60377 );
nor U117911 ( n27259, n27074, n27232 );
nor U117912 ( n27251, n27063, n27232 );
nor U117913 ( n60402, n60215, n60377 );
nor U117914 ( n60394, n60204, n60377 );
nor U117915 ( n34993, n34329, n34962 );
nor U117916 ( n69733, n69081, n69702 );
nor U117917 ( n34969, n34296, n34962 );
nor U117918 ( n35003, n34340, n34962 );
nor U117919 ( n35011, n34351, n34962 );
nor U117920 ( n35019, n34372, n34962 );
nor U117921 ( n69709, n69048, n69702 );
nor U117922 ( n69749, n69103, n69702 );
nor U117923 ( n69757, n69124, n69702 );
nor U117924 ( n69741, n69092, n69702 );
nor U117925 ( n34985, n34318, n34962 );
nor U117926 ( n34977, n34307, n34962 );
nor U117927 ( n69717, n69059, n69702 );
nor U117928 ( n69725, n69070, n69702 );
nor U117929 ( n48315, n74442, n48130 );
nor U117930 ( n34512, n34329, n34477 );
nor U117931 ( n69260, n69081, n69227 );
nor U117932 ( n34486, n34296, n34477 );
nor U117933 ( n34520, n34340, n34477 );
nor U117934 ( n34528, n34351, n34477 );
nor U117935 ( n34544, n34372, n34477 );
nor U117936 ( n69236, n69048, n69227 );
nor U117937 ( n69276, n69103, n69227 );
nor U117938 ( n69292, n69124, n69227 );
nor U117939 ( n69268, n69092, n69227 );
nor U117940 ( n34504, n34318, n34477 );
nor U117941 ( n34494, n34307, n34477 );
nor U117942 ( n69244, n69059, n69227 );
nor U117943 ( n69252, n69070, n69227 );
nor U117944 ( n63143, n63070, n74848 );
nor U117945 ( n63195, n63070, n74805 );
nor U117946 ( n63362, n63070, n74687 );
nor U117947 ( n29380, n29303, n74849 );
nor U117948 ( n29432, n29303, n74804 );
nor U117949 ( n29533, n29303, n74688 );
nor U117950 ( n22061, n21988, n74850 );
nor U117951 ( n22214, n21988, n74689 );
nor U117952 ( n22113, n21988, n74806 );
nor U117953 ( n55171, n55098, n74851 );
nor U117954 ( n55328, n55098, n74690 );
nor U117955 ( n21977, n21988, n75186 );
nor U117956 ( n55223, n55098, n74807 );
nor U117957 ( n29292, n29303, n75185 );
nor U117958 ( n63059, n63070, n75188 );
nor U117959 ( n55087, n55098, n75187 );
and U117960 ( n49461, n51662, n76325 );
nor U117961 ( n51662, n51663, n51664 );
nor U117962 ( n51664, n7850, n7457 );
nor U117963 ( n51663, n51666, n51667 );
nor U117964 ( n51661, n49461, n74132 );
nand U117965 ( n46789, n46741, n46331 );
nand U117966 ( n33080, n33033, n32630 );
nand U117967 ( n67836, n67788, n67395 );
nand U117968 ( n25833, n25785, n25390 );
nand U117969 ( n58971, n58923, n58527 );
nor U117970 ( n67830, n67835, n67836 );
nor U117971 ( n33074, n33079, n33080 );
nor U117972 ( n46783, n46788, n46789 );
nor U117973 ( n25827, n25832, n25833 );
nor U117974 ( n58965, n58970, n58971 );
nor U117975 ( n15162, n74435, n5208 );
nor U117976 ( n21114, n15162, n15053 );
not U117977 ( n5208, n15389 );
nand U117978 ( n42682, n42683, n42433 );
nand U117979 ( n42683, n900, n42432 );
nor U117980 ( n42679, n42680, n42681 );
nor U117981 ( n42680, n42684, n42685 );
nor U117982 ( n42681, n897, n42682 );
nand U117983 ( n42685, n42686, n42432 );
nor U117984 ( n47895, n47896, n47884 );
nor U117985 ( n47896, n47897, n43348 );
nor U117986 ( n14668, n14669, n14654 );
nor U117987 ( n14669, n14670, n9402 );
xor U117988 ( n68461, n74452, n68369 );
xor U117989 ( n47440, n74443, n47337 );
xor U117990 ( n26460, n74453, n26368 );
xor U117991 ( n59599, n74454, n59507 );
xor U117992 ( n33705, n74455, n33613 );
xor U117993 ( n14090, n74461, n13969 );
nand U117994 ( n34228, n34269, n34270 );
nand U117995 ( n34270, P1_P3_STATE2_REG_3_, n74591 );
nor U117996 ( n34269, n34223, n34271 );
nor U117997 ( n34271, n189, n29193 );
nand U117998 ( n26983, n27024, n27025 );
nand U117999 ( n27025, P1_P2_STATE2_REG_3_, n74592 );
nor U118000 ( n27024, n26978, n27026 );
nor U118001 ( n27026, n152, n21876 );
nand U118002 ( n68982, n69021, n69022 );
nand U118003 ( n69022, P2_P3_STATE2_REG_3_, n74593 );
nor U118004 ( n69021, n68977, n69023 );
nor U118005 ( n69023, n460, n62911 );
nand U118006 ( n60126, n60165, n60166 );
nand U118007 ( n60166, P2_P2_STATE2_REG_3_, n74594 );
nor U118008 ( n60165, n60118, n60167 );
nor U118009 ( n60167, n424, n54967 );
nor U118010 ( n63037, n75179, n63041 );
nor U118011 ( n29270, n75180, n29274 );
nor U118012 ( n21953, n75178, n21957 );
nor U118013 ( n55065, n75177, n55069 );
nand U118014 ( n47974, n48013, n48014 );
nand U118015 ( n48014, n76176, n74648 );
nor U118016 ( n48013, n47969, n48015 );
nor U118017 ( n48015, n494, n42402 );
nand U118018 ( n14752, n14807, n14808 );
nand U118019 ( n14808, n76186, n74649 );
nor U118020 ( n14807, n14745, n14809 );
nor U118021 ( n14809, n223, n8319 );
and U118022 ( n34267, n34228, n34268 );
and U118023 ( n27022, n26983, n27023 );
and U118024 ( n69019, n68982, n69020 );
and U118025 ( n60163, n60126, n60164 );
nor U118026 ( n62610, n74827, n76234 );
nor U118027 ( n62695, n74925, n76233 );
nor U118028 ( n62707, n74969, n76233 );
nor U118029 ( n62622, n74882, n76234 );
nor U118030 ( n62719, n73295, n76233 );
nor U118031 ( n62723, n75000, n76233 );
nor U118032 ( n62614, n74837, n76234 );
nor U118033 ( n62626, n74898, n76234 );
nor U118034 ( n62699, n74938, n76233 );
nor U118035 ( n62711, n74990, n76233 );
nor U118036 ( n62790, n73316, n76233 );
nor U118037 ( n62794, n75063, n76233 );
nor U118038 ( n62598, n74788, n76234 );
nor U118039 ( n62534, n74747, n76234 );
nor U118040 ( n62618, n73247, n76234 );
nor U118041 ( n62691, n73261, n76233 );
nor U118042 ( n62703, n73275, n76233 );
nor U118043 ( n62715, n73290, n76233 );
nor U118044 ( n62530, n73198, n76234 );
nor U118045 ( n62606, n73233, n76234 );
nor U118046 ( n62594, n74743, n76234 );
nor U118047 ( n62727, n75300, n76233 );
nor U118048 ( n62590, n73214, n76234 );
nor U118049 ( n62602, n74798, n76234 );
nand U118050 ( n12987, n12992, n12993 );
nand U118051 ( n12992, n12732, n74653 );
and U118052 ( n48011, n47974, n48012 );
and U118053 ( n14804, n14752, n14805 );
nor U118054 ( n28368, n28296, n73908 );
nor U118055 ( n61645, n61518, n73909 );
nor U118056 ( n35521, n35522, n74002 );
nor U118057 ( n28295, n28296, n73661 );
nor U118058 ( n70249, n70250, n73659 );
nor U118059 ( n28382, n28296, n74058 );
nor U118060 ( n61659, n61518, n74057 );
nor U118061 ( n61517, n61518, n73660 );
nand U118062 ( n60072, n6543, n60062 );
nand U118063 ( n26932, n3910, n26922 );
nand U118064 ( n34177, n3067, n34167 );
nand U118065 ( n68931, n5668, n68921 );
nor U118066 ( n35564, n35522, n74262 );
nor U118067 ( n35572, n35522, n74304 );
nor U118068 ( n35548, n35522, n74107 );
nor U118069 ( n35556, n35522, n74224 );
nor U118070 ( n35539, n35522, n74048 );
nor U118071 ( n28325, n28296, n73748 );
nor U118072 ( n28340, n28296, n73759 );
nor U118073 ( n70267, n70250, n73746 );
nor U118074 ( n70276, n70250, n73758 );
nor U118075 ( n70300, n70250, n74056 );
nor U118076 ( n70292, n70250, n73907 );
nor U118077 ( n61562, n61518, n73760 );
nor U118078 ( n70284, n70250, n73840 );
nor U118079 ( n61547, n61518, n73747 );
nor U118080 ( n61533, n61518, n73634 );
nor U118081 ( n28311, n28296, n73635 );
nor U118082 ( n61576, n61518, n73842 );
nor U118083 ( n28354, n28296, n73841 );
nor U118084 ( n35531, n35522, n73969 );
nor U118085 ( n70259, n70250, n73628 );
nor U118086 ( n29095, n74970, n76502 );
nor U118087 ( n29079, n74926, n76502 );
nor U118088 ( n29067, n74883, n76503 );
nor U118089 ( n29055, n74828, n76503 );
nor U118090 ( n29107, n73294, n76502 );
nor U118091 ( n29111, n74999, n76502 );
nor U118092 ( n29099, n74991, n76502 );
nor U118093 ( n29083, n74939, n76502 );
nor U118094 ( n29071, n74899, n76503 );
nor U118095 ( n29059, n74838, n76503 );
nor U118096 ( n29119, n73317, n76502 );
nor U118097 ( n29123, n75064, n76502 );
nor U118098 ( n34276, n34282, n34283 );
nor U118099 ( n69028, n69034, n69035 );
nor U118100 ( n54794, n74860, n76303 );
nor U118101 ( n54833, n74951, n76302 );
nor U118102 ( n54845, n74995, n76302 );
nor U118103 ( n54806, n74904, n76303 );
nor U118104 ( n54857, n73308, n76302 );
nor U118105 ( n29039, n74789, n76503 );
nor U118106 ( n29027, n74748, n76503 );
nor U118107 ( n29103, n73291, n76502 );
nor U118108 ( n29091, n73276, n76502 );
nor U118109 ( n29075, n73262, n76502 );
nor U118110 ( n29063, n73248, n76503 );
nor U118111 ( n29051, n73234, n76503 );
nor U118112 ( n29035, n74744, n76503 );
nor U118113 ( n29023, n73199, n76503 );
not U118114 ( n1788, n45750 );
not U118115 ( n2904, n38147 );
nor U118116 ( n54861, n75014, n76302 );
nor U118117 ( n29115, n75301, n76502 );
nor U118118 ( n54798, n74868, n76303 );
nor U118119 ( n54825, n74914, n76303 );
nor U118120 ( n54837, n74958, n76302 );
nor U118121 ( n54849, n75005, n76302 );
nor U118122 ( n54884, n73391, n76302 );
nor U118123 ( n56323, n75326, n56330 );
nor U118124 ( n29031, n73215, n76503 );
nor U118125 ( n29047, n74799, n76503 );
nor U118126 ( n54888, n75237, n76302 );
nor U118127 ( n54782, n74811, n76303 );
nor U118128 ( n54766, n75965, n76303 );
nor U118129 ( n54802, n73253, n76303 );
nor U118130 ( n54829, n73267, n76302 );
nor U118131 ( n54841, n73280, n76302 );
nor U118132 ( n54853, n73304, n76302 );
nor U118133 ( n54790, n73239, n76303 );
nor U118134 ( n54747, n73206, n76303 );
nor U118135 ( n54778, n74769, n76303 );
nor U118136 ( n54880, n75302, n76302 );
nor U118137 ( n54770, n73221, n76303 );
nor U118138 ( n54786, n74815, n76303 );
nor U118139 ( n42672, n898, n42673 );
not U118140 ( n898, n42675 );
nand U118141 ( n42673, n42674, n42425 );
nand U118142 ( n42674, n902, n42424 );
nor U118143 ( n62514, n72960, n76234 );
nor U118144 ( n62518, n74640, n76234 );
nor U118145 ( n62522, n74693, n76233 );
nand U118146 ( n3971, n34877, n34878 );
nor U118147 ( n34878, n34879, n34880 );
nor U118148 ( n34877, n34885, n34886 );
nand U118149 ( n34880, n34881, n34882 );
nand U118150 ( n10706, n69619, n69620 );
nor U118151 ( n69620, n69621, n69622 );
nor U118152 ( n69619, n69627, n69628 );
nand U118153 ( n69622, n69623, n69624 );
nor U118154 ( n62510, n74619, n76233 );
nor U118155 ( n62506, n72959, n76233 );
nor U118156 ( n62526, n74709, n76234 );
nor U118157 ( n28396, n28296, n74178 );
nor U118158 ( n61677, n61518, n74179 );
nor U118159 ( n35579, n35522, n74341 );
nor U118160 ( n70307, n70250, n74177 );
nor U118161 ( n29007, n72961, n76503 );
nor U118162 ( n27283, n27107, n27232 );
nor U118163 ( n27231, n27039, n27232 );
nor U118164 ( n60426, n60251, n60377 );
nor U118165 ( n60376, n60180, n60377 );
nor U118166 ( n29011, n74641, n76503 );
nor U118167 ( n29015, n74694, n76502 );
nor U118168 ( n34956, n34283, n34962 );
nor U118169 ( n69696, n69035, n69702 );
nor U118170 ( n69632, n69479, n6047 );
nor U118171 ( n69640, n69488, n6047 );
nor U118172 ( n69648, n69497, n6047 );
nor U118173 ( n69672, n69524, n6047 );
nor U118174 ( n69664, n69515, n6047 );
nor U118175 ( n69621, n69468, n6047 );
nor U118176 ( n34890, n34735, n3432 );
nor U118177 ( n34924, n34771, n3432 );
nor U118178 ( n34932, n34780, n3432 );
nor U118179 ( n34908, n34753, n3432 );
nor U118180 ( n34879, n34724, n3432 );
nor U118181 ( n34898, n34744, n3432 );
nor U118182 ( n34940, n34796, n3432 );
nor U118183 ( n34916, n34762, n3432 );
nor U118184 ( n69680, n69540, n6047 );
nor U118185 ( n69656, n69506, n6047 );
nor U118186 ( n29003, n74620, n76502 );
nor U118187 ( n28995, n72958, n76502 );
nor U118188 ( n54731, n72964, n76302 );
nor U118189 ( n29019, n74710, n76503 );
nor U118190 ( n21755, n74905, n76562 );
nor U118191 ( n23202, n23209, n75327 );
nor U118192 ( n21743, n74861, n76562 );
nor U118193 ( n21781, n74996, n76561 );
nor U118194 ( n21767, n74952, n76561 );
nor U118195 ( n21793, n73309, n76561 );
nor U118196 ( n21797, n75015, n76561 );
nor U118197 ( n21809, n75238, n76561 );
nor U118198 ( n21747, n74869, n76562 );
nor U118199 ( n21759, n74915, n76562 );
nor U118200 ( n21785, n75006, n76561 );
nor U118201 ( n21773, n74959, n76561 );
nor U118202 ( n21731, n74812, n76562 );
nor U118203 ( n54735, n74672, n76302 );
nor U118204 ( n21719, n75967, n76562 );
nor U118205 ( n21805, n73392, n76561 );
nor U118206 ( n54739, n74726, n76303 );
nor U118207 ( n21751, n73254, n76562 );
nor U118208 ( n21763, n73268, n76561 );
nor U118209 ( n21789, n73305, n76561 );
nor U118210 ( n21777, n73281, n76561 );
nor U118211 ( n21739, n73240, n76562 );
nor U118212 ( n21727, n74770, n76562 );
nor U118213 ( n21715, n73207, n76562 );
nor U118214 ( n21801, n75303, n76561 );
nor U118215 ( n21723, n73222, n76562 );
nor U118216 ( n21735, n74816, n76562 );
nor U118217 ( n70025, n69479, n70016 );
nor U118218 ( n69714, n69479, n69705 );
nor U118219 ( n70033, n69488, n70016 );
nor U118220 ( n69722, n69488, n69705 );
nor U118221 ( n70041, n69497, n70016 );
nor U118222 ( n69730, n69497, n69705 );
nor U118223 ( n70065, n69524, n70016 );
nor U118224 ( n69754, n69524, n69705 );
nor U118225 ( n70057, n69515, n70016 );
nor U118226 ( n69746, n69515, n69705 );
nor U118227 ( n70170, n69468, n70171 );
nor U118228 ( n70093, n69468, n70094 );
nor U118229 ( n70015, n69468, n70016 );
nor U118230 ( n69939, n69468, n69940 );
nor U118231 ( n69861, n69468, n69862 );
nor U118232 ( n69783, n69468, n69784 );
nor U118233 ( n69704, n69468, n69705 );
nor U118234 ( n69552, n69468, n69553 );
nor U118235 ( n69467, n69468, n69469 );
nor U118236 ( n34476, n34283, n34477 );
nor U118237 ( n69226, n69035, n69227 );
nor U118238 ( n35291, n34735, n35282 );
nor U118239 ( n34974, n34735, n34965 );
nor U118240 ( n35325, n34771, n35282 );
nor U118241 ( n35008, n34771, n34965 );
nor U118242 ( n35333, n34780, n35282 );
nor U118243 ( n35016, n34780, n34965 );
nor U118244 ( n35309, n34753, n35282 );
nor U118245 ( n34990, n34753, n34965 );
nor U118246 ( n35440, n34724, n35441 );
nor U118247 ( n35361, n34724, n35362 );
nor U118248 ( n35281, n34724, n35282 );
nor U118249 ( n35203, n34724, n35204 );
nor U118250 ( n35125, n34724, n35126 );
nor U118251 ( n35045, n34724, n35046 );
nor U118252 ( n34964, n34724, n34965 );
nor U118253 ( n34808, n34724, n34809 );
nor U118254 ( n34723, n34724, n34725 );
nor U118255 ( n35299, n34744, n35282 );
nor U118256 ( n34982, n34744, n34965 );
nor U118257 ( n35349, n34796, n35282 );
nor U118258 ( n35032, n34796, n34965 );
nor U118259 ( n35317, n34762, n35282 );
nor U118260 ( n34998, n34762, n34965 );
nor U118261 ( n70081, n69540, n70016 );
nor U118262 ( n69770, n69540, n69705 );
nor U118263 ( n70049, n69506, n70016 );
nor U118264 ( n69738, n69506, n69705 );
nor U118265 ( n54727, n74655, n76303 );
nor U118266 ( n54723, n72962, n76303 );
nor U118267 ( n54743, n74728, n76302 );
not U118268 ( n5834, n68552 );
not U118269 ( n7622, n47531 );
not U118270 ( n4063, n26551 );
not U118271 ( n6695, n59693 );
nor U118272 ( n68626, n5819, n68628 );
nor U118273 ( n68628, n68629, n5834 );
nor U118274 ( n26625, n4050, n26627 );
nor U118275 ( n26627, n26628, n4063 );
nor U118276 ( n59767, n6683, n59769 );
nor U118277 ( n59769, n59770, n6695 );
nor U118278 ( n47605, n7607, n47607 );
nor U118279 ( n47607, n47608, n7622 );
not U118280 ( n4968, n14204 );
not U118281 ( n3235, n33796 );
nor U118282 ( n33870, n3220, n33872 );
nor U118283 ( n33872, n33873, n3235 );
nor U118284 ( n14297, n4953, n14299 );
nor U118285 ( n14299, n14300, n4968 );
nand U118286 ( n60065, P2_P2_STATE2_REG_3_, n60062 );
nand U118287 ( n26925, P1_P2_STATE2_REG_3_, n26922 );
nand U118288 ( n34170, P1_P3_STATE2_REG_3_, n34167 );
nand U118289 ( n68924, P2_P3_STATE2_REG_3_, n68921 );
nand U118290 ( n12827, n12732, n72970 );
xnor U118291 ( n67176, n68530, n68457 );
xnor U118292 ( n46212, n47509, n47436 );
xnor U118293 ( n25278, n26529, n26456 );
xnor U118294 ( n58414, n59671, n59595 );
xnor U118295 ( n32520, n33774, n33701 );
xnor U118296 ( n12585, n14177, n14085 );
nor U118297 ( n68630, n68629, n68631 );
nor U118298 ( n68631, n5819, n68552 );
nor U118299 ( n26629, n26628, n26630 );
nor U118300 ( n26630, n4050, n26551 );
nor U118301 ( n59771, n59770, n59772 );
nor U118302 ( n59772, n6683, n59693 );
nor U118303 ( n47609, n47608, n47610 );
nor U118304 ( n47610, n7607, n47531 );
nor U118305 ( n33874, n33873, n33875 );
nor U118306 ( n33875, n3220, n33796 );
nor U118307 ( n14302, n14300, n14303 );
nor U118308 ( n14303, n4953, n14204 );
nor U118309 ( n34284, n34288, n34289 );
nor U118310 ( n69036, n69040, n69041 );
nor U118311 ( n34297, n34288, n34300 );
nor U118312 ( n34341, n34288, n34344 );
nor U118313 ( n34352, n34288, n34355 );
nor U118314 ( n34375, n34288, n34379 );
nor U118315 ( n34319, n34288, n34322 );
nor U118316 ( n34330, n34288, n34333 );
nor U118317 ( n34308, n34288, n34311 );
nor U118318 ( n69049, n69040, n69052 );
nor U118319 ( n69060, n69040, n69063 );
nor U118320 ( n69071, n69040, n69074 );
nor U118321 ( n69104, n69040, n69107 );
nor U118322 ( n69127, n69040, n69131 );
nor U118323 ( n69093, n69040, n69096 );
nor U118324 ( n69082, n69040, n69085 );
nor U118325 ( n21707, n74727, n76562 );
nor U118326 ( n21695, n74656, n76561 );
nor U118327 ( n21699, n72965, n76561 );
nor U118328 ( n21691, n72963, n76562 );
nor U118329 ( n21703, n74673, n76562 );
nor U118330 ( n21711, n74729, n76561 );
nor U118331 ( n27552, n4287, n26969 );
nor U118332 ( n34797, n3449, n34214 );
nor U118333 ( n69541, n6064, n68968 );
nor U118334 ( n60704, n6919, n60109 );
nor U118335 ( n69311, n69052, n69304 );
nor U118336 ( n69231, n69052, n69224 );
nor U118337 ( n69149, n69052, n69142 );
nor U118338 ( n70262, n69063, n70247 );
nor U118339 ( n69319, n69063, n69304 );
nor U118340 ( n69239, n69063, n69224 );
nor U118341 ( n69157, n69063, n69142 );
nor U118342 ( n70270, n69074, n70247 );
nor U118343 ( n69327, n69074, n69304 );
nor U118344 ( n69247, n69074, n69224 );
nor U118345 ( n69165, n69074, n69142 );
nor U118346 ( n70295, n69107, n70247 );
nor U118347 ( n69351, n69107, n69304 );
nor U118348 ( n69271, n69107, n69224 );
nor U118349 ( n69189, n69107, n69142 );
nor U118350 ( n69359, n69131, n69304 );
nor U118351 ( n69279, n69131, n69224 );
nor U118352 ( n69197, n69131, n69142 );
nor U118353 ( n70287, n69096, n70247 );
nor U118354 ( n69343, n69096, n69304 );
nor U118355 ( n69263, n69096, n69224 );
nor U118356 ( n69181, n69096, n69142 );
nor U118357 ( n70279, n69085, n70247 );
nor U118358 ( n69335, n69085, n69304 );
nor U118359 ( n69255, n69085, n69224 );
nor U118360 ( n69173, n69085, n69142 );
nor U118361 ( n69298, n69041, n69304 );
nor U118362 ( n69218, n69041, n69224 );
nor U118363 ( n69136, n69041, n69142 );
nor U118364 ( n70238, n69041, n70247 );
nor U118365 ( n70303, n69131, n70247 );
nor U118366 ( n70254, n69052, n70247 );
nor U118367 ( n34563, n34300, n34556 );
nor U118368 ( n34481, n34300, n34474 );
nor U118369 ( n34399, n34300, n34390 );
nor U118370 ( n35559, n34344, n35519 );
nor U118371 ( n34597, n34344, n34556 );
nor U118372 ( n34515, n34344, n34474 );
nor U118373 ( n34431, n34344, n34390 );
nor U118374 ( n35567, n34355, n35519 );
nor U118375 ( n34605, n34355, n34556 );
nor U118376 ( n34523, n34355, n34474 );
nor U118377 ( n34439, n34355, n34390 );
nor U118378 ( n34613, n34379, n34556 );
nor U118379 ( n34531, n34379, n34474 );
nor U118380 ( n34447, n34379, n34390 );
nor U118381 ( n35542, n34322, n35519 );
nor U118382 ( n34579, n34322, n34556 );
nor U118383 ( n34499, n34322, n34474 );
nor U118384 ( n34415, n34322, n34390 );
nor U118385 ( n35551, n34333, n35519 );
nor U118386 ( n34587, n34333, n34556 );
nor U118387 ( n34507, n34333, n34474 );
nor U118388 ( n34423, n34333, n34390 );
nor U118389 ( n34550, n34289, n34556 );
nor U118390 ( n34468, n34289, n34474 );
nor U118391 ( n34384, n34289, n34390 );
nor U118392 ( n35534, n34311, n35519 );
nor U118393 ( n34571, n34311, n34556 );
nor U118394 ( n34489, n34311, n34474 );
nor U118395 ( n34407, n34311, n34390 );
nor U118396 ( n35510, n34289, n35519 );
nor U118397 ( n35575, n34379, n35519 );
nor U118398 ( n35526, n34300, n35519 );
nor U118399 ( n60078, n60065, n60079 );
nor U118400 ( n26938, n26925, n26939 );
nor U118401 ( n34183, n34170, n34184 );
nor U118402 ( n68937, n68924, n68938 );
nor U118403 ( n69637, n69052, n69629 );
nor U118404 ( n69645, n69063, n69629 );
nor U118405 ( n69653, n69074, n69629 );
nor U118406 ( n69677, n69107, n69629 );
nor U118407 ( n69693, n69131, n69629 );
nor U118408 ( n69669, n69096, n69629 );
nor U118409 ( n69661, n69085, n69629 );
nor U118410 ( n69628, n69041, n69629 );
nor U118411 ( n34895, n34300, n34887 );
nor U118412 ( n34929, n34344, n34887 );
nor U118413 ( n34937, n34355, n34887 );
nor U118414 ( n34953, n34379, n34887 );
nor U118415 ( n34913, n34322, n34887 );
nor U118416 ( n34921, n34333, n34887 );
nor U118417 ( n34886, n34289, n34887 );
nor U118418 ( n34903, n34311, n34887 );
nor U118419 ( n69385, n69041, n69388 );
nor U118420 ( n34639, n34289, n34642 );
nor U118421 ( n69395, n69052, n69388 );
nor U118422 ( n69403, n69063, n69388 );
nor U118423 ( n69411, n69074, n69388 );
nor U118424 ( n69435, n69107, n69388 );
nor U118425 ( n69454, n69131, n69388 );
nor U118426 ( n69427, n69096, n69388 );
nor U118427 ( n69419, n69085, n69388 );
nor U118428 ( n34649, n34300, n34642 );
nor U118429 ( n34681, n34344, n34642 );
nor U118430 ( n34689, n34355, n34642 );
nor U118431 ( n34710, n34379, n34642 );
nor U118432 ( n34665, n34322, n34642 );
nor U118433 ( n34673, n34333, n34642 );
nor U118434 ( n34657, n34311, n34642 );
nor U118435 ( n60070, n60071, n60072 );
nor U118436 ( n60071, n60073, n60074 );
nor U118437 ( n60073, n60075, n74424 );
nor U118438 ( n26930, n26931, n26932 );
nor U118439 ( n26931, n26933, n26934 );
nor U118440 ( n26933, n26935, n74423 );
nor U118441 ( n34175, n34176, n34177 );
nor U118442 ( n34176, n34178, n34179 );
nor U118443 ( n34178, n34180, n74426 );
nor U118444 ( n68929, n68930, n68931 );
nor U118445 ( n68930, n68932, n68933 );
nor U118446 ( n68932, n68934, n74425 );
nand U118447 ( n34881, n34884, n88 );
not U118448 ( n88, n34287 );
nand U118449 ( n69623, n69626, n353 );
not U118450 ( n353, n69039 );
nand U118451 ( n14402, n14304, n4954 );
xor U118452 ( n18715, n20929, n15273 );
nand U118453 ( n60076, n6925, n60062 );
nand U118454 ( n26936, n4293, n26922 );
nand U118455 ( n34181, n3455, n34167 );
nand U118456 ( n68935, n6070, n68921 );
and U118457 ( n27310, n27378, n4268 );
and U118458 ( n27378, n26955, n4287 );
and U118459 ( n34555, n34623, n3430 );
and U118460 ( n34623, n34200, n3449 );
and U118461 ( n60453, n60526, n6900 );
and U118462 ( n60526, n60095, n6919 );
and U118463 ( n69303, n69369, n6045 );
and U118464 ( n69369, n68954, n6064 );
and U118465 ( n63216, n75864, n63218 );
or U118466 ( n75864, n63219, n63220 );
and U118467 ( n29453, n75865, n29455 );
or U118468 ( n75865, n29456, n29457 );
and U118469 ( n22134, n75866, n22136 );
or U118470 ( n75866, n22137, n22138 );
and U118471 ( n55244, n75867, n55246 );
or U118472 ( n75867, n55247, n55248 );
nor U118473 ( n8668, n5273, n8637 );
nor U118474 ( n42728, n7928, n42703 );
nor U118475 ( n31658, n75278, n31646 );
nor U118476 ( n31662, n74731, n31646 );
nor U118477 ( n31666, n75280, n31646 );
nor U118478 ( n31670, n74676, n31646 );
nor U118479 ( n31678, n75252, n31646 );
nor U118480 ( n31682, n75281, n31646 );
nor U118481 ( n31698, n74540, n31646 );
nor U118482 ( n31710, n75286, n31646 );
nor U118483 ( n31706, n73135, n31646 );
nor U118484 ( n31714, n72957, n31646 );
nor U118485 ( n31702, n75279, n31646 );
nor U118486 ( n31690, n75282, n31646 );
nor U118487 ( n31686, n74582, n31646 );
nor U118488 ( n31654, n74778, n31646 );
nor U118489 ( n31718, n74488, n31646 );
nor U118490 ( n31674, n74629, n31646 );
nor U118491 ( n8703, n5273, n8704 );
nor U118492 ( n8704, n8705, n8707 );
nor U118493 ( n8705, n8708, n8709 );
nor U118494 ( n42760, n7928, n42761 );
nor U118495 ( n42761, n42762, n42763 );
nor U118496 ( n42762, n42764, n42765 );
nand U118497 ( n28408, n74423, n27459 );
nand U118498 ( n61717, n74424, n60608 );
nand U118499 ( n70317, n74425, n69448 );
nand U118500 ( n35589, n74426, n34704 );
nor U118501 ( n31752, n75311, n31756 );
nor U118502 ( n31736, n75296, n31756 );
nor U118503 ( n31732, n75297, n31756 );
nor U118504 ( n31740, n75298, n31756 );
nor U118505 ( n31727, n75288, n31756 );
nand U118506 ( n27227, n27290, n76517 );
nor U118507 ( n27290, n27291, n27292 );
and U118508 ( n27292, n27232, P1_P2_STATE2_REG_3_ );
nor U118509 ( n27291, n27293, n27294 );
nand U118510 ( n60372, n60433, n76259 );
nor U118511 ( n60433, n60434, n60435 );
and U118512 ( n60435, n60377, P2_P2_STATE2_REG_3_ );
nor U118513 ( n60434, n60436, n60437 );
nand U118514 ( n34472, n34535, n76461 );
nor U118515 ( n34535, n34536, n34537 );
and U118516 ( n34537, n34477, P1_P3_STATE2_REG_3_ );
nor U118517 ( n34536, n34538, n34539 );
nand U118518 ( n69222, n69283, n76193 );
nor U118519 ( n69283, n69284, n69285 );
and U118520 ( n69285, n69227, P2_P3_STATE2_REG_3_ );
nor U118521 ( n69284, n69286, n69287 );
nand U118522 ( n11244, n11245, n10120 );
nor U118523 ( n42671, n42675, n42676 );
nand U118524 ( n42676, n42677, n42424 );
nand U118525 ( n34280, n34362, n76461 );
nor U118526 ( n34362, n34363, n34364 );
and U118527 ( n34364, n34282, P1_P3_STATE2_REG_3_ );
nor U118528 ( n34363, n34365, n34366 );
nand U118529 ( n69032, n69114, n76193 );
nor U118530 ( n69114, n69115, n69116 );
and U118531 ( n69116, n69034, P2_P3_STATE2_REG_3_ );
nor U118532 ( n69115, n69117, n69118 );
nand U118533 ( n27035, n27117, n76517 );
nor U118534 ( n27117, n27118, n27119 );
and U118535 ( n27119, n27038, P1_P2_STATE2_REG_3_ );
nor U118536 ( n27118, n27120, n27121 );
nand U118537 ( n60176, n60261, n76259 );
nor U118538 ( n60261, n60262, n60263 );
and U118539 ( n60263, n60179, P2_P2_STATE2_REG_3_ );
nor U118540 ( n60262, n60264, n60265 );
nand U118541 ( n15609, n15693, n76591 );
nor U118542 ( n15693, n15694, n15695 );
nor U118543 ( n15695, n5194, n4813 );
nor U118544 ( n15694, n15697, n15692 );
nor U118545 ( n35432, n34287, n35438 );
nor U118546 ( n35353, n34287, n35359 );
nor U118547 ( n35195, n34287, n35201 );
nor U118548 ( n35117, n34287, n35123 );
nor U118549 ( n35037, n34287, n35043 );
nor U118550 ( n34800, n34287, n34806 );
nor U118551 ( n34715, n34287, n34721 );
nor U118552 ( n69853, n69039, n69859 );
nor U118553 ( n69544, n69039, n69550 );
nor U118554 ( n69459, n69039, n69465 );
nor U118555 ( n70162, n69039, n70168 );
nor U118556 ( n70085, n69039, n70091 );
nor U118557 ( n69931, n69039, n69937 );
nor U118558 ( n69775, n69039, n69781 );
nor U118559 ( n60112, n73137, n60062 );
nor U118560 ( n26972, n73136, n26922 );
nor U118561 ( n34217, n73138, n34167 );
nor U118562 ( n68971, n73139, n68921 );
nor U118563 ( n31809, n75316, n31756 );
nor U118564 ( n31805, n75317, n31756 );
nor U118565 ( n31801, n75318, n31756 );
nor U118566 ( n31793, n75319, n31756 );
nor U118567 ( n31785, n75320, n31756 );
nor U118568 ( n31773, n75312, n31756 );
nor U118569 ( n31769, n75313, n31756 );
nor U118570 ( n31777, n75314, n31756 );
nor U118571 ( n31781, n75315, n31756 );
nor U118572 ( n31816, n75363, n31756 );
nor U118573 ( n31797, n75321, n31756 );
nor U118574 ( n48523, n74442, n7855 );
nand U118575 ( n46926, n47063, n47064 );
nor U118576 ( n47063, n74734, n47011 );
nand U118577 ( n47497, n47583, n7879 );
nor U118578 ( n47583, n74400, n73071 );
nand U118579 ( n46711, n46816, n46817 );
nor U118580 ( n46816, n74524, n46818 );
nor U118581 ( n46591, n46695, n46711 );
nor U118582 ( n47311, n47497, n75934 );
nand U118583 ( n46450, n46590, n46591 );
nor U118584 ( n46590, n74881, n46592 );
nor U118585 ( n46817, n46926, n46927 );
nand U118586 ( n46432, n46448, n46449 );
nor U118587 ( n46449, n74930, n73220 );
nor U118588 ( n46448, n74919, n46450 );
and U118589 ( n47064, n47169, n47170 );
nor U118590 ( n47170, n73078, n74659 );
nor U118591 ( n47169, n73178, n47171 );
nor U118592 ( n27301, n74423, n4294 );
nor U118593 ( n34546, n74426, n3457 );
nor U118594 ( n60444, n74424, n6927 );
nor U118595 ( n69294, n74425, n6072 );
nor U118596 ( n28413, n27301, n27219 );
nor U118597 ( n35594, n34546, n34464 );
nor U118598 ( n61722, n60444, n60364 );
nor U118599 ( n70322, n69294, n69214 );
not U118600 ( n4294, n27459 );
not U118601 ( n3457, n34704 );
not U118602 ( n6927, n60608 );
not U118603 ( n6072, n69448 );
and U118604 ( n34389, n34457, n34179 );
nor U118605 ( n34457, n34214, n34458 );
and U118606 ( n69141, n69207, n68933 );
nor U118607 ( n69207, n68968, n69208 );
and U118608 ( n27146, n27212, n26934 );
nor U118609 ( n27212, n26969, n27213 );
and U118610 ( n60288, n60357, n60074 );
nor U118611 ( n60357, n60109, n60358 );
not U118612 ( n2903, n38163 );
nand U118613 ( n34892, n34884, n90 );
not U118614 ( n90, n34299 );
nand U118615 ( n34926, n34884, n98 );
not U118616 ( n98, n34343 );
nand U118617 ( n34934, n34884, n100 );
not U118618 ( n100, n34354 );
nand U118619 ( n34942, n34884, n102 );
not U118620 ( n102, n34377 );
nand U118621 ( n34910, n34884, n94 );
not U118622 ( n94, n34321 );
nand U118623 ( n34918, n34884, n96 );
not U118624 ( n96, n34332 );
nand U118625 ( n34900, n34884, n92 );
not U118626 ( n92, n34310 );
nand U118627 ( n69634, n69626, n355 );
not U118628 ( n355, n69051 );
nand U118629 ( n69642, n69626, n358 );
not U118630 ( n358, n69062 );
nand U118631 ( n69650, n69626, n360 );
not U118632 ( n360, n69073 );
nand U118633 ( n69674, n69626, n368 );
not U118634 ( n368, n69106 );
nand U118635 ( n69682, n69626, n370 );
not U118636 ( n370, n69129 );
nand U118637 ( n69666, n69626, n365 );
not U118638 ( n365, n69095 );
nand U118639 ( n69658, n69626, n363 );
not U118640 ( n363, n69084 );
nor U118641 ( n14692, n15167, n15058 );
nand U118642 ( n14733, n14717, n15062 );
xnor U118643 ( n14177, n75941, n14144 );
nor U118644 ( n47939, n7413, n47942 );
nor U118645 ( n47942, n47943, n47944 );
nor U118646 ( n47944, n7415, n7838 );
nor U118647 ( n47943, n47946, n47918 );
nand U118648 ( n15511, n47937, n47938 );
nor U118649 ( n47937, n47949, n47950 );
nor U118650 ( n47938, n47939, n47940 );
nor U118651 ( n47949, n7457, n47951 );
xnor U118652 ( n68530, n75937, n68504 );
xnor U118653 ( n47509, n75934, n47483 );
xnor U118654 ( n26529, n75938, n26503 );
xnor U118655 ( n59671, n75939, n59642 );
xnor U118656 ( n33774, n75940, n33748 );
nand U118657 ( n42426, n42427, n42428 );
nand U118658 ( n42427, n42430, n42431 );
nand U118659 ( n42428, n42429, n900 );
nand U118660 ( n42430, n42432, n42433 );
xor U118661 ( n68627, n74408, n68546 );
xor U118662 ( n26626, n74409, n26545 );
xor U118663 ( n59768, n74410, n59687 );
xor U118664 ( n47606, n74400, n47525 );
xor U118665 ( n33871, n74412, n33790 );
xor U118666 ( n14298, n74429, n14197 );
nor U118667 ( n63338, n6140, n63339 );
nor U118668 ( n63339, n63340, n6168 );
not U118669 ( n6168, n63341 );
nor U118670 ( n63340, n63342, n63343 );
nor U118671 ( n29509, n3525, n29510 );
nor U118672 ( n29510, n29511, n3553 );
not U118673 ( n3553, n29512 );
nor U118674 ( n29511, n29513, n29514 );
nor U118675 ( n22190, n4363, n22191 );
nor U118676 ( n22191, n22192, n4390 );
not U118677 ( n4390, n22193 );
nor U118678 ( n22192, n22194, n22195 );
nor U118679 ( n55304, n6995, n55305 );
nor U118680 ( n55305, n55306, n7023 );
not U118681 ( n7023, n55307 );
nor U118682 ( n55306, n55308, n55309 );
nand U118683 ( n68696, n68632, n5820 );
nand U118684 ( n47675, n47611, n7608 );
nand U118685 ( n26695, n26631, n4052 );
nand U118686 ( n59837, n59773, n6684 );
nand U118687 ( n33940, n33876, n3222 );
not U118688 ( n3503, n32961 );
nand U118689 ( n41977, n842, n41908 );
not U118690 ( n2978, n31722 );
nand U118691 ( n67200, n68708, n68709 );
nand U118692 ( n68708, n5835, n68712 );
nand U118693 ( n68709, n68710, n68671 );
nand U118694 ( n68710, n5818, n68535 );
nand U118695 ( n46248, n47687, n47688 );
nand U118696 ( n47687, n7623, n47691 );
nand U118697 ( n47688, n47689, n47650 );
nand U118698 ( n47689, n7605, n47514 );
nand U118699 ( n25302, n26707, n26708 );
nand U118700 ( n26707, n4064, n26711 );
nand U118701 ( n26708, n26709, n26670 );
nand U118702 ( n26709, n4049, n26534 );
nand U118703 ( n58441, n59849, n59850 );
nand U118704 ( n59849, n6697, n59853 );
nand U118705 ( n59850, n59851, n59812 );
nand U118706 ( n59851, n6682, n59676 );
nand U118707 ( n32544, n33952, n33953 );
nand U118708 ( n33952, n3236, n33956 );
nand U118709 ( n33953, n33954, n33915 );
nand U118710 ( n33954, n3219, n33779 );
nand U118711 ( n42420, n42421, n902 );
xor U118712 ( n42421, n74281, n893 );
nor U118713 ( n35445, n34299, n35438 );
nor U118714 ( n35366, n34299, n35359 );
nor U118715 ( n35210, n34299, n35201 );
nor U118716 ( n35130, n34299, n35123 );
nor U118717 ( n35050, n34299, n35043 );
nor U118718 ( n34815, n34299, n34806 );
nor U118719 ( n34729, n34299, n34721 );
nor U118720 ( n35400, n34343, n35359 );
nor U118721 ( n35242, n34343, n35201 );
nor U118722 ( n35162, n34343, n35123 );
nor U118723 ( n35082, n34343, n35043 );
nor U118724 ( n34847, n34343, n34806 );
nor U118725 ( n34765, n34343, n34721 );
nor U118726 ( n35477, n34343, n35438 );
nor U118727 ( n35408, n34354, n35359 );
nor U118728 ( n35250, n34354, n35201 );
nor U118729 ( n35170, n34354, n35123 );
nor U118730 ( n35090, n34354, n35043 );
nor U118731 ( n34855, n34354, n34806 );
nor U118732 ( n34774, n34354, n34721 );
nor U118733 ( n35485, n34354, n35438 );
nor U118734 ( n35495, n34377, n35438 );
nor U118735 ( n35416, n34377, n35359 );
nor U118736 ( n35258, n34377, n35201 );
nor U118737 ( n35178, n34377, n35123 );
nor U118738 ( n35100, n34377, n35043 );
nor U118739 ( n34863, n34377, n34806 );
nor U118740 ( n34783, n34377, n34721 );
nor U118741 ( n35461, n34321, n35438 );
nor U118742 ( n35382, n34321, n35359 );
nor U118743 ( n35226, n34321, n35201 );
nor U118744 ( n35146, n34321, n35123 );
nor U118745 ( n35066, n34321, n35043 );
nor U118746 ( n34831, n34321, n34806 );
nor U118747 ( n34747, n34321, n34721 );
nor U118748 ( n35469, n34332, n35438 );
nor U118749 ( n35390, n34332, n35359 );
nor U118750 ( n35234, n34332, n35201 );
nor U118751 ( n35154, n34332, n35123 );
nor U118752 ( n35074, n34332, n35043 );
nor U118753 ( n34839, n34332, n34806 );
nor U118754 ( n34756, n34332, n34721 );
nor U118755 ( n35374, n34310, n35359 );
nor U118756 ( n35218, n34310, n35201 );
nor U118757 ( n35138, n34310, n35123 );
nor U118758 ( n35058, n34310, n35043 );
nor U118759 ( n34823, n34310, n34806 );
nor U118760 ( n34738, n34310, n34721 );
nor U118761 ( n70175, n69051, n70168 );
nor U118762 ( n70098, n69051, n70091 );
nor U118763 ( n69944, n69051, n69937 );
nor U118764 ( n69866, n69051, n69859 );
nor U118765 ( n69788, n69051, n69781 );
nor U118766 ( n69557, n69051, n69550 );
nor U118767 ( n69473, n69051, n69465 );
nor U118768 ( n70106, n69062, n70091 );
nor U118769 ( n69952, n69062, n69937 );
nor U118770 ( n69874, n69062, n69859 );
nor U118771 ( n69796, n69062, n69781 );
nor U118772 ( n69565, n69062, n69550 );
nor U118773 ( n69482, n69062, n69465 );
nor U118774 ( n70191, n69073, n70168 );
nor U118775 ( n70114, n69073, n70091 );
nor U118776 ( n69960, n69073, n69937 );
nor U118777 ( n69882, n69073, n69859 );
nor U118778 ( n69804, n69073, n69781 );
nor U118779 ( n69573, n69073, n69550 );
nor U118780 ( n69491, n69073, n69465 );
nor U118781 ( n70138, n69106, n70091 );
nor U118782 ( n69984, n69106, n69937 );
nor U118783 ( n69906, n69106, n69859 );
nor U118784 ( n69828, n69106, n69781 );
nor U118785 ( n69597, n69106, n69550 );
nor U118786 ( n69518, n69106, n69465 );
nor U118787 ( n70215, n69106, n70168 );
nor U118788 ( n70223, n69129, n70168 );
nor U118789 ( n70146, n69129, n70091 );
nor U118790 ( n69992, n69129, n69937 );
nor U118791 ( n69914, n69129, n69859 );
nor U118792 ( n69836, n69129, n69781 );
nor U118793 ( n69605, n69129, n69550 );
nor U118794 ( n69527, n69129, n69465 );
nor U118795 ( n70130, n69095, n70091 );
nor U118796 ( n69976, n69095, n69937 );
nor U118797 ( n69898, n69095, n69859 );
nor U118798 ( n69820, n69095, n69781 );
nor U118799 ( n69589, n69095, n69550 );
nor U118800 ( n69509, n69095, n69465 );
nor U118801 ( n70207, n69095, n70168 );
nor U118802 ( n70199, n69084, n70168 );
nor U118803 ( n70122, n69084, n70091 );
nor U118804 ( n69968, n69084, n69937 );
nor U118805 ( n69890, n69084, n69859 );
nor U118806 ( n69812, n69084, n69781 );
nor U118807 ( n69581, n69084, n69550 );
nor U118808 ( n69500, n69084, n69465 );
nor U118809 ( n70183, n69062, n70168 );
nor U118810 ( n35453, n34310, n35438 );
nor U118811 ( n49554, n49461, n73640 );
nor U118812 ( n49599, n49461, n73808 );
nor U118813 ( n49524, n49461, n73611 );
nor U118814 ( n49460, n49461, n73556 );
nor U118815 ( n49495, n49461, n73552 );
nor U118816 ( n49627, n49461, n73882 );
nor U118817 ( n49657, n49461, n73968 );
xor U118818 ( n28412, n28408, n27384 );
xor U118819 ( n70321, n70317, n69375 );
xor U118820 ( n35593, n35589, n34629 );
xor U118821 ( n61721, n61717, n60532 );
nand U118822 ( n60084, n60062, n60085 );
nand U118823 ( n60085, P2_P2_STATE2_REG_3_, n60086 );
nand U118824 ( n26944, n26922, n26945 );
nand U118825 ( n26945, P1_P2_STATE2_REG_3_, n26946 );
nand U118826 ( n34189, n34167, n34190 );
nand U118827 ( n34190, P1_P3_STATE2_REG_3_, n34191 );
nand U118828 ( n68943, n68921, n68944 );
nand U118829 ( n68944, P2_P3_STATE2_REG_3_, n68945 );
nand U118830 ( n68621, n68538, n74408 );
nand U118831 ( n26620, n26537, n74409 );
nand U118832 ( n59762, n59679, n74410 );
nand U118833 ( n47600, n47517, n74400 );
nand U118834 ( n33865, n33782, n74412 );
nand U118835 ( n14290, n14187, n74429 );
nand U118836 ( n31624, n31619, n74591 );
nand U118837 ( n27638, n27699, n76517 );
nor U118838 ( n27699, n27700, n27701 );
nor U118839 ( n27701, n4284, n76916 );
nor U118840 ( n27700, n27702, n27703 );
nand U118841 ( n34883, n34944, n76461 );
nor U118842 ( n34944, n34945, n34946 );
nor U118843 ( n34946, n3447, n76918 );
nor U118844 ( n34945, n34947, n34948 );
nand U118845 ( n69625, n69684, n76193 );
nor U118846 ( n69684, n69685, n69686 );
nor U118847 ( n69686, n6062, n76914 );
nor U118848 ( n69685, n69687, n69688 );
nand U118849 ( n60791, n60850, n76259 );
nor U118850 ( n60850, n60851, n60852 );
nor U118851 ( n60852, n6917, n76912 );
nor U118852 ( n60851, n60853, n60854 );
not U118853 ( n3822, n24460 );
nand U118854 ( n43413, n43421, n8089 );
nor U118855 ( n43421, n75071, n73310 );
nand U118856 ( n30144, n30152, n3674 );
nor U118857 ( n30152, n75072, n73311 );
nand U118858 ( n64157, n64165, n6308 );
nor U118859 ( n64165, n75073, n73312 );
nand U118860 ( n22819, n22827, n4568 );
nor U118861 ( n22827, n75074, n73313 );
nand U118862 ( n55933, n55941, n7200 );
nor U118863 ( n55941, n75076, n73314 );
not U118864 ( n3688, n30381 );
not U118865 ( n4582, n23052 );
not U118866 ( n6322, n64544 );
not U118867 ( n7214, n56175 );
not U118868 ( n8103, n43702 );
nand U118869 ( n30364, n30366, n3688 );
nor U118870 ( n30366, n74568, n73144 );
nand U118871 ( n23035, n23037, n4582 );
nor U118872 ( n23037, n74572, n73145 );
nand U118873 ( n64483, n64485, n6322 );
nor U118874 ( n64485, n74570, n73146 );
nand U118875 ( n56154, n56156, n7214 );
nor U118876 ( n56156, n74573, n73147 );
nand U118877 ( n43685, n43687, n8103 );
nor U118878 ( n43687, n74571, n73142 );
nand U118879 ( n43471, n43473, n8090 );
nor U118880 ( n43473, n75021, n73298 );
nand U118881 ( n43490, n43492, n8092 );
nor U118882 ( n43492, n74978, n73282 );
nand U118883 ( n43509, n43511, n8093 );
nor U118884 ( n43511, n74932, n73269 );
nand U118885 ( n43528, n43530, n8094 );
nor U118886 ( n43530, n74892, n73255 );
nand U118887 ( n43547, n43549, n8095 );
nor U118888 ( n43549, n74831, n73241 );
nand U118889 ( n43579, n43581, n8097 );
nor U118890 ( n43581, n74795, n73226 );
nand U118891 ( n30169, n30171, n3675 );
nor U118892 ( n30171, n75022, n73299 );
nand U118893 ( n30188, n30190, n3677 );
nor U118894 ( n30190, n74979, n73283 );
nand U118895 ( n30211, n30213, n3678 );
nor U118896 ( n30213, n74933, n73270 );
nand U118897 ( n30230, n30232, n3679 );
nor U118898 ( n30232, n74893, n73256 );
nand U118899 ( n30249, n30251, n3680 );
nor U118900 ( n30251, n74832, n73242 );
nand U118901 ( n30268, n30270, n3682 );
nor U118902 ( n30270, n74792, n73227 );
nand U118903 ( n30287, n30289, n3683 );
nor U118904 ( n30289, n74762, n73208 );
nand U118905 ( n30310, n30312, n3684 );
nor U118906 ( n30312, n74719, n73200 );
nand U118907 ( n64182, n64184, n6309 );
nor U118908 ( n64184, n75023, n73300 );
nand U118909 ( n64254, n64256, n6310 );
nor U118910 ( n64256, n74980, n73284 );
nand U118911 ( n64273, n64275, n6312 );
nor U118912 ( n64275, n74934, n73271 );
nand U118913 ( n64292, n64294, n6313 );
nor U118914 ( n64294, n74894, n73257 );
nand U118915 ( n64311, n64313, n6314 );
nor U118916 ( n64313, n74833, n73243 );
nand U118917 ( n64330, n64332, n6315 );
nor U118918 ( n64332, n74793, n73228 );
nand U118919 ( n64410, n64412, n6317 );
nor U118920 ( n64412, n74763, n73209 );
nand U118921 ( n64429, n64431, n6318 );
nor U118922 ( n64431, n74720, n73201 );
nand U118923 ( n30329, n30331, n3685 );
nor U118924 ( n30331, n74664, n73170 );
nand U118925 ( n30347, n30349, n3687 );
nor U118926 ( n30349, n74601, n73152 );
nand U118927 ( n22844, n22846, n4569 );
nor U118928 ( n22846, n75024, n73301 );
nand U118929 ( n22863, n22865, n4570 );
nor U118930 ( n22865, n74982, n73285 );
nand U118931 ( n22884, n22886, n4572 );
nor U118932 ( n22886, n74936, n73272 );
nand U118933 ( n22903, n22905, n4573 );
nor U118934 ( n22905, n74896, n73258 );
nand U118935 ( n22922, n22924, n4574 );
nor U118936 ( n22924, n74835, n73244 );
nand U118937 ( n22941, n22943, n4575 );
nor U118938 ( n22943, n74796, n73229 );
nand U118939 ( n22960, n22962, n4577 );
nor U118940 ( n22962, n74766, n73210 );
nand U118941 ( n22981, n22983, n4578 );
nor U118942 ( n22983, n74723, n73202 );
nand U118943 ( n23000, n23002, n4579 );
nor U118944 ( n23002, n74668, n73171 );
nand U118945 ( n23018, n23020, n4580 );
nor U118946 ( n23020, n74605, n73153 );
nand U118947 ( n64448, n64450, n6319 );
nor U118948 ( n64450, n74666, n73172 );
nand U118949 ( n64466, n64468, n6320 );
nor U118950 ( n64468, n74603, n73154 );
nand U118951 ( n55961, n55963, n7202 );
nor U118952 ( n55963, n75026, n73302 );
nand U118953 ( n55980, n55982, n7203 );
nor U118954 ( n55982, n74983, n73286 );
nand U118955 ( n55999, n56001, n7204 );
nor U118956 ( n56001, n74937, n73273 );
nand U118957 ( n56018, n56020, n7205 );
nor U118958 ( n56020, n74897, n73259 );
nand U118959 ( n56037, n56039, n7207 );
nor U118960 ( n56039, n74836, n73245 );
nand U118961 ( n56059, n56061, n7208 );
nor U118962 ( n56061, n74797, n73230 );
nand U118963 ( n56078, n56080, n7209 );
nor U118964 ( n56080, n74767, n73211 );
nand U118965 ( n56097, n56099, n7210 );
nor U118966 ( n56099, n74724, n73203 );
nand U118967 ( n56116, n56118, n7212 );
nor U118968 ( n56118, n74669, n73173 );
nand U118969 ( n56134, n56136, n7213 );
nor U118970 ( n56136, n74606, n73155 );
nand U118971 ( n43598, n43600, n8098 );
nor U118972 ( n43600, n74765, n73212 );
nand U118973 ( n43617, n43619, n8099 );
nor U118974 ( n43619, n74722, n73204 );
nand U118975 ( n43636, n43638, n8100 );
nor U118976 ( n43638, n74667, n73174 );
nand U118977 ( n43654, n43656, n8102 );
nor U118978 ( n43656, n74604, n73156 );
nand U118979 ( n47012, n47100, n47101 );
nor U118980 ( n47100, n72948, n74734 );
nand U118981 ( n47132, n47221, n47222 );
nor U118982 ( n47221, n74659, n73178 );
nand U118983 ( n47270, n47408, n47409 );
nor U118984 ( n47408, n75934, n74443 );
nor U118985 ( n47409, n7873, n74400 );
nor U118986 ( n46980, n47012, n74427 );
nand U118987 ( n46491, n46498, n7870 );
nor U118988 ( n46498, n46499, n74919 );
nor U118989 ( n47222, n47270, n73065 );
nor U118990 ( n47101, n47132, n73078 );
nand U118991 ( n46627, n46630, n7872 );
nor U118992 ( n46630, n73148, n46592 );
nand U118993 ( n46725, n46740, n46741 );
nor U118994 ( n46740, n74524, n46734 );
nand U118995 ( n9483, n9493, n5434 );
nor U118996 ( n9493, n75075, n73315 );
not U118997 ( n5448, n9775 );
nand U118998 ( n9750, n9753, n5448 );
nor U118999 ( n9753, n74569, n73143 );
nand U119000 ( n9514, n9517, n5435 );
nor U119001 ( n9517, n75025, n73303 );
nand U119002 ( n9538, n9540, n5437 );
nor U119003 ( n9540, n74981, n73287 );
nand U119004 ( n9562, n9564, n5438 );
nor U119005 ( n9564, n74935, n73274 );
nand U119006 ( n9585, n9587, n5439 );
nor U119007 ( n9587, n74895, n73260 );
nand U119008 ( n9608, n9610, n5440 );
nor U119009 ( n9610, n74834, n73246 );
nand U119010 ( n9659, n9662, n5443 );
nor U119011 ( n9662, n74764, n73213 );
nand U119012 ( n9683, n9685, n5444 );
nor U119013 ( n9685, n74721, n73205 );
nand U119014 ( n9707, n9709, n5445 );
nor U119015 ( n9709, n74665, n73175 );
nand U119016 ( n9729, n9732, n5447 );
nor U119017 ( n9732, n74602, n73157 );
nand U119018 ( n9632, n9634, n5442 );
nor U119019 ( n9634, n74794, n73231 );
nand U119020 ( n13579, n13690, n13692 );
nor U119021 ( n13690, n73116, n74735 );
nand U119022 ( n13730, n13833, n13834 );
nor U119023 ( n13833, n74658, n73176 );
nand U119024 ( n13893, n14065, n14067 );
nor U119025 ( n14065, n75941, n74461 );
nor U119026 ( n14067, n5219, n74429 );
nor U119027 ( n13539, n13579, n74476 );
nand U119028 ( n12944, n12950, n5217 );
nor U119029 ( n12950, n74886, n12952 );
nor U119030 ( n13834, n13893, n73090 );
nor U119031 ( n13692, n13730, n73109 );
nand U119032 ( n13098, n13102, n5218 );
nor U119033 ( n13102, n73158, n13052 );
nand U119034 ( n13237, n13257, n13258 );
nor U119035 ( n13257, n74599, n13247 );
not U119036 ( n1785, n46220 );
and U119037 ( n12755, n5215, n12778 );
not U119038 ( n2902, n38182 );
nor U119039 ( n43333, n72962, n42617 );
nand U119040 ( n13487, n13637, n13638 );
nor U119041 ( n13637, n74735, n13578 );
nand U119042 ( n14162, n14269, n5225 );
nor U119043 ( n14269, n74429, n73079 );
nand U119044 ( n13219, n13348, n13349 );
nor U119045 ( n13348, n74599, n13350 );
nor U119046 ( n13050, n13197, n13219 );
nor U119047 ( n13944, n14162, n75941 );
nand U119048 ( n12898, n13049, n13050 );
nor U119049 ( n13049, n74653, n13052 );
nor U119050 ( n13349, n13487, n13488 );
and U119051 ( n13638, n13777, n13778 );
nor U119052 ( n13778, n73109, n74658 );
nor U119053 ( n13777, n73176, n13779 );
nand U119054 ( n13889, n14160, n5225 );
nor U119055 ( n14160, n74429, n75941 );
nand U119056 ( n13002, n13155, n13157 );
nor U119057 ( n13155, n74625, n13158 );
nand U119058 ( n13312, n13429, n13430 );
nor U119059 ( n13430, n74818, n73117 );
nor U119060 ( n13429, n74823, n13432 );
nor U119061 ( n13157, n13310, n13312 );
or U119062 ( n13310, n74847, n13313 );
nand U119063 ( n13432, n13577, n5223 );
nor U119064 ( n13577, n74468, n13578 );
nand U119065 ( n13643, n13737, n5224 );
nor U119066 ( n13737, n73176, n13738 );
nor U119067 ( n12838, n13000, n13002 );
or U119068 ( n13000, n74920, n12952 );
nand U119069 ( n12822, n12838, n12839 );
nand U119070 ( n13880, n13887, n13888 );
nor U119071 ( n13887, n74658, n13889 );
nand U119072 ( n47267, n47496, n7879 );
nor U119073 ( n47496, n74400, n75934 );
nor U119074 ( n42345, n42346, n42347 );
nor U119075 ( n42346, n42350, n42351 );
nor U119076 ( n42347, n907, n42348 );
nand U119077 ( n42351, n42352, n42309 );
nand U119078 ( n46787, n46888, n46889 );
nor U119079 ( n46889, n73118, n74417 );
nor U119080 ( n46888, n74822, n46890 );
nand U119081 ( n46536, n46666, n46667 );
nor U119082 ( n46666, n74585, n46668 );
nor U119083 ( n46667, n46786, n46787 );
or U119084 ( n46786, n74841, n46788 );
nand U119085 ( n46890, n47010, n7877 );
nor U119086 ( n47010, n73099, n47011 );
nand U119087 ( n47068, n47137, n7878 );
nor U119088 ( n47137, n73178, n47138 );
nand U119089 ( n42310, n42353, n42354 );
nand U119090 ( n42354, n42256, n42257 );
nor U119091 ( n46410, n46535, n46536 );
or U119092 ( n46535, n73159, n46499 );
nand U119093 ( n46392, n46409, n46410 );
nor U119094 ( n46409, n74919, n46369 );
nand U119095 ( n47260, n47265, n47266 );
nor U119096 ( n47265, n74659, n47267 );
nand U119097 ( n42348, n42349, n42308 );
nand U119098 ( n42349, n910, n42309 );
nand U119099 ( n30112, n30125, n30126 );
nor U119100 ( n30126, n75181, n73387 );
nand U119101 ( n64125, n64138, n64139 );
nor U119102 ( n64139, n75182, n73388 );
nand U119103 ( n22787, n22800, n22801 );
nor U119104 ( n22801, n75183, n73386 );
nand U119105 ( n55901, n55914, n55915 );
nor U119106 ( n55915, n75184, n73389 );
nor U119107 ( n30125, n75171, n30144 );
nor U119108 ( n64138, n75172, n64157 );
nor U119109 ( n22800, n75173, n22819 );
nor U119110 ( n55914, n75174, n55933 );
nor U119111 ( n9384, n72963, n8559 );
not U119112 ( n5579, n66162 );
nand U119113 ( n43381, n43394, n43395 );
nor U119114 ( n43395, n75190, n73385 );
nand U119115 ( n9443, n9459, n9460 );
nor U119116 ( n9460, n75189, n73384 );
nor U119117 ( n43394, n75175, n43413 );
nor U119118 ( n9459, n75176, n9483 );
nand U119119 ( n12759, n12778, n5215 );
not U119120 ( n6454, n57586 );
nand U119121 ( n33218, n33337, n33338 );
nor U119122 ( n33337, n73115, n33287 );
nand U119123 ( n33762, n33848, n3475 );
nor U119124 ( n33848, n74412, n73077 );
nand U119125 ( n32749, n32876, n32877 );
nor U119126 ( n32876, n74671, n32878 );
nand U119127 ( n33002, n33107, n33108 );
nor U119128 ( n33107, n74635, n33109 );
nor U119129 ( n32877, n32985, n33002 );
nor U119130 ( n33587, n33762, n75940 );
nor U119131 ( n33108, n33218, n33219 );
nand U119132 ( n32731, n32747, n32748 );
nor U119133 ( n32748, n74961, n73232 );
nor U119134 ( n32747, n74948, n32749 );
and U119135 ( n33338, n33449, n33450 );
nor U119136 ( n33450, n73114, n74696 );
nor U119137 ( n33449, n73197, n33451 );
nand U119138 ( n67973, n68094, n68095 );
nor U119139 ( n68094, n74758, n68046 );
nand U119140 ( n25970, n26091, n26092 );
nor U119141 ( n26091, n74759, n26043 );
nand U119142 ( n59108, n59232, n59233 );
nor U119143 ( n59232, n74760, n59184 );
nand U119144 ( n68518, n68604, n6090 );
nor U119145 ( n68604, n74408, n73076 );
nand U119146 ( n26517, n26603, n4313 );
nor U119147 ( n26603, n74409, n73075 );
nand U119148 ( n59656, n59745, n6945 );
nor U119149 ( n59745, n74410, n73074 );
nand U119150 ( n67514, n67637, n67638 );
nor U119151 ( n67637, n74916, n67639 );
nand U119152 ( n67758, n67863, n67864 );
nor U119153 ( n67863, n74546, n67865 );
nand U119154 ( n25509, n25632, n25633 );
nor U119155 ( n25632, n74917, n25634 );
nand U119156 ( n25753, n25860, n25861 );
nor U119157 ( n25860, n74547, n25862 );
nand U119158 ( n58646, n58769, n58770 );
nor U119159 ( n58769, n74918, n58771 );
nand U119160 ( n58893, n58998, n58999 );
nor U119161 ( n58998, n74548, n59000 );
nor U119162 ( n67638, n67742, n67758 );
nor U119163 ( n25633, n25737, n25753 );
nor U119164 ( n58770, n58877, n58893 );
nor U119165 ( n68343, n68518, n75937 );
nor U119166 ( n26342, n26517, n75938 );
nor U119167 ( n59481, n59656, n75939 );
nor U119168 ( n67864, n67973, n67974 );
nor U119169 ( n25861, n25970, n25971 );
nor U119170 ( n58999, n59108, n59109 );
nand U119171 ( n25491, n25507, n25508 );
nor U119172 ( n25508, n74960, n73224 );
nor U119173 ( n25507, n74949, n25509 );
nand U119174 ( n67496, n67512, n67513 );
nor U119175 ( n67513, n74962, n73223 );
nor U119176 ( n67512, n74947, n67514 );
nand U119177 ( n58628, n58644, n58645 );
nor U119178 ( n58645, n74963, n73225 );
nor U119179 ( n58644, n74950, n58646 );
and U119180 ( n68095, n68200, n68201 );
nor U119181 ( n68201, n73084, n74695 );
nor U119182 ( n68200, n73187, n68202 );
and U119183 ( n26092, n26199, n26200 );
nor U119184 ( n26200, n73085, n74697 );
nor U119185 ( n26199, n73188, n26201 );
and U119186 ( n59233, n59338, n59339 );
nor U119187 ( n59339, n73086, n74698 );
nor U119188 ( n59338, n73189, n59340 );
not U119189 ( n7879, n47577 );
not U119190 ( n7873, n47660 );
not U119191 ( n5219, n14365 );
nor U119192 ( n57441, n56380, n74490 );
nor U119193 ( n24318, n23256, n74491 );
nor U119194 ( n31614, n30577, n74488 );
nor U119195 ( n65900, n64736, n74487 );
not U119196 ( n7793, n44508 );
not U119197 ( n5138, n10713 );
not U119198 ( n3390, n31129 );
not U119199 ( n6005, n65383 );
nor U119200 ( n30831, n74351, n30832 );
nor U119201 ( n10334, n74375, n10335 );
nor U119202 ( n65033, n74202, n65034 );
nor U119203 ( n44191, n74148, n44192 );
nand U119204 ( n30827, n30828, n30829 );
nor U119205 ( n30828, n30834, n30835 );
nor U119206 ( n30829, n30830, n30831 );
nor U119207 ( n30834, n74353, n30837 );
nand U119208 ( n10329, n10330, n10332 );
nor U119209 ( n10330, n10338, n10339 );
nor U119210 ( n10332, n10333, n10334 );
nor U119211 ( n10338, n74373, n10342 );
nand U119212 ( n65029, n65030, n65031 );
nor U119213 ( n65030, n65036, n65037 );
nor U119214 ( n65031, n65032, n65033 );
nor U119215 ( n65036, n74208, n65039 );
nand U119216 ( n44187, n44188, n44189 );
nor U119217 ( n44188, n44194, n44195 );
nor U119218 ( n44189, n44190, n44191 );
nor U119219 ( n44194, n74158, n44197 );
not U119220 ( n4228, n23837 );
not U119221 ( n6860, n56961 );
nor U119222 ( n23524, n74203, n23525 );
nor U119223 ( n56646, n74204, n56647 );
nand U119224 ( n23520, n23521, n23522 );
nor U119225 ( n23521, n23527, n23528 );
nor U119226 ( n23522, n23523, n23524 );
nor U119227 ( n23527, n74209, n23530 );
nand U119228 ( n56642, n56643, n56644 );
nor U119229 ( n56643, n56649, n56650 );
nor U119230 ( n56644, n56645, n56646 );
nor U119231 ( n56649, n74210, n56652 );
nor U119232 ( n30830, n74355, n30833 );
nor U119233 ( n10333, n74377, n10337 );
nor U119234 ( n65032, n74214, n65035 );
nor U119235 ( n44190, n74160, n44193 );
nor U119236 ( n23523, n74215, n23526 );
nor U119237 ( n56645, n74216, n56648 );
nor U119238 ( n30835, n74348, n30836 );
nor U119239 ( n10339, n74368, n10340 );
nor U119240 ( n65037, n74192, n65038 );
nor U119241 ( n44195, n74145, n44196 );
not U119242 ( n3797, n23824 );
nand U119243 ( n63378, n63385, n63386 );
nor U119244 ( n63386, n63387, n63388 );
nor U119245 ( n63385, n63389, n63390 );
nand U119246 ( n63387, n73037, n73460 );
nand U119247 ( n63390, n73489, n73043 );
nor U119248 ( n23528, n74193, n23529 );
nor U119249 ( n56650, n74194, n56651 );
nor U119250 ( n29160, n74591, n29164 );
nand U119251 ( n29164, n29165, n29163 );
nand U119252 ( n29165, n29172, n29173 );
nor U119253 ( n29172, n29176, n74662 );
nand U119254 ( n29163, n29166, n29167 );
nand U119255 ( n29167, n29168, n74591 );
nor U119256 ( n29166, n29144, n3068 );
nand U119257 ( n29168, n29169, n29170 );
nor U119258 ( n62882, n74593, n62886 );
nand U119259 ( n62886, n62887, n62885 );
nand U119260 ( n62887, n62894, n62895 );
nor U119261 ( n62894, n62898, n74660 );
nor U119262 ( n54938, n74594, n54942 );
nand U119263 ( n54942, n54943, n54941 );
nand U119264 ( n54943, n54950, n54951 );
nor U119265 ( n54950, n54954, n74661 );
nor U119266 ( n21847, n74592, n21851 );
nand U119267 ( n21851, n21852, n21850 );
nand U119268 ( n21852, n21859, n21860 );
nor U119269 ( n21859, n21863, n74663 );
nand U119270 ( n62885, n62888, n62889 );
nand U119271 ( n62889, n62890, n74593 );
nor U119272 ( n62888, n62811, n5669 );
nand U119273 ( n62890, n62891, n62892 );
nand U119274 ( n54941, n54944, n54945 );
nand U119275 ( n54945, n54946, n74594 );
nor U119276 ( n54944, n54905, n6544 );
nand U119277 ( n54946, n54947, n54948 );
nand U119278 ( n21850, n21853, n21854 );
nand U119279 ( n21854, n21855, n74592 );
nor U119280 ( n21853, n21829, n3912 );
nand U119281 ( n21855, n21856, n21857 );
nor U119282 ( n15397, n74435, n5200 );
nor U119283 ( n42373, n74648, n42377 );
nand U119284 ( n42377, n42378, n42376 );
nand U119285 ( n42378, n42385, n42386 );
nor U119286 ( n42385, n42389, n73190 );
nand U119287 ( n42376, n42379, n42380 );
nand U119288 ( n42380, n42381, n74648 );
nor U119289 ( n42379, n42323, n7454 );
nand U119290 ( n42381, n42382, n42383 );
nor U119291 ( n8758, n5274, n8759 );
nor U119292 ( n8759, n8760, n5299 );
not U119293 ( n5299, n8762 );
nor U119294 ( n8760, n8763, n8764 );
nor U119295 ( n42804, n7929, n42805 );
nor U119296 ( n42805, n42806, n7954 );
not U119297 ( n7954, n42807 );
nor U119298 ( n42806, n42808, n42809 );
nand U119299 ( n42301, n42339, n42340 );
nand U119300 ( n42340, n42246, n42247 );
nor U119301 ( n42333, n908, n42334 );
not U119302 ( n908, n42336 );
nand U119303 ( n42334, n42335, n42303 );
nand U119304 ( n42335, n912, n42302 );
nor U119305 ( n13261, n75035, n60062 );
nor U119306 ( n6526, n75033, n26922 );
nor U119307 ( n4281, n75032, n34167 );
nor U119308 ( n11016, n75034, n68921 );
nand U119309 ( n8287, n8290, n8292 );
nand U119310 ( n8292, n8293, n74649 );
nor U119311 ( n8290, n8263, n4810 );
nand U119312 ( n8293, n8294, n8295 );
nor U119313 ( n8283, n74649, n8288 );
nand U119314 ( n8288, n8289, n8287 );
nand U119315 ( n8289, n8298, n8299 );
nor U119316 ( n8298, n8303, n73191 );
nand U119317 ( n42419, n42422, n42423 );
nand U119318 ( n42422, n42424, n42425 );
nand U119319 ( n63388, n73466, n73036 );
nand U119320 ( n63396, n73031, n73444 );
nand U119321 ( n63395, n73033, n73454 );
not U119322 ( n5253, n13158 );
nand U119323 ( n63389, n73476, n73040 );
nand U119324 ( n63402, n73048, n73507 );
nor U119325 ( n30841, n74341, n30842 );
nor U119326 ( n10347, n74361, n10348 );
nor U119327 ( n65043, n74177, n65044 );
nor U119328 ( n44201, n74132, n44202 );
nand U119329 ( n30826, n30838, n30839 );
nor U119330 ( n30838, n30844, n30845 );
nor U119331 ( n30839, n30840, n30841 );
nor U119332 ( n30844, n74347, n30847 );
nand U119333 ( n10328, n10343, n10344 );
nor U119334 ( n10343, n10350, n10352 );
nor U119335 ( n10344, n10345, n10347 );
nor U119336 ( n10350, n74370, n10354 );
nand U119337 ( n65028, n65040, n65041 );
nor U119338 ( n65040, n65046, n65047 );
nor U119339 ( n65041, n65042, n65043 );
nor U119340 ( n65046, n74189, n65049 );
nand U119341 ( n44186, n44198, n44199 );
nor U119342 ( n44198, n44204, n44205 );
nor U119343 ( n44199, n44200, n44201 );
nor U119344 ( n44204, n74144, n44207 );
nor U119345 ( n23534, n74178, n23535 );
nor U119346 ( n56656, n74179, n56657 );
nand U119347 ( n23519, n23531, n23532 );
nor U119348 ( n23531, n23537, n23538 );
nor U119349 ( n23532, n23533, n23534 );
nor U119350 ( n23537, n74190, n23540 );
nand U119351 ( n56641, n56653, n56654 );
nor U119352 ( n56653, n56659, n56660 );
nor U119353 ( n56654, n56655, n56656 );
nor U119354 ( n56659, n74191, n56662 );
nand U119355 ( n44203, n44539, n44507 );
nor U119356 ( n44539, n7793, n44511 );
nand U119357 ( n10349, n10752, n10712 );
nor U119358 ( n10752, n5138, n10717 );
nand U119359 ( n30843, n31160, n31128 );
nor U119360 ( n31160, n3390, n31132 );
nand U119361 ( n65045, n65414, n65382 );
nor U119362 ( n65414, n6005, n65386 );
nor U119363 ( n30840, n74350, n30843 );
nor U119364 ( n10345, n74376, n10349 );
nor U119365 ( n65042, n74199, n65045 );
nor U119366 ( n44200, n74147, n44203 );
nand U119367 ( n12615, n14388, n14389 );
nand U119368 ( n14388, n4969, n14393 );
nand U119369 ( n14389, n14390, n14353 );
nand U119370 ( n14390, n4952, n14183 );
nand U119371 ( n23536, n23868, n23836 );
nor U119372 ( n23868, n4228, n23840 );
nand U119373 ( n56658, n56992, n56960 );
nor U119374 ( n56992, n6860, n56964 );
nor U119375 ( n23533, n74200, n23536 );
nor U119376 ( n56655, n74201, n56658 );
nand U119377 ( n44206, n44542, n44507 );
nor U119378 ( n44542, n7793, n44515 );
nand U119379 ( n10353, n10755, n10712 );
nor U119380 ( n10755, n5138, n10722 );
nand U119381 ( n30846, n31163, n31128 );
nor U119382 ( n31163, n3390, n31136 );
nand U119383 ( n65048, n65417, n65382 );
nor U119384 ( n65417, n6005, n65390 );
nor U119385 ( n30845, n74340, n30846 );
nor U119386 ( n10352, n74362, n10353 );
nor U119387 ( n65047, n74174, n65048 );
nor U119388 ( n44205, n74133, n44206 );
nand U119389 ( n23539, n23871, n23836 );
nor U119390 ( n23871, n4228, n23844 );
nand U119391 ( n56661, n56995, n56960 );
nor U119392 ( n56995, n6860, n56968 );
nor U119393 ( n23538, n74175, n23539 );
nor U119394 ( n56660, n74176, n56661 );
nor U119395 ( n48142, n47935, n74442 );
nand U119396 ( n68047, n68131, n68132 );
nor U119397 ( n68131, n72950, n74758 );
nand U119398 ( n33288, n33379, n33380 );
nor U119399 ( n33379, n74755, n73115 );
nand U119400 ( n26044, n26128, n26129 );
nor U119401 ( n26128, n72951, n74759 );
nand U119402 ( n59185, n59269, n59270 );
nor U119403 ( n59269, n72952, n74760 );
nand U119404 ( n68163, n68252, n68253 );
nor U119405 ( n68252, n74695, n73187 );
nand U119406 ( n33413, n33497, n33498 );
nor U119407 ( n33497, n74696, n73197 );
nand U119408 ( n26162, n26251, n26252 );
nor U119409 ( n26251, n74697, n73188 );
nand U119410 ( n59301, n59390, n59391 );
nor U119411 ( n59390, n74698, n73189 );
nand U119412 ( n68301, n68440, n68441 );
nor U119413 ( n68440, n75937, n74452 );
nor U119414 ( n68441, n6083, n74408 );
nand U119415 ( n33545, n33684, n33685 );
nor U119416 ( n33684, n75940, n74455 );
nor U119417 ( n33685, n3468, n74412 );
nand U119418 ( n26300, n26439, n26440 );
nor U119419 ( n26439, n75938, n74453 );
nor U119420 ( n26440, n4305, n74409 );
nand U119421 ( n59439, n59578, n59579 );
nor U119422 ( n59578, n75939, n74454 );
nor U119423 ( n59579, n6938, n74410 );
nor U119424 ( n33256, n33288, n74458 );
nor U119425 ( n68015, n68047, n74438 );
nor U119426 ( n26012, n26044, n74439 );
nor U119427 ( n59150, n59185, n74440 );
nand U119428 ( n25549, n25556, n4303 );
nor U119429 ( n25556, n25557, n74949 );
nand U119430 ( n58686, n58693, n6935 );
nor U119431 ( n58693, n58694, n74950 );
nand U119432 ( n32789, n32796, n3465 );
nor U119433 ( n32796, n32797, n74948 );
nand U119434 ( n67554, n67561, n6080 );
nor U119435 ( n67561, n67562, n74947 );
nor U119436 ( n68253, n68301, n73066 );
nor U119437 ( n26252, n26300, n73067 );
nor U119438 ( n59391, n59439, n73068 );
nor U119439 ( n33498, n33545, n73088 );
nor U119440 ( n68132, n68163, n73084 );
nor U119441 ( n26129, n26162, n73085 );
nor U119442 ( n59270, n59301, n73086 );
nor U119443 ( n33380, n33413, n73114 );
nand U119444 ( n25669, n25672, n4304 );
nor U119445 ( n25672, n73150, n25634 );
nand U119446 ( n58809, n58812, n6937 );
nor U119447 ( n58812, n73151, n58771 );
nand U119448 ( n32913, n32916, n3467 );
nor U119449 ( n32916, n73167, n32878 );
nand U119450 ( n67674, n67677, n6082 );
nor U119451 ( n67677, n73149, n67639 );
nand U119452 ( n25769, n25784, n25785 );
nor U119453 ( n25784, n74547, n25778 );
nand U119454 ( n58907, n58922, n58923 );
nor U119455 ( n58922, n74548, n58916 );
nand U119456 ( n33016, n33032, n33033 );
nor U119457 ( n33032, n74635, n33024 );
nand U119458 ( n67772, n67787, n67788 );
nor U119459 ( n67787, n74546, n67781 );
nor U119460 ( n42332, n42336, n42337 );
nand U119461 ( n42337, n42338, n42302 );
nand U119462 ( n42338, n42301, n42303 );
nor U119463 ( n45145, n852, n45077 );
not U119464 ( n852, n45010 );
not U119465 ( n1784, n46549 );
not U119466 ( n2900, n38195 );
not U119467 ( n5225, n14262 );
not U119468 ( n850, n45018 );
nand U119469 ( n22477, n22564, n22565 );
nor U119470 ( n22564, n74710, n73199 );
nor U119471 ( n22565, n22566, n74694 );
nand U119472 ( n22566, n22633, n22634 );
nor U119473 ( n22633, n72961, n74641 );
nor U119474 ( n22634, n72958, n74620 );
nand U119475 ( n55592, n55677, n55678 );
nor U119476 ( n55677, n74709, n73198 );
nor U119477 ( n55678, n55679, n74693 );
nand U119478 ( n55679, n55746, n55747 );
nor U119479 ( n55746, n72960, n74640 );
nor U119480 ( n55747, n72959, n74619 );
nand U119481 ( n22233, n22324, n22325 );
nor U119482 ( n22324, n74838, n73248 );
nor U119483 ( n22325, n22326, n74828 );
nand U119484 ( n22326, n22406, n22407 );
nor U119485 ( n22406, n74799, n73234 );
nor U119486 ( n22407, n22408, n74789 );
nand U119487 ( n55345, n55436, n55437 );
nor U119488 ( n55436, n74837, n73247 );
nor U119489 ( n55437, n55438, n74827 );
nand U119490 ( n55438, n55518, n55519 );
nor U119491 ( n55518, n74798, n73233 );
nor U119492 ( n55519, n55520, n74788 );
nand U119493 ( n22170, n22231, n22232 );
nor U119494 ( n22231, n74899, n73262 );
nor U119495 ( n22232, n22233, n74883 );
nand U119496 ( n22079, n22168, n22169 );
nor U119497 ( n22168, n74939, n73276 );
nor U119498 ( n22169, n22170, n74926 );
nand U119499 ( n55284, n55343, n55344 );
nor U119500 ( n55343, n74898, n73261 );
nor U119501 ( n55344, n55345, n74882 );
nand U119502 ( n55189, n55282, n55283 );
nor U119503 ( n55282, n74938, n73275 );
nor U119504 ( n55283, n55284, n74925 );
xor U119505 ( n21948, n75178, n21949 );
nand U119506 ( n21949, n21946, n21947 );
xor U119507 ( n55060, n75177, n55061 );
nand U119508 ( n55061, n55058, n55059 );
nand U119509 ( n22075, n22077, n22078 );
nor U119510 ( n22077, n74991, n73291 );
nor U119511 ( n22078, n22079, n74970 );
nand U119512 ( n55185, n55187, n55188 );
nor U119513 ( n55187, n74990, n73290 );
nor U119514 ( n55188, n55189, n74969 );
nand U119515 ( n21998, n4643, n22001 );
nand U119516 ( n55108, n7275, n55111 );
nand U119517 ( n22408, n22475, n22476 );
nor U119518 ( n22475, n74748, n73215 );
nor U119519 ( n22476, n22477, n74744 );
nand U119520 ( n55520, n55590, n55591 );
nor U119521 ( n55590, n74747, n73214 );
nor U119522 ( n55591, n55592, n74743 );
nand U119523 ( n63758, n63843, n63844 );
nor U119524 ( n63843, n74711, n72966 );
nor U119525 ( n63844, n63845, n73193 );
nand U119526 ( n63845, n63912, n63913 );
nor U119527 ( n63912, n73168, n74642 );
nor U119528 ( n63913, n73163, n74621 );
nand U119529 ( n29798, n29887, n29888 );
nor U119530 ( n29887, n74712, n72967 );
nor U119531 ( n29888, n29889, n73194 );
nand U119532 ( n29889, n29956, n29957 );
nor U119533 ( n29956, n73169, n74643 );
nor U119534 ( n29957, n73164, n74622 );
nand U119535 ( n63252, n63451, n63452 );
nor U119536 ( n63451, n74900, n73263 );
nor U119537 ( n63452, n63453, n74884 );
nand U119538 ( n63453, n63544, n63545 );
nor U119539 ( n63544, n74840, n73249 );
nor U119540 ( n63545, n63546, n74830 );
nand U119541 ( n63546, n63626, n63627 );
nor U119542 ( n63626, n74800, n73236 );
nor U119543 ( n63627, n63628, n74790 );
nand U119544 ( n29489, n29548, n29549 );
nor U119545 ( n29548, n74901, n73264 );
nor U119546 ( n29549, n29550, n74885 );
nand U119547 ( n29550, n29645, n29646 );
nor U119548 ( n29645, n74839, n73250 );
nor U119549 ( n29646, n29647, n74829 );
nand U119550 ( n29647, n29727, n29728 );
nor U119551 ( n29727, n74801, n73235 );
nor U119552 ( n29728, n29729, n74791 );
nand U119553 ( n63161, n63250, n63251 );
nor U119554 ( n63250, n74944, n73277 );
nor U119555 ( n63251, n63252, n74928 );
nand U119556 ( n29398, n29487, n29488 );
nor U119557 ( n29487, n74945, n73278 );
nor U119558 ( n29488, n29489, n74929 );
xor U119559 ( n63032, n75179, n63033 );
nand U119560 ( n63033, n63030, n63031 );
xor U119561 ( n29265, n75180, n29266 );
nand U119562 ( n29266, n29263, n29264 );
nand U119563 ( n63157, n63159, n63160 );
nor U119564 ( n63159, n74993, n73292 );
nor U119565 ( n63160, n63161, n74987 );
nand U119566 ( n29394, n29396, n29397 );
nor U119567 ( n29396, n74994, n73293 );
nor U119568 ( n29397, n29398, n74988 );
nand U119569 ( n63080, n6383, n63083 );
nand U119570 ( n29317, n3749, n29320 );
nand U119571 ( n63628, n63756, n63757 );
nor U119572 ( n63756, n74749, n73216 );
nor U119573 ( n63757, n63758, n74745 );
nand U119574 ( n29729, n29796, n29797 );
nor U119575 ( n29796, n74750, n73217 );
nor U119576 ( n29797, n29798, n74746 );
nor U119577 ( n42259, n73911, n42260 );
xor U119578 ( n42260, n42251, n42256 );
nand U119579 ( n42253, n42254, n42255 );
nand U119580 ( n42255, n913, n42256 );
nor U119581 ( n42254, n42258, n42259 );
not U119582 ( n913, n42257 );
xor U119583 ( n12619, n14353, n14393 );
nand U119584 ( n8285, n73191, n74685 );
xor U119585 ( n67203, n68671, n68712 );
xor U119586 ( n46251, n47650, n47691 );
nand U119587 ( n9432, n21121, n76188 );
nor U119588 ( n21121, n74649, n8285 );
xor U119589 ( n25305, n26670, n26711 );
xor U119590 ( n58444, n59812, n59853 );
xor U119591 ( n32547, n33915, n33956 );
nor U119592 ( n47266, n74443, n73065 );
not U119593 ( n3475, n33842 );
not U119594 ( n6090, n68598 );
not U119595 ( n4313, n26597 );
not U119596 ( n6945, n59739 );
not U119597 ( n849, n45007 );
nand U119598 ( n45011, n849, n74415 );
nand U119599 ( n68299, n68517, n6090 );
nor U119600 ( n68517, n74408, n75937 );
nand U119601 ( n33543, n33761, n3475 );
nor U119602 ( n33761, n74412, n75940 );
nand U119603 ( n26298, n26516, n4313 );
nor U119604 ( n26516, n74409, n75938 );
nand U119605 ( n59437, n59655, n6945 );
nor U119606 ( n59655, n74410, n75939 );
nand U119607 ( n67598, n67713, n67714 );
nor U119608 ( n67713, n74595, n67715 );
nand U119609 ( n32833, n32959, n32960 );
nor U119610 ( n32959, n74652, n32961 );
nand U119611 ( n25593, n25708, n25709 );
nor U119612 ( n25708, n74596, n25710 );
nand U119613 ( n58730, n58848, n58849 );
nor U119614 ( n58848, n74597, n58850 );
nand U119615 ( n67834, n67935, n67936 );
nor U119616 ( n67936, n73130, n74431 );
nor U119617 ( n67935, n74852, n67937 );
nand U119618 ( n33078, n33172, n33173 );
nor U119619 ( n33173, n74845, n73160 );
nor U119620 ( n33172, n74855, n33174 );
nand U119621 ( n25831, n25932, n25933 );
nor U119622 ( n25933, n73131, n74432 );
nor U119623 ( n25932, n74853, n25934 );
nand U119624 ( n58969, n59070, n59071 );
nor U119625 ( n59071, n73132, n74433 );
nor U119626 ( n59070, n74854, n59072 );
nor U119627 ( n67714, n67833, n67834 );
or U119628 ( n67833, n74872, n67835 );
nor U119629 ( n32960, n33077, n33078 );
or U119630 ( n33077, n74879, n33079 );
nor U119631 ( n25709, n25830, n25831 );
or U119632 ( n25830, n74873, n25832 );
nor U119633 ( n58849, n58968, n58969 );
or U119634 ( n58968, n74874, n58970 );
not U119635 ( n6083, n68681 );
not U119636 ( n3468, n33925 );
not U119637 ( n4305, n26680 );
not U119638 ( n6938, n59822 );
nand U119639 ( n67937, n68045, n6088 );
nor U119640 ( n68045, n73104, n68046 );
nand U119641 ( n33174, n33286, n3473 );
nor U119642 ( n33286, n74460, n33287 );
nand U119643 ( n25934, n26042, n4310 );
nor U119644 ( n26042, n73105, n26043 );
nand U119645 ( n59072, n59183, n6943 );
nor U119646 ( n59183, n73106, n59184 );
nand U119647 ( n68099, n68168, n6089 );
nor U119648 ( n68168, n73187, n68169 );
nand U119649 ( n33342, n33418, n3474 );
nor U119650 ( n33418, n73197, n33419 );
nand U119651 ( n26096, n26167, n4312 );
nor U119652 ( n26167, n73188, n26168 );
nand U119653 ( n59237, n59306, n6944 );
nor U119654 ( n59306, n73189, n59307 );
nand U119655 ( n67456, n67473, n67474 );
nor U119656 ( n67473, n74947, n67433 );
nand U119657 ( n32691, n32708, n32709 );
nor U119658 ( n32708, n74948, n32668 );
nand U119659 ( n25451, n25468, n25469 );
nor U119660 ( n25468, n74949, n25428 );
nand U119661 ( n58588, n58605, n58606 );
nor U119662 ( n58605, n74950, n58565 );
nand U119663 ( n68291, n68297, n68298 );
nor U119664 ( n68297, n74695, n68299 );
nand U119665 ( n33535, n33541, n33542 );
nor U119666 ( n33541, n74696, n33543 );
nand U119667 ( n26290, n26296, n26297 );
nor U119668 ( n26296, n74697, n26298 );
nand U119669 ( n59429, n59435, n59436 );
nor U119670 ( n59435, n74698, n59437 );
nand U119671 ( n45019, n849, n74416 );
nand U119672 ( n9059, n9165, n9167 );
nor U119673 ( n9165, n74729, n73207 );
nor U119674 ( n9167, n9168, n74727 );
nand U119675 ( n9168, n9252, n9253 );
nor U119676 ( n9252, n72965, n74673 );
nor U119677 ( n9253, n72963, n74656 );
nand U119678 ( n43059, n43144, n43145 );
nor U119679 ( n43144, n74728, n73206 );
nor U119680 ( n43145, n43146, n74726 );
nand U119681 ( n43146, n43213, n43214 );
nor U119682 ( n43213, n72964, n74672 );
nor U119683 ( n43214, n72962, n74655 );
nand U119684 ( n8678, n8752, n8753 );
nor U119685 ( n8752, n74915, n73268 );
nor U119686 ( n8753, n8754, n74905 );
nand U119687 ( n42801, n42892, n42893 );
nor U119688 ( n42892, n74868, n73253 );
nor U119689 ( n42893, n42894, n74860 );
nand U119690 ( n8754, n8868, n8869 );
nor U119691 ( n8868, n74869, n73254 );
nor U119692 ( n8869, n8870, n74861 );
nand U119693 ( n8870, n8970, n8972 );
nor U119694 ( n8970, n74816, n73240 );
nor U119695 ( n8972, n8973, n74812 );
nand U119696 ( n42736, n42799, n42800 );
nor U119697 ( n42799, n74914, n73267 );
nor U119698 ( n42800, n42801, n74904 );
nand U119699 ( n42894, n42988, n42989 );
nor U119700 ( n42988, n74815, n73239 );
nor U119701 ( n42989, n42990, n74811 );
nand U119702 ( n42621, n42734, n42735 );
nor U119703 ( n42734, n74958, n73280 );
nor U119704 ( n42735, n42736, n74951 );
nand U119705 ( n8564, n8675, n8677 );
nor U119706 ( n8675, n74959, n73281 );
nor U119707 ( n8677, n8678, n74952 );
nand U119708 ( n42616, n42619, n42620 );
nor U119709 ( n42619, n75005, n73304 );
nor U119710 ( n42620, n42621, n74995 );
nand U119711 ( n8558, n8562, n8563 );
nor U119712 ( n8562, n75006, n73305 );
nor U119713 ( n8563, n8564, n74996 );
nand U119714 ( n8973, n9057, n9058 );
nor U119715 ( n9057, n75967, n73222 );
nor U119716 ( n9058, n9059, n74770 );
nand U119717 ( n42990, n43057, n43058 );
nor U119718 ( n43057, n75965, n73221 );
nor U119719 ( n43058, n43059, n74769 );
and U119720 ( n42537, n8164, n42543 );
and U119721 ( n8460, n5510, n8468 );
nor U119722 ( n27462, n74423, n4287 );
nor U119723 ( n60611, n74424, n6919 );
and U119724 ( n21946, n4643, n22001 );
and U119725 ( n55058, n7275, n55111 );
nor U119726 ( n69451, n74425, n6064 );
nor U119727 ( n34707, n74426, n3449 );
nand U119728 ( n42375, n73190, n74686 );
nand U119729 ( n43372, n54104, n76178 );
nor U119730 ( n54104, n74648, n42375 );
and U119731 ( n63030, n6383, n63083 );
and U119732 ( n29263, n3749, n29320 );
xor U119733 ( n16717, n16726, n73430 );
xor U119734 ( n42250, n42251, n42246 );
nor U119735 ( n42244, n42248, n42249 );
nor U119736 ( n42248, n42246, n42252 );
nor U119737 ( n42249, n73910, n42250 );
nand U119738 ( n42252, n42251, n73910 );
nor U119739 ( n44522, n44507, n44508 );
nor U119740 ( n31143, n31128, n31129 );
nor U119741 ( n65397, n65382, n65383 );
nor U119742 ( n30819, n74339, n30820 );
nor U119743 ( n65021, n74171, n65022 );
nor U119744 ( n44179, n74130, n44180 );
nand U119745 ( n30804, n30816, n30817 );
nor U119746 ( n30816, n30822, n30823 );
nor U119747 ( n30817, n30818, n30819 );
nor U119748 ( n30822, n74343, n30825 );
nand U119749 ( n65006, n65018, n65019 );
nor U119750 ( n65018, n65024, n65025 );
nor U119751 ( n65019, n65020, n65021 );
nor U119752 ( n65024, n74180, n65027 );
nand U119753 ( n44164, n44176, n44177 );
nor U119754 ( n44176, n44182, n44183 );
nor U119755 ( n44177, n44178, n44179 );
nor U119756 ( n44182, n74135, n44185 );
nor U119757 ( n23851, n23836, n23837 );
nor U119758 ( n56975, n56960, n56961 );
nor U119759 ( n23512, n74172, n23513 );
nor U119760 ( n56634, n74173, n56635 );
nand U119761 ( n23497, n23509, n23510 );
nor U119762 ( n23509, n23515, n23516 );
nor U119763 ( n23510, n23511, n23512 );
nor U119764 ( n23515, n74182, n23518 );
nand U119765 ( n56619, n56631, n56632 );
nor U119766 ( n56631, n56637, n56638 );
nor U119767 ( n56632, n56633, n56634 );
nor U119768 ( n56637, n74183, n56640 );
nor U119769 ( n30818, n74345, n30821 );
nor U119770 ( n65020, n74186, n65023 );
nor U119771 ( n44178, n74141, n44181 );
nor U119772 ( n23511, n74187, n23514 );
nor U119773 ( n56633, n74188, n56636 );
nor U119774 ( n30823, n74338, n30824 );
nor U119775 ( n65025, n74167, n65026 );
nor U119776 ( n44183, n74106, n44184 );
nor U119777 ( n23516, n74168, n23517 );
nor U119778 ( n56638, n74169, n56639 );
not U119779 ( n7343, n43348 );
nor U119780 ( n10730, n10712, n10713 );
nor U119781 ( n10319, n74359, n10320 );
nand U119782 ( n10300, n10315, n10317 );
nor U119783 ( n10315, n10323, n10324 );
nor U119784 ( n10317, n10318, n10319 );
nor U119785 ( n10323, n74364, n10327 );
nor U119786 ( n10318, n74367, n10322 );
nand U119787 ( n11573, n11574, n622 );
nor U119788 ( n10324, n74357, n10325 );
not U119789 ( n2899, n38211 );
nor U119790 ( n27214, n4293, n74423 );
nor U119791 ( n60359, n6925, n74424 );
nor U119792 ( n34459, n3455, n74426 );
nor U119793 ( n69209, n6070, n74425 );
not U119794 ( n1783, n46937 );
not U119795 ( n4711, n9402 );
nor U119796 ( n44544, n73511, n7817 );
nor U119797 ( n10758, n73527, n5162 );
nor U119798 ( n31165, n73526, n3414 );
nor U119799 ( n65419, n73515, n6029 );
nor U119800 ( n23873, n73516, n4252 );
nor U119801 ( n56997, n73517, n6884 );
nand U119802 ( n14640, n4813, n73191 );
and U119803 ( n9433, n74649, n8264 );
and U119804 ( n63457, n75868, n63459 );
or U119805 ( n75868, n63460, n63461 );
and U119806 ( n29554, n75869, n29556 );
or U119807 ( n75869, n29557, n29558 );
and U119808 ( n22237, n75870, n22239 );
or U119809 ( n75870, n22240, n22241 );
and U119810 ( n55349, n75871, n55351 );
or U119811 ( n75871, n55352, n55353 );
nand U119812 ( n23503, n23835, n23836 );
nor U119813 ( n23835, n23837, n23838 );
nand U119814 ( n56625, n56959, n56960 );
nor U119815 ( n56959, n56961, n56962 );
nor U119816 ( n23500, n23501, n23502 );
nor U119817 ( n23501, n74212, n23504 );
nor U119818 ( n23502, n74196, n23503 );
nor U119819 ( n56622, n56623, n56624 );
nor U119820 ( n56623, n74213, n56626 );
nor U119821 ( n56624, n74197, n56625 );
xor U119822 ( n37983, n74483, n38038 );
nand U119823 ( n44170, n44506, n44507 );
nor U119824 ( n44506, n44508, n44509 );
nand U119825 ( n10308, n10710, n10712 );
nor U119826 ( n10710, n10713, n10714 );
nand U119827 ( n30810, n31127, n31128 );
nor U119828 ( n31127, n31129, n31130 );
nand U119829 ( n65012, n65381, n65382 );
nor U119830 ( n65381, n65383, n65384 );
nor U119831 ( n30807, n30808, n30809 );
nor U119832 ( n30808, n74354, n30811 );
nor U119833 ( n30809, n74349, n30810 );
nor U119834 ( n10304, n10305, n10307 );
nor U119835 ( n10305, n74374, n10309 );
nor U119836 ( n10307, n74369, n10308 );
nor U119837 ( n65009, n65010, n65011 );
nor U119838 ( n65010, n74211, n65013 );
nor U119839 ( n65011, n74195, n65012 );
nor U119840 ( n44167, n44168, n44169 );
nor U119841 ( n44168, n74159, n44171 );
nor U119842 ( n44169, n74146, n44170 );
nand U119843 ( n23507, n23843, n23836 );
nor U119844 ( n23843, n23837, n23844 );
nand U119845 ( n56629, n56967, n56960 );
nor U119846 ( n56967, n56961, n56968 );
nor U119847 ( n23499, n23505, n23506 );
nor U119848 ( n23505, n74206, n23508 );
nor U119849 ( n23506, n74184, n23507 );
nor U119850 ( n56621, n56627, n56628 );
nor U119851 ( n56627, n74207, n56630 );
nor U119852 ( n56628, n74185, n56629 );
xor U119853 ( n38043, n74482, n38038 );
nor U119854 ( n42827, n7930, n42808 );
nor U119855 ( n8787, n5275, n8763 );
nand U119856 ( n44174, n44514, n44507 );
nor U119857 ( n44514, n44508, n44515 );
nand U119858 ( n10313, n10720, n10712 );
nor U119859 ( n10720, n10713, n10722 );
nand U119860 ( n30814, n31135, n31128 );
nor U119861 ( n31135, n31129, n31136 );
nand U119862 ( n65016, n65389, n65382 );
nor U119863 ( n65389, n65383, n65390 );
nor U119864 ( n30806, n30812, n30813 );
nor U119865 ( n30812, n74352, n30815 );
nor U119866 ( n30813, n74344, n30814 );
nor U119867 ( n10303, n10310, n10312 );
nor U119868 ( n10310, n74365, n10314 );
nor U119869 ( n10312, n74363, n10313 );
nor U119870 ( n65008, n65014, n65015 );
nor U119871 ( n65014, n74205, n65017 );
nor U119872 ( n65015, n74181, n65016 );
nor U119873 ( n44166, n44172, n44173 );
nor U119874 ( n44172, n74151, n44175 );
nor U119875 ( n44173, n74138, n44174 );
nor U119876 ( n54900, n54905, n54906 );
nor U119877 ( n21824, n21829, n21830 );
nor U119878 ( n29139, n29144, n29145 );
nor U119879 ( n62806, n62811, n62812 );
nor U119880 ( n46954, n73099, n74417 );
nand U119881 ( n44171, n44510, n44507 );
nor U119882 ( n44510, n44508, n44511 );
nand U119883 ( n30811, n31131, n31128 );
nor U119884 ( n31131, n31129, n31132 );
nand U119885 ( n65013, n65385, n65382 );
nor U119886 ( n65385, n65383, n65386 );
nand U119887 ( n26968, n26955, n27213 );
nand U119888 ( n34213, n34200, n34458 );
nand U119889 ( n68967, n68954, n69208 );
nand U119890 ( n60108, n60095, n60358 );
nand U119891 ( n23504, n23839, n23836 );
nor U119892 ( n23839, n23837, n23840 );
nand U119893 ( n56626, n56963, n56960 );
nor U119894 ( n56963, n56961, n56964 );
nor U119895 ( n42318, n42323, n42324 );
nand U119896 ( n47873, n7457, n73190 );
and U119897 ( n43373, n74648, n42324 );
nand U119898 ( n10309, n10715, n10712 );
nor U119899 ( n10715, n10713, n10717 );
nand U119900 ( n44175, n44516, n44507 );
nor U119901 ( n44516, n44508, n44517 );
nand U119902 ( n30815, n31137, n31128 );
nor U119903 ( n31137, n31129, n31138 );
nand U119904 ( n65017, n65391, n65382 );
nor U119905 ( n65391, n65383, n65392 );
nand U119906 ( n23508, n23845, n23836 );
nor U119907 ( n23845, n23837, n23846 );
nand U119908 ( n56630, n56969, n56960 );
nor U119909 ( n56969, n56961, n56970 );
nand U119910 ( n10314, n10723, n10712 );
nor U119911 ( n10723, n10713, n10724 );
nor U119912 ( n8257, n8263, n8264 );
nand U119913 ( n10475, n10530, n10532 );
nor U119914 ( n10530, n74909, n73266 );
nand U119915 ( n9907, n9968, n9969 );
nor U119916 ( n9968, n75085, n73321 );
nand U119917 ( n10068, n10132, n10133 );
nor U119918 ( n10132, n75013, n73307 );
nand U119919 ( n10245, n10369, n10370 );
nor U119920 ( n10369, n74966, n73289 );
nand U119921 ( n43807, n43891, n43892 );
nor U119922 ( n43891, n75084, n73320 );
nand U119923 ( n44304, n44348, n44349 );
nor U119924 ( n44348, n74908, n73265 );
nand U119925 ( n43982, n44029, n44030 );
nor U119926 ( n44029, n75012, n73306 );
nand U119927 ( n44120, n44219, n44220 );
nor U119928 ( n44219, n74965, n73288 );
nand U119929 ( n44447, n44491, n44492 );
nor U119930 ( n44491, n73251, n74865 );
nand U119931 ( n10637, n10692, n10693 );
nor U119932 ( n10692, n73252, n74864 );
nand U119933 ( n11002, n11050, n11052 );
nor U119934 ( n11050, n73219, n74756 );
nand U119935 ( n11152, n11222, n11223 );
nor U119936 ( n11222, n73196, n74705 );
nand U119937 ( n44734, n44773, n44774 );
nor U119938 ( n44773, n73218, n74757 );
nand U119939 ( n10852, n10900, n10902 );
nor U119940 ( n10900, n73238, n74802 );
nand U119941 ( n11254, n11265, n11267 );
nor U119942 ( n11265, n73166, n74630 );
nand U119943 ( n44868, n44924, n44925 );
nor U119944 ( n44924, n73195, n74704 );
nand U119945 ( n44945, n44954, n44955 );
nor U119946 ( n44954, n73165, n74631 );
nand U119947 ( n44614, n44653, n44654 );
nor U119948 ( n44653, n73237, n74803 );
nor U119949 ( n10532, n10637, n74903 );
nor U119950 ( n9969, n10068, n75062 );
nor U119951 ( n10133, n10245, n75002 );
nor U119952 ( n10370, n10475, n74954 );
nor U119953 ( n43892, n43982, n75061 );
nor U119954 ( n44349, n44447, n74902 );
nor U119955 ( n44030, n44120, n75001 );
nor U119956 ( n44220, n44304, n74953 );
nor U119957 ( n11052, n11152, n74739 );
nor U119958 ( n11223, n11254, n74682 );
nor U119959 ( n44774, n44868, n74738 );
nor U119960 ( n10902, n11002, n74787 );
nor U119961 ( n44925, n44945, n74681 );
nor U119962 ( n44654, n44734, n74786 );
nor U119963 ( n44492, n44614, n74842 );
nor U119964 ( n10693, n10852, n74843 );
nor U119965 ( n14958, n15062, n74435 );
nor U119966 ( n54197, n73511, n73052 );
nor U119967 ( n35699, n73526, n73059 );
nor U119968 ( n28520, n73516, n73055 );
nor U119969 ( n70425, n73515, n73053 );
nor U119970 ( n61825, n73517, n73054 );
nor U119971 ( n13888, n74461, n73090 );
nor U119972 ( n11267, n73162, n74608 );
nor U119973 ( n44955, n73161, n74609 );
nand U119974 ( n8776, n14719, n14720 );
nor U119975 ( n14719, n14737, n14738 );
nor U119976 ( n14720, n14722, n14723 );
nor U119977 ( n14737, n4813, n14739 );
nand U119978 ( n61685, n61692, n61693 );
nor U119979 ( n61693, n61694, n61695 );
nor U119980 ( n61692, n61696, n61697 );
nand U119981 ( n61694, n73061, n73821 );
nand U119982 ( n61697, n73027, n73472 );
not U119983 ( n853, n45083 );
nor U119984 ( n33542, n74455, n73088 );
nor U119985 ( n68298, n74452, n73066 );
nor U119986 ( n26297, n74453, n73067 );
nor U119987 ( n59436, n74454, n73068 );
nor U119988 ( n30771, n3397, n30801 );
nor U119989 ( n10259, n5144, n10297 );
nor U119990 ( n64973, n6012, n65003 );
nor U119991 ( n44131, n7799, n44161 );
nor U119992 ( n30783, n3395, n73526 );
nor U119993 ( n10274, n5143, n73527 );
nor U119994 ( n64985, n6010, n73515 );
nor U119995 ( n44143, n7798, n73511 );
nor U119996 ( n30780, n74008, n30464 );
nor U119997 ( n10270, n74038, n9873 );
nor U119998 ( n64982, n73676, n64623 );
nor U119999 ( n44140, n73562, n43780 );
nand U120000 ( n10252, n10268, n10269 );
nor U120001 ( n10268, n10275, n10277 );
nor U120002 ( n10269, n10270, n10272 );
nor U120003 ( n10275, n74026, n9868 );
nand U120004 ( n30765, n30778, n30779 );
nor U120005 ( n30778, n30784, n30785 );
nor U120006 ( n30779, n30780, n30781 );
nor U120007 ( n30784, n74003, n30460 );
nand U120008 ( n64967, n64980, n64981 );
nor U120009 ( n64980, n64986, n64987 );
nor U120010 ( n64981, n64982, n64983 );
nor U120011 ( n64986, n73665, n64619 );
nand U120012 ( n44125, n44138, n44139 );
nor U120013 ( n44138, n44144, n44145 );
nor U120014 ( n44139, n44140, n44141 );
nor U120015 ( n44144, n73557, n43776 );
nand U120016 ( n62884, n74660, n73183 );
nand U120017 ( n29162, n74662, n73182 );
nand U120018 ( n54940, n74661, n73180 );
nand U120019 ( n21849, n74663, n73181 );
xnor U120020 ( n67330, n68769, n68700 );
xor U120021 ( n68769, n75054, n68701 );
xnor U120022 ( n32565, n34013, n33944 );
xor U120023 ( n34013, n75055, n33945 );
xnor U120024 ( n25323, n26770, n26699 );
xor U120025 ( n26770, n75056, n26700 );
xnor U120026 ( n58462, n59910, n59841 );
xor U120027 ( n59910, n75057, n59842 );
xnor U120028 ( n46269, n47748, n47679 );
xor U120029 ( n47748, n75058, n47680 );
xnor U120030 ( n12642, n14484, n14407 );
xor U120031 ( n14484, n75059, n14408 );
nand U120032 ( n61703, n73069, n74385 );
nor U120033 ( n30785, n73987, n30461 );
nor U120034 ( n10277, n74005, n9869 );
nor U120035 ( n64987, n73643, n64620 );
nor U120036 ( n44145, n73553, n43777 );
nor U120037 ( n23464, n4234, n23494 );
nor U120038 ( n56586, n6867, n56616 );
nor U120039 ( n23476, n4233, n73516 );
nor U120040 ( n56598, n6865, n73517 );
nor U120041 ( n23473, n73683, n23133 );
nor U120042 ( n56595, n73682, n56254 );
nand U120043 ( n23458, n23471, n23472 );
nor U120044 ( n23471, n23477, n23478 );
nor U120045 ( n23472, n23473, n23474 );
nor U120046 ( n23477, n73669, n23129 );
nand U120047 ( n56580, n56593, n56594 );
nor U120048 ( n56593, n56599, n56600 );
nor U120049 ( n56594, n56595, n56596 );
nor U120050 ( n56599, n73668, n56250 );
nor U120051 ( n23478, n73641, n23130 );
nor U120052 ( n56600, n73642, n56251 );
nand U120053 ( n61695, n73056, n73528 );
nor U120054 ( n42258, n42256, n42261 );
nand U120055 ( n42261, n42251, n73911 );
nand U120056 ( n61702, n73095, n74434 );
nand U120057 ( n8294, n4813, n74685 );
nand U120058 ( n61696, n73045, n73498 );
not U120059 ( n7802, n44902 );
not U120060 ( n3399, n31517 );
not U120061 ( n4237, n24223 );
not U120062 ( n6014, n65767 );
not U120063 ( n6869, n57345 );
nand U120064 ( n61709, n73124, n74493 );
xor U120065 ( n45140, n74474, n847 );
not U120066 ( n847, n45270 );
nand U120067 ( n42540, n8164, n42543 );
nand U120068 ( n8464, n5510, n8468 );
nand U120069 ( n42382, n7457, n74686 );
nor U120070 ( n27127, n27213, n74423 );
nor U120071 ( n34371, n34458, n74426 );
nor U120072 ( n69123, n69208, n74425 );
nor U120073 ( n60271, n60358, n74424 );
nor U120074 ( n30727, n73959, n30464 );
nor U120075 ( n10208, n73986, n9873 );
nor U120076 ( n64933, n73596, n64623 );
nor U120077 ( n44090, n73545, n43780 );
nand U120078 ( n30717, n30725, n30726 );
nor U120079 ( n30725, n30729, n30730 );
nor U120080 ( n30726, n30727, n30728 );
nor U120081 ( n30729, n73952, n30460 );
nand U120082 ( n10195, n10205, n10207 );
nor U120083 ( n10205, n10210, n10212 );
nor U120084 ( n10207, n10208, n10209 );
nor U120085 ( n10210, n73979, n9868 );
nand U120086 ( n64923, n64931, n64932 );
nor U120087 ( n64931, n64935, n64936 );
nor U120088 ( n64932, n64933, n64934 );
nor U120089 ( n64935, n73585, n64619 );
nand U120090 ( n44080, n44088, n44089 );
nor U120091 ( n44088, n44092, n44093 );
nor U120092 ( n44089, n44090, n44091 );
nor U120093 ( n44092, n73537, n43776 );
not U120094 ( n498, n42384 );
nor U120095 ( n23417, n73620, n23133 );
nor U120096 ( n56539, n73619, n56254 );
nand U120097 ( n23407, n23415, n23416 );
nor U120098 ( n23415, n23419, n23420 );
nor U120099 ( n23416, n23417, n23418 );
nor U120100 ( n23419, n73601, n23129 );
nand U120101 ( n56529, n56537, n56538 );
nor U120102 ( n56537, n56541, n56542 );
nor U120103 ( n56538, n56539, n56540 );
nor U120104 ( n56541, n73600, n56250 );
nor U120105 ( n30730, n73949, n30461 );
nor U120106 ( n10212, n73964, n9869 );
nor U120107 ( n64936, n73564, n64620 );
nor U120108 ( n44093, n73534, n43777 );
not U120109 ( n882, n43559 );
nor U120110 ( n23420, n73569, n23130 );
nor U120111 ( n56542, n73568, n56251 );
not U120112 ( n2898, n38227 );
not U120113 ( n227, n8297 );
not U120114 ( n5147, n11194 );
nor U120115 ( n8314, n8319, n8320 );
xnor U120116 ( n12637, n14460, n14483 );
xor U120117 ( n14483, n75059, n11304 );
xnor U120118 ( n67326, n68750, n68768 );
xor U120119 ( n68768, n75054, n65893 );
xnor U120120 ( n46265, n47729, n47747 );
xor U120121 ( n47747, n75058, n44985 );
xnor U120122 ( n25319, n26749, n26769 );
xor U120123 ( n26769, n75056, n24311 );
xnor U120124 ( n58458, n59891, n59909 );
xor U120125 ( n59909, n75057, n57434 );
xnor U120126 ( n32561, n33994, n34012 );
xor U120127 ( n34012, n75055, n31607 );
nand U120128 ( n12658, n14460, n14587 );
nand U120129 ( n14587, n4978, n73079 );
nand U120130 ( n25329, n26749, n26851 );
nand U120131 ( n26851, n4069, n73075 );
nand U120132 ( n58468, n59891, n59991 );
nand U120133 ( n59991, n6702, n73074 );
nand U120134 ( n46275, n47729, n47830 );
nand U120135 ( n47830, n7632, n73071 );
nand U120136 ( n32571, n33994, n34096 );
nand U120137 ( n34096, n3244, n73077 );
nand U120138 ( n67336, n68750, n68850 );
nand U120139 ( n68850, n5844, n73076 );
not U120140 ( n887, n42957 );
nor U120141 ( n29189, n29193, n29194 );
nor U120142 ( n21872, n21876, n21877 );
nor U120143 ( n62907, n62911, n62912 );
nor U120144 ( n54963, n54967, n54968 );
nor U120145 ( n21214, n73527, n73060 );
nor U120146 ( n4936, n31619, n73436 );
nor U120147 ( n13916, n75427, n57446 );
nor U120148 ( n11671, n73429, n65905 );
nor U120149 ( n7181, n24323, n75428 );
nor U120150 ( n42398, n42402, n42403 );
nand U120151 ( n11630, n11632, n11633 );
nor U120152 ( n67989, n73104, n74431 );
nor U120153 ( n25986, n73105, n74432 );
nor U120154 ( n59124, n73106, n74433 );
nor U120155 ( n30792, n73526, n30771 );
nor U120156 ( n10285, n73527, n10259 );
nor U120157 ( n64994, n73515, n64973 );
nor U120158 ( n44152, n73511, n44131 );
nor U120159 ( n30790, n74018, n30452 );
nor U120160 ( n10283, n74061, n9858 );
nor U120161 ( n64992, n73702, n64611 );
nor U120162 ( n44150, n73574, n43768 );
nand U120163 ( n30787, n30788, n30789 );
nor U120164 ( n30788, n30793, n30794 );
nor U120165 ( n30789, n30790, n30791 );
nor U120166 ( n30793, n74014, n30448 );
nand U120167 ( n10279, n10280, n10282 );
nor U120168 ( n10280, n10287, n10288 );
nor U120169 ( n10282, n10283, n10284 );
nor U120170 ( n10287, n74059, n9853 );
nand U120171 ( n64989, n64990, n64991 );
nor U120172 ( n64990, n64995, n64996 );
nor U120173 ( n64991, n64992, n64993 );
nor U120174 ( n64995, n73695, n64607 );
nand U120175 ( n44147, n44148, n44149 );
nor U120176 ( n44148, n44153, n44154 );
nor U120177 ( n44149, n44150, n44151 );
nor U120178 ( n44153, n73571, n43764 );
nor U120179 ( n42901, n7932, n42902 );
nor U120180 ( n42902, n42903, n42904 );
nor U120181 ( n42903, n42905, n42906 );
nor U120182 ( n8879, n5277, n8880 );
nor U120183 ( n8880, n8882, n8883 );
nor U120184 ( n8882, n8884, n8885 );
nor U120185 ( n30794, n74007, n30449 );
nor U120186 ( n10288, n74037, n9854 );
nor U120187 ( n64996, n73675, n64608 );
nor U120188 ( n44154, n73561, n43765 );
nor U120189 ( n23485, n73516, n23464 );
nor U120190 ( n56607, n73517, n56586 );
nor U120191 ( n23483, n73704, n23121 );
nor U120192 ( n56605, n73703, n56242 );
nand U120193 ( n23480, n23481, n23482 );
nor U120194 ( n23481, n23486, n23487 );
nor U120195 ( n23482, n23483, n23484 );
nor U120196 ( n23486, n73697, n23117 );
nand U120197 ( n56602, n56603, n56604 );
nor U120198 ( n56603, n56608, n56609 );
nor U120199 ( n56604, n56605, n56606 );
nor U120200 ( n56608, n73696, n56238 );
nor U120201 ( n33234, n74460, n73160 );
not U120202 ( n1780, n47958 );
not U120203 ( n2897, n38243 );
nor U120204 ( n23487, n73680, n23118 );
nor U120205 ( n56609, n73679, n56239 );
and U120206 ( n27715, n27788, n27135 );
and U120207 ( n60866, n60936, n60279 );
and U120208 ( n34960, n35029, n34380 );
and U120209 ( n69700, n69767, n69132 );
nor U120210 ( n23484, n73691, n23122 );
nor U120211 ( n56606, n73690, n56243 );
nor U120212 ( n30791, n74011, n30453 );
nor U120213 ( n10284, n74045, n9859 );
nor U120214 ( n64993, n73687, n64612 );
nor U120215 ( n44151, n73567, n43769 );
and U120216 ( n27882, n27788, n27297 );
and U120217 ( n61029, n60936, n60440 );
and U120218 ( n35121, n35029, n34542 );
and U120219 ( n69857, n69767, n69290 );
nand U120220 ( n30443, n30772, n3395 );
nand U120221 ( n9847, n10260, n5143 );
nand U120222 ( n64602, n64974, n6010 );
nand U120223 ( n43759, n44132, n7798 );
nor U120224 ( n30796, n30797, n30798 );
nor U120225 ( n30797, n74010, n30442 );
nor U120226 ( n30798, n74002, n30443 );
nor U120227 ( n10290, n10292, n10293 );
nor U120228 ( n10292, n74043, n9845 );
nor U120229 ( n10293, n74019, n9847 );
nor U120230 ( n64998, n64999, n65000 );
nor U120231 ( n64999, n73686, n64601 );
nor U120232 ( n65000, n73659, n64602 );
nor U120233 ( n44156, n44157, n44158 );
nor U120234 ( n44157, n73565, n43758 );
nor U120235 ( n44158, n73556, n43759 );
nand U120236 ( n30442, n30773, n3395 );
nand U120237 ( n9845, n10262, n5143 );
nand U120238 ( n64601, n64975, n6010 );
nand U120239 ( n43758, n44133, n7798 );
nand U120240 ( n23112, n23465, n4233 );
nand U120241 ( n56233, n56587, n6865 );
nor U120242 ( n23489, n23490, n23491 );
nor U120243 ( n23490, n73689, n23111 );
nor U120244 ( n23491, n73661, n23112 );
nor U120245 ( n56611, n56612, n56613 );
nor U120246 ( n56612, n73688, n56232 );
nor U120247 ( n56613, n73660, n56233 );
nand U120248 ( n30439, n30776, n3395 );
nand U120249 ( n9842, n10265, n5143 );
nand U120250 ( n64598, n64978, n6010 );
nand U120251 ( n43755, n44136, n7798 );
nor U120252 ( n30795, n30799, n30800 );
nor U120253 ( n30799, n74006, n30438 );
nor U120254 ( n30800, n74000, n30439 );
nor U120255 ( n10289, n10294, n10295 );
nor U120256 ( n10294, n74035, n9840 );
nor U120257 ( n10295, n74016, n9842 );
nor U120258 ( n64997, n65001, n65002 );
nor U120259 ( n65001, n73674, n64597 );
nor U120260 ( n65002, n73652, n64598 );
nor U120261 ( n44155, n44159, n44160 );
nor U120262 ( n44159, n73560, n43754 );
nor U120263 ( n44160, n73554, n43755 );
nand U120264 ( n23111, n23466, n4233 );
nand U120265 ( n56232, n56588, n6865 );
nand U120266 ( n30438, n30777, n3395 );
nand U120267 ( n9840, n10267, n5143 );
nand U120268 ( n64597, n64979, n6010 );
nand U120269 ( n43754, n44137, n7798 );
nand U120270 ( n23108, n23469, n4233 );
nand U120271 ( n56229, n56591, n6865 );
nor U120272 ( n23488, n23492, n23493 );
nor U120273 ( n23492, n73678, n23107 );
nor U120274 ( n23493, n73654, n23108 );
nor U120275 ( n56610, n56614, n56615 );
nor U120276 ( n56614, n73677, n56228 );
nor U120277 ( n56615, n73653, n56229 );
nand U120278 ( n42245, n914, n42246 );
not U120279 ( n914, n42247 );
nand U120280 ( n23107, n23470, n4233 );
nand U120281 ( n56228, n56592, n6865 );
and U120282 ( n28040, n28111, n27135 );
and U120283 ( n61199, n61266, n60279 );
and U120284 ( n35277, n35346, n34380 );
and U120285 ( n70011, n70078, n69132 );
and U120286 ( n28203, n28111, n27297 );
and U120287 ( n61367, n61266, n60440 );
and U120288 ( n70166, n70078, n69290 );
and U120289 ( n35436, n35346, n34542 );
nand U120290 ( n27217, n3909, n26954 );
not U120291 ( n3909, n27124 );
nand U120292 ( n60362, n6542, n60094 );
not U120293 ( n6542, n60268 );
nand U120294 ( n34462, n3065, n34199 );
not U120295 ( n3065, n34369 );
nand U120296 ( n69212, n5667, n68953 );
not U120297 ( n5667, n69121 );
nor U120298 ( n34378, n3064, n34704 );
not U120299 ( n3064, n34462 );
nor U120300 ( n27134, n3908, n27459 );
not U120301 ( n3908, n27217 );
nor U120302 ( n69130, n5665, n69448 );
not U120303 ( n5665, n69212 );
nor U120304 ( n60278, n6540, n60608 );
not U120305 ( n6540, n60362 );
nand U120306 ( n26965, n3912, n74888 );
nand U120307 ( n68964, n5669, n74889 );
nand U120308 ( n34210, n3068, n74887 );
nand U120309 ( n60105, n6544, n74890 );
not U120310 ( n6165, n63514 );
not U120311 ( n3550, n29615 );
not U120312 ( n4388, n22294 );
not U120313 ( n7020, n55406 );
nor U120314 ( n30735, n73965, n30452 );
nor U120315 ( n10218, n73995, n9858 );
nor U120316 ( n64941, n73621, n64611 );
nor U120317 ( n44098, n73550, n43768 );
nand U120318 ( n30732, n30733, n30734 );
nor U120319 ( n30733, n30737, n30738 );
nor U120320 ( n30734, n30735, n30736 );
nor U120321 ( n30737, n73960, n30448 );
nand U120322 ( n64938, n64939, n64940 );
nor U120323 ( n64939, n64943, n64944 );
nor U120324 ( n64940, n64941, n64942 );
nor U120325 ( n64943, n73602, n64607 );
nand U120326 ( n44095, n44096, n44097 );
nor U120327 ( n44096, n44100, n44101 );
nor U120328 ( n44097, n44098, n44099 );
nor U120329 ( n44100, n73546, n43764 );
nand U120330 ( n10214, n10215, n10217 );
nor U120331 ( n10215, n10220, n10222 );
nor U120332 ( n10217, n10218, n10219 );
nor U120333 ( n10220, n73988, n9853 );
nor U120334 ( n30684, n74034, n30464 );
nor U120335 ( n10152, n74097, n9873 );
nor U120336 ( n64890, n73728, n64623 );
nor U120337 ( n44045, n73584, n43780 );
nand U120338 ( n10139, n10149, n10150 );
nor U120339 ( n10149, n10154, n10155 );
nor U120340 ( n10150, n10152, n10153 );
nor U120341 ( n10154, n74072, n9868 );
nand U120342 ( n30674, n30682, n30683 );
nor U120343 ( n30682, n30686, n30687 );
nor U120344 ( n30683, n30684, n30685 );
nor U120345 ( n30686, n74022, n30460 );
nand U120346 ( n64880, n64888, n64889 );
nor U120347 ( n64888, n64892, n64893 );
nor U120348 ( n64889, n64890, n64891 );
nor U120349 ( n64892, n73707, n64619 );
nand U120350 ( n44035, n44043, n44044 );
nor U120351 ( n44043, n44047, n44048 );
nor U120352 ( n44044, n44045, n44046 );
nor U120353 ( n44047, n73575, n43776 );
nor U120354 ( n23373, n73730, n23133 );
nor U120355 ( n56497, n73729, n56254 );
nand U120356 ( n23363, n23371, n23372 );
nor U120357 ( n23371, n23375, n23376 );
nor U120358 ( n23372, n23373, n23374 );
nor U120359 ( n23375, n73709, n23129 );
nand U120360 ( n56487, n56495, n56496 );
nor U120361 ( n56495, n56499, n56500 );
nor U120362 ( n56496, n56497, n56498 );
nor U120363 ( n56499, n73708, n56250 );
nor U120364 ( n23425, n73632, n23121 );
nor U120365 ( n56547, n73631, n56242 );
nand U120366 ( n23422, n23423, n23424 );
nor U120367 ( n23423, n23427, n23428 );
nor U120368 ( n23424, n23425, n23426 );
nor U120369 ( n23427, n73623, n23117 );
nand U120370 ( n56544, n56545, n56546 );
nor U120371 ( n56545, n56549, n56550 );
nor U120372 ( n56546, n56547, n56548 );
nor U120373 ( n56549, n73622, n56238 );
nor U120374 ( n30738, n73956, n30449 );
nor U120375 ( n10222, n73983, n9854 );
nor U120376 ( n64944, n73592, n64608 );
nor U120377 ( n44101, n73541, n43765 );
nor U120378 ( n30687, n74012, n30461 );
nor U120379 ( n10155, n74046, n9869 );
nor U120380 ( n64893, n73666, n64620 );
nor U120381 ( n44048, n73558, n43777 );
nor U120382 ( n23376, n73671, n23130 );
nor U120383 ( n56500, n73670, n56251 );
nor U120384 ( n23428, n73614, n23118 );
nor U120385 ( n56550, n73613, n56239 );
nand U120386 ( n66978, n67070, n67071 );
nor U120387 ( n67071, n74502, n73100 );
nor U120388 ( n67070, n74526, n67072 );
nand U120389 ( n67072, n67131, n67132 );
nor U120390 ( n67131, n74479, n73091 );
nand U120391 ( n32339, n32407, n32408 );
nor U120392 ( n32408, n74503, n73102 );
nor U120393 ( n32407, n74527, n32409 );
nand U120394 ( n32409, n32475, n32476 );
nor U120395 ( n32475, n74478, n73093 );
nand U120396 ( n25174, n25233, n25234 );
nor U120397 ( n25233, n74480, n73094 );
nand U120398 ( n25102, n25172, n25173 );
nor U120399 ( n25173, n74504, n73103 );
nor U120400 ( n25172, n74528, n25174 );
nand U120401 ( n58310, n58369, n58370 );
nor U120402 ( n58369, n74481, n73092 );
nand U120403 ( n58240, n58308, n58309 );
nor U120404 ( n58309, n74505, n73101 );
nor U120405 ( n58308, n74529, n58310 );
nand U120406 ( n66798, n66846, n6185 );
nor U120407 ( n66846, n66847, n74563 );
nand U120408 ( n66934, n66976, n66977 );
nor U120409 ( n66977, n73110, n74558 );
nor U120410 ( n66976, n74463, n66978 );
nand U120411 ( n32152, n32200, n3570 );
nor U120412 ( n32200, n32201, n74564 );
nand U120413 ( n32295, n32337, n32338 );
nor U120414 ( n32338, n73112, n74557 );
nor U120415 ( n32337, n74465, n32339 );
nand U120416 ( n24920, n24970, n4408 );
nor U120417 ( n24970, n24971, n74565 );
nand U120418 ( n25058, n25100, n25101 );
nor U120419 ( n25101, n73113, n74559 );
nor U120420 ( n25100, n74466, n25102 );
nand U120421 ( n58057, n58105, n7040 );
nor U120422 ( n58105, n58106, n74566 );
nand U120423 ( n58193, n58238, n58239 );
nor U120424 ( n58239, n73111, n74560 );
nor U120425 ( n58238, n74464, n58240 );
nand U120426 ( n66599, n66660, n6183 );
nor U120427 ( n66660, n74751, n66661 );
nand U120428 ( n66678, n66783, n6184 );
nor U120429 ( n66783, n66784, n74940 );
nand U120430 ( n31996, n32057, n3568 );
nor U120431 ( n32057, n74752, n32058 );
nand U120432 ( n32075, n32137, n3569 );
nor U120433 ( n32137, n32138, n74941 );
nand U120434 ( n24764, n24825, n4405 );
nor U120435 ( n24825, n74753, n24826 );
nand U120436 ( n24843, n24905, n4407 );
nor U120437 ( n24905, n24906, n74942 );
nand U120438 ( n57898, n57959, n7038 );
nor U120439 ( n57959, n74754, n57960 );
nand U120440 ( n24676, n24746, n4404 );
nor U120441 ( n24746, n75043, n24747 );
nand U120442 ( n57977, n58042, n7039 );
nor U120443 ( n58042, n58043, n74943 );
nand U120444 ( n31888, n31978, n3567 );
nor U120445 ( n31978, n75044, n31979 );
nand U120446 ( n66511, n66581, n6182 );
nor U120447 ( n66581, n75045, n66582 );
nand U120448 ( n57810, n57880, n7037 );
nor U120449 ( n57880, n75046, n57881 );
nor U120450 ( n67132, n74700, n73080 );
nor U120451 ( n32476, n74699, n73082 );
nor U120452 ( n25234, n74701, n73083 );
nor U120453 ( n58370, n74702, n73081 );
nand U120454 ( n24644, n24656, n4403 );
nor U120455 ( n24656, n74910, n24657 );
nand U120456 ( n57780, n57792, n7035 );
nor U120457 ( n57792, n74911, n57793 );
nand U120458 ( n31858, n31870, n3565 );
nor U120459 ( n31870, n74912, n31871 );
nand U120460 ( n66481, n66493, n6180 );
nor U120461 ( n66493, n74913, n66494 );
not U120462 ( n6185, n66870 );
not U120463 ( n3570, n32232 );
not U120464 ( n4408, n24994 );
not U120465 ( n7040, n58129 );
nor U120466 ( n70855, n72927, n8208 );
nor U120467 ( n62418, n74636, n8208 );
nor U120468 ( n62483, n62418, n8208 );
nor U120469 ( n70864, n70855, n8208 );
nand U120470 ( n10161, n70856, n70857 );
nor U120471 ( n70856, n70866, n70867 );
nor U120472 ( n70857, n70858, n70859 );
nor U120473 ( n70866, n72927, n70842 );
nand U120474 ( n12406, n62475, n62476 );
nor U120475 ( n62475, n62485, n62486 );
nor U120476 ( n62476, n62477, n62478 );
nor U120477 ( n62485, n74636, n62405 );
nor U120478 ( n30736, n73962, n30453 );
nor U120479 ( n10219, n73991, n9859 );
nor U120480 ( n64942, n73610, n64612 );
nor U120481 ( n44099, n73548, n43769 );
nor U120482 ( n30740, n30741, n30742 );
nor U120483 ( n30741, n73963, n30442 );
nor U120484 ( n30742, n73969, n30443 );
nor U120485 ( n10224, n10225, n10227 );
nor U120486 ( n10225, n73992, n9845 );
nor U120487 ( n10227, n73998, n9847 );
nor U120488 ( n64946, n64947, n64948 );
nor U120489 ( n64947, n73612, n64601 );
nor U120490 ( n64948, n73628, n64602 );
nor U120491 ( n44103, n44104, n44105 );
nor U120492 ( n44104, n73549, n43758 );
nor U120493 ( n44105, n73552, n43759 );
nor U120494 ( n23426, n73627, n23122 );
nor U120495 ( n56548, n73626, n56243 );
nor U120496 ( n23430, n23431, n23432 );
nor U120497 ( n23431, n73630, n23111 );
nor U120498 ( n23432, n73635, n23112 );
nor U120499 ( n56552, n56553, n56554 );
nor U120500 ( n56553, n73629, n56232 );
nor U120501 ( n56554, n73634, n56233 );
nor U120502 ( n30739, n30743, n30744 );
nor U120503 ( n30743, n73958, n30438 );
nor U120504 ( n30744, n73953, n30439 );
nor U120505 ( n10223, n10228, n10229 );
nor U120506 ( n10228, n73985, n9840 );
nor U120507 ( n10229, n73980, n9842 );
nor U120508 ( n64945, n64949, n64950 );
nor U120509 ( n64949, n73595, n64597 );
nor U120510 ( n64950, n73588, n64598 );
nor U120511 ( n44102, n44106, n44107 );
nor U120512 ( n44106, n73543, n43754 );
nor U120513 ( n44107, n73538, n43755 );
nor U120514 ( n23429, n23433, n23434 );
nor U120515 ( n23433, n73618, n23107 );
nor U120516 ( n23434, n73605, n23108 );
nor U120517 ( n56551, n56555, n56556 );
nor U120518 ( n56555, n73617, n56228 );
nor U120519 ( n56556, n73604, n56229 );
xor U120520 ( n37954, n74420, n37955 );
nand U120521 ( n12408, n12409, n843 );
nand U120522 ( n30475, n30771, n30772 );
nand U120523 ( n9887, n10259, n10260 );
nand U120524 ( n64634, n64973, n64974 );
nand U120525 ( n43791, n44131, n44132 );
nor U120526 ( n30770, n74009, n30475 );
nor U120527 ( n10258, n74039, n9887 );
nor U120528 ( n64972, n73681, n64634 );
nor U120529 ( n44130, n73563, n43791 );
nand U120530 ( n30766, n30767, n30768 );
nor U120531 ( n30767, n30774, n30775 );
nor U120532 ( n30768, n30769, n30770 );
nor U120533 ( n30774, n74013, n30470 );
nand U120534 ( n10253, n10254, n10255 );
nor U120535 ( n10254, n10263, n10264 );
nor U120536 ( n10255, n10257, n10258 );
nor U120537 ( n10263, n74052, n9880 );
nand U120538 ( n64968, n64969, n64970 );
nor U120539 ( n64969, n64976, n64977 );
nor U120540 ( n64970, n64971, n64972 );
nor U120541 ( n64976, n73692, n64629 );
nand U120542 ( n44126, n44127, n44128 );
nor U120543 ( n44127, n44134, n44135 );
nor U120544 ( n44128, n44129, n44130 );
nor U120545 ( n44134, n73570, n43786 );
nor U120546 ( n30781, n74001, n30465 );
nor U120547 ( n10272, n74017, n9874 );
nor U120548 ( n64983, n73655, n64624 );
nor U120549 ( n44141, n73555, n43781 );
nand U120550 ( n30474, n30771, n30773 );
nand U120551 ( n9885, n10259, n10262 );
nand U120552 ( n64633, n64973, n64975 );
nand U120553 ( n43790, n44131, n44133 );
nor U120554 ( n30769, n74015, n30474 );
nor U120555 ( n10257, n74060, n9885 );
nor U120556 ( n64971, n73698, n64633 );
nor U120557 ( n44129, n73572, n43790 );
nand U120558 ( n23144, n23464, n23465 );
nand U120559 ( n56265, n56586, n56587 );
nor U120560 ( n23463, n73685, n23144 );
nor U120561 ( n56585, n73684, n56265 );
nand U120562 ( n23459, n23460, n23461 );
nor U120563 ( n23460, n23467, n23468 );
nor U120564 ( n23461, n23462, n23463 );
nor U120565 ( n23467, n73694, n23139 );
nand U120566 ( n56581, n56582, n56583 );
nor U120567 ( n56582, n56589, n56590 );
nor U120568 ( n56583, n56584, n56585 );
nor U120569 ( n56589, n73693, n56260 );
nor U120570 ( n23474, n73658, n23134 );
nor U120571 ( n56596, n73657, n56255 );
nand U120572 ( n12401, n62487, n62488 );
nor U120573 ( n62487, n62496, n62497 );
nor U120574 ( n62488, n76235, n62489 );
nor U120575 ( n62496, n74636, n62502 );
nand U120576 ( n30471, n30771, n30776 );
nand U120577 ( n9882, n10259, n10265 );
nand U120578 ( n64630, n64973, n64978 );
nand U120579 ( n43787, n44131, n44136 );
nor U120580 ( n30775, n74004, n30471 );
nor U120581 ( n10264, n74031, n9882 );
nor U120582 ( n64977, n73667, n64630 );
nor U120583 ( n44135, n73559, n43787 );
nand U120584 ( n23143, n23464, n23466 );
nand U120585 ( n56264, n56586, n56588 );
nor U120586 ( n23462, n73700, n23143 );
nor U120587 ( n56584, n73699, n56264 );
nand U120588 ( n30470, n30771, n30777 );
nand U120589 ( n9880, n10259, n10267 );
nand U120590 ( n64629, n64973, n64979 );
nand U120591 ( n43786, n44131, n44137 );
nand U120592 ( n23140, n23464, n23469 );
nand U120593 ( n56261, n56586, n56591 );
nor U120594 ( n23468, n73673, n23140 );
nor U120595 ( n56590, n73672, n56261 );
nand U120596 ( n23139, n23464, n23470 );
nand U120597 ( n56260, n56586, n56592 );
nor U120598 ( n30638, n74126, n30464 );
nor U120599 ( n10087, n74154, n9873 );
nor U120600 ( n64844, n73773, n64623 );
nor U120601 ( n43997, n73648, n43780 );
nand U120602 ( n10074, n10084, n10085 );
nor U120603 ( n10084, n10089, n10090 );
nor U120604 ( n10085, n10087, n10088 );
nor U120605 ( n10089, n74149, n9868 );
nand U120606 ( n30628, n30636, n30637 );
nor U120607 ( n30636, n30640, n30641 );
nor U120608 ( n30637, n30638, n30639 );
nor U120609 ( n30640, n74121, n30460 );
nand U120610 ( n64834, n64842, n64843 );
nor U120611 ( n64842, n64846, n64847 );
nor U120612 ( n64843, n64844, n64845 );
nor U120613 ( n64846, n73761, n64619 );
nand U120614 ( n43987, n43995, n43996 );
nor U120615 ( n43995, n43999, n44000 );
nor U120616 ( n43996, n43997, n43998 );
nor U120617 ( n43999, n73644, n43776 );
nor U120618 ( n23324, n73774, n23133 );
nor U120619 ( n56448, n73775, n56254 );
nand U120620 ( n23314, n23322, n23323 );
nor U120621 ( n23322, n23326, n23327 );
nor U120622 ( n23323, n23324, n23325 );
nor U120623 ( n23326, n73763, n23129 );
nand U120624 ( n56438, n56446, n56447 );
nor U120625 ( n56446, n56450, n56451 );
nor U120626 ( n56447, n56448, n56449 );
nor U120627 ( n56450, n73764, n56250 );
nor U120628 ( n30641, n74063, n30461 );
nor U120629 ( n10090, n74128, n9869 );
nor U120630 ( n64847, n73749, n64620 );
nor U120631 ( n44000, n73636, n43777 );
nor U120632 ( n23327, n73750, n23130 );
nor U120633 ( n56451, n73751, n56251 );
and U120634 ( n27561, n27297, n27467 );
and U120635 ( n60711, n60440, n60616 );
and U120636 ( n34804, n34542, n34712 );
and U120637 ( n69548, n69290, n69456 );
nor U120638 ( n13507, n74468, n73117 );
nor U120639 ( n54709, n54710, n74684 );
nor U120640 ( n54710, n54711, n54712 );
nor U120641 ( n54711, n54717, n54718 );
nor U120642 ( n54712, n54713, n8208 );
nor U120643 ( n21670, n21671, n74713 );
nor U120644 ( n21671, n21672, n21673 );
nor U120645 ( n21672, n21678, n21679 );
nor U120646 ( n21673, n21674, n8208 );
nor U120647 ( n36154, n36155, n73192 );
nor U120648 ( n36155, n36156, n36157 );
nor U120649 ( n36156, n36162, n36163 );
nor U120650 ( n36157, n36158, n8208 );
nor U120651 ( n28981, n28982, n74691 );
nor U120652 ( n28982, n28983, n28984 );
nor U120653 ( n28983, n28989, n28990 );
nor U120654 ( n28984, n28985, n8208 );
nand U120655 ( n12362, n12453, n12454 );
nor U120656 ( n12454, n74506, n73097 );
nor U120657 ( n12453, n74541, n12455 );
nand U120658 ( n12455, n12529, n12530 );
nor U120659 ( n12529, n74484, n73087 );
nand U120660 ( n12125, n12185, n5319 );
nor U120661 ( n12185, n12187, n74512 );
nand U120662 ( n12307, n12359, n12360 );
nor U120663 ( n12360, n73107, n74577 );
nor U120664 ( n12359, n74450, n12362 );
nand U120665 ( n11838, n11910, n5315 );
nor U120666 ( n11910, n74808, n11912 );
nand U120667 ( n11938, n12002, n5317 );
nor U120668 ( n12002, n74997, n12003 );
nand U120669 ( n12024, n12102, n5318 );
nor U120670 ( n12102, n12103, n74956 );
nor U120671 ( n12530, n74718, n73072 );
nand U120672 ( n11797, n11812, n5314 );
nor U120673 ( n11812, n75170, n11813 );
not U120674 ( n5319, n12228 );
not U120675 ( n2895, n38259 );
nand U120676 ( n46038, n46106, n46107 );
nor U120677 ( n46107, n74500, n73098 );
nor U120678 ( n46106, n74522, n46108 );
nand U120679 ( n46108, n46167, n46168 );
nor U120680 ( n46167, n74473, n73089 );
nand U120681 ( n45847, n45895, n7974 );
nor U120682 ( n45895, n45896, n74515 );
nand U120683 ( n45983, n46036, n46037 );
nor U120684 ( n46037, n73108, n74554 );
nor U120685 ( n46036, n74451, n46038 );
nand U120686 ( n45586, n45657, n7970 );
nor U120687 ( n45657, n74810, n45658 );
nand U120688 ( n45675, n45734, n7972 );
nor U120689 ( n45734, n74998, n45735 );
nand U120690 ( n45770, n45832, n7973 );
nor U120691 ( n45832, n45833, n74957 );
nor U120692 ( n30722, n73957, n30475 );
nor U120693 ( n10202, n73984, n9887 );
nor U120694 ( n64928, n73594, n64634 );
nor U120695 ( n44085, n73542, n43791 );
nor U120696 ( n46168, n74717, n73073 );
nand U120697 ( n45556, n45568, n7969 );
nor U120698 ( n45568, n75077, n45569 );
nand U120699 ( n30718, n30719, n30720 );
nor U120700 ( n30719, n30723, n30724 );
nor U120701 ( n30720, n30721, n30722 );
nor U120702 ( n30723, n73955, n30470 );
nand U120703 ( n10197, n10198, n10199 );
nor U120704 ( n10198, n10203, n10204 );
nor U120705 ( n10199, n10200, n10202 );
nor U120706 ( n10203, n73982, n9880 );
nand U120707 ( n64924, n64925, n64926 );
nor U120708 ( n64925, n64929, n64930 );
nor U120709 ( n64926, n64927, n64928 );
nor U120710 ( n64929, n73590, n64629 );
nand U120711 ( n44081, n44082, n44083 );
nor U120712 ( n44082, n44086, n44087 );
nor U120713 ( n44083, n44084, n44085 );
nor U120714 ( n44086, n73540, n43786 );
not U120715 ( n7974, n45919 );
nor U120716 ( n30728, n73954, n30465 );
nor U120717 ( n10209, n73981, n9874 );
nor U120718 ( n64934, n73589, n64624 );
nor U120719 ( n44091, n73539, n43781 );
nor U120720 ( n30721, n73961, n30474 );
nor U120721 ( n10200, n73989, n9885 );
nor U120722 ( n64927, n73603, n64633 );
nor U120723 ( n44084, n73547, n43790 );
nand U120724 ( n62415, n62416, n62417 );
nand U120725 ( n62417, n62418, n73184 );
nand U120726 ( n62416, n76300, n75228 );
nand U120727 ( n12411, n62407, n62408 );
nor U120728 ( n62408, n62409, n62410 );
nor U120729 ( n62407, n62414, n62415 );
nor U120730 ( n62409, n61915, n54949 );
nor U120731 ( n56534, n73615, n56265 );
not U120732 ( n76300, n76301 );
nor U120733 ( n23412, n73616, n23144 );
nand U120734 ( n23408, n23409, n23410 );
nor U120735 ( n23409, n23413, n23414 );
nor U120736 ( n23410, n23411, n23412 );
nor U120737 ( n23413, n73609, n23139 );
nand U120738 ( n56530, n56531, n56532 );
nor U120739 ( n56531, n56535, n56536 );
nor U120740 ( n56532, n56533, n56534 );
nor U120741 ( n56535, n73608, n56260 );
not U120742 ( n76299, n76301 );
nor U120743 ( n23418, n73607, n23134 );
nor U120744 ( n56540, n73606, n56255 );
nor U120745 ( n23411, n73625, n23143 );
nor U120746 ( n56533, n73624, n56264 );
nor U120747 ( n30724, n73951, n30471 );
nor U120748 ( n10204, n73978, n9882 );
nor U120749 ( n64930, n73583, n64630 );
nor U120750 ( n44087, n73536, n43787 );
nand U120751 ( n62480, n76301, n74636 );
not U120752 ( n7900, n46818 );
nor U120753 ( n23414, n73598, n23140 );
nor U120754 ( n56536, n73597, n56261 );
nor U120755 ( n62486, n76299, n54949 );
not U120756 ( n76372, n76373 );
nand U120757 ( n14656, n54679, n54680 );
nor U120758 ( n54680, n54681, n54682 );
nor U120759 ( n54679, n54686, n54687 );
nor U120760 ( n54681, n54287, n42384 );
not U120761 ( n76371, n76373 );
nor U120762 ( n47917, n47919, n47920 );
nor U120763 ( n47919, n47921, n74442 );
nor U120764 ( n47909, n7413, n47913 );
nor U120765 ( n47913, n47914, n47915 );
nor U120766 ( n47915, n47916, n7415 );
nor U120767 ( n47914, n47917, n47918 );
nand U120768 ( n15521, n47906, n47907 );
nand U120769 ( n47907, n47908, n7394 );
nor U120770 ( n47906, n47909, n47910 );
not U120771 ( n7394, n47904 );
or U120772 ( n36123, n73192, n35789 );
not U120773 ( n76554, n76555 );
nand U120774 ( n5676, n28951, n28952 );
nor U120775 ( n28952, n28953, n28954 );
nor U120776 ( n28951, n28958, n28959 );
nor U120777 ( n28953, n28610, n21858 );
nand U120778 ( n28968, n76555, n74651 );
not U120779 ( n76553, n76555 );
nor U120780 ( n54703, n76371, n42384 );
nand U120781 ( n14651, n54691, n54692 );
nor U120782 ( n54692, n54693, n54694 );
nor U120783 ( n54691, n54702, n54703 );
nor U120784 ( n54693, n75253, n54701 );
nor U120785 ( n28975, n76553, n21858 );
nand U120786 ( n54696, n76373, n74650 );
nand U120787 ( n5671, n28963, n28964 );
nor U120788 ( n28964, n28965, n28966 );
nor U120789 ( n28963, n28974, n28975 );
nor U120790 ( n28965, n75254, n28973 );
not U120791 ( n76644, n76645 );
nand U120792 ( n7921, n21641, n21642 );
nor U120793 ( n21642, n21643, n21644 );
nor U120794 ( n21641, n21648, n21649 );
nor U120795 ( n21643, n21304, n8297 );
not U120796 ( n76643, n76645 );
nor U120797 ( n63554, n63555, n63556 );
nor U120798 ( n63555, n63557, n63558 );
nor U120799 ( n29655, n29656, n29657 );
nor U120800 ( n29656, n29658, n29659 );
nor U120801 ( n22334, n22335, n22336 );
nor U120802 ( n22335, n22337, n22338 );
nor U120803 ( n55446, n55447, n55448 );
nor U120804 ( n55447, n55449, n55450 );
xor U120805 ( n44391, n74428, n859 );
not U120806 ( n859, n44395 );
or U120807 ( n21640, n74713, n21304 );
or U120808 ( n54662, n74684, n54287 );
or U120809 ( n28950, n74691, n28610 );
nor U120810 ( n21664, n76643, n8297 );
nand U120811 ( n7916, n21653, n21654 );
nor U120812 ( n21654, n21655, n21656 );
nor U120813 ( n21653, n21663, n21664 );
nor U120814 ( n21655, n75255, n21662 );
nand U120815 ( n21658, n76645, n74670 );
nor U120816 ( n23384, n73721, n23118 );
nor U120817 ( n56508, n73720, n56239 );
nand U120818 ( n23378, n23379, n23380 );
nor U120819 ( n23380, n23381, n23382 );
nor U120820 ( n23379, n23383, n23384 );
nor U120821 ( n23381, n73745, n23121 );
nand U120822 ( n56502, n56503, n56504 );
nor U120823 ( n56504, n56505, n56506 );
nor U120824 ( n56503, n56507, n56508 );
nor U120825 ( n56505, n73744, n56242 );
nor U120826 ( n30695, n74030, n30449 );
nor U120827 ( n10165, n74088, n9854 );
nor U120828 ( n64901, n73719, n64608 );
nor U120829 ( n44056, n73580, n43765 );
nand U120830 ( n30689, n30690, n30691 );
nor U120831 ( n30691, n30692, n30693 );
nor U120832 ( n30690, n30694, n30695 );
nor U120833 ( n30693, n74042, n30453 );
nand U120834 ( n10158, n10159, n10160 );
nor U120835 ( n10160, n10162, n10163 );
nor U120836 ( n10159, n10164, n10165 );
nor U120837 ( n10163, n74100, n9859 );
nand U120838 ( n64895, n64896, n64897 );
nor U120839 ( n64897, n64898, n64899 );
nor U120840 ( n64896, n64900, n64901 );
nor U120841 ( n64899, n73737, n64612 );
nand U120842 ( n44050, n44051, n44052 );
nor U120843 ( n44052, n44053, n44054 );
nor U120844 ( n44051, n44055, n44056 );
nor U120845 ( n44054, n73591, n43769 );
buf U120846 ( n76478, n76479 );
nand U120847 ( n28966, n28967, n76508 );
nand U120848 ( n28967, n28969, n28970 );
nor U120849 ( n28969, n73179, n74691 );
nor U120850 ( n28970, n28971, n28972 );
or U120851 ( n70843, n73186, n70515 );
nand U120852 ( n54694, n54695, n76308 );
nand U120853 ( n54695, n54697, n54698 );
nor U120854 ( n54697, n73177, n74684 );
nor U120855 ( n54698, n54699, n54700 );
nor U120856 ( n23382, n73739, n23122 );
nor U120857 ( n56506, n73738, n56243 );
nor U120858 ( n30692, n74047, n30452 );
nor U120859 ( n10162, n74103, n9858 );
nor U120860 ( n64898, n73743, n64611 );
nor U120861 ( n44053, n73599, n43768 );
nor U120862 ( n30694, n74036, n30448 );
nor U120863 ( n10164, n74098, n9853 );
nor U120864 ( n64900, n73731, n64607 );
nor U120865 ( n44055, n73586, n43764 );
nor U120866 ( n23383, n73733, n23117 );
nor U120867 ( n56507, n73732, n56238 );
or U120868 ( n62406, n74683, n61915 );
nor U120869 ( n23386, n23387, n23388 );
nor U120870 ( n23387, n73742, n23111 );
nor U120871 ( n23388, n73748, n23112 );
nor U120872 ( n56510, n56511, n56512 );
nor U120873 ( n56511, n73741, n56232 );
nor U120874 ( n56512, n73747, n56233 );
nor U120875 ( n30697, n30698, n30699 );
nor U120876 ( n30698, n74044, n30442 );
nor U120877 ( n30699, n74048, n30443 );
nor U120878 ( n10168, n10169, n10170 );
nor U120879 ( n10169, n74101, n9845 );
nor U120880 ( n10170, n74111, n9847 );
nor U120881 ( n64903, n64904, n64905 );
nor U120882 ( n64904, n73740, n64601 );
nor U120883 ( n64905, n73746, n64602 );
nor U120884 ( n44058, n44059, n44060 );
nor U120885 ( n44059, n73593, n43758 );
nor U120886 ( n44060, n73611, n43759 );
nand U120887 ( n21656, n21657, n76567 );
nand U120888 ( n21657, n21647, n21659 );
nor U120889 ( n21659, n21660, n21661 );
nor U120890 ( n21661, n227, n21652 );
not U120891 ( n3794, n38139 );
nor U120892 ( n23385, n23389, n23390 );
nor U120893 ( n23389, n73727, n23107 );
nor U120894 ( n23390, n73713, n23108 );
nor U120895 ( n56509, n56513, n56514 );
nor U120896 ( n56513, n73726, n56228 );
nor U120897 ( n56514, n73712, n56229 );
nand U120898 ( n10156, n70868, n70869 );
nor U120899 ( n70868, n70877, n70878 );
nor U120900 ( n70869, n5582, n70870 );
nor U120901 ( n70877, n72927, n70886 );
nor U120902 ( n30696, n30700, n30701 );
nor U120903 ( n30700, n74033, n30438 );
nor U120904 ( n30701, n74023, n30439 );
nor U120905 ( n10167, n10172, n10173 );
nor U120906 ( n10172, n74093, n9840 );
nor U120907 ( n10173, n74082, n9842 );
nor U120908 ( n64902, n64906, n64907 );
nor U120909 ( n64906, n73725, n64597 );
nor U120910 ( n64907, n73710, n64598 );
nor U120911 ( n44057, n44061, n44062 );
nor U120912 ( n44061, n73582, n43754 );
nor U120913 ( n44062, n73576, n43755 );
not U120914 ( n1972, n37930 );
not U120915 ( n2894, n38275 );
nor U120916 ( n8919, n5278, n8884 );
nor U120917 ( n42933, n7933, n42905 );
nor U120918 ( n47932, n47933, n47918 );
xor U120919 ( n47933, n47934, n47935 );
nand U120920 ( n47927, n47928, n47929 );
nand U120921 ( n47929, n7857, n47930 );
nor U120922 ( n47928, n47931, n47932 );
nor U120923 ( n47931, n47926, n47936 );
not U120924 ( n1778, n48202 );
nand U120925 ( n62405, n74683, n73184 );
nand U120926 ( n70842, n73186, n74657 );
not U120927 ( n897, n42684 );
not U120928 ( n907, n42350 );
not U120929 ( n3910, n26954 );
nor U120930 ( n30646, n74142, n30452 );
nor U120931 ( n10097, n74164, n9858 );
nor U120932 ( n64852, n73794, n64611 );
nor U120933 ( n44005, n73664, n43768 );
nand U120934 ( n30643, n30644, n30645 );
nor U120935 ( n30644, n30648, n30649 );
nor U120936 ( n30645, n30646, n30647 );
nor U120937 ( n30648, n74136, n30448 );
nand U120938 ( n10093, n10094, n10095 );
nor U120939 ( n10094, n10099, n10100 );
nor U120940 ( n10095, n10097, n10098 );
nor U120941 ( n10099, n74162, n9853 );
nand U120942 ( n64849, n64850, n64851 );
nor U120943 ( n64850, n64854, n64855 );
nor U120944 ( n64851, n64852, n64853 );
nor U120945 ( n64854, n73788, n64607 );
nand U120946 ( n44002, n44003, n44004 );
nor U120947 ( n44003, n44007, n44008 );
nor U120948 ( n44004, n44005, n44006 );
nor U120949 ( n44007, n73662, n43764 );
nand U120950 ( n28949, n74691, n73179 );
nand U120951 ( n36122, n73192, n74654 );
nor U120952 ( n30595, n74230, n30464 );
nor U120953 ( n10038, n74248, n9873 );
nor U120954 ( n64754, n73855, n64623 );
nor U120955 ( n43954, n73813, n43780 );
nor U120956 ( n30649, n74125, n30449 );
nor U120957 ( n10100, n74153, n9854 );
nor U120958 ( n64855, n73768, n64608 );
nor U120959 ( n44008, n73647, n43765 );
nand U120960 ( n10028, n10036, n10037 );
nor U120961 ( n10036, n10040, n10041 );
nor U120962 ( n10037, n10038, n10039 );
nor U120963 ( n10040, n74244, n9868 );
nand U120964 ( n30585, n30593, n30594 );
nor U120965 ( n30593, n30597, n30598 );
nor U120966 ( n30594, n30595, n30596 );
nor U120967 ( n30597, n74226, n30460 );
nand U120968 ( n64744, n64752, n64753 );
nor U120969 ( n64752, n64756, n64757 );
nor U120970 ( n64753, n64754, n64755 );
nor U120971 ( n64756, n73843, n64619 );
nand U120972 ( n43944, n43952, n43953 );
nor U120973 ( n43952, n43956, n43957 );
nor U120974 ( n43953, n43954, n43955 );
nor U120975 ( n43956, n73809, n43776 );
nor U120976 ( n23332, n73795, n23121 );
nor U120977 ( n56456, n73796, n56242 );
nor U120978 ( n23335, n73771, n23118 );
nor U120979 ( n56459, n73772, n56239 );
nand U120980 ( n23329, n23330, n23331 );
nor U120981 ( n23330, n23334, n23335 );
nor U120982 ( n23331, n23332, n23333 );
nor U120983 ( n23334, n73789, n23117 );
nand U120984 ( n56453, n56454, n56455 );
nor U120985 ( n56454, n56458, n56459 );
nor U120986 ( n56455, n56456, n56457 );
nor U120987 ( n56458, n73790, n56238 );
xnor U120988 ( n43431, n74381, n880 );
nand U120989 ( n54661, n74684, n73177 );
nor U120990 ( n23274, n73856, n23133 );
nor U120991 ( n56398, n73857, n56254 );
nand U120992 ( n23264, n23272, n23273 );
nor U120993 ( n23272, n23276, n23277 );
nor U120994 ( n23273, n23274, n23275 );
nor U120995 ( n23276, n73845, n23129 );
nand U120996 ( n56388, n56396, n56397 );
nor U120997 ( n56396, n56400, n56401 );
nor U120998 ( n56397, n56398, n56399 );
nor U120999 ( n56400, n73846, n56250 );
nor U121000 ( n30598, n74221, n30461 );
nor U121001 ( n10041, n74232, n9869 );
nor U121002 ( n64757, n73830, n64620 );
nor U121003 ( n43957, n73805, n43777 );
xnor U121004 ( n43444, n74380, n880 );
not U121005 ( n6543, n60094 );
nor U121006 ( n23277, n73831, n23130 );
nor U121007 ( n56401, n73832, n56251 );
nor U121008 ( n30647, n74131, n30453 );
nor U121009 ( n10098, n74157, n9859 );
nor U121010 ( n64853, n73782, n64612 );
nor U121011 ( n23333, n73783, n23122 );
nor U121012 ( n44006, n73651, n43769 );
nor U121013 ( n56457, n73784, n56243 );
nor U121014 ( n70867, n76646, n62893 );
nor U121015 ( n36148, n76500, n29171 );
nand U121016 ( n3426, n36136, n36137 );
nor U121017 ( n36137, n36138, n36139 );
nor U121018 ( n36136, n36147, n36148 );
nor U121019 ( n36138, n75256, n36146 );
nor U121020 ( n30651, n30652, n30653 );
nor U121021 ( n30652, n74129, n30442 );
nor U121022 ( n30653, n74107, n30443 );
nor U121023 ( n10103, n10104, n10105 );
nor U121024 ( n10104, n74156, n9845 );
nor U121025 ( n10105, n74143, n9847 );
nor U121026 ( n64857, n64858, n64859 );
nor U121027 ( n64858, n73779, n64601 );
nor U121028 ( n64859, n73758, n64602 );
nor U121029 ( n44010, n44011, n44012 );
nor U121030 ( n44011, n73650, n43758 );
nor U121031 ( n44012, n73640, n43759 );
nor U121032 ( n23337, n23338, n23339 );
nor U121033 ( n23338, n73780, n23111 );
nor U121034 ( n23339, n73759, n23112 );
nor U121035 ( n56461, n56462, n56463 );
nor U121036 ( n56462, n73781, n56232 );
nor U121037 ( n56463, n73760, n56233 );
buf U121038 ( n76613, n76609 );
nand U121039 ( n21639, n74713, n73185 );
nor U121040 ( n30650, n30654, n30655 );
nor U121041 ( n30654, n74124, n30438 );
nor U121042 ( n30655, n74102, n30439 );
nor U121043 ( n10102, n10107, n10108 );
nor U121044 ( n10107, n74152, n9840 );
nor U121045 ( n10108, n74139, n9842 );
nor U121046 ( n64856, n64860, n64861 );
nor U121047 ( n64860, n73767, n64597 );
nor U121048 ( n64861, n73752, n64598 );
nor U121049 ( n44009, n44013, n44014 );
nor U121050 ( n44013, n73646, n43754 );
nor U121051 ( n44014, n73638, n43755 );
nor U121052 ( n36382, n76920, n75247 );
nor U121053 ( n36614, n76920, n72953 );
nor U121054 ( n37081, n76920, n72944 );
nor U121055 ( n36731, n76920, n72941 );
nor U121056 ( n36763, n76920, n72938 );
nor U121057 ( n36288, n76920, n72930 );
nor U121058 ( n36590, n76920, n74123 );
nor U121059 ( n36668, n76920, n72932 );
nor U121060 ( n36798, n76920, n72956 );
nor U121061 ( n36573, n76920, n72947 );
nor U121062 ( n36323, n76920, n72945 );
nor U121063 ( n36533, n76920, n72940 );
nor U121064 ( n36356, n76920, n72933 );
nor U121065 ( n36463, n76920, n72934 );
nor U121066 ( n36818, n76920, n74198 );
nor U121067 ( n23336, n23340, n23341 );
nor U121068 ( n23340, n73769, n23107 );
nor U121069 ( n23341, n73753, n23108 );
nor U121070 ( n56460, n56464, n56465 );
nor U121071 ( n56464, n73770, n56228 );
nor U121072 ( n56465, n73754, n56229 );
nor U121073 ( n30679, n74032, n30475 );
nor U121074 ( n10145, n74089, n9887 );
nor U121075 ( n64885, n73722, n64634 );
nor U121076 ( n44040, n73581, n43791 );
nand U121077 ( n30675, n30676, n30677 );
nor U121078 ( n30676, n30680, n30681 );
nor U121079 ( n30677, n30678, n30679 );
nor U121080 ( n30680, n74025, n30470 );
nand U121081 ( n10140, n10142, n10143 );
nor U121082 ( n10142, n10147, n10148 );
nor U121083 ( n10143, n10144, n10145 );
nor U121084 ( n10147, n74085, n9880 );
nand U121085 ( n64881, n64882, n64883 );
nor U121086 ( n64882, n64886, n64887 );
nor U121087 ( n64883, n64884, n64885 );
nor U121088 ( n64886, n73711, n64629 );
nand U121089 ( n44036, n44037, n44038 );
nor U121090 ( n44037, n44041, n44042 );
nor U121091 ( n44038, n44039, n44040 );
nor U121092 ( n44041, n73578, n43786 );
nor U121093 ( n23368, n73724, n23144 );
nor U121094 ( n56492, n73723, n56265 );
nand U121095 ( n23364, n23365, n23366 );
nor U121096 ( n23365, n23369, n23370 );
nor U121097 ( n23366, n23367, n23368 );
nor U121098 ( n23369, n73718, n23139 );
nand U121099 ( n56488, n56489, n56490 );
nor U121100 ( n56489, n56493, n56494 );
nor U121101 ( n56490, n56491, n56492 );
nor U121102 ( n56493, n73717, n56260 );
nor U121103 ( n30685, n74024, n30465 );
nor U121104 ( n10153, n74084, n9874 );
nor U121105 ( n64891, n73714, n64624 );
nor U121106 ( n44046, n73577, n43781 );
nor U121107 ( n23374, n73716, n23134 );
nor U121108 ( n56498, n73715, n56255 );
nand U121109 ( n70852, n70853, n70854 );
nand U121110 ( n70854, n70855, n74657 );
nand U121111 ( n70853, n76646, n75227 );
nand U121112 ( n10166, n70844, n70845 );
nor U121113 ( n70845, n70846, n70847 );
nor U121114 ( n70844, n70851, n70852 );
nor U121115 ( n70846, n70515, n62893 );
not U121116 ( n76646, n76647 );
nor U121117 ( n30678, n74040, n30474 );
nor U121118 ( n10144, n74099, n9885 );
nor U121119 ( n64884, n73734, n64633 );
nor U121120 ( n44039, n73587, n43790 );
nor U121121 ( n23367, n73736, n23143 );
nor U121122 ( n56491, n73735, n56264 );
nor U121123 ( n30681, n74021, n30471 );
nor U121124 ( n10148, n74071, n9882 );
nor U121125 ( n64887, n73701, n64630 );
nor U121126 ( n44042, n73573, n43787 );
nor U121127 ( n23370, n73706, n23140 );
nor U121128 ( n56494, n73705, n56261 );
nor U121129 ( n62477, n75228, n62484 );
or U121130 ( n62484, n74683, n62418 );
nor U121131 ( n70858, n75227, n70865 );
or U121132 ( n70865, n73186, n70855 );
nor U121133 ( n36650, n76920, n74062 );
nand U121134 ( n3431, n36124, n36125 );
nor U121135 ( n36125, n36126, n36127 );
nor U121136 ( n36124, n36131, n36132 );
nor U121137 ( n36126, n35789, n29171 );
not U121138 ( n76500, n76501 );
nor U121139 ( n30548, n74269, n30464 );
nor U121140 ( n9990, n74291, n9873 );
nor U121141 ( n64707, n73924, n64623 );
nor U121142 ( n43909, n73887, n43780 );
nand U121143 ( n30538, n30546, n30547 );
nor U121144 ( n30546, n30550, n30551 );
nor U121145 ( n30547, n30548, n30549 );
nor U121146 ( n30550, n74264, n30460 );
nand U121147 ( n9978, n9988, n9989 );
nor U121148 ( n9988, n9993, n9994 );
nor U121149 ( n9989, n9990, n9992 );
nor U121150 ( n9993, n74284, n9868 );
nand U121151 ( n64697, n64705, n64706 );
nor U121152 ( n64705, n64709, n64710 );
nor U121153 ( n64706, n64707, n64708 );
nor U121154 ( n64709, n73912, n64619 );
nand U121155 ( n43899, n43907, n43908 );
nor U121156 ( n43907, n43911, n43912 );
nor U121157 ( n43908, n43909, n43910 );
nor U121158 ( n43911, n73883, n43776 );
not U121159 ( n3497, n33109 );
nor U121160 ( n23228, n73925, n23133 );
nor U121161 ( n56349, n73926, n56254 );
nor U121162 ( n30551, n74258, n30461 );
nor U121163 ( n9994, n74280, n9869 );
nor U121164 ( n64710, n73898, n64620 );
nor U121165 ( n43912, n73867, n43777 );
nand U121166 ( n23218, n23226, n23227 );
nor U121167 ( n23226, n23230, n23231 );
nor U121168 ( n23227, n23228, n23229 );
nor U121169 ( n23230, n73914, n23129 );
nand U121170 ( n56339, n56347, n56348 );
nor U121171 ( n56347, n56351, n56352 );
nor U121172 ( n56348, n56349, n56350 );
nor U121173 ( n56351, n73915, n56250 );
nor U121174 ( n23231, n73899, n23130 );
nor U121175 ( n56352, n73900, n56251 );
nor U121176 ( n3446, n76497, n75105 );
nor U121177 ( n3451, n76497, n73361 );
nor U121178 ( n3456, n76497, n75153 );
nor U121179 ( n3461, n76497, n73371 );
nor U121180 ( n3466, n76497, n75111 );
nor U121181 ( n3471, n76497, n73341 );
nor U121182 ( n3476, n76497, n75147 );
and U121183 ( n42307, n42308, n42309 );
nor U121184 ( n3481, n76497, n73369 );
nor U121185 ( n3486, n76497, n75099 );
nor U121186 ( n3491, n76497, n73333 );
nor U121187 ( n3496, n76497, n75088 );
nor U121188 ( n3501, n76497, n73330 );
nor U121189 ( n3506, n76497, n75117 );
nor U121190 ( n3511, n76497, n73347 );
nor U121191 ( n3516, n76497, n75141 );
nor U121192 ( n3521, n76497, n73367 );
nor U121193 ( n3526, n76496, n75165 );
nor U121194 ( n3531, n76497, n73383 );
nor U121195 ( n3536, n76496, n75129 );
nor U121196 ( n3541, n76496, n73355 );
nor U121197 ( n3546, n76496, n75159 );
nor U121198 ( n3551, n76496, n73377 );
nor U121199 ( n3556, n76496, n75089 );
nor U121200 ( n3561, n76496, n73331 );
nor U121201 ( n3566, n76496, n75123 );
nor U121202 ( n3571, n76496, n73349 );
nor U121203 ( n3576, n76496, n75079 );
nor U121204 ( n3581, n76496, n73323 );
nor U121205 ( n3586, n76496, n73335 );
nor U121206 ( n3591, n76496, n75135 );
nor U121207 ( n66510, n66494, n66511 );
nor U121208 ( n31887, n31871, n31888 );
nor U121209 ( n24675, n24657, n24676 );
nor U121210 ( n57809, n57793, n57810 );
nor U121211 ( n45585, n45569, n45586 );
nor U121212 ( n7936, n76640, n75109 );
nor U121213 ( n7941, n76640, n73365 );
nor U121214 ( n7946, n76640, n75157 );
nor U121215 ( n7951, n76640, n73375 );
nor U121216 ( n7956, n76640, n75115 );
nor U121217 ( n7961, n76640, n73345 );
nor U121218 ( n7966, n76640, n75151 );
nor U121219 ( n14671, n76368, n75106 );
nor U121220 ( n14676, n76368, n73362 );
nor U121221 ( n14681, n76368, n75154 );
nor U121222 ( n14686, n76368, n73372 );
nor U121223 ( n14691, n76368, n75112 );
nor U121224 ( n14696, n76368, n73342 );
nor U121225 ( n14701, n76368, n75148 );
nor U121226 ( n5691, n76550, n75107 );
nor U121227 ( n5696, n76550, n73363 );
nor U121228 ( n5701, n76550, n75155 );
nor U121229 ( n5706, n76550, n73373 );
nor U121230 ( n5711, n76550, n75113 );
nor U121231 ( n5716, n76550, n73343 );
nor U121232 ( n5721, n76550, n75149 );
nor U121233 ( n7971, n76640, n72994 );
nor U121234 ( n7976, n76640, n75103 );
nor U121235 ( n7981, n76640, n72982 );
nor U121236 ( n7986, n76640, n75096 );
nor U121237 ( n7991, n76640, n72977 );
nor U121238 ( n7996, n76640, n75121 );
nor U121239 ( n8001, n76640, n72986 );
nor U121240 ( n8006, n76640, n75145 );
nor U121241 ( n8011, n76640, n72990 );
nor U121242 ( n8016, n76639, n75169 );
nor U121243 ( n8021, n76640, n72998 );
nor U121244 ( n8026, n76639, n75133 );
nor U121245 ( n8031, n76639, n73359 );
nor U121246 ( n8036, n76639, n75163 );
nor U121247 ( n8041, n76639, n73381 );
nor U121248 ( n8046, n76639, n75097 );
nor U121249 ( n8051, n76639, n72978 );
nor U121250 ( n8056, n76639, n75127 );
nor U121251 ( n8061, n76639, n73353 );
nor U121252 ( n8066, n76639, n75083 );
nor U121253 ( n8071, n76639, n73327 );
nor U121254 ( n8076, n76639, n73339 );
nor U121255 ( n8081, n76639, n75139 );
nor U121256 ( n14706, n76368, n72991 );
nor U121257 ( n14711, n76368, n75101 );
nor U121258 ( n14716, n76368, n72980 );
nor U121259 ( n14721, n76368, n75090 );
nor U121260 ( n14726, n76368, n72971 );
nor U121261 ( n14731, n76368, n75118 );
nor U121262 ( n14736, n76368, n72983 );
nor U121263 ( n14741, n76368, n75142 );
nor U121264 ( n14746, n76368, n72987 );
nor U121265 ( n14751, n76367, n75166 );
nor U121266 ( n14756, n76368, n72995 );
nor U121267 ( n14761, n76367, n75130 );
nor U121268 ( n14766, n76367, n73356 );
nor U121269 ( n14771, n76367, n75160 );
nor U121270 ( n14776, n76367, n73378 );
nor U121271 ( n14781, n76367, n75091 );
nor U121272 ( n14786, n76367, n72972 );
nor U121273 ( n14791, n76367, n75124 );
nor U121274 ( n14796, n76367, n73350 );
nor U121275 ( n14801, n76367, n75080 );
nor U121276 ( n14806, n76367, n73324 );
nor U121277 ( n14811, n76367, n73336 );
nor U121278 ( n14816, n76367, n75136 );
nor U121279 ( n5726, n76550, n72992 );
nor U121280 ( n5731, n76550, n75102 );
nor U121281 ( n5736, n76550, n72981 );
nor U121282 ( n5741, n76550, n75092 );
nor U121283 ( n5746, n76550, n72973 );
nor U121284 ( n5751, n76550, n75119 );
nor U121285 ( n5756, n76550, n72984 );
nor U121286 ( n5761, n76550, n75143 );
nor U121287 ( n5766, n76550, n72988 );
nor U121288 ( n5771, n76549, n75167 );
nor U121289 ( n5776, n76550, n72996 );
nor U121290 ( n5781, n76549, n75131 );
nor U121291 ( n5786, n76549, n73357 );
nor U121292 ( n5791, n76549, n75161 );
nor U121293 ( n5796, n76549, n73379 );
nor U121294 ( n5801, n76549, n75093 );
nor U121295 ( n5806, n76549, n72974 );
nor U121296 ( n5811, n76549, n75125 );
nor U121297 ( n5816, n76549, n73351 );
nor U121298 ( n5821, n76549, n75081 );
nor U121299 ( n5826, n76549, n73325 );
nor U121300 ( n5831, n76549, n73337 );
nor U121301 ( n5836, n76549, n75137 );
nor U121302 ( n30633, n74127, n30475 );
nor U121303 ( n10080, n74155, n9887 );
nor U121304 ( n64839, n73776, n64634 );
nor U121305 ( n43992, n73649, n43791 );
nand U121306 ( n30629, n30630, n30631 );
nor U121307 ( n30630, n30634, n30635 );
nor U121308 ( n30631, n30632, n30633 );
nor U121309 ( n30634, n74134, n30470 );
nand U121310 ( n10075, n10077, n10078 );
nor U121311 ( n10077, n10082, n10083 );
nor U121312 ( n10078, n10079, n10080 );
nor U121313 ( n10082, n74161, n9880 );
nand U121314 ( n64835, n64836, n64837 );
nor U121315 ( n64836, n64840, n64841 );
nor U121316 ( n64837, n64838, n64839 );
nor U121317 ( n64840, n73785, n64629 );
nand U121318 ( n43988, n43989, n43990 );
nor U121319 ( n43989, n43993, n43994 );
nor U121320 ( n43990, n43991, n43992 );
nor U121321 ( n43993, n73656, n43786 );
nor U121322 ( n30639, n74104, n30465 );
nor U121323 ( n10088, n74140, n9874 );
nor U121324 ( n64845, n73755, n64624 );
nor U121325 ( n43998, n73639, n43781 );
nor U121326 ( n30632, n74137, n30474 );
nor U121327 ( n10079, n74163, n9885 );
nor U121328 ( n64838, n73791, n64633 );
nor U121329 ( n43991, n73663, n43790 );
nor U121330 ( n23319, n73777, n23144 );
nor U121331 ( n56443, n73778, n56265 );
nand U121332 ( n23315, n23316, n23317 );
nor U121333 ( n23316, n23320, n23321 );
nor U121334 ( n23317, n23318, n23319 );
nor U121335 ( n23320, n73786, n23139 );
nand U121336 ( n56439, n56440, n56441 );
nor U121337 ( n56440, n56444, n56445 );
nor U121338 ( n56441, n56442, n56443 );
nor U121339 ( n56444, n73787, n56260 );
nor U121340 ( n23325, n73756, n23134 );
nor U121341 ( n56449, n73757, n56255 );
nor U121342 ( n23318, n73792, n23143 );
nor U121343 ( n56442, n73793, n56264 );
not U121344 ( n6112, n67865 );
not U121345 ( n4334, n25862 );
not U121346 ( n6967, n59000 );
nor U121347 ( n30635, n74122, n30471 );
nor U121348 ( n10083, n74150, n9882 );
nor U121349 ( n64841, n73762, n64630 );
nor U121350 ( n43994, n73645, n43787 );
nor U121351 ( n23321, n73765, n23140 );
nor U121352 ( n56445, n73766, n56261 );
nor U121353 ( n8955, n8958, n8959 );
nor U121354 ( n42976, n42978, n42979 );
nor U121355 ( n10181, n76230, n75104 );
nor U121356 ( n10186, n76230, n73360 );
nor U121357 ( n10191, n76230, n75152 );
nor U121358 ( n10196, n76230, n73370 );
nor U121359 ( n10201, n76230, n75110 );
nor U121360 ( n10206, n76230, n73340 );
nor U121361 ( n10211, n76230, n75146 );
nor U121362 ( n10216, n76230, n73368 );
nor U121363 ( n10221, n76230, n75098 );
nor U121364 ( n10226, n76230, n73332 );
nor U121365 ( n10231, n76230, n75086 );
nor U121366 ( n10236, n76230, n73328 );
nor U121367 ( n10241, n76230, n75116 );
nor U121368 ( n10246, n76230, n73346 );
nor U121369 ( n10251, n76230, n75140 );
nor U121370 ( n10256, n76230, n73366 );
nor U121371 ( n10261, n76229, n75164 );
nor U121372 ( n10266, n76230, n73382 );
nor U121373 ( n10271, n76229, n75128 );
nor U121374 ( n10276, n76229, n73354 );
nor U121375 ( n10281, n76229, n75158 );
nor U121376 ( n10286, n76229, n73376 );
nor U121377 ( n10291, n76229, n75087 );
nor U121378 ( n10296, n76229, n73329 );
nor U121379 ( n10301, n76229, n75122 );
nor U121380 ( n10306, n76229, n73348 );
nor U121381 ( n10311, n76229, n75078 );
nor U121382 ( n10316, n76229, n73322 );
nor U121383 ( n10321, n76229, n73334 );
nor U121384 ( n10326, n76229, n75134 );
nand U121385 ( n60096, P2_P2_STATE2_REG_3_, n74517 );
nand U121386 ( n26956, P1_P2_STATE2_REG_3_, n74516 );
nand U121387 ( n34201, P1_P3_STATE2_REG_3_, n74513 );
nand U121388 ( n68955, P2_P3_STATE2_REG_3_, n74514 );
nor U121389 ( n60088, n60091, n60092 );
nor U121390 ( n60092, n60093, n60094 );
nor U121391 ( n60091, n60086, n60096 );
xor U121392 ( n60093, n60095, n6919 );
nor U121393 ( n26948, n26951, n26952 );
nor U121394 ( n26952, n26953, n26954 );
nor U121395 ( n26951, n26946, n26956 );
xor U121396 ( n26953, n26955, n4287 );
nor U121397 ( n34193, n34196, n34197 );
nor U121398 ( n34197, n34198, n34199 );
nor U121399 ( n34196, n34191, n34201 );
xor U121400 ( n34198, n34200, n3449 );
nor U121401 ( n68947, n68950, n68951 );
nor U121402 ( n68951, n68952, n68953 );
nor U121403 ( n68950, n68945, n68955 );
xor U121404 ( n68952, n68954, n6064 );
nor U121405 ( n12426, n76296, n75108 );
nor U121406 ( n12431, n76296, n73364 );
nor U121407 ( n12436, n76296, n75156 );
nor U121408 ( n12441, n76296, n73374 );
nor U121409 ( n12446, n76296, n75114 );
nor U121410 ( n12451, n76296, n73344 );
nor U121411 ( n12456, n76296, n75150 );
not U121412 ( n1930, n37816 );
not U121413 ( n1950, n37872 );
nor U121414 ( n31151, n74011, n30832 );
nor U121415 ( n44530, n73567, n44192 );
nor U121416 ( n65405, n73687, n65034 );
nand U121417 ( n31147, n31148, n31149 );
nor U121418 ( n31148, n31153, n31154 );
nor U121419 ( n31149, n31150, n31151 );
nor U121420 ( n31153, n74014, n30837 );
nand U121421 ( n44526, n44527, n44528 );
nor U121422 ( n44527, n44532, n44533 );
nor U121423 ( n44528, n44529, n44530 );
nor U121424 ( n44532, n73571, n44197 );
nand U121425 ( n65401, n65402, n65403 );
nor U121426 ( n65402, n65407, n65408 );
nor U121427 ( n65403, n65404, n65405 );
nor U121428 ( n65407, n73695, n65039 );
not U121429 ( n5247, n13350 );
not U121430 ( n3067, n34199 );
not U121431 ( n5668, n68953 );
nor U121432 ( n12461, n76296, n72993 );
nor U121433 ( n12466, n76296, n75100 );
nor U121434 ( n12471, n76296, n72979 );
nor U121435 ( n12476, n76296, n75094 );
nor U121436 ( n12481, n76296, n72975 );
nor U121437 ( n12486, n76296, n75120 );
nor U121438 ( n12491, n76296, n72985 );
nor U121439 ( n12496, n76296, n75144 );
nor U121440 ( n12501, n76296, n72989 );
nor U121441 ( n12506, n76295, n75168 );
nor U121442 ( n12511, n76296, n72997 );
nor U121443 ( n12516, n76295, n75132 );
nor U121444 ( n12521, n76295, n73358 );
nor U121445 ( n12526, n76295, n75162 );
nor U121446 ( n12531, n76295, n73380 );
nor U121447 ( n12536, n76295, n75095 );
nor U121448 ( n12541, n76295, n72976 );
nor U121449 ( n12546, n76295, n75126 );
nor U121450 ( n12551, n76295, n73352 );
nor U121451 ( n12556, n76295, n75082 );
nor U121452 ( n12561, n76295, n73326 );
nor U121453 ( n12566, n76295, n73338 );
nor U121454 ( n12571, n76295, n75138 );
nor U121455 ( n23285, n73853, n23118 );
nor U121456 ( n56409, n73854, n56239 );
nand U121457 ( n23279, n23280, n23281 );
nor U121458 ( n23281, n23282, n23283 );
nor U121459 ( n23280, n23284, n23285 );
nor U121460 ( n23282, n73878, n23121 );
nand U121461 ( n56403, n56404, n56405 );
nor U121462 ( n56405, n56406, n56407 );
nor U121463 ( n56404, n56408, n56409 );
nor U121464 ( n56406, n73879, n56242 );
nor U121465 ( n30606, n74229, n30449 );
nor U121466 ( n10049, n74247, n9854 );
nor U121467 ( n64765, n73850, n64608 );
nor U121468 ( n43965, n73812, n43765 );
nand U121469 ( n30600, n30601, n30602 );
nor U121470 ( n30602, n30603, n30604 );
nor U121471 ( n30601, n30605, n30606 );
nor U121472 ( n30603, n74242, n30452 );
nand U121473 ( n10043, n10044, n10045 );
nor U121474 ( n10045, n10046, n10047 );
nor U121475 ( n10044, n10048, n10049 );
nor U121476 ( n10046, n74255, n9858 );
nand U121477 ( n64759, n64760, n64761 );
nor U121478 ( n64761, n64762, n64763 );
nor U121479 ( n64760, n64764, n64765 );
nor U121480 ( n64762, n73877, n64611 );
nand U121481 ( n43959, n43960, n43961 );
nor U121482 ( n43961, n43962, n43963 );
nor U121483 ( n43960, n43964, n43965 );
nor U121484 ( n43962, n73820, n43768 );
not U121485 ( n5294, n8957 );
not U121486 ( n7949, n42977 );
nor U121487 ( n31154, n74007, n30836 );
nor U121488 ( n44533, n73561, n44196 );
nor U121489 ( n65408, n73675, n65038 );
nor U121490 ( n23283, n73865, n23122 );
nor U121491 ( n56407, n73866, n56243 );
nor U121492 ( n30604, n74235, n30453 );
nor U121493 ( n10047, n74251, n9859 );
nor U121494 ( n64763, n73864, n64612 );
nor U121495 ( n43963, n73816, n43769 );
nor U121496 ( n31094, n73962, n30832 );
nor U121497 ( n30882, n74312, n30832 );
nor U121498 ( n30924, n74272, n30832 );
nor U121499 ( n30967, n74235, n30832 );
nor U121500 ( n10559, n74157, n10335 );
nor U121501 ( n10614, n74100, n10335 );
nor U121502 ( n10453, n74294, n10335 );
nor U121503 ( n10398, n74331, n10335 );
nor U121504 ( n44371, n73651, n44192 );
nor U121505 ( n44429, n73591, n44192 );
nor U121506 ( n44242, n73977, n44192 );
nor U121507 ( n44286, n73890, n44192 );
nor U121508 ( n44471, n73548, n44192 );
nor U121509 ( n10667, n73991, n10335 );
nor U121510 ( n65084, n74094, n65034 );
nor U121511 ( n65126, n73933, n65034 );
nor U121512 ( n65169, n73864, n65034 );
nor U121513 ( n65211, n73782, n65034 );
nor U121514 ( n65254, n73737, n65034 );
nor U121515 ( n31009, n74131, n30832 );
nor U121516 ( n31052, n74042, n30832 );
nor U121517 ( n65296, n73610, n65034 );
nand U121518 ( n31090, n31091, n31092 );
nor U121519 ( n31091, n31095, n31096 );
nor U121520 ( n31092, n31093, n31094 );
nor U121521 ( n31095, n73960, n30837 );
nand U121522 ( n30878, n30879, n30880 );
nor U121523 ( n30879, n30883, n30884 );
nor U121524 ( n30880, n30881, n30882 );
nor U121525 ( n30883, n74315, n30837 );
nand U121526 ( n30920, n30921, n30922 );
nor U121527 ( n30921, n30925, n30926 );
nor U121528 ( n30922, n30923, n30924 );
nor U121529 ( n30925, n74276, n30837 );
nand U121530 ( n30963, n30964, n30965 );
nor U121531 ( n30964, n30968, n30969 );
nor U121532 ( n30965, n30966, n30967 );
nor U121533 ( n30968, n74238, n30837 );
nand U121534 ( n10554, n10555, n10557 );
nor U121535 ( n10555, n10560, n10562 );
nor U121536 ( n10557, n10558, n10559 );
nor U121537 ( n10560, n74162, n10342 );
nand U121538 ( n10609, n10610, n10612 );
nor U121539 ( n10610, n10615, n10617 );
nor U121540 ( n10612, n10613, n10614 );
nor U121541 ( n10615, n74098, n10342 );
nand U121542 ( n10448, n10449, n10450 );
nor U121543 ( n10449, n10454, n10455 );
nor U121544 ( n10450, n10452, n10453 );
nor U121545 ( n10454, n74292, n10342 );
nand U121546 ( n10393, n10394, n10395 );
nor U121547 ( n10394, n10399, n10400 );
nor U121548 ( n10395, n10397, n10398 );
nor U121549 ( n10399, n74329, n10342 );
nand U121550 ( n44367, n44368, n44369 );
nor U121551 ( n44368, n44372, n44373 );
nor U121552 ( n44369, n44370, n44371 );
nor U121553 ( n44372, n73662, n44197 );
nand U121554 ( n44425, n44426, n44427 );
nor U121555 ( n44426, n44430, n44431 );
nor U121556 ( n44427, n44428, n44429 );
nor U121557 ( n44430, n73586, n44197 );
nand U121558 ( n44238, n44239, n44240 );
nor U121559 ( n44239, n44243, n44244 );
nor U121560 ( n44240, n44241, n44242 );
nor U121561 ( n44243, n73993, n44197 );
nand U121562 ( n44282, n44283, n44284 );
nor U121563 ( n44283, n44287, n44288 );
nor U121564 ( n44284, n44285, n44286 );
nor U121565 ( n44287, n73892, n44197 );
nand U121566 ( n44467, n44468, n44469 );
nor U121567 ( n44468, n44472, n44473 );
nor U121568 ( n44469, n44470, n44471 );
nor U121569 ( n44472, n73546, n44197 );
nand U121570 ( n10662, n10663, n10664 );
nor U121571 ( n10663, n10668, n10669 );
nor U121572 ( n10664, n10665, n10667 );
nor U121573 ( n10668, n73988, n10342 );
nand U121574 ( n65080, n65081, n65082 );
nor U121575 ( n65081, n65085, n65086 );
nor U121576 ( n65082, n65083, n65084 );
nor U121577 ( n65085, n74112, n65039 );
nand U121578 ( n65122, n65123, n65124 );
nor U121579 ( n65123, n65127, n65128 );
nor U121580 ( n65124, n65125, n65126 );
nor U121581 ( n65127, n73939, n65039 );
nand U121582 ( n65165, n65166, n65167 );
nor U121583 ( n65166, n65170, n65171 );
nor U121584 ( n65167, n65168, n65169 );
nor U121585 ( n65170, n73871, n65039 );
nand U121586 ( n65207, n65208, n65209 );
nor U121587 ( n65208, n65212, n65213 );
nor U121588 ( n65209, n65210, n65211 );
nor U121589 ( n65212, n73788, n65039 );
nand U121590 ( n65250, n65251, n65252 );
nor U121591 ( n65251, n65255, n65256 );
nor U121592 ( n65252, n65253, n65254 );
nor U121593 ( n65255, n73731, n65039 );
nand U121594 ( n31005, n31006, n31007 );
nor U121595 ( n31006, n31010, n31011 );
nor U121596 ( n31007, n31008, n31009 );
nor U121597 ( n31010, n74136, n30837 );
nand U121598 ( n31048, n31049, n31050 );
nor U121599 ( n31049, n31053, n31054 );
nor U121600 ( n31050, n31051, n31052 );
nor U121601 ( n31053, n74036, n30837 );
nand U121602 ( n65292, n65293, n65294 );
nor U121603 ( n65293, n65297, n65298 );
nor U121604 ( n65294, n65295, n65296 );
nor U121605 ( n65297, n73602, n65039 );
not U121606 ( n1777, n48331 );
nand U121607 ( n42300, n42302, n42303 );
not U121608 ( n2893, n38294 );
nor U121609 ( n31093, n73965, n30833 );
nor U121610 ( n30881, n74317, n30833 );
nor U121611 ( n30923, n74278, n30833 );
nor U121612 ( n30966, n74242, n30833 );
nor U121613 ( n10558, n74164, n10337 );
nor U121614 ( n10613, n74103, n10337 );
nor U121615 ( n10452, n74296, n10337 );
nor U121616 ( n10397, n74334, n10337 );
nor U121617 ( n44370, n73664, n44193 );
nor U121618 ( n44428, n73599, n44193 );
nor U121619 ( n44241, n73996, n44193 );
nor U121620 ( n44285, n73894, n44193 );
nor U121621 ( n44470, n73550, n44193 );
nor U121622 ( n10665, n73995, n10337 );
nor U121623 ( n65083, n74118, n65035 );
nor U121624 ( n65125, n73945, n65035 );
nor U121625 ( n65168, n73877, n65035 );
nor U121626 ( n65210, n73794, n65035 );
nor U121627 ( n65253, n73743, n65035 );
nor U121628 ( n31008, n74142, n30833 );
nor U121629 ( n31051, n74047, n30833 );
nor U121630 ( n65295, n73621, n65035 );
nor U121631 ( n10740, n74045, n10335 );
nand U121632 ( n10735, n10737, n10738 );
nor U121633 ( n10737, n10743, n10744 );
nor U121634 ( n10738, n10739, n10740 );
nor U121635 ( n10743, n74059, n10342 );
nor U121636 ( n10509, n74251, n10335 );
nor U121637 ( n44331, n73816, n44192 );
nand U121638 ( n10504, n10505, n10507 );
nor U121639 ( n10505, n10510, n10512 );
nor U121640 ( n10507, n10508, n10509 );
nor U121641 ( n10510, n74253, n10342 );
nand U121642 ( n44327, n44328, n44329 );
nor U121643 ( n44328, n44332, n44333 );
nor U121644 ( n44329, n44330, n44331 );
nor U121645 ( n44332, n73818, n44197 );
nor U121646 ( n31150, n74018, n30833 );
nor U121647 ( n44529, n73574, n44193 );
nor U121648 ( n10739, n74061, n10337 );
nor U121649 ( n65404, n73702, n65035 );
nor U121650 ( n31096, n73956, n30836 );
nor U121651 ( n30884, n74308, n30836 );
nor U121652 ( n30926, n74268, n30836 );
nor U121653 ( n30969, n74229, n30836 );
nor U121654 ( n10562, n74153, n10340 );
nor U121655 ( n10617, n74088, n10340 );
nor U121656 ( n10455, n74288, n10340 );
nor U121657 ( n10400, n74325, n10340 );
nor U121658 ( n44373, n73647, n44196 );
nor U121659 ( n44431, n73580, n44196 );
nor U121660 ( n44244, n73973, n44196 );
nor U121661 ( n44288, n73886, n44196 );
nor U121662 ( n44473, n73541, n44196 );
nor U121663 ( n10669, n73983, n10340 );
nor U121664 ( n65086, n74074, n65038 );
nor U121665 ( n65128, n73919, n65038 );
nor U121666 ( n65171, n73850, n65038 );
nor U121667 ( n65213, n73768, n65038 );
nor U121668 ( n65256, n73719, n65038 );
nor U121669 ( n31011, n74125, n30836 );
nor U121670 ( n31054, n74030, n30836 );
nor U121671 ( n65298, n73592, n65038 );
nor U121672 ( n23666, n73865, n23525 );
nor U121673 ( n23710, n73783, n23525 );
nor U121674 ( n23755, n73739, n23525 );
nor U121675 ( n23621, n73934, n23525 );
nor U121676 ( n23577, n74096, n23525 );
nor U121677 ( n56743, n73935, n56647 );
nor U121678 ( n56788, n73866, n56647 );
nor U121679 ( n56699, n74095, n56647 );
nor U121680 ( n56832, n73784, n56647 );
nor U121681 ( n56877, n73738, n56647 );
nor U121682 ( n23799, n73627, n23525 );
nor U121683 ( n56924, n73626, n56647 );
nand U121684 ( n23662, n23663, n23664 );
nor U121685 ( n23663, n23667, n23668 );
nor U121686 ( n23664, n23665, n23666 );
nor U121687 ( n23667, n73872, n23530 );
nand U121688 ( n23706, n23707, n23708 );
nor U121689 ( n23707, n23711, n23712 );
nor U121690 ( n23708, n23709, n23710 );
nor U121691 ( n23711, n73789, n23530 );
nand U121692 ( n23751, n23752, n23753 );
nor U121693 ( n23752, n23756, n23757 );
nor U121694 ( n23753, n23754, n23755 );
nor U121695 ( n23756, n73733, n23530 );
nand U121696 ( n23617, n23618, n23619 );
nor U121697 ( n23618, n23622, n23623 );
nor U121698 ( n23619, n23620, n23621 );
nor U121699 ( n23622, n73940, n23530 );
nand U121700 ( n23573, n23574, n23575 );
nor U121701 ( n23574, n23578, n23579 );
nor U121702 ( n23575, n23576, n23577 );
nor U121703 ( n23578, n74114, n23530 );
nand U121704 ( n56739, n56740, n56741 );
nor U121705 ( n56740, n56744, n56745 );
nor U121706 ( n56741, n56742, n56743 );
nor U121707 ( n56744, n73941, n56652 );
nand U121708 ( n56784, n56785, n56786 );
nor U121709 ( n56785, n56789, n56790 );
nor U121710 ( n56786, n56787, n56788 );
nor U121711 ( n56789, n73873, n56652 );
nand U121712 ( n56695, n56696, n56697 );
nor U121713 ( n56696, n56700, n56701 );
nor U121714 ( n56697, n56698, n56699 );
nor U121715 ( n56700, n74113, n56652 );
nand U121716 ( n56828, n56829, n56830 );
nor U121717 ( n56829, n56833, n56834 );
nor U121718 ( n56830, n56831, n56832 );
nor U121719 ( n56833, n73790, n56652 );
nand U121720 ( n56873, n56874, n56875 );
nor U121721 ( n56874, n56878, n56879 );
nor U121722 ( n56875, n56876, n56877 );
nor U121723 ( n56878, n73732, n56652 );
nand U121724 ( n23795, n23796, n23797 );
nor U121725 ( n23796, n23800, n23801 );
nor U121726 ( n23797, n23798, n23799 );
nor U121727 ( n23800, n73623, n23530 );
nand U121728 ( n56920, n56921, n56922 );
nor U121729 ( n56921, n56925, n56926 );
nor U121730 ( n56922, n56923, n56924 );
nor U121731 ( n56925, n73622, n56652 );
nor U121732 ( n10508, n74255, n10337 );
nor U121733 ( n44330, n73820, n44193 );
nor U121734 ( n10744, n74037, n10340 );
xor U121735 ( n42429, n74282, n893 );
nor U121736 ( n23284, n73872, n23117 );
nor U121737 ( n56408, n73873, n56238 );
nor U121738 ( n30605, n74238, n30448 );
nor U121739 ( n10048, n74253, n9853 );
nor U121740 ( n64764, n73871, n64607 );
nor U121741 ( n43964, n73818, n43764 );
nor U121742 ( n10512, n74247, n10340 );
nor U121743 ( n44333, n73812, n44196 );
nor U121744 ( n23668, n73853, n23529 );
nor U121745 ( n23712, n73771, n23529 );
nor U121746 ( n23757, n73721, n23529 );
nor U121747 ( n23623, n73922, n23529 );
nor U121748 ( n23579, n74078, n23529 );
nor U121749 ( n56745, n73923, n56651 );
nor U121750 ( n56790, n73854, n56651 );
nor U121751 ( n56701, n74077, n56651 );
nor U121752 ( n56834, n73772, n56651 );
nor U121753 ( n56879, n73720, n56651 );
nor U121754 ( n23801, n73614, n23529 );
nor U121755 ( n56926, n73613, n56651 );
nor U121756 ( n23287, n23288, n23289 );
nor U121757 ( n23288, n73862, n23111 );
nor U121758 ( n23289, n73841, n23112 );
nor U121759 ( n56411, n56412, n56413 );
nor U121760 ( n56412, n73863, n56232 );
nor U121761 ( n56413, n73842, n56233 );
nor U121762 ( n30608, n30609, n30610 );
nor U121763 ( n30609, n74233, n30442 );
nor U121764 ( n30610, n74224, n30443 );
nor U121765 ( n10051, n10052, n10053 );
nor U121766 ( n10052, n74250, n9845 );
nor U121767 ( n10053, n74243, n9847 );
nor U121768 ( n64767, n64768, n64769 );
nor U121769 ( n64768, n73861, n64601 );
nor U121770 ( n64769, n73840, n64602 );
nor U121771 ( n43967, n43968, n43969 );
nor U121772 ( n43968, n73815, n43758 );
nor U121773 ( n43969, n73808, n43759 );
nor U121774 ( n23665, n73878, n23526 );
nor U121775 ( n23709, n73795, n23526 );
nor U121776 ( n23754, n73745, n23526 );
nor U121777 ( n23620, n73946, n23526 );
nor U121778 ( n23576, n74120, n23526 );
nor U121779 ( n56742, n73947, n56648 );
nor U121780 ( n56787, n73879, n56648 );
nor U121781 ( n56698, n74119, n56648 );
nor U121782 ( n56831, n73796, n56648 );
nor U121783 ( n56876, n73744, n56648 );
nor U121784 ( n23798, n73632, n23526 );
nor U121785 ( n56923, n73631, n56648 );
nor U121786 ( n54700, n498, n54690 );
nor U121787 ( n28972, n167, n28962 );
nor U121788 ( n36145, n200, n36135 );
nand U121789 ( n36139, n36140, n76124 );
nand U121790 ( n36140, n36142, n36143 );
nor U121791 ( n36142, n74654, n73192 );
nor U121792 ( n36143, n36144, n36145 );
nor U121793 ( n23286, n23290, n23291 );
nor U121794 ( n23290, n73851, n23107 );
nor U121795 ( n23291, n73835, n23108 );
nor U121796 ( n56410, n56414, n56415 );
nor U121797 ( n56414, n73852, n56228 );
nor U121798 ( n56415, n73836, n56229 );
nor U121799 ( n30607, n30611, n30612 );
nor U121800 ( n30611, n74228, n30438 );
nor U121801 ( n30612, n74222, n30439 );
nor U121802 ( n10050, n10054, n10055 );
nor U121803 ( n10054, n74246, n9840 );
nor U121804 ( n10055, n74240, n9842 );
nor U121805 ( n64766, n64770, n64771 );
nor U121806 ( n64770, n73849, n64597 );
nor U121807 ( n64771, n73834, n64598 );
nor U121808 ( n43966, n43970, n43971 );
nor U121809 ( n43970, n73811, n43754 );
nor U121810 ( n43971, n73806, n43755 );
nand U121811 ( n42210, n42211, n42212 );
nor U121812 ( n14713, n14714, n14715 );
xor U121813 ( n14714, n14717, n5200 );
nand U121814 ( n14707, n14708, n14709 );
nand U121815 ( n14709, n5202, n14710 );
nor U121816 ( n14708, n14712, n14713 );
nor U121817 ( n14712, n14705, n14718 );
nand U121818 ( n30074, n74887, n29171 );
nor U121819 ( n63614, n63616, n63617 );
nor U121820 ( n29715, n29717, n29718 );
nor U121821 ( n22394, n22396, n22397 );
nor U121822 ( n55506, n55508, n55509 );
nand U121823 ( n64091, n74889, n62893 );
nor U121824 ( n31158, n74002, n30842 );
nor U121825 ( n44537, n73556, n44202 );
nor U121826 ( n65412, n73659, n65044 );
nand U121827 ( n31146, n31155, n31156 );
nor U121828 ( n31155, n31161, n31162 );
nor U121829 ( n31156, n31157, n31158 );
nor U121830 ( n31161, n74006, n30847 );
nand U121831 ( n44525, n44534, n44535 );
nor U121832 ( n44534, n44540, n44541 );
nor U121833 ( n44535, n44536, n44537 );
nor U121834 ( n44540, n73560, n44207 );
nand U121835 ( n65400, n65409, n65410 );
nor U121836 ( n65409, n65415, n65416 );
nor U121837 ( n65410, n65411, n65412 );
nor U121838 ( n65415, n73674, n65049 );
and U121839 ( n14747, n74649, n21107 );
nand U121840 ( n21107, n21108, n14759 );
nand U121841 ( n21108, n14812, n8285 );
and U121842 ( n47970, n74648, n54092 );
nand U121843 ( n54092, n54093, n47980 );
nand U121844 ( n54093, n48017, n42375 );
xor U121845 ( n42311, n74219, n42299 );
xor U121846 ( n37896, n74399, n37897 );
nor U121847 ( n31100, n73969, n30842 );
nor U121848 ( n30888, n74304, n30842 );
nor U121849 ( n30930, n74262, n30842 );
nor U121850 ( n30973, n74224, n30842 );
nor U121851 ( n10567, n74143, n10348 );
nor U121852 ( n10622, n74111, n10348 );
nor U121853 ( n10460, n74297, n10348 );
nor U121854 ( n10405, n74333, n10348 );
nor U121855 ( n44377, n73640, n44202 );
nor U121856 ( n44435, n73611, n44202 );
nor U121857 ( n44248, n73968, n44202 );
nor U121858 ( n44292, n73882, n44202 );
nor U121859 ( n44477, n73552, n44202 );
nor U121860 ( n10674, n73998, n10348 );
nor U121861 ( n65090, n74056, n65044 );
nor U121862 ( n65132, n73907, n65044 );
nor U121863 ( n65175, n73840, n65044 );
nor U121864 ( n65217, n73758, n65044 );
nor U121865 ( n65260, n73746, n65044 );
nor U121866 ( n31015, n74107, n30842 );
nor U121867 ( n31058, n74048, n30842 );
nor U121868 ( n65302, n73628, n65044 );
nand U121869 ( n31089, n31097, n31098 );
nor U121870 ( n31097, n31101, n31102 );
nor U121871 ( n31098, n31099, n31100 );
nor U121872 ( n31101, n73958, n30847 );
nand U121873 ( n30877, n30885, n30886 );
nor U121874 ( n30885, n30889, n30890 );
nor U121875 ( n30886, n30887, n30888 );
nor U121876 ( n30889, n74307, n30847 );
nand U121877 ( n30919, n30927, n30928 );
nor U121878 ( n30927, n30931, n30932 );
nor U121879 ( n30928, n30929, n30930 );
nor U121880 ( n30931, n74267, n30847 );
nand U121881 ( n30962, n30970, n30971 );
nor U121882 ( n30970, n30974, n30975 );
nor U121883 ( n30971, n30972, n30973 );
nor U121884 ( n30974, n74228, n30847 );
nand U121885 ( n10553, n10563, n10564 );
nor U121886 ( n10563, n10568, n10569 );
nor U121887 ( n10564, n10565, n10567 );
nor U121888 ( n10568, n74152, n10354 );
nand U121889 ( n10608, n10618, n10619 );
nor U121890 ( n10618, n10623, n10624 );
nor U121891 ( n10619, n10620, n10622 );
nor U121892 ( n10623, n74093, n10354 );
nand U121893 ( n10447, n10457, n10458 );
nor U121894 ( n10457, n10462, n10463 );
nor U121895 ( n10458, n10459, n10460 );
nor U121896 ( n10462, n74290, n10354 );
nand U121897 ( n10392, n10402, n10403 );
nor U121898 ( n10402, n10407, n10408 );
nor U121899 ( n10403, n10404, n10405 );
nor U121900 ( n10407, n74327, n10354 );
nand U121901 ( n44366, n44374, n44375 );
nor U121902 ( n44374, n44378, n44379 );
nor U121903 ( n44375, n44376, n44377 );
nor U121904 ( n44378, n73646, n44207 );
nand U121905 ( n44424, n44432, n44433 );
nor U121906 ( n44432, n44436, n44437 );
nor U121907 ( n44433, n44434, n44435 );
nor U121908 ( n44436, n73582, n44207 );
nand U121909 ( n44237, n44245, n44246 );
nor U121910 ( n44245, n44249, n44250 );
nor U121911 ( n44246, n44247, n44248 );
nor U121912 ( n44249, n73972, n44207 );
nand U121913 ( n44281, n44289, n44290 );
nor U121914 ( n44289, n44293, n44294 );
nor U121915 ( n44290, n44291, n44292 );
nor U121916 ( n44293, n73885, n44207 );
nand U121917 ( n44466, n44474, n44475 );
nor U121918 ( n44474, n44478, n44479 );
nor U121919 ( n44475, n44476, n44477 );
nor U121920 ( n44478, n73543, n44207 );
nand U121921 ( n10660, n10670, n10672 );
nor U121922 ( n10670, n10675, n10677 );
nor U121923 ( n10672, n10673, n10674 );
nor U121924 ( n10675, n73985, n10354 );
nand U121925 ( n65079, n65087, n65088 );
nor U121926 ( n65087, n65091, n65092 );
nor U121927 ( n65088, n65089, n65090 );
nor U121928 ( n65091, n74073, n65049 );
nand U121929 ( n65121, n65129, n65130 );
nor U121930 ( n65129, n65133, n65134 );
nor U121931 ( n65130, n65131, n65132 );
nor U121932 ( n65133, n73918, n65049 );
nand U121933 ( n65164, n65172, n65173 );
nor U121934 ( n65172, n65176, n65177 );
nor U121935 ( n65173, n65174, n65175 );
nor U121936 ( n65176, n73849, n65049 );
nand U121937 ( n65206, n65214, n65215 );
nor U121938 ( n65214, n65218, n65219 );
nor U121939 ( n65215, n65216, n65217 );
nor U121940 ( n65218, n73767, n65049 );
nand U121941 ( n65249, n65257, n65258 );
nor U121942 ( n65257, n65261, n65262 );
nor U121943 ( n65258, n65259, n65260 );
nor U121944 ( n65261, n73725, n65049 );
nand U121945 ( n31004, n31012, n31013 );
nor U121946 ( n31012, n31016, n31017 );
nor U121947 ( n31013, n31014, n31015 );
nor U121948 ( n31016, n74124, n30847 );
nand U121949 ( n31047, n31055, n31056 );
nor U121950 ( n31055, n31059, n31060 );
nor U121951 ( n31056, n31057, n31058 );
nor U121952 ( n31059, n74033, n30847 );
nand U121953 ( n65291, n65299, n65300 );
nor U121954 ( n65299, n65303, n65304 );
nor U121955 ( n65300, n65301, n65302 );
nor U121956 ( n65303, n73595, n65049 );
nor U121957 ( n31162, n74000, n30846 );
nor U121958 ( n44541, n73554, n44206 );
nor U121959 ( n65416, n73652, n65048 );
nor U121960 ( n31099, n73963, n30843 );
nor U121961 ( n30887, n74311, n30843 );
nor U121962 ( n30929, n74271, n30843 );
nor U121963 ( n30972, n74233, n30843 );
nor U121964 ( n10565, n74156, n10349 );
nor U121965 ( n10620, n74101, n10349 );
nor U121966 ( n10459, n74295, n10349 );
nor U121967 ( n10404, n74332, n10349 );
nor U121968 ( n44376, n73650, n44203 );
nor U121969 ( n44434, n73593, n44203 );
nor U121970 ( n44247, n73976, n44203 );
nor U121971 ( n44291, n73889, n44203 );
nor U121972 ( n44476, n73549, n44203 );
nor U121973 ( n10673, n73992, n10349 );
nor U121974 ( n65089, n74090, n65045 );
nor U121975 ( n65131, n73930, n65045 );
nor U121976 ( n65174, n73861, n65045 );
nor U121977 ( n65216, n73779, n65045 );
nor U121978 ( n65259, n73740, n65045 );
nor U121979 ( n31014, n74129, n30843 );
nor U121980 ( n31057, n74044, n30843 );
nor U121981 ( n65301, n73612, n65045 );
nor U121982 ( n10749, n74019, n10348 );
nor U121983 ( n8983, n5279, n8958 );
nor U121984 ( n42998, n7934, n42978 );
nand U121985 ( n10734, n10745, n10747 );
nor U121986 ( n10745, n10753, n10754 );
nor U121987 ( n10747, n10748, n10749 );
nor U121988 ( n10753, n74035, n10354 );
nor U121989 ( n10517, n74243, n10348 );
nor U121990 ( n44337, n73808, n44202 );
nand U121991 ( n10503, n10513, n10514 );
nor U121992 ( n10513, n10518, n10519 );
nor U121993 ( n10514, n10515, n10517 );
nor U121994 ( n10518, n74246, n10354 );
nand U121995 ( n44326, n44334, n44335 );
nor U121996 ( n44334, n44338, n44339 );
nor U121997 ( n44335, n44336, n44337 );
nor U121998 ( n44338, n73811, n44207 );
nor U121999 ( n31157, n74010, n30843 );
nor U122000 ( n30890, n74302, n30846 );
nor U122001 ( n30932, n74260, n30846 );
nor U122002 ( n30975, n74222, n30846 );
nor U122003 ( n10569, n74139, n10353 );
nor U122004 ( n10624, n74082, n10353 );
nor U122005 ( n10463, n74285, n10353 );
nor U122006 ( n10408, n74322, n10353 );
nor U122007 ( n44379, n73638, n44206 );
nor U122008 ( n44437, n73576, n44206 );
nor U122009 ( n44250, n73966, n44206 );
nor U122010 ( n44294, n73880, n44206 );
nor U122011 ( n44479, n73538, n44206 );
nor U122012 ( n10677, n73980, n10353 );
nor U122013 ( n65092, n74049, n65048 );
nor U122014 ( n65134, n73901, n65048 );
nor U122015 ( n65177, n73834, n65048 );
nor U122016 ( n65219, n73752, n65048 );
nor U122017 ( n65262, n73710, n65048 );
nor U122018 ( n31017, n74102, n30846 );
nor U122019 ( n31060, n74023, n30846 );
nor U122020 ( n65304, n73588, n65048 );
nor U122021 ( n44536, n73565, n44203 );
nor U122022 ( n10748, n74043, n10349 );
nor U122023 ( n65411, n73686, n65045 );
nor U122024 ( n31102, n73953, n30846 );
nor U122025 ( n10515, n74250, n10349 );
nor U122026 ( n44336, n73815, n44203 );
nor U122027 ( n10754, n74016, n10353 );
nor U122028 ( n30559, n74268, n30449 );
nor U122029 ( n10004, n74288, n9854 );
nor U122030 ( n64718, n73919, n64608 );
nor U122031 ( n43920, n73886, n43765 );
nand U122032 ( n30553, n30554, n30555 );
nor U122033 ( n30555, n30556, n30557 );
nor U122034 ( n30554, n30558, n30559 );
nor U122035 ( n30556, n74278, n30452 );
nand U122036 ( n9997, n9998, n9999 );
nor U122037 ( n9999, n10000, n10002 );
nor U122038 ( n9998, n10003, n10004 );
nor U122039 ( n10000, n74296, n9858 );
nand U122040 ( n64712, n64713, n64714 );
nor U122041 ( n64714, n64715, n64716 );
nor U122042 ( n64713, n64717, n64718 );
nor U122043 ( n64715, n73945, n64611 );
nand U122044 ( n43914, n43915, n43916 );
nor U122045 ( n43916, n43917, n43918 );
nor U122046 ( n43915, n43919, n43920 );
nor U122047 ( n43917, n73894, n43768 );
nor U122048 ( n10519, n74240, n10353 );
nor U122049 ( n23672, n73841, n23535 );
nor U122050 ( n23716, n73759, n23535 );
nor U122051 ( n23761, n73748, n23535 );
nor U122052 ( n23627, n73908, n23535 );
nor U122053 ( n23583, n74058, n23535 );
nor U122054 ( n44339, n73806, n44206 );
nor U122055 ( n56749, n73909, n56657 );
nor U122056 ( n56794, n73842, n56657 );
nor U122057 ( n56705, n74057, n56657 );
nor U122058 ( n56838, n73760, n56657 );
nor U122059 ( n56883, n73747, n56657 );
nor U122060 ( n23805, n73635, n23535 );
nor U122061 ( n56930, n73634, n56657 );
nor U122062 ( n23239, n73922, n23118 );
nor U122063 ( n56360, n73923, n56239 );
nand U122064 ( n23661, n23669, n23670 );
nor U122065 ( n23669, n23673, n23674 );
nor U122066 ( n23670, n23671, n23672 );
nor U122067 ( n23673, n73851, n23540 );
nand U122068 ( n23705, n23713, n23714 );
nor U122069 ( n23713, n23717, n23718 );
nor U122070 ( n23714, n23715, n23716 );
nor U122071 ( n23717, n73769, n23540 );
nand U122072 ( n23750, n23758, n23759 );
nor U122073 ( n23758, n23762, n23763 );
nor U122074 ( n23759, n23760, n23761 );
nor U122075 ( n23762, n73727, n23540 );
nand U122076 ( n23616, n23624, n23625 );
nor U122077 ( n23624, n23628, n23629 );
nor U122078 ( n23625, n23626, n23627 );
nor U122079 ( n23628, n73920, n23540 );
nand U122080 ( n23572, n23580, n23581 );
nor U122081 ( n23580, n23584, n23585 );
nor U122082 ( n23581, n23582, n23583 );
nor U122083 ( n23584, n74076, n23540 );
nand U122084 ( n56738, n56746, n56747 );
nor U122085 ( n56746, n56750, n56751 );
nor U122086 ( n56747, n56748, n56749 );
nor U122087 ( n56750, n73921, n56662 );
nand U122088 ( n56783, n56791, n56792 );
nor U122089 ( n56791, n56795, n56796 );
nor U122090 ( n56792, n56793, n56794 );
nor U122091 ( n56795, n73852, n56662 );
nand U122092 ( n56694, n56702, n56703 );
nor U122093 ( n56702, n56706, n56707 );
nor U122094 ( n56703, n56704, n56705 );
nor U122095 ( n56706, n74075, n56662 );
nand U122096 ( n56827, n56835, n56836 );
nor U122097 ( n56835, n56839, n56840 );
nor U122098 ( n56836, n56837, n56838 );
nor U122099 ( n56839, n73770, n56662 );
nand U122100 ( n56872, n56880, n56881 );
nor U122101 ( n56880, n56884, n56885 );
nor U122102 ( n56881, n56882, n56883 );
nor U122103 ( n56884, n73726, n56662 );
nand U122104 ( n23794, n23802, n23803 );
nor U122105 ( n23802, n23806, n23807 );
nor U122106 ( n23803, n23804, n23805 );
nor U122107 ( n23806, n73618, n23540 );
nand U122108 ( n56919, n56927, n56928 );
nor U122109 ( n56927, n56931, n56932 );
nor U122110 ( n56928, n56929, n56930 );
nor U122111 ( n56931, n73617, n56662 );
nand U122112 ( n23233, n23234, n23235 );
nor U122113 ( n23235, n23236, n23237 );
nor U122114 ( n23234, n23238, n23239 );
nor U122115 ( n23236, n73946, n23121 );
nand U122116 ( n56354, n56355, n56356 );
nor U122117 ( n56356, n56357, n56358 );
nor U122118 ( n56355, n56359, n56360 );
nor U122119 ( n56357, n73947, n56242 );
nor U122120 ( n30557, n74272, n30453 );
nor U122121 ( n10002, n74294, n9859 );
nor U122122 ( n64716, n73933, n64612 );
nor U122123 ( n43918, n73890, n43769 );
nor U122124 ( n23237, n73934, n23122 );
nor U122125 ( n56358, n73935, n56243 );
nor U122126 ( n23674, n73835, n23539 );
nor U122127 ( n23718, n73753, n23539 );
nor U122128 ( n23763, n73713, n23539 );
nor U122129 ( n23629, n73902, n23539 );
nor U122130 ( n23585, n74051, n23539 );
nor U122131 ( n56751, n73903, n56661 );
nor U122132 ( n56796, n73836, n56661 );
nor U122133 ( n56707, n74050, n56661 );
nor U122134 ( n56840, n73754, n56661 );
nor U122135 ( n56885, n73712, n56661 );
nor U122136 ( n23807, n73605, n23539 );
nor U122137 ( n56932, n73604, n56661 );
nor U122138 ( n23671, n73862, n23536 );
nor U122139 ( n23715, n73780, n23536 );
nor U122140 ( n23760, n73742, n23536 );
nor U122141 ( n23626, n73931, n23536 );
nor U122142 ( n23582, n74092, n23536 );
nor U122143 ( n56748, n73932, n56658 );
nor U122144 ( n56793, n73863, n56658 );
nor U122145 ( n56704, n74091, n56658 );
nor U122146 ( n56837, n73781, n56658 );
nor U122147 ( n56882, n73741, n56658 );
nor U122148 ( n23804, n73630, n23536 );
nor U122149 ( n56929, n73629, n56658 );
not U122150 ( n6162, n63615 );
not U122151 ( n3547, n29716 );
not U122152 ( n4384, n22395 );
not U122153 ( n7017, n55507 );
xor U122154 ( n37844, n74372, n37841 );
nor U122155 ( n30505, n74309, n30464 );
nor U122156 ( n9929, n74328, n9873 );
nor U122157 ( n64664, n74079, n64623 );
nor U122158 ( n43825, n73974, n43780 );
nand U122159 ( n30495, n30503, n30504 );
nor U122160 ( n30503, n30507, n30508 );
nor U122161 ( n30504, n30505, n30506 );
nor U122162 ( n30507, n74305, n30460 );
nand U122163 ( n9917, n9927, n9928 );
nor U122164 ( n9927, n9932, n9933 );
nor U122165 ( n9928, n9929, n9930 );
nor U122166 ( n9932, n74321, n9868 );
nand U122167 ( n64654, n64662, n64663 );
nor U122168 ( n64662, n64666, n64667 );
nor U122169 ( n64663, n64664, n64665 );
nor U122170 ( n64666, n74065, n64619 );
nand U122171 ( n43815, n43823, n43824 );
nor U122172 ( n43823, n43827, n43828 );
nor U122173 ( n43824, n43825, n43826 );
nor U122174 ( n43827, n73970, n43776 );
nor U122175 ( n23181, n74081, n23133 );
nor U122176 ( n56302, n74080, n56254 );
nand U122177 ( n23171, n23179, n23180 );
nor U122178 ( n23179, n23183, n23184 );
nor U122179 ( n23180, n23181, n23182 );
nor U122180 ( n23183, n74068, n23129 );
nand U122181 ( n56292, n56300, n56301 );
nor U122182 ( n56300, n56304, n56305 );
nor U122183 ( n56301, n56302, n56303 );
nor U122184 ( n56304, n74067, n56250 );
xor U122185 ( n37705, n73804, n37706 );
nor U122186 ( n30558, n74276, n30448 );
nor U122187 ( n10003, n74292, n9853 );
nor U122188 ( n64717, n73939, n64607 );
nor U122189 ( n43919, n73892, n43764 );
nor U122190 ( n30508, n74299, n30461 );
nor U122191 ( n9933, n74319, n9869 );
nor U122192 ( n64667, n74027, n64620 );
nor U122193 ( n43828, n73950, n43777 );
nor U122194 ( n23238, n73940, n23117 );
nor U122195 ( n56359, n73941, n56238 );
nor U122196 ( n23184, n74029, n23130 );
nor U122197 ( n56305, n74028, n56251 );
nor U122198 ( n23859, n73691, n23525 );
nor U122199 ( n56983, n73690, n56647 );
nand U122200 ( n23855, n23856, n23857 );
nor U122201 ( n23856, n23861, n23862 );
nor U122202 ( n23857, n23858, n23859 );
nor U122203 ( n23861, n73697, n23530 );
nand U122204 ( n56979, n56980, n56981 );
nor U122205 ( n56980, n56985, n56986 );
nor U122206 ( n56981, n56982, n56983 );
nor U122207 ( n56985, n73696, n56652 );
xnor U122208 ( n37707, n37708, n37709 );
xor U122209 ( n37709, n73802, n37706 );
nor U122210 ( n23858, n73704, n23526 );
nor U122211 ( n56982, n73703, n56648 );
nor U122212 ( n30561, n30562, n30563 );
nor U122213 ( n30562, n74271, n30442 );
nor U122214 ( n30563, n74262, n30443 );
nor U122215 ( n10006, n10007, n10008 );
nor U122216 ( n10007, n74295, n9845 );
nor U122217 ( n10008, n74297, n9847 );
nor U122218 ( n64720, n64721, n64722 );
nor U122219 ( n64721, n73930, n64601 );
nor U122220 ( n64722, n73907, n64602 );
nor U122221 ( n43922, n43923, n43924 );
nor U122222 ( n43923, n73889, n43758 );
nor U122223 ( n43924, n73882, n43759 );
nor U122224 ( n23241, n23242, n23243 );
nor U122225 ( n23242, n73931, n23111 );
nor U122226 ( n23243, n73908, n23112 );
nor U122227 ( n56362, n56363, n56364 );
nor U122228 ( n56363, n73932, n56232 );
nor U122229 ( n56364, n73909, n56233 );
nor U122230 ( n23862, n73680, n23529 );
nor U122231 ( n56986, n73679, n56651 );
nor U122232 ( n30560, n30564, n30565 );
nor U122233 ( n30564, n74267, n30438 );
nor U122234 ( n30565, n74260, n30439 );
nor U122235 ( n10005, n10009, n10010 );
nor U122236 ( n10009, n74290, n9840 );
nor U122237 ( n10010, n74285, n9842 );
nor U122238 ( n64719, n64723, n64724 );
nor U122239 ( n64723, n73918, n64597 );
nor U122240 ( n64724, n73901, n64598 );
nor U122241 ( n43921, n43925, n43926 );
nor U122242 ( n43925, n73885, n43754 );
nor U122243 ( n43926, n73880, n43755 );
nor U122244 ( n23240, n23244, n23245 );
nor U122245 ( n23244, n73920, n23107 );
nor U122246 ( n23245, n73902, n23108 );
nor U122247 ( n56361, n56365, n56366 );
nor U122248 ( n56365, n73921, n56228 );
nor U122249 ( n56366, n73903, n56229 );
nor U122250 ( n14685, n14687, n14688 );
nor U122251 ( n14687, n14689, n14690 );
nor U122252 ( n14689, n14692, n74435 );
nand U122253 ( n8786, n14682, n14683 );
nor U122254 ( n14682, n14694, n14695 );
nor U122255 ( n14683, n14684, n14685 );
nor U122256 ( n14695, n14679, n14697 );
nor U122257 ( n31142, n74001, n30820 );
nor U122258 ( n44521, n73555, n44180 );
nor U122259 ( n10729, n74017, n10320 );
nor U122260 ( n65396, n73655, n65022 );
nand U122261 ( n31121, n31139, n31140 );
nor U122262 ( n31139, n31144, n31145 );
nor U122263 ( n31140, n31141, n31142 );
nor U122264 ( n31144, n74003, n30825 );
nand U122265 ( n44500, n44518, n44519 );
nor U122266 ( n44518, n44523, n44524 );
nor U122267 ( n44519, n44520, n44521 );
nor U122268 ( n44523, n73557, n44185 );
nand U122269 ( n10703, n10725, n10727 );
nor U122270 ( n10725, n10732, n10733 );
nor U122271 ( n10727, n10728, n10729 );
nor U122272 ( n10732, n74026, n10327 );
nand U122273 ( n65375, n65393, n65394 );
nor U122274 ( n65393, n65398, n65399 );
nor U122275 ( n65394, n65395, n65396 );
nor U122276 ( n65398, n73665, n65027 );
nor U122277 ( n30590, n74231, n30475 );
nor U122278 ( n10033, n74249, n9887 );
nor U122279 ( n64749, n73858, n64634 );
nor U122280 ( n43949, n73814, n43791 );
nand U122281 ( n30586, n30587, n30588 );
nor U122282 ( n30587, n30591, n30592 );
nor U122283 ( n30588, n30589, n30590 );
nor U122284 ( n30591, n74237, n30470 );
nand U122285 ( n10029, n10030, n10031 );
nor U122286 ( n10030, n10034, n10035 );
nor U122287 ( n10031, n10032, n10033 );
nor U122288 ( n10034, n74252, n9880 );
nand U122289 ( n64745, n64746, n64747 );
nor U122290 ( n64746, n64750, n64751 );
nor U122291 ( n64747, n64748, n64749 );
nor U122292 ( n64750, n73868, n64629 );
nand U122293 ( n43945, n43946, n43947 );
nor U122294 ( n43946, n43950, n43951 );
nor U122295 ( n43947, n43948, n43949 );
nor U122296 ( n43950, n73817, n43786 );
nor U122297 ( n30596, n74223, n30465 );
nor U122298 ( n10039, n74241, n9874 );
nor U122299 ( n64755, n73837, n64624 );
nor U122300 ( n43955, n73807, n43781 );
nand U122301 ( n62502, n8209, n74683 );
nand U122302 ( n70886, n8209, n73186 );
nor U122303 ( n30589, n74239, n30474 );
nor U122304 ( n10032, n74254, n9885 );
nor U122305 ( n64748, n73874, n64633 );
nor U122306 ( n43948, n73819, n43790 );
nor U122307 ( n23269, n73859, n23144 );
nor U122308 ( n56393, n73860, n56265 );
nand U122309 ( n23265, n23266, n23267 );
nor U122310 ( n23266, n23270, n23271 );
nor U122311 ( n23267, n23268, n23269 );
nor U122312 ( n23270, n73869, n23139 );
nand U122313 ( n56389, n56390, n56391 );
nor U122314 ( n56390, n56394, n56395 );
nor U122315 ( n56391, n56392, n56393 );
nor U122316 ( n56394, n73870, n56260 );
nor U122317 ( n23275, n73838, n23134 );
nor U122318 ( n56399, n73839, n56255 );
nor U122319 ( n31145, n73987, n30824 );
nor U122320 ( n44524, n73553, n44184 );
nor U122321 ( n10733, n74005, n10325 );
nor U122322 ( n65399, n73643, n65026 );
nor U122323 ( n23268, n73875, n23143 );
nor U122324 ( n56392, n73876, n56264 );
nor U122325 ( n45674, n45658, n45675 );
nor U122326 ( n30592, n74227, n30471 );
nor U122327 ( n10035, n74245, n9882 );
nor U122328 ( n64751, n73844, n64630 );
nor U122329 ( n43951, n73810, n43787 );
nor U122330 ( n11937, n11912, n11938 );
nor U122331 ( n66598, n66582, n66599 );
nor U122332 ( n31995, n31979, n31996 );
nor U122333 ( n24763, n24747, n24764 );
nor U122334 ( n57897, n57881, n57898 );
nor U122335 ( n31086, n73954, n30820 );
nor U122336 ( n30874, n74303, n30820 );
nor U122337 ( n30916, n74261, n30820 );
nor U122338 ( n30959, n74223, n30820 );
nor U122339 ( n10549, n74140, n10320 );
nor U122340 ( n10604, n74084, n10320 );
nor U122341 ( n10443, n74286, n10320 );
nor U122342 ( n10388, n74323, n10320 );
nor U122343 ( n44363, n73639, n44180 );
nor U122344 ( n44421, n73577, n44180 );
nor U122345 ( n44234, n73967, n44180 );
nor U122346 ( n44278, n73881, n44180 );
nor U122347 ( n44463, n73539, n44180 );
nor U122348 ( n10657, n73981, n10320 );
nor U122349 ( n65076, n74053, n65022 );
nor U122350 ( n65118, n73904, n65022 );
nor U122351 ( n65161, n73837, n65022 );
nor U122352 ( n65203, n73755, n65022 );
nor U122353 ( n65246, n73714, n65022 );
nor U122354 ( n31001, n74104, n30820 );
nor U122355 ( n31044, n74024, n30820 );
nor U122356 ( n65288, n73589, n65022 );
nor U122357 ( n23271, n73847, n23140 );
nor U122358 ( n56395, n73848, n56261 );
nand U122359 ( n31075, n31083, n31084 );
nor U122360 ( n31083, n31087, n31088 );
nor U122361 ( n31084, n31085, n31086 );
nor U122362 ( n31087, n73952, n30825 );
nand U122363 ( n30863, n30871, n30872 );
nor U122364 ( n30871, n30875, n30876 );
nor U122365 ( n30872, n30873, n30874 );
nor U122366 ( n30875, n74305, n30825 );
nand U122367 ( n30905, n30913, n30914 );
nor U122368 ( n30913, n30917, n30918 );
nor U122369 ( n30914, n30915, n30916 );
nor U122370 ( n30917, n74264, n30825 );
nand U122371 ( n30948, n30956, n30957 );
nor U122372 ( n30956, n30960, n30961 );
nor U122373 ( n30957, n30958, n30959 );
nor U122374 ( n30960, n74226, n30825 );
nand U122375 ( n10535, n10545, n10547 );
nor U122376 ( n10545, n10550, n10552 );
nor U122377 ( n10547, n10548, n10549 );
nor U122378 ( n10550, n74149, n10327 );
nand U122379 ( n10590, n10600, n10602 );
nor U122380 ( n10600, n10605, n10607 );
nor U122381 ( n10602, n10603, n10604 );
nor U122382 ( n10605, n74072, n10327 );
nand U122383 ( n10429, n10439, n10440 );
nor U122384 ( n10439, n10444, n10445 );
nor U122385 ( n10440, n10442, n10443 );
nor U122386 ( n10444, n74284, n10327 );
nand U122387 ( n10374, n10384, n10385 );
nor U122388 ( n10384, n10389, n10390 );
nor U122389 ( n10385, n10387, n10388 );
nor U122390 ( n10389, n74321, n10327 );
nand U122391 ( n44352, n44360, n44361 );
nor U122392 ( n44360, n44364, n44365 );
nor U122393 ( n44361, n44362, n44363 );
nor U122394 ( n44364, n73644, n44185 );
nand U122395 ( n44410, n44418, n44419 );
nor U122396 ( n44418, n44422, n44423 );
nor U122397 ( n44419, n44420, n44421 );
nor U122398 ( n44422, n73575, n44185 );
nand U122399 ( n44223, n44231, n44232 );
nor U122400 ( n44231, n44235, n44236 );
nor U122401 ( n44232, n44233, n44234 );
nor U122402 ( n44235, n73970, n44185 );
nand U122403 ( n44267, n44275, n44276 );
nor U122404 ( n44275, n44279, n44280 );
nor U122405 ( n44276, n44277, n44278 );
nor U122406 ( n44279, n73883, n44185 );
nand U122407 ( n44452, n44460, n44461 );
nor U122408 ( n44460, n44464, n44465 );
nor U122409 ( n44461, n44462, n44463 );
nor U122410 ( n44464, n73537, n44185 );
nand U122411 ( n10643, n10653, n10654 );
nor U122412 ( n10653, n10658, n10659 );
nor U122413 ( n10654, n10655, n10657 );
nor U122414 ( n10658, n73979, n10327 );
nand U122415 ( n65065, n65073, n65074 );
nor U122416 ( n65073, n65077, n65078 );
nor U122417 ( n65074, n65075, n65076 );
nor U122418 ( n65077, n74065, n65027 );
nand U122419 ( n65107, n65115, n65116 );
nor U122420 ( n65115, n65119, n65120 );
nor U122421 ( n65116, n65117, n65118 );
nor U122422 ( n65119, n73912, n65027 );
nand U122423 ( n65150, n65158, n65159 );
nor U122424 ( n65158, n65162, n65163 );
nor U122425 ( n65159, n65160, n65161 );
nor U122426 ( n65162, n73843, n65027 );
nand U122427 ( n65192, n65200, n65201 );
nor U122428 ( n65200, n65204, n65205 );
nor U122429 ( n65201, n65202, n65203 );
nor U122430 ( n65204, n73761, n65027 );
nand U122431 ( n65235, n65243, n65244 );
nor U122432 ( n65243, n65247, n65248 );
nor U122433 ( n65244, n65245, n65246 );
nor U122434 ( n65247, n73707, n65027 );
nand U122435 ( n30990, n30998, n30999 );
nor U122436 ( n30998, n31002, n31003 );
nor U122437 ( n30999, n31000, n31001 );
nor U122438 ( n31002, n74121, n30825 );
nand U122439 ( n31033, n31041, n31042 );
nor U122440 ( n31041, n31045, n31046 );
nor U122441 ( n31042, n31043, n31044 );
nor U122442 ( n31045, n74022, n30825 );
nand U122443 ( n65277, n65285, n65286 );
nor U122444 ( n65285, n65289, n65290 );
nor U122445 ( n65286, n65287, n65288 );
nor U122446 ( n65289, n73585, n65027 );
nor U122447 ( n23658, n73838, n23513 );
nor U122448 ( n23702, n73756, n23513 );
nor U122449 ( n23747, n73716, n23513 );
nor U122450 ( n23613, n73905, n23513 );
nor U122451 ( n23569, n74055, n23513 );
nor U122452 ( n56735, n73906, n56635 );
nor U122453 ( n56780, n73839, n56635 );
nor U122454 ( n56691, n74054, n56635 );
nor U122455 ( n56824, n73757, n56635 );
nor U122456 ( n56869, n73715, n56635 );
nor U122457 ( n23791, n73607, n23513 );
nor U122458 ( n56916, n73606, n56635 );
nand U122459 ( n23647, n23655, n23656 );
nor U122460 ( n23655, n23659, n23660 );
nor U122461 ( n23656, n23657, n23658 );
nor U122462 ( n23659, n73845, n23518 );
nand U122463 ( n23691, n23699, n23700 );
nor U122464 ( n23699, n23703, n23704 );
nor U122465 ( n23700, n23701, n23702 );
nor U122466 ( n23703, n73763, n23518 );
nand U122467 ( n23736, n23744, n23745 );
nor U122468 ( n23744, n23748, n23749 );
nor U122469 ( n23745, n23746, n23747 );
nor U122470 ( n23748, n73709, n23518 );
nand U122471 ( n23602, n23610, n23611 );
nor U122472 ( n23610, n23614, n23615 );
nor U122473 ( n23611, n23612, n23613 );
nor U122474 ( n23614, n73914, n23518 );
nand U122475 ( n23558, n23566, n23567 );
nor U122476 ( n23566, n23570, n23571 );
nor U122477 ( n23567, n23568, n23569 );
nor U122478 ( n23570, n74068, n23518 );
nand U122479 ( n56724, n56732, n56733 );
nor U122480 ( n56732, n56736, n56737 );
nor U122481 ( n56733, n56734, n56735 );
nor U122482 ( n56736, n73915, n56640 );
nand U122483 ( n56769, n56777, n56778 );
nor U122484 ( n56777, n56781, n56782 );
nor U122485 ( n56778, n56779, n56780 );
nor U122486 ( n56781, n73846, n56640 );
nand U122487 ( n56680, n56688, n56689 );
nor U122488 ( n56688, n56692, n56693 );
nor U122489 ( n56689, n56690, n56691 );
nor U122490 ( n56692, n74067, n56640 );
nand U122491 ( n56813, n56821, n56822 );
nor U122492 ( n56821, n56825, n56826 );
nor U122493 ( n56822, n56823, n56824 );
nor U122494 ( n56825, n73764, n56640 );
nand U122495 ( n56858, n56866, n56867 );
nor U122496 ( n56866, n56870, n56871 );
nor U122497 ( n56867, n56868, n56869 );
nor U122498 ( n56870, n73708, n56640 );
nand U122499 ( n23780, n23788, n23789 );
nor U122500 ( n23788, n23792, n23793 );
nor U122501 ( n23789, n23790, n23791 );
nor U122502 ( n23792, n73601, n23518 );
nand U122503 ( n56905, n56913, n56914 );
nor U122504 ( n56913, n56917, n56918 );
nor U122505 ( n56914, n56915, n56916 );
nor U122506 ( n56917, n73600, n56640 );
nor U122507 ( n31088, n73949, n30824 );
nor U122508 ( n30876, n74299, n30824 );
nor U122509 ( n30918, n74258, n30824 );
nor U122510 ( n30961, n74221, n30824 );
nor U122511 ( n10552, n74128, n10325 );
nor U122512 ( n10607, n74046, n10325 );
nor U122513 ( n10445, n74280, n10325 );
nor U122514 ( n10390, n74319, n10325 );
nor U122515 ( n44365, n73636, n44184 );
nor U122516 ( n44423, n73558, n44184 );
nor U122517 ( n44236, n73950, n44184 );
nor U122518 ( n44280, n73867, n44184 );
nor U122519 ( n44465, n73534, n44184 );
nor U122520 ( n10659, n73964, n10325 );
nor U122521 ( n65078, n74027, n65026 );
nor U122522 ( n65120, n73898, n65026 );
nor U122523 ( n65163, n73830, n65026 );
nor U122524 ( n65205, n73749, n65026 );
nor U122525 ( n65248, n73666, n65026 );
nor U122526 ( n31003, n74063, n30824 );
nor U122527 ( n31046, n74012, n30824 );
nor U122528 ( n65290, n73564, n65026 );
nor U122529 ( n23866, n73661, n23535 );
nor U122530 ( n56990, n73660, n56657 );
nor U122531 ( n31141, n74008, n30821 );
nor U122532 ( n44520, n73562, n44181 );
nor U122533 ( n10728, n74038, n10322 );
nor U122534 ( n65395, n73676, n65023 );
nor U122535 ( n10499, n74241, n10320 );
nor U122536 ( n44323, n73807, n44180 );
nand U122537 ( n10485, n10495, n10497 );
nor U122538 ( n10495, n10500, n10502 );
nor U122539 ( n10497, n10498, n10499 );
nor U122540 ( n10500, n74244, n10327 );
nand U122541 ( n44312, n44320, n44321 );
nor U122542 ( n44320, n44324, n44325 );
nor U122543 ( n44321, n44322, n44323 );
nor U122544 ( n44324, n73809, n44185 );
nand U122545 ( n23854, n23863, n23864 );
nor U122546 ( n23863, n23869, n23870 );
nor U122547 ( n23864, n23865, n23866 );
nor U122548 ( n23869, n73678, n23540 );
nand U122549 ( n56978, n56987, n56988 );
nor U122550 ( n56987, n56993, n56994 );
nor U122551 ( n56988, n56989, n56990 );
nor U122552 ( n56993, n73677, n56662 );
nor U122553 ( n31124, n31125, n31126 );
nor U122554 ( n31125, n74015, n30811 );
nor U122555 ( n31126, n74009, n30810 );
nor U122556 ( n44503, n44504, n44505 );
nor U122557 ( n44504, n73572, n44171 );
nor U122558 ( n44505, n73563, n44170 );
nor U122559 ( n10707, n10708, n10709 );
nor U122560 ( n10708, n74060, n10309 );
nor U122561 ( n10709, n74039, n10308 );
nor U122562 ( n65378, n65379, n65380 );
nor U122563 ( n65379, n73698, n65013 );
nor U122564 ( n65380, n73681, n65012 );
nor U122565 ( n23865, n73689, n23536 );
nor U122566 ( n56989, n73688, n56658 );
nor U122567 ( n23660, n73831, n23517 );
nor U122568 ( n23704, n73750, n23517 );
nor U122569 ( n23749, n73671, n23517 );
nor U122570 ( n23615, n73899, n23517 );
nor U122571 ( n23571, n74029, n23517 );
nor U122572 ( n56737, n73900, n56639 );
nor U122573 ( n56782, n73832, n56639 );
nor U122574 ( n56693, n74028, n56639 );
nor U122575 ( n56826, n73751, n56639 );
nor U122576 ( n56871, n73670, n56639 );
nor U122577 ( n23793, n73569, n23517 );
nor U122578 ( n56918, n73568, n56639 );
nor U122579 ( n23870, n73654, n23539 );
nor U122580 ( n56994, n73653, n56661 );
nor U122581 ( n10502, n74232, n10325 );
nor U122582 ( n44325, n73805, n44184 );
nor U122583 ( n31123, n31133, n31134 );
nor U122584 ( n31133, n74013, n30815 );
nor U122585 ( n31134, n74004, n30814 );
nor U122586 ( n44502, n44512, n44513 );
nor U122587 ( n44512, n73570, n44175 );
nor U122588 ( n44513, n73559, n44174 );
nor U122589 ( n10705, n10718, n10719 );
nor U122590 ( n10718, n74052, n10314 );
nor U122591 ( n10719, n74031, n10313 );
nor U122592 ( n65377, n65387, n65388 );
nor U122593 ( n65387, n73692, n65017 );
nor U122594 ( n65388, n73667, n65016 );
nor U122595 ( n31085, n73959, n30821 );
nor U122596 ( n30873, n74309, n30821 );
nor U122597 ( n30915, n74269, n30821 );
nor U122598 ( n30958, n74230, n30821 );
nor U122599 ( n10548, n74154, n10322 );
nor U122600 ( n10603, n74097, n10322 );
nor U122601 ( n10442, n74291, n10322 );
nor U122602 ( n10387, n74328, n10322 );
nor U122603 ( n44362, n73648, n44181 );
nor U122604 ( n44420, n73584, n44181 );
nor U122605 ( n44233, n73974, n44181 );
nor U122606 ( n44277, n73887, n44181 );
nor U122607 ( n44462, n73545, n44181 );
nor U122608 ( n10655, n73986, n10322 );
nor U122609 ( n65075, n74079, n65023 );
nor U122610 ( n65117, n73924, n65023 );
nor U122611 ( n65160, n73855, n65023 );
nor U122612 ( n65202, n73773, n65023 );
nor U122613 ( n65245, n73728, n65023 );
nor U122614 ( n31000, n74126, n30821 );
nor U122615 ( n31043, n74034, n30821 );
nor U122616 ( n65287, n73596, n65023 );
nand U122617 ( n21686, n21687, n76557 );
nor U122618 ( n31078, n31079, n31080 );
nor U122619 ( n31079, n73961, n30811 );
nor U122620 ( n31080, n73957, n30810 );
nor U122621 ( n30866, n30867, n30868 );
nor U122622 ( n30867, n74316, n30811 );
nor U122623 ( n30868, n74310, n30810 );
nor U122624 ( n30908, n30909, n30910 );
nor U122625 ( n30909, n74277, n30811 );
nor U122626 ( n30910, n74270, n30810 );
nor U122627 ( n30951, n30952, n30953 );
nor U122628 ( n30952, n74239, n30811 );
nor U122629 ( n30953, n74231, n30810 );
nor U122630 ( n10539, n10540, n10542 );
nor U122631 ( n10540, n74163, n10309 );
nor U122632 ( n10542, n74155, n10308 );
nor U122633 ( n10594, n10595, n10597 );
nor U122634 ( n10595, n74099, n10309 );
nor U122635 ( n10597, n74089, n10308 );
nor U122636 ( n10433, n10434, n10435 );
nor U122637 ( n10434, n74293, n10309 );
nor U122638 ( n10435, n74289, n10308 );
nor U122639 ( n10378, n10379, n10380 );
nor U122640 ( n10379, n74330, n10309 );
nor U122641 ( n10380, n74326, n10308 );
nor U122642 ( n44355, n44356, n44357 );
nor U122643 ( n44356, n73663, n44171 );
nor U122644 ( n44357, n73649, n44170 );
nor U122645 ( n44413, n44414, n44415 );
nor U122646 ( n44414, n73587, n44171 );
nor U122647 ( n44415, n73581, n44170 );
nor U122648 ( n44226, n44227, n44228 );
nor U122649 ( n44227, n73994, n44171 );
nor U122650 ( n44228, n73975, n44170 );
nor U122651 ( n44270, n44271, n44272 );
nor U122652 ( n44271, n73893, n44171 );
nor U122653 ( n44272, n73888, n44170 );
nor U122654 ( n44455, n44456, n44457 );
nor U122655 ( n44456, n73547, n44171 );
nor U122656 ( n44457, n73542, n44170 );
nor U122657 ( n10647, n10648, n10649 );
nor U122658 ( n10648, n73989, n10309 );
nor U122659 ( n10649, n73984, n10308 );
nor U122660 ( n65068, n65069, n65070 );
nor U122661 ( n65069, n74115, n65013 );
nor U122662 ( n65070, n74083, n65012 );
nor U122663 ( n65110, n65111, n65112 );
nor U122664 ( n65111, n73942, n65013 );
nor U122665 ( n65112, n73927, n65012 );
nor U122666 ( n65153, n65154, n65155 );
nor U122667 ( n65154, n73874, n65013 );
nor U122668 ( n65155, n73858, n65012 );
nor U122669 ( n65195, n65196, n65197 );
nor U122670 ( n65196, n73791, n65013 );
nor U122671 ( n65197, n73776, n65012 );
nor U122672 ( n65238, n65239, n65240 );
nor U122673 ( n65239, n73734, n65013 );
nor U122674 ( n65240, n73722, n65012 );
nor U122675 ( n30993, n30994, n30995 );
nor U122676 ( n30994, n74137, n30811 );
nor U122677 ( n30995, n74127, n30810 );
nor U122678 ( n31036, n31037, n31038 );
nor U122679 ( n31037, n74040, n30811 );
nor U122680 ( n31038, n74032, n30810 );
nor U122681 ( n65280, n65281, n65282 );
nor U122682 ( n65281, n73603, n65013 );
nor U122683 ( n65282, n73594, n65012 );
nor U122684 ( n23657, n73856, n23514 );
nor U122685 ( n23701, n73774, n23514 );
nor U122686 ( n23746, n73730, n23514 );
nor U122687 ( n23612, n73925, n23514 );
nor U122688 ( n23568, n74081, n23514 );
nor U122689 ( n56734, n73926, n56636 );
nor U122690 ( n56779, n73857, n56636 );
nor U122691 ( n56690, n74080, n56636 );
nor U122692 ( n56823, n73775, n56636 );
nor U122693 ( n56868, n73729, n56636 );
nor U122694 ( n23790, n73620, n23514 );
nor U122695 ( n56915, n73619, n56636 );
nor U122696 ( n23650, n23651, n23652 );
nor U122697 ( n23651, n73875, n23504 );
nor U122698 ( n23652, n73859, n23503 );
nor U122699 ( n23694, n23695, n23696 );
nor U122700 ( n23695, n73792, n23504 );
nor U122701 ( n23696, n73777, n23503 );
nor U122702 ( n23739, n23740, n23741 );
nor U122703 ( n23740, n73736, n23504 );
nor U122704 ( n23741, n73724, n23503 );
nor U122705 ( n23605, n23606, n23607 );
nor U122706 ( n23606, n73943, n23504 );
nor U122707 ( n23607, n73928, n23503 );
nor U122708 ( n23561, n23562, n23563 );
nor U122709 ( n23562, n74117, n23504 );
nor U122710 ( n23563, n74087, n23503 );
nor U122711 ( n56727, n56728, n56729 );
nor U122712 ( n56728, n73944, n56626 );
nor U122713 ( n56729, n73929, n56625 );
nor U122714 ( n56772, n56773, n56774 );
nor U122715 ( n56773, n73876, n56626 );
nor U122716 ( n56774, n73860, n56625 );
nor U122717 ( n56683, n56684, n56685 );
nor U122718 ( n56684, n74116, n56626 );
nor U122719 ( n56685, n74086, n56625 );
nor U122720 ( n56816, n56817, n56818 );
nor U122721 ( n56817, n73793, n56626 );
nor U122722 ( n56818, n73778, n56625 );
nor U122723 ( n56861, n56862, n56863 );
nor U122724 ( n56862, n73735, n56626 );
nor U122725 ( n56863, n73723, n56625 );
nor U122726 ( n23783, n23784, n23785 );
nor U122727 ( n23784, n73625, n23504 );
nor U122728 ( n23785, n73616, n23503 );
nor U122729 ( n56908, n56909, n56910 );
nor U122730 ( n56909, n73624, n56626 );
nor U122731 ( n56910, n73615, n56625 );
nor U122732 ( n10498, n74248, n10322 );
nor U122733 ( n44322, n73813, n44181 );
nor U122734 ( n31077, n31081, n31082 );
nor U122735 ( n31081, n73955, n30815 );
nor U122736 ( n31082, n73951, n30814 );
nor U122737 ( n30865, n30869, n30870 );
nor U122738 ( n30869, n74313, n30815 );
nor U122739 ( n30870, n74306, n30814 );
nor U122740 ( n30907, n30911, n30912 );
nor U122741 ( n30911, n74275, n30815 );
nor U122742 ( n30912, n74265, n30814 );
nor U122743 ( n30950, n30954, n30955 );
nor U122744 ( n30954, n74237, n30815 );
nor U122745 ( n30955, n74227, n30814 );
nor U122746 ( n10538, n10543, n10544 );
nor U122747 ( n10543, n74161, n10314 );
nor U122748 ( n10544, n74150, n10313 );
nor U122749 ( n10593, n10598, n10599 );
nor U122750 ( n10598, n74085, n10314 );
nor U122751 ( n10599, n74071, n10313 );
nor U122752 ( n10432, n10437, n10438 );
nor U122753 ( n10437, n74287, n10314 );
nor U122754 ( n10438, n74283, n10313 );
nor U122755 ( n10377, n10382, n10383 );
nor U122756 ( n10382, n74324, n10314 );
nor U122757 ( n10383, n74320, n10313 );
nor U122758 ( n44354, n44358, n44359 );
nor U122759 ( n44358, n73656, n44175 );
nor U122760 ( n44359, n73645, n44174 );
nor U122761 ( n44412, n44416, n44417 );
nor U122762 ( n44416, n73578, n44175 );
nor U122763 ( n44417, n73573, n44174 );
nor U122764 ( n44225, n44229, n44230 );
nor U122765 ( n44229, n73990, n44175 );
nor U122766 ( n44230, n73971, n44174 );
nor U122767 ( n44269, n44273, n44274 );
nor U122768 ( n44273, n73891, n44175 );
nor U122769 ( n44274, n73884, n44174 );
nor U122770 ( n44454, n44458, n44459 );
nor U122771 ( n44458, n73540, n44175 );
nor U122772 ( n44459, n73536, n44174 );
nor U122773 ( n10645, n10650, n10652 );
nor U122774 ( n10650, n73982, n10314 );
nor U122775 ( n10652, n73978, n10313 );
nor U122776 ( n65067, n65071, n65072 );
nor U122777 ( n65071, n74108, n65017 );
nor U122778 ( n65072, n74066, n65016 );
nor U122779 ( n65109, n65113, n65114 );
nor U122780 ( n65113, n73936, n65017 );
nor U122781 ( n65114, n73913, n65016 );
nor U122782 ( n65152, n65156, n65157 );
nor U122783 ( n65156, n73868, n65017 );
nor U122784 ( n65157, n73844, n65016 );
nor U122785 ( n65194, n65198, n65199 );
nor U122786 ( n65198, n73785, n65017 );
nor U122787 ( n65199, n73762, n65016 );
nor U122788 ( n65237, n65241, n65242 );
nor U122789 ( n65241, n73711, n65017 );
nor U122790 ( n65242, n73701, n65016 );
nor U122791 ( n30992, n30996, n30997 );
nor U122792 ( n30996, n74134, n30815 );
nor U122793 ( n30997, n74122, n30814 );
nor U122794 ( n31035, n31039, n31040 );
nor U122795 ( n31039, n74025, n30815 );
nor U122796 ( n31040, n74021, n30814 );
nor U122797 ( n65279, n65283, n65284 );
nor U122798 ( n65283, n73590, n65017 );
nor U122799 ( n65284, n73583, n65016 );
nor U122800 ( n10489, n10490, n10492 );
nor U122801 ( n10490, n74254, n10309 );
nor U122802 ( n10492, n74249, n10308 );
nor U122803 ( n44315, n44316, n44317 );
nor U122804 ( n44316, n73819, n44171 );
nor U122805 ( n44317, n73814, n44170 );
nor U122806 ( n23649, n23653, n23654 );
nor U122807 ( n23653, n73869, n23508 );
nor U122808 ( n23654, n73847, n23507 );
nor U122809 ( n23693, n23697, n23698 );
nor U122810 ( n23697, n73786, n23508 );
nor U122811 ( n23698, n73765, n23507 );
nor U122812 ( n23738, n23742, n23743 );
nor U122813 ( n23742, n73718, n23508 );
nor U122814 ( n23743, n73706, n23507 );
nor U122815 ( n23604, n23608, n23609 );
nor U122816 ( n23608, n73937, n23508 );
nor U122817 ( n23609, n73916, n23507 );
nor U122818 ( n23560, n23564, n23565 );
nor U122819 ( n23564, n74110, n23508 );
nor U122820 ( n23565, n74070, n23507 );
nor U122821 ( n56726, n56730, n56731 );
nor U122822 ( n56730, n73938, n56630 );
nor U122823 ( n56731, n73917, n56629 );
nor U122824 ( n56771, n56775, n56776 );
nor U122825 ( n56775, n73870, n56630 );
nor U122826 ( n56776, n73848, n56629 );
nor U122827 ( n56682, n56686, n56687 );
nor U122828 ( n56686, n74109, n56630 );
nor U122829 ( n56687, n74069, n56629 );
nor U122830 ( n56815, n56819, n56820 );
nor U122831 ( n56819, n73787, n56630 );
nor U122832 ( n56820, n73766, n56629 );
nor U122833 ( n56860, n56864, n56865 );
nor U122834 ( n56864, n73717, n56630 );
nor U122835 ( n56865, n73705, n56629 );
nor U122836 ( n23782, n23786, n23787 );
nor U122837 ( n23786, n73609, n23508 );
nor U122838 ( n23787, n73598, n23507 );
nor U122839 ( n56907, n56911, n56912 );
nor U122840 ( n56911, n73608, n56630 );
nor U122841 ( n56912, n73597, n56629 );
nor U122842 ( n10488, n10493, n10494 );
nor U122843 ( n10493, n74252, n10314 );
nor U122844 ( n10494, n74245, n10313 );
nor U122845 ( n44314, n44318, n44319 );
nor U122846 ( n44318, n73817, n44175 );
nor U122847 ( n44319, n73810, n44174 );
nand U122848 ( n32421, n32422, n76464 );
nor U122849 ( n30543, n74270, n30475 );
nor U122850 ( n9984, n74289, n9887 );
nor U122851 ( n64702, n73927, n64634 );
nor U122852 ( n43904, n73888, n43791 );
nand U122853 ( n30539, n30540, n30541 );
nor U122854 ( n30540, n30544, n30545 );
nor U122855 ( n30541, n30542, n30543 );
nor U122856 ( n30544, n74275, n30470 );
nand U122857 ( n9979, n9980, n9982 );
nor U122858 ( n9980, n9985, n9987 );
nor U122859 ( n9982, n9983, n9984 );
nor U122860 ( n9985, n74287, n9880 );
nand U122861 ( n64698, n64699, n64700 );
nor U122862 ( n64699, n64703, n64704 );
nor U122863 ( n64700, n64701, n64702 );
nor U122864 ( n64703, n73936, n64629 );
nand U122865 ( n43900, n43901, n43902 );
nor U122866 ( n43901, n43905, n43906 );
nor U122867 ( n43902, n43903, n43904 );
nor U122868 ( n43905, n73891, n43786 );
nor U122869 ( n30549, n74261, n30465 );
nor U122870 ( n9992, n74286, n9874 );
nor U122871 ( n64708, n73904, n64624 );
nor U122872 ( n43910, n73881, n43781 );
nor U122873 ( n30542, n74277, n30474 );
nor U122874 ( n9983, n74293, n9885 );
nor U122875 ( n64701, n73942, n64633 );
nor U122876 ( n43903, n73893, n43790 );
nor U122877 ( n23223, n73928, n23144 );
nor U122878 ( n56344, n73929, n56265 );
nand U122879 ( n23219, n23220, n23221 );
nor U122880 ( n23220, n23224, n23225 );
nor U122881 ( n23221, n23222, n23223 );
nor U122882 ( n23224, n73937, n23139 );
nand U122883 ( n56340, n56341, n56342 );
nor U122884 ( n56341, n56345, n56346 );
nor U122885 ( n56342, n56343, n56344 );
nor U122886 ( n56345, n73938, n56260 );
or U122887 ( n30457, n75872, n75873 );
nor U122888 ( n75872, n30461, n74338 );
nor U122889 ( n75873, n30460, n74343 );
or U122890 ( n9864, n75874, n75875 );
nor U122891 ( n75874, n9869, n74357 );
nor U122892 ( n75875, n9868, n74364 );
or U122893 ( n64616, n75876, n75877 );
nor U122894 ( n75876, n64620, n74167 );
nor U122895 ( n75877, n64619, n74180 );
or U122896 ( n43773, n75878, n75879 );
nor U122897 ( n75878, n43777, n74106 );
nor U122898 ( n75879, n43776, n74135 );
nor U122899 ( n23229, n73905, n23134 );
nor U122900 ( n56350, n73906, n56255 );
nor U122901 ( n23222, n73943, n23143 );
nor U122902 ( n56343, n73944, n56264 );
or U122903 ( n9863, n75880, n75881 );
nor U122904 ( n75880, n9874, n74359 );
nor U122905 ( n75881, n9873, n74367 );
or U122906 ( n30456, n75882, n75883 );
nor U122907 ( n75882, n30465, n74339 );
nor U122908 ( n75883, n30464, n74345 );
or U122909 ( n64615, n75884, n75885 );
nor U122910 ( n75884, n64624, n74171 );
nor U122911 ( n75885, n64623, n74186 );
or U122912 ( n43772, n75886, n75887 );
nor U122913 ( n75886, n43781, n74130 );
nor U122914 ( n75887, n43780, n74141 );
nor U122915 ( n30545, n74265, n30471 );
nor U122916 ( n9987, n74283, n9882 );
nor U122917 ( n64704, n73913, n64630 );
nor U122918 ( n43906, n73884, n43787 );
or U122919 ( n23126, n75888, n75889 );
nor U122920 ( n75888, n23130, n74168 );
nor U122921 ( n75889, n23129, n74182 );
or U122922 ( n56247, n75890, n75891 );
nor U122923 ( n75890, n56251, n74169 );
nor U122924 ( n75891, n56250, n74183 );
or U122925 ( n23125, n75892, n75893 );
nor U122926 ( n75892, n23134, n74172 );
nor U122927 ( n75893, n23133, n74187 );
or U122928 ( n56246, n75894, n75895 );
nor U122929 ( n75894, n56255, n74173 );
nor U122930 ( n75895, n56254, n74188 );
nor U122931 ( n23225, n73916, n23140 );
nor U122932 ( n56346, n73917, n56261 );
nand U122933 ( n15904, n15822, n15910 );
nand U122934 ( n15910, n15804, n15053 );
nor U122935 ( n30516, n74308, n30449 );
nor U122936 ( n9943, n74325, n9854 );
nor U122937 ( n64675, n74074, n64608 );
nor U122938 ( n43836, n73973, n43765 );
nand U122939 ( n30510, n30511, n30512 );
nor U122940 ( n30512, n30513, n30514 );
nor U122941 ( n30511, n30515, n30516 );
nor U122942 ( n30513, n74317, n30452 );
nand U122943 ( n9935, n9937, n9938 );
nor U122944 ( n9938, n9939, n9940 );
nor U122945 ( n9937, n9942, n9943 );
nor U122946 ( n9939, n74334, n9858 );
nand U122947 ( n64669, n64670, n64671 );
nor U122948 ( n64671, n64672, n64673 );
nor U122949 ( n64670, n64674, n64675 );
nor U122950 ( n64672, n74118, n64611 );
nand U122951 ( n43830, n43831, n43832 );
nor U122952 ( n43832, n43833, n43834 );
nor U122953 ( n43831, n43835, n43836 );
nor U122954 ( n43833, n73996, n43768 );
nor U122955 ( n23192, n74078, n23118 );
nor U122956 ( n56313, n74077, n56239 );
nand U122957 ( n23186, n23187, n23188 );
nor U122958 ( n23188, n23189, n23190 );
nor U122959 ( n23187, n23191, n23192 );
nor U122960 ( n23189, n74120, n23121 );
nand U122961 ( n56307, n56308, n56309 );
nor U122962 ( n56309, n56310, n56311 );
nor U122963 ( n56308, n56312, n56313 );
nor U122964 ( n56310, n74119, n56242 );
nor U122965 ( n30514, n74312, n30453 );
nor U122966 ( n9940, n74331, n9859 );
nor U122967 ( n64673, n74094, n64612 );
nor U122968 ( n43834, n73977, n43769 );
nor U122969 ( n23190, n74096, n23122 );
nor U122970 ( n56311, n74095, n56243 );
nand U122971 ( n15492, n15407, n15498 );
nand U122972 ( n15498, n15053, n5192 );
nand U122973 ( n54707, n8209, n74684 );
nand U122974 ( n21668, n8209, n74713 );
nand U122975 ( n28979, n8209, n74691 );
nand U122976 ( n36152, n8209, n73192 );
nor U122977 ( n23850, n73658, n23513 );
nor U122978 ( n56974, n73657, n56635 );
nand U122979 ( n23829, n23847, n23848 );
nor U122980 ( n23847, n23852, n23853 );
nor U122981 ( n23848, n23849, n23850 );
nor U122982 ( n23852, n73669, n23518 );
nand U122983 ( n56953, n56971, n56972 );
nor U122984 ( n56971, n56976, n56977 );
nor U122985 ( n56972, n56973, n56974 );
nor U122986 ( n56976, n73668, n56640 );
nor U122987 ( n30515, n74315, n30448 );
nor U122988 ( n9942, n74329, n9853 );
nor U122989 ( n64674, n74112, n64607 );
nor U122990 ( n43835, n73993, n43764 );
nor U122991 ( n23191, n74114, n23117 );
nor U122992 ( n56312, n74113, n56238 );
nor U122993 ( n23853, n73641, n23517 );
nor U122994 ( n56977, n73642, n56639 );
nand U122995 ( n48973, n48892, n48978 );
nand U122996 ( n48978, n48878, n48233 );
nor U122997 ( n30518, n30519, n30520 );
nor U122998 ( n30519, n74311, n30442 );
nor U122999 ( n30520, n74304, n30443 );
nor U123000 ( n9945, n9947, n9948 );
nor U123001 ( n9947, n74332, n9845 );
nor U123002 ( n9948, n74333, n9847 );
nor U123003 ( n64677, n64678, n64679 );
nor U123004 ( n64678, n74090, n64601 );
nor U123005 ( n64679, n74056, n64602 );
nor U123006 ( n43838, n43839, n43840 );
nor U123007 ( n43839, n73976, n43758 );
nor U123008 ( n43840, n73968, n43759 );
nor U123009 ( n23194, n23195, n23196 );
nor U123010 ( n23195, n74092, n23111 );
nor U123011 ( n23196, n74058, n23112 );
nor U123012 ( n56315, n56316, n56317 );
nor U123013 ( n56316, n74091, n56232 );
nor U123014 ( n56317, n74057, n56233 );
nor U123015 ( n30517, n30521, n30522 );
nor U123016 ( n30521, n74307, n30438 );
nor U123017 ( n30522, n74302, n30439 );
nor U123018 ( n9944, n9949, n9950 );
nor U123019 ( n9949, n74327, n9840 );
nor U123020 ( n9950, n74322, n9842 );
nor U123021 ( n64676, n64680, n64681 );
nor U123022 ( n64680, n74073, n64597 );
nor U123023 ( n64681, n74049, n64598 );
nor U123024 ( n43837, n43841, n43842 );
nor U123025 ( n43841, n73972, n43754 );
nor U123026 ( n43842, n73966, n43755 );
nor U123027 ( n70962, n73263, n70876 );
nor U123028 ( n70958, n74900, n70876 );
nor U123029 ( n70954, n74884, n70876 );
nor U123030 ( n70950, n73249, n70876 );
nor U123031 ( n70946, n74840, n70876 );
nor U123032 ( n70942, n74830, n70876 );
nor U123033 ( n70938, n73236, n70876 );
nor U123034 ( n70934, n74800, n70876 );
nor U123035 ( n70930, n74790, n70876 );
nor U123036 ( n70926, n74745, n70876 );
nor U123037 ( n70922, n73216, n70876 );
nor U123038 ( n70918, n74749, n70876 );
nor U123039 ( n70914, n72966, n70876 );
nor U123040 ( n70910, n74711, n70876 );
nor U123041 ( n70906, n73193, n70876 );
nor U123042 ( n70902, n74642, n70876 );
nor U123043 ( n70898, n73168, n70876 );
nor U123044 ( n70894, n74621, n70876 );
nor U123045 ( n70890, n73163, n70876 );
nand U123046 ( n48608, n48531, n48613 );
nand U123047 ( n48613, n48233, n7847 );
nor U123048 ( n23193, n23197, n23198 );
nor U123049 ( n23197, n74076, n23107 );
nor U123050 ( n23198, n74051, n23108 );
nor U123051 ( n56314, n56318, n56319 );
nor U123052 ( n56318, n74075, n56228 );
nor U123053 ( n56319, n74050, n56229 );
nor U123054 ( n23849, n73683, n23514 );
nor U123055 ( n56973, n73682, n56636 );
nor U123056 ( n23832, n23833, n23834 );
nor U123057 ( n23833, n73700, n23504 );
nor U123058 ( n23834, n73685, n23503 );
nor U123059 ( n56956, n56957, n56958 );
nor U123060 ( n56957, n73699, n56626 );
nor U123061 ( n56958, n73684, n56625 );
not U123062 ( n1774, n48566 );
nor U123063 ( n40785, n76925, n75248 );
nor U123064 ( n41007, n76925, n72954 );
nor U123065 ( n41450, n76925, n72943 );
nor U123066 ( n41115, n76925, n72939 );
nor U123067 ( n41146, n76925, n72937 );
nor U123068 ( n41055, n76925, n72931 );
nor U123069 ( n40692, n76925, n72929 );
nor U123070 ( n40985, n76925, n74170 );
nor U123071 ( n41179, n76925, n72955 );
nor U123072 ( n40968, n76925, n72946 );
nor U123073 ( n40728, n76925, n72949 );
nor U123074 ( n40931, n76925, n72942 );
nor U123075 ( n40761, n76925, n72935 );
nor U123076 ( n40865, n76925, n72936 );
nor U123077 ( n41199, n76925, n74256 );
nor U123078 ( n23831, n23841, n23842 );
nor U123079 ( n23841, n73694, n23508 );
nor U123080 ( n23842, n73673, n23507 );
nor U123081 ( n56955, n56965, n56966 );
nor U123082 ( n56965, n73693, n56630 );
nor U123083 ( n56966, n73672, n56629 );
nor U123084 ( n36247, n73264, n36167 );
nor U123085 ( n36243, n74901, n36167 );
nor U123086 ( n36239, n74885, n36167 );
nor U123087 ( n36235, n73250, n36167 );
nor U123088 ( n36231, n74839, n36167 );
nor U123089 ( n36227, n74829, n36167 );
nor U123090 ( n36223, n73235, n36167 );
nor U123091 ( n36217, n74801, n36167 );
nor U123092 ( n36213, n74791, n36167 );
nor U123093 ( n36209, n74746, n36167 );
nor U123094 ( n36205, n73217, n36167 );
nor U123095 ( n36201, n74750, n36167 );
nor U123096 ( n36197, n72967, n36167 );
nor U123097 ( n36193, n74712, n36167 );
nor U123098 ( n36189, n73194, n36167 );
nor U123099 ( n36185, n74643, n36167 );
nor U123100 ( n36181, n73169, n36167 );
nor U123101 ( n36175, n74622, n36167 );
nor U123102 ( n36171, n73164, n36167 );
nor U123103 ( n14849, n14823, n14854 );
nor U123104 ( n48047, n48026, n48051 );
not U123105 ( n2890, n38332 );
or U123106 ( n54708, n73177, n54699 );
or U123107 ( n28980, n73179, n28971 );
or U123108 ( n36153, n74654, n36144 );
or U123109 ( n21669, n73185, n21660 );
and U123110 ( n16220, n15273, n15272 );
nand U123111 ( n49337, n49276, n49342 );
nand U123112 ( n49342, n49247, n48233 );
nor U123113 ( n41037, n76925, n74064 );
nor U123114 ( n14863, n14823, n14868 );
nor U123115 ( n48058, n48026, n48062 );
nor U123116 ( n14835, n14823, n14840 );
nor U123117 ( n48036, n48026, n48040 );
nor U123118 ( n11165, n11169, n5147 );
nor U123119 ( n44879, n44882, n7802 );
nor U123120 ( n31494, n31497, n3399 );
nor U123121 ( n65744, n65747, n6014 );
nor U123122 ( n31189, n74341, n31190 );
nor U123123 ( n31246, n74304, n31190 );
nor U123124 ( n31290, n74262, n31190 );
nor U123125 ( n31331, n74224, n31190 );
nor U123126 ( n31371, n74107, n31190 );
nor U123127 ( n10864, n74333, n10797 );
nor U123128 ( n10914, n74297, n10797 );
nor U123129 ( n10965, n74243, n10797 );
nor U123130 ( n11014, n74143, n10797 );
nor U123131 ( n11064, n74111, n10797 );
nor U123132 ( n11115, n73998, n10797 );
nor U123133 ( n11164, n74019, n10797 );
nor U123134 ( n65500, n74056, n65444 );
nor U123135 ( n65540, n73907, n65444 );
nor U123136 ( n65581, n73840, n65444 );
nor U123137 ( n65621, n73758, n65444 );
nor U123138 ( n44664, n73882, n44570 );
nor U123139 ( n44705, n73808, n44570 );
nor U123140 ( n44744, n73640, n44570 );
nor U123141 ( n44784, n73611, n44570 );
nor U123142 ( n44878, n73556, n44570 );
nor U123143 ( n44825, n73552, n44570 );
nor U123144 ( n44624, n73968, n44570 );
nor U123145 ( n10795, n74361, n10797 );
nor U123146 ( n65443, n74177, n65444 );
nor U123147 ( n44569, n74132, n44570 );
nor U123148 ( n31412, n74048, n31190 );
nor U123149 ( n31452, n73969, n31190 );
nor U123150 ( n31493, n74002, n31190 );
nor U123151 ( n65662, n73746, n65444 );
nor U123152 ( n65702, n73628, n65444 );
nor U123153 ( n65743, n73659, n65444 );
nand U123154 ( n31185, n31186, n31187 );
nor U123155 ( n31186, n31192, n31193 );
nor U123156 ( n31187, n31188, n31189 );
nor U123157 ( n31192, n74347, n31195 );
nand U123158 ( n31242, n31243, n31244 );
nor U123159 ( n31243, n31247, n31248 );
nor U123160 ( n31244, n31245, n31246 );
nor U123161 ( n31247, n74307, n31195 );
nand U123162 ( n31286, n31287, n31288 );
nor U123163 ( n31287, n31291, n31292 );
nor U123164 ( n31288, n31289, n31290 );
nor U123165 ( n31291, n74267, n31195 );
nand U123166 ( n31327, n31328, n31329 );
nor U123167 ( n31328, n31332, n31333 );
nor U123168 ( n31329, n31330, n31331 );
nor U123169 ( n31332, n74228, n31195 );
nand U123170 ( n31367, n31368, n31369 );
nor U123171 ( n31368, n31372, n31373 );
nor U123172 ( n31369, n31370, n31371 );
nor U123173 ( n31372, n74124, n31195 );
nand U123174 ( n10859, n10860, n10862 );
nor U123175 ( n10860, n10865, n10867 );
nor U123176 ( n10862, n10863, n10864 );
nor U123177 ( n10865, n74327, n10803 );
nand U123178 ( n10909, n10910, n10912 );
nor U123179 ( n10910, n10915, n10917 );
nor U123180 ( n10912, n10913, n10914 );
nor U123181 ( n10915, n74290, n10803 );
nand U123182 ( n10960, n10962, n10963 );
nor U123183 ( n10962, n10967, n10968 );
nor U123184 ( n10963, n10964, n10965 );
nor U123185 ( n10967, n74246, n10803 );
nand U123186 ( n11009, n11010, n11012 );
nor U123187 ( n11010, n11015, n11017 );
nor U123188 ( n11012, n11013, n11014 );
nor U123189 ( n11015, n74152, n10803 );
nand U123190 ( n11059, n11060, n11062 );
nor U123191 ( n11060, n11065, n11067 );
nor U123192 ( n11062, n11063, n11064 );
nor U123193 ( n11065, n74093, n10803 );
nand U123194 ( n11110, n11112, n11113 );
nor U123195 ( n11112, n11117, n11118 );
nor U123196 ( n11113, n11114, n11115 );
nor U123197 ( n11117, n73985, n10803 );
nand U123198 ( n11159, n11160, n11162 );
nor U123199 ( n11160, n11167, n11168 );
nor U123200 ( n11162, n11163, n11164 );
nor U123201 ( n11167, n74035, n10803 );
nand U123202 ( n65496, n65497, n65498 );
nor U123203 ( n65497, n65501, n65502 );
nor U123204 ( n65498, n65499, n65500 );
nor U123205 ( n65501, n74073, n65449 );
nand U123206 ( n65536, n65537, n65538 );
nor U123207 ( n65537, n65541, n65542 );
nor U123208 ( n65538, n65539, n65540 );
nor U123209 ( n65541, n73918, n65449 );
nand U123210 ( n65577, n65578, n65579 );
nor U123211 ( n65578, n65582, n65583 );
nor U123212 ( n65579, n65580, n65581 );
nor U123213 ( n65582, n73849, n65449 );
nand U123214 ( n65617, n65618, n65619 );
nor U123215 ( n65618, n65622, n65623 );
nor U123216 ( n65619, n65620, n65621 );
nor U123217 ( n65622, n73767, n65449 );
nand U123218 ( n44660, n44661, n44662 );
nor U123219 ( n44661, n44665, n44666 );
nor U123220 ( n44662, n44663, n44664 );
nor U123221 ( n44665, n73885, n44575 );
nand U123222 ( n44701, n44702, n44703 );
nor U123223 ( n44702, n44706, n44707 );
nor U123224 ( n44703, n44704, n44705 );
nor U123225 ( n44706, n73811, n44575 );
nand U123226 ( n44740, n44741, n44742 );
nor U123227 ( n44741, n44745, n44746 );
nor U123228 ( n44742, n44743, n44744 );
nor U123229 ( n44745, n73646, n44575 );
nand U123230 ( n44780, n44781, n44782 );
nor U123231 ( n44781, n44785, n44786 );
nor U123232 ( n44782, n44783, n44784 );
nor U123233 ( n44785, n73582, n44575 );
nand U123234 ( n44874, n44875, n44876 );
nor U123235 ( n44875, n44880, n44881 );
nor U123236 ( n44876, n44877, n44878 );
nor U123237 ( n44880, n73560, n44575 );
nand U123238 ( n44821, n44822, n44823 );
nor U123239 ( n44822, n44826, n44827 );
nor U123240 ( n44823, n44824, n44825 );
nor U123241 ( n44826, n73543, n44575 );
nand U123242 ( n44620, n44621, n44622 );
nor U123243 ( n44621, n44625, n44626 );
nor U123244 ( n44622, n44623, n44624 );
nor U123245 ( n44625, n73972, n44575 );
nand U123246 ( n10790, n10792, n10793 );
nor U123247 ( n10792, n10799, n10800 );
nor U123248 ( n10793, n10794, n10795 );
nor U123249 ( n10799, n74370, n10803 );
nand U123250 ( n65439, n65440, n65441 );
nor U123251 ( n65440, n65446, n65447 );
nor U123252 ( n65441, n65442, n65443 );
nor U123253 ( n65446, n74189, n65449 );
nand U123254 ( n44565, n44566, n44567 );
nor U123255 ( n44566, n44572, n44573 );
nor U123256 ( n44567, n44568, n44569 );
nor U123257 ( n44572, n74144, n44575 );
nand U123258 ( n31408, n31409, n31410 );
nor U123259 ( n31409, n31413, n31414 );
nor U123260 ( n31410, n31411, n31412 );
nor U123261 ( n31413, n74033, n31195 );
nand U123262 ( n31448, n31449, n31450 );
nor U123263 ( n31449, n31453, n31454 );
nor U123264 ( n31450, n31451, n31452 );
nor U123265 ( n31453, n73958, n31195 );
nand U123266 ( n31489, n31490, n31491 );
nor U123267 ( n31490, n31495, n31496 );
nor U123268 ( n31491, n31492, n31493 );
nor U123269 ( n31495, n74006, n31195 );
nand U123270 ( n65658, n65659, n65660 );
nor U123271 ( n65659, n65663, n65664 );
nor U123272 ( n65660, n65661, n65662 );
nor U123273 ( n65663, n73725, n65449 );
nand U123274 ( n65698, n65699, n65700 );
nor U123275 ( n65699, n65703, n65704 );
nor U123276 ( n65700, n65701, n65702 );
nor U123277 ( n65703, n73595, n65449 );
nand U123278 ( n65739, n65740, n65741 );
nor U123279 ( n65740, n65745, n65746 );
nor U123280 ( n65741, n65742, n65743 );
nor U123281 ( n65745, n73674, n65449 );
nor U123282 ( n14877, n14823, n14882 );
nor U123283 ( n48083, n48026, n48087 );
nand U123284 ( n48226, n48155, n48232 );
nand U123285 ( n48232, n48233, n48131 );
nor U123286 ( n14890, n14823, n14895 );
nor U123287 ( n48094, n48026, n48098 );
nor U123288 ( n31193, n74340, n31194 );
nor U123289 ( n31248, n74302, n31194 );
nor U123290 ( n31292, n74260, n31194 );
nor U123291 ( n31333, n74222, n31194 );
nor U123292 ( n31373, n74102, n31194 );
nor U123293 ( n10867, n74322, n10802 );
nor U123294 ( n10917, n74285, n10802 );
nor U123295 ( n10968, n74240, n10802 );
nor U123296 ( n11017, n74139, n10802 );
nor U123297 ( n11067, n74082, n10802 );
nor U123298 ( n11118, n73980, n10802 );
nor U123299 ( n11168, n74016, n10802 );
nor U123300 ( n65502, n74049, n65448 );
nor U123301 ( n65542, n73901, n65448 );
nor U123302 ( n65583, n73834, n65448 );
nor U123303 ( n65623, n73752, n65448 );
nor U123304 ( n44666, n73880, n44574 );
nor U123305 ( n44707, n73806, n44574 );
nor U123306 ( n44746, n73638, n44574 );
nor U123307 ( n44786, n73576, n44574 );
nor U123308 ( n44881, n73554, n44574 );
nor U123309 ( n44827, n73538, n44574 );
nor U123310 ( n44626, n73966, n44574 );
nor U123311 ( n10800, n74362, n10802 );
nor U123312 ( n65447, n74174, n65448 );
nor U123313 ( n44573, n74133, n44574 );
nor U123314 ( n31414, n74023, n31194 );
nor U123315 ( n31454, n73953, n31194 );
nor U123316 ( n31496, n74000, n31194 );
nor U123317 ( n65664, n73710, n65448 );
nor U123318 ( n65704, n73588, n65448 );
nor U123319 ( n65746, n73652, n65448 );
nor U123320 ( n14815, n14823, n14824 );
nor U123321 ( n48020, n48026, n48027 );
nor U123322 ( n14904, n14823, n14909 );
nor U123323 ( n48105, n48026, n48109 );
not U123324 ( n1834, n10118 );
nand U123325 ( n47980, n76175, n74626 );
nand U123326 ( n14759, n76185, n74646 );
and U123327 ( n49247, n48413, n48412 );
nor U123328 ( n31188, n74350, n31191 );
nor U123329 ( n31245, n74311, n31191 );
nor U123330 ( n31289, n74271, n31191 );
nor U123331 ( n31330, n74233, n31191 );
nor U123332 ( n31370, n74129, n31191 );
nor U123333 ( n10863, n74332, n10798 );
nor U123334 ( n10913, n74295, n10798 );
nor U123335 ( n10964, n74250, n10798 );
nor U123336 ( n11013, n74156, n10798 );
nor U123337 ( n11063, n74101, n10798 );
nor U123338 ( n11114, n73992, n10798 );
nor U123339 ( n11163, n74043, n10798 );
nor U123340 ( n65499, n74090, n65445 );
nor U123341 ( n65539, n73930, n65445 );
nor U123342 ( n65580, n73861, n65445 );
nor U123343 ( n65620, n73779, n65445 );
nor U123344 ( n44663, n73889, n44571 );
nor U123345 ( n44704, n73815, n44571 );
nor U123346 ( n44743, n73650, n44571 );
nor U123347 ( n44783, n73593, n44571 );
nor U123348 ( n44877, n73565, n44571 );
nor U123349 ( n44824, n73549, n44571 );
nor U123350 ( n44623, n73976, n44571 );
nor U123351 ( n10794, n74376, n10798 );
nor U123352 ( n65442, n74199, n65445 );
nor U123353 ( n44568, n74147, n44571 );
nor U123354 ( n31411, n74044, n31191 );
nor U123355 ( n31451, n73963, n31191 );
nor U123356 ( n31492, n74010, n31191 );
nor U123357 ( n65661, n73740, n65445 );
nor U123358 ( n65701, n73612, n65445 );
nor U123359 ( n65742, n73686, n65445 );
nand U123360 ( n48227, n7452, n47918 );
not U123361 ( n7452, n48133 );
nand U123362 ( n47945, n7454, n74907 );
nand U123363 ( n43346, n74907, n42384 );
nand U123364 ( n22753, n74888, n21858 );
nand U123365 ( n55867, n74890, n54949 );
not U123366 ( n7413, n47901 );
nand U123367 ( n15045, n4808, n14715 );
not U123368 ( n4808, n14947 );
nand U123369 ( n14729, n4810, n74906 );
nor U123370 ( n14955, n4807, n15389 );
not U123371 ( n4807, n15045 );
nor U123372 ( n30432, n30444, n30445 );
nand U123373 ( n30444, n30450, n30451 );
nand U123374 ( n30445, n30446, n30447 );
or U123375 ( n30450, n30453, n74351 );
nor U123376 ( n9833, n9848, n9849 );
nand U123377 ( n9848, n9855, n9857 );
nand U123378 ( n9849, n9850, n9852 );
or U123379 ( n9855, n9859, n74375 );
nor U123380 ( n64591, n64603, n64604 );
nand U123381 ( n64603, n64609, n64610 );
nand U123382 ( n64604, n64605, n64606 );
or U123383 ( n64609, n64612, n74202 );
nor U123384 ( n43748, n43760, n43761 );
nand U123385 ( n43760, n43766, n43767 );
nand U123386 ( n43761, n43762, n43763 );
or U123387 ( n43766, n43769, n74148 );
or U123388 ( n30447, n30448, n74353 );
or U123389 ( n9852, n9853, n74373 );
or U123390 ( n64606, n64607, n74208 );
or U123391 ( n43763, n43764, n74158 );
nor U123392 ( n23101, n23113, n23114 );
nand U123393 ( n23113, n23119, n23120 );
nand U123394 ( n23114, n23115, n23116 );
or U123395 ( n23119, n23122, n74203 );
nor U123396 ( n56222, n56234, n56235 );
nand U123397 ( n56234, n56240, n56241 );
nand U123398 ( n56235, n56236, n56237 );
or U123399 ( n56240, n56243, n74204 );
or U123400 ( n23116, n23117, n74209 );
or U123401 ( n56237, n56238, n74210 );
nor U123402 ( n30433, n30434, n30435 );
nand U123403 ( n30434, n30440, n30441 );
nand U123404 ( n30435, n30436, n30437 );
or U123405 ( n30440, n30443, n74341 );
nor U123406 ( n9834, n9835, n9837 );
nand U123407 ( n9835, n9843, n9844 );
nand U123408 ( n9837, n9838, n9839 );
or U123409 ( n9843, n9847, n74361 );
nor U123410 ( n64592, n64593, n64594 );
nand U123411 ( n64593, n64599, n64600 );
nand U123412 ( n64594, n64595, n64596 );
or U123413 ( n64599, n64602, n74177 );
nor U123414 ( n43749, n43750, n43751 );
nand U123415 ( n43750, n43756, n43757 );
nand U123416 ( n43751, n43752, n43753 );
or U123417 ( n43756, n43759, n74132 );
or U123418 ( n30437, n30438, n74347 );
or U123419 ( n9839, n9840, n74370 );
or U123420 ( n64596, n64597, n74189 );
or U123421 ( n43753, n43754, n74144 );
nand U123422 ( n9399, n74906, n8297 );
or U123423 ( n30446, n30449, n74348 );
or U123424 ( n9850, n9854, n74368 );
or U123425 ( n64605, n64608, n74192 );
or U123426 ( n43762, n43765, n74145 );
nor U123427 ( n23102, n23103, n23104 );
nand U123428 ( n23103, n23109, n23110 );
nand U123429 ( n23104, n23105, n23106 );
or U123430 ( n23109, n23112, n74178 );
nor U123431 ( n56223, n56224, n56225 );
nand U123432 ( n56224, n56230, n56231 );
nand U123433 ( n56225, n56226, n56227 );
or U123434 ( n56230, n56233, n74179 );
or U123435 ( n23106, n23107, n74190 );
or U123436 ( n56227, n56228, n74191 );
nor U123437 ( n66677, n66661, n66678 );
nor U123438 ( n32074, n32058, n32075 );
nor U123439 ( n24842, n24826, n24843 );
nor U123440 ( n57976, n57960, n57977 );
or U123441 ( n23115, n23118, n74193 );
or U123442 ( n56236, n56239, n74194 );
nor U123443 ( n12023, n12003, n12024 );
nor U123444 ( n45769, n45735, n45770 );
or U123445 ( n30436, n30439, n74340 );
or U123446 ( n9838, n9842, n74362 );
or U123447 ( n64595, n64598, n74174 );
or U123448 ( n43752, n43755, n74133 );
not U123449 ( n5582, n70876 );
or U123450 ( n23105, n23108, n74175 );
or U123451 ( n56226, n56229, n74176 );
or U123452 ( n30451, n30452, n74355 );
or U123453 ( n9857, n9858, n74377 );
or U123454 ( n64610, n64611, n74214 );
or U123455 ( n43767, n43768, n74160 );
nand U123456 ( n44580, n44887, n7802 );
nor U123457 ( n44887, n44882, n43330 );
nand U123458 ( n31200, n31502, n3399 );
nor U123459 ( n31502, n31497, n30059 );
nand U123460 ( n65454, n65752, n6014 );
nor U123461 ( n65752, n65747, n64076 );
nor U123462 ( n31199, n74351, n31200 );
nor U123463 ( n31252, n74312, n31200 );
nor U123464 ( n31296, n74272, n31200 );
nor U123465 ( n31337, n74235, n31200 );
nor U123466 ( n31377, n74131, n31200 );
nor U123467 ( n10872, n74331, n10809 );
nor U123468 ( n10922, n74294, n10809 );
nor U123469 ( n10973, n74251, n10809 );
nor U123470 ( n11022, n74157, n10809 );
nor U123471 ( n11072, n74100, n10809 );
nor U123472 ( n11123, n73991, n10809 );
nor U123473 ( n11174, n74045, n10809 );
nor U123474 ( n65506, n74094, n65454 );
nor U123475 ( n65546, n73933, n65454 );
nor U123476 ( n65587, n73864, n65454 );
nor U123477 ( n65627, n73782, n65454 );
nor U123478 ( n44670, n73890, n44580 );
nor U123479 ( n44711, n73816, n44580 );
nor U123480 ( n44750, n73651, n44580 );
nor U123481 ( n44790, n73591, n44580 );
nor U123482 ( n44886, n73567, n44580 );
nor U123483 ( n44831, n73548, n44580 );
nor U123484 ( n44630, n73977, n44580 );
nor U123485 ( n10808, n74375, n10809 );
nor U123486 ( n65453, n74202, n65454 );
nor U123487 ( n44579, n74148, n44580 );
nor U123488 ( n31418, n74042, n31200 );
nor U123489 ( n31458, n73962, n31200 );
nor U123490 ( n31501, n74011, n31200 );
nor U123491 ( n65668, n73737, n65454 );
nor U123492 ( n65708, n73610, n65454 );
nor U123493 ( n65751, n73687, n65454 );
nand U123494 ( n10809, n11175, n5147 );
nor U123495 ( n11175, n11169, n9380 );
nand U123496 ( n31184, n31196, n31197 );
nor U123497 ( n31196, n31202, n31203 );
nor U123498 ( n31197, n31198, n31199 );
nor U123499 ( n31202, n74353, n31205 );
nand U123500 ( n31241, n31249, n31250 );
nor U123501 ( n31249, n31253, n31254 );
nor U123502 ( n31250, n31251, n31252 );
nor U123503 ( n31253, n74315, n31205 );
nand U123504 ( n31285, n31293, n31294 );
nor U123505 ( n31293, n31297, n31298 );
nor U123506 ( n31294, n31295, n31296 );
nor U123507 ( n31297, n74276, n31205 );
nand U123508 ( n31326, n31334, n31335 );
nor U123509 ( n31334, n31338, n31339 );
nor U123510 ( n31335, n31336, n31337 );
nor U123511 ( n31338, n74238, n31205 );
nand U123512 ( n31366, n31374, n31375 );
nor U123513 ( n31374, n31378, n31379 );
nor U123514 ( n31375, n31376, n31377 );
nor U123515 ( n31378, n74136, n31205 );
nand U123516 ( n10858, n10868, n10869 );
nor U123517 ( n10868, n10873, n10874 );
nor U123518 ( n10869, n10870, n10872 );
nor U123519 ( n10873, n74329, n10815 );
nand U123520 ( n10908, n10918, n10919 );
nor U123521 ( n10918, n10923, n10924 );
nor U123522 ( n10919, n10920, n10922 );
nor U123523 ( n10923, n74292, n10815 );
nand U123524 ( n10959, n10969, n10970 );
nor U123525 ( n10969, n10974, n10975 );
nor U123526 ( n10970, n10972, n10973 );
nor U123527 ( n10974, n74253, n10815 );
nand U123528 ( n11008, n11018, n11019 );
nor U123529 ( n11018, n11023, n11024 );
nor U123530 ( n11019, n11020, n11022 );
nor U123531 ( n11023, n74162, n10815 );
nand U123532 ( n11058, n11068, n11069 );
nor U123533 ( n11068, n11073, n11074 );
nor U123534 ( n11069, n11070, n11072 );
nor U123535 ( n11073, n74098, n10815 );
nand U123536 ( n11109, n11119, n11120 );
nor U123537 ( n11119, n11124, n11125 );
nor U123538 ( n11120, n11122, n11123 );
nor U123539 ( n11124, n73988, n10815 );
nand U123540 ( n11158, n11170, n11172 );
nor U123541 ( n11170, n11179, n11180 );
nor U123542 ( n11172, n11173, n11174 );
nor U123543 ( n11179, n74059, n10815 );
nand U123544 ( n65495, n65503, n65504 );
nor U123545 ( n65503, n65507, n65508 );
nor U123546 ( n65504, n65505, n65506 );
nor U123547 ( n65507, n74112, n65459 );
nand U123548 ( n65535, n65543, n65544 );
nor U123549 ( n65543, n65547, n65548 );
nor U123550 ( n65544, n65545, n65546 );
nor U123551 ( n65547, n73939, n65459 );
nand U123552 ( n65576, n65584, n65585 );
nor U123553 ( n65584, n65588, n65589 );
nor U123554 ( n65585, n65586, n65587 );
nor U123555 ( n65588, n73871, n65459 );
nand U123556 ( n65616, n65624, n65625 );
nor U123557 ( n65624, n65628, n65629 );
nor U123558 ( n65625, n65626, n65627 );
nor U123559 ( n65628, n73788, n65459 );
nand U123560 ( n44659, n44667, n44668 );
nor U123561 ( n44667, n44671, n44672 );
nor U123562 ( n44668, n44669, n44670 );
nor U123563 ( n44671, n73892, n44585 );
nand U123564 ( n44700, n44708, n44709 );
nor U123565 ( n44708, n44712, n44713 );
nor U123566 ( n44709, n44710, n44711 );
nor U123567 ( n44712, n73818, n44585 );
nand U123568 ( n44739, n44747, n44748 );
nor U123569 ( n44747, n44751, n44752 );
nor U123570 ( n44748, n44749, n44750 );
nor U123571 ( n44751, n73662, n44585 );
nand U123572 ( n44779, n44787, n44788 );
nor U123573 ( n44787, n44791, n44792 );
nor U123574 ( n44788, n44789, n44790 );
nor U123575 ( n44791, n73586, n44585 );
nand U123576 ( n44873, n44883, n44884 );
nor U123577 ( n44883, n44890, n44891 );
nor U123578 ( n44884, n44885, n44886 );
nor U123579 ( n44890, n73571, n44585 );
nand U123580 ( n44820, n44828, n44829 );
nor U123581 ( n44828, n44832, n44833 );
nor U123582 ( n44829, n44830, n44831 );
nor U123583 ( n44832, n73546, n44585 );
nand U123584 ( n44619, n44627, n44628 );
nor U123585 ( n44627, n44631, n44632 );
nor U123586 ( n44628, n44629, n44630 );
nor U123587 ( n44631, n73993, n44585 );
nand U123588 ( n10789, n10804, n10805 );
nor U123589 ( n10804, n10812, n10813 );
nor U123590 ( n10805, n10807, n10808 );
nor U123591 ( n10812, n74373, n10815 );
nand U123592 ( n65438, n65450, n65451 );
nor U123593 ( n65450, n65456, n65457 );
nor U123594 ( n65451, n65452, n65453 );
nor U123595 ( n65456, n74208, n65459 );
nand U123596 ( n44564, n44576, n44577 );
nor U123597 ( n44576, n44582, n44583 );
nor U123598 ( n44577, n44578, n44579 );
nor U123599 ( n44582, n74158, n44585 );
nand U123600 ( n31407, n31415, n31416 );
nor U123601 ( n31415, n31419, n31420 );
nor U123602 ( n31416, n31417, n31418 );
nor U123603 ( n31419, n74036, n31205 );
nand U123604 ( n31447, n31455, n31456 );
nor U123605 ( n31455, n31459, n31460 );
nor U123606 ( n31456, n31457, n31458 );
nor U123607 ( n31459, n73960, n31205 );
nand U123608 ( n31488, n31498, n31499 );
nor U123609 ( n31498, n31505, n31506 );
nor U123610 ( n31499, n31500, n31501 );
nor U123611 ( n31505, n74014, n31205 );
nand U123612 ( n65657, n65665, n65666 );
nor U123613 ( n65665, n65669, n65670 );
nor U123614 ( n65666, n65667, n65668 );
nor U123615 ( n65669, n73731, n65459 );
nand U123616 ( n65697, n65705, n65706 );
nor U123617 ( n65705, n65709, n65710 );
nor U123618 ( n65706, n65707, n65708 );
nor U123619 ( n65709, n73602, n65459 );
nand U123620 ( n65738, n65748, n65749 );
nor U123621 ( n65748, n65755, n65756 );
nor U123622 ( n65749, n65750, n65751 );
nor U123623 ( n65755, n73695, n65459 );
or U123624 ( n23120, n23121, n74215 );
or U123625 ( n56241, n56242, n74216 );
nor U123626 ( n47902, n47905, n74442 );
nor U123627 ( n47905, n7413, n46293 );
nor U123628 ( n12857, n72970, n74886 );
nor U123629 ( n57322, n57325, n6869 );
nor U123630 ( n24200, n24203, n4237 );
nor U123631 ( n23894, n74178, n23895 );
nor U123632 ( n57018, n74179, n57019 );
nand U123633 ( n23890, n23891, n23892 );
nor U123634 ( n23891, n23897, n23898 );
nor U123635 ( n23892, n23893, n23894 );
nor U123636 ( n23897, n74190, n23900 );
nand U123637 ( n57014, n57015, n57016 );
nor U123638 ( n57015, n57021, n57022 );
nor U123639 ( n57016, n57017, n57018 );
nor U123640 ( n57021, n74191, n57024 );
or U123641 ( n30441, n30442, n74350 );
or U123642 ( n9844, n9845, n74376 );
or U123643 ( n64600, n64601, n74199 );
or U123644 ( n43757, n43758, n74147 );
nand U123645 ( n10814, n11182, n5147 );
nor U123646 ( n11182, n11169, n9382 );
nand U123647 ( n44584, n44892, n7802 );
nor U123648 ( n44892, n44882, n43331 );
nand U123649 ( n31204, n31507, n3399 );
nor U123650 ( n31507, n31497, n30060 );
nand U123651 ( n65458, n65757, n6014 );
nor U123652 ( n65757, n65747, n64077 );
nor U123653 ( n14944, n15272, n15273 );
nor U123654 ( n31203, n74348, n31204 );
nor U123655 ( n31254, n74308, n31204 );
nor U123656 ( n31298, n74268, n31204 );
nor U123657 ( n31339, n74229, n31204 );
nor U123658 ( n31379, n74125, n31204 );
nor U123659 ( n10874, n74325, n10814 );
nor U123660 ( n10924, n74288, n10814 );
nor U123661 ( n10975, n74247, n10814 );
nor U123662 ( n11024, n74153, n10814 );
nor U123663 ( n11074, n74088, n10814 );
nor U123664 ( n11125, n73983, n10814 );
nor U123665 ( n11180, n74037, n10814 );
nor U123666 ( n65508, n74074, n65458 );
nor U123667 ( n65548, n73919, n65458 );
nor U123668 ( n65589, n73850, n65458 );
nor U123669 ( n65629, n73768, n65458 );
nor U123670 ( n44672, n73886, n44584 );
nor U123671 ( n44713, n73812, n44584 );
nor U123672 ( n44752, n73647, n44584 );
nor U123673 ( n44792, n73580, n44584 );
nor U123674 ( n44891, n73561, n44584 );
nor U123675 ( n44833, n73541, n44584 );
nor U123676 ( n44632, n73973, n44584 );
nor U123677 ( n10813, n74368, n10814 );
nor U123678 ( n65457, n74192, n65458 );
nor U123679 ( n44583, n74145, n44584 );
nor U123680 ( n31420, n74030, n31204 );
nor U123681 ( n31460, n73956, n31204 );
nor U123682 ( n31506, n74007, n31204 );
nor U123683 ( n65670, n73719, n65458 );
nor U123684 ( n65710, n73592, n65458 );
nor U123685 ( n65756, n73675, n65458 );
nand U123686 ( n15044, n14974, n15052 );
nand U123687 ( n15052, n15053, n14944 );
or U123688 ( n23110, n23111, n74200 );
or U123689 ( n56231, n56232, n74201 );
nand U123690 ( n15154, n15078, n15160 );
nand U123691 ( n15160, n15162, n14944 );
not U123692 ( n4769, n14675 );
nor U123693 ( n23898, n74175, n23899 );
nor U123694 ( n57022, n74176, n57023 );
nor U123695 ( n30500, n74310, n30475 );
nor U123696 ( n9923, n74326, n9887 );
nor U123697 ( n64659, n74083, n64634 );
nor U123698 ( n43820, n73975, n43791 );
nand U123699 ( n30496, n30497, n30498 );
nor U123700 ( n30497, n30501, n30502 );
nor U123701 ( n30498, n30499, n30500 );
nor U123702 ( n30501, n74313, n30470 );
nand U123703 ( n9918, n9919, n9920 );
nor U123704 ( n9919, n9924, n9925 );
nor U123705 ( n9920, n9922, n9923 );
nor U123706 ( n9924, n74324, n9880 );
nand U123707 ( n64655, n64656, n64657 );
nor U123708 ( n64656, n64660, n64661 );
nor U123709 ( n64657, n64658, n64659 );
nor U123710 ( n64660, n74108, n64629 );
nand U123711 ( n43816, n43817, n43818 );
nor U123712 ( n43817, n43821, n43822 );
nor U123713 ( n43818, n43819, n43820 );
nor U123714 ( n43821, n73990, n43786 );
nor U123715 ( n30506, n74303, n30465 );
nor U123716 ( n9930, n74323, n9874 );
nor U123717 ( n23176, n74087, n23144 );
nor U123718 ( n64665, n74053, n64624 );
nor U123719 ( n43826, n73967, n43781 );
nor U123720 ( n56297, n74086, n56265 );
nand U123721 ( n23172, n23173, n23174 );
nor U123722 ( n23173, n23177, n23178 );
nor U123723 ( n23174, n23175, n23176 );
nor U123724 ( n23177, n74110, n23139 );
nand U123725 ( n56293, n56294, n56295 );
nor U123726 ( n56294, n56298, n56299 );
nor U123727 ( n56295, n56296, n56297 );
nor U123728 ( n56298, n74109, n56260 );
not U123729 ( n2980, n36167 );
nor U123730 ( n30499, n74316, n30474 );
nor U123731 ( n9922, n74330, n9885 );
nor U123732 ( n64658, n74115, n64633 );
nor U123733 ( n43819, n73994, n43790 );
nor U123734 ( n23182, n74055, n23134 );
nor U123735 ( n56303, n74054, n56255 );
nor U123736 ( n23175, n74117, n23143 );
nor U123737 ( n56296, n74116, n56264 );
nor U123738 ( n31198, n74355, n31201 );
nor U123739 ( n31251, n74317, n31201 );
nor U123740 ( n31295, n74278, n31201 );
nor U123741 ( n31336, n74242, n31201 );
nor U123742 ( n31376, n74142, n31201 );
nor U123743 ( n10870, n74334, n10810 );
nor U123744 ( n10920, n74296, n10810 );
nor U123745 ( n10972, n74255, n10810 );
nor U123746 ( n11020, n74164, n10810 );
nor U123747 ( n11070, n74103, n10810 );
nor U123748 ( n11122, n73995, n10810 );
nor U123749 ( n11173, n74061, n10810 );
nor U123750 ( n65505, n74118, n65455 );
nor U123751 ( n65545, n73945, n65455 );
nor U123752 ( n65586, n73877, n65455 );
nor U123753 ( n65626, n73794, n65455 );
nor U123754 ( n44669, n73894, n44581 );
nor U123755 ( n44710, n73820, n44581 );
nor U123756 ( n44749, n73664, n44581 );
nor U123757 ( n44789, n73599, n44581 );
nor U123758 ( n44885, n73574, n44581 );
nor U123759 ( n44830, n73550, n44581 );
nor U123760 ( n44629, n73996, n44581 );
nor U123761 ( n10807, n74377, n10810 );
nor U123762 ( n65452, n74214, n65455 );
nor U123763 ( n44578, n74160, n44581 );
nor U123764 ( n31417, n74047, n31201 );
nor U123765 ( n31457, n73965, n31201 );
nor U123766 ( n31500, n74018, n31201 );
nor U123767 ( n65667, n73743, n65455 );
nor U123768 ( n65707, n73621, n65455 );
nor U123769 ( n65750, n73702, n65455 );
nand U123770 ( n44581, n44888, n7802 );
nor U123771 ( n44888, n44882, n44889 );
nand U123772 ( n31201, n31503, n3399 );
nor U123773 ( n31503, n31497, n31504 );
nand U123774 ( n65455, n65753, n6014 );
nor U123775 ( n65753, n65747, n65754 );
nand U123776 ( n10810, n11177, n5147 );
nor U123777 ( n11177, n11169, n11178 );
nor U123778 ( n30502, n74306, n30471 );
nor U123779 ( n9925, n74320, n9882 );
nor U123780 ( n64661, n74066, n64630 );
nor U123781 ( n43822, n73971, n43787 );
nor U123782 ( n14677, n14680, n74435 );
nor U123783 ( n14680, n4769, n12680 );
nand U123784 ( n16321, n16237, n16327 );
nand U123785 ( n16327, n16220, n15053 );
nor U123786 ( n23178, n74070, n23140 );
nor U123787 ( n56299, n74069, n56261 );
nor U123788 ( n23893, n74200, n23896 );
nor U123789 ( n57017, n74201, n57020 );
nand U123790 ( n10815, n11183, n5147 );
nor U123791 ( n11183, n11169, n11184 );
nand U123792 ( n44585, n44893, n7802 );
nor U123793 ( n44893, n44882, n44894 );
nand U123794 ( n31205, n31508, n3399 );
nor U123795 ( n31508, n31497, n31509 );
nand U123796 ( n65459, n65758, n6014 );
nor U123797 ( n65758, n65747, n65759 );
nor U123798 ( n23996, n73908, n23895 );
nor U123799 ( n24037, n73841, n23895 );
nor U123800 ( n24077, n73759, n23895 );
nor U123801 ( n57078, n74057, n57019 );
nor U123802 ( n57118, n73909, n57019 );
nor U123803 ( n57159, n73842, n57019 );
nor U123804 ( n57199, n73760, n57019 );
nor U123805 ( n23956, n74058, n23895 );
nor U123806 ( n57240, n73747, n57019 );
nor U123807 ( n57280, n73634, n57019 );
nor U123808 ( n57321, n73660, n57019 );
nor U123809 ( n24118, n73748, n23895 );
nor U123810 ( n24158, n73635, n23895 );
nor U123811 ( n24199, n73661, n23895 );
nand U123812 ( n23992, n23993, n23994 );
nor U123813 ( n23993, n23997, n23998 );
nor U123814 ( n23994, n23995, n23996 );
nor U123815 ( n23997, n73920, n23900 );
nand U123816 ( n24033, n24034, n24035 );
nor U123817 ( n24034, n24038, n24039 );
nor U123818 ( n24035, n24036, n24037 );
nor U123819 ( n24038, n73851, n23900 );
nand U123820 ( n24073, n24074, n24075 );
nor U123821 ( n24074, n24078, n24079 );
nor U123822 ( n24075, n24076, n24077 );
nor U123823 ( n24078, n73769, n23900 );
nand U123824 ( n57074, n57075, n57076 );
nor U123825 ( n57075, n57079, n57080 );
nor U123826 ( n57076, n57077, n57078 );
nor U123827 ( n57079, n74075, n57024 );
nand U123828 ( n57114, n57115, n57116 );
nor U123829 ( n57115, n57119, n57120 );
nor U123830 ( n57116, n57117, n57118 );
nor U123831 ( n57119, n73921, n57024 );
nand U123832 ( n57155, n57156, n57157 );
nor U123833 ( n57156, n57160, n57161 );
nor U123834 ( n57157, n57158, n57159 );
nor U123835 ( n57160, n73852, n57024 );
nand U123836 ( n57195, n57196, n57197 );
nor U123837 ( n57196, n57200, n57201 );
nor U123838 ( n57197, n57198, n57199 );
nor U123839 ( n57200, n73770, n57024 );
nand U123840 ( n23952, n23953, n23954 );
nor U123841 ( n23953, n23957, n23958 );
nor U123842 ( n23954, n23955, n23956 );
nor U123843 ( n23957, n74076, n23900 );
nand U123844 ( n57236, n57237, n57238 );
nor U123845 ( n57237, n57241, n57242 );
nor U123846 ( n57238, n57239, n57240 );
nor U123847 ( n57241, n73726, n57024 );
nand U123848 ( n57276, n57277, n57278 );
nor U123849 ( n57277, n57281, n57282 );
nor U123850 ( n57278, n57279, n57280 );
nor U123851 ( n57281, n73617, n57024 );
nand U123852 ( n57317, n57318, n57319 );
nor U123853 ( n57318, n57323, n57324 );
nor U123854 ( n57319, n57320, n57321 );
nor U123855 ( n57323, n73677, n57024 );
nand U123856 ( n24114, n24115, n24116 );
nor U123857 ( n24115, n24119, n24120 );
nor U123858 ( n24116, n24117, n24118 );
nor U123859 ( n24119, n73727, n23900 );
nand U123860 ( n24154, n24155, n24156 );
nor U123861 ( n24155, n24159, n24160 );
nor U123862 ( n24156, n24157, n24158 );
nor U123863 ( n24159, n73618, n23900 );
nand U123864 ( n24195, n24196, n24197 );
nor U123865 ( n24196, n24201, n24202 );
nor U123866 ( n24197, n24198, n24199 );
nor U123867 ( n24201, n73678, n23900 );
nor U123868 ( n15388, n15389, n15390 );
nor U123869 ( n23998, n73902, n23899 );
nor U123870 ( n24039, n73835, n23899 );
nor U123871 ( n24079, n73753, n23899 );
nor U123872 ( n57080, n74050, n57023 );
nor U123873 ( n57120, n73903, n57023 );
nor U123874 ( n57161, n73836, n57023 );
nor U123875 ( n57201, n73754, n57023 );
nor U123876 ( n23958, n74051, n23899 );
nor U123877 ( n57242, n73712, n57023 );
nor U123878 ( n57282, n73604, n57023 );
nor U123879 ( n57324, n73653, n57023 );
nor U123880 ( n24120, n73713, n23899 );
nor U123881 ( n24160, n73605, n23899 );
nor U123882 ( n24202, n73654, n23899 );
nor U123883 ( n48131, n48412, n48413 );
nand U123884 ( n48309, n48253, n48314 );
nand U123885 ( n48314, n48315, n48131 );
nor U123886 ( n23995, n73931, n23896 );
nor U123887 ( n24036, n73862, n23896 );
nor U123888 ( n24076, n73780, n23896 );
nor U123889 ( n57077, n74091, n57020 );
nor U123890 ( n57117, n73932, n57020 );
nor U123891 ( n57158, n73863, n57020 );
nor U123892 ( n57198, n73781, n57020 );
nor U123893 ( n23955, n74092, n23896 );
nor U123894 ( n57239, n73741, n57020 );
nor U123895 ( n57279, n73629, n57020 );
nor U123896 ( n57320, n73688, n57020 );
nor U123897 ( n24117, n73742, n23896 );
nor U123898 ( n24157, n73630, n23896 );
nor U123899 ( n24198, n73689, n23896 );
nand U123900 ( n57029, n57330, n6869 );
nor U123901 ( n57330, n57325, n55852 );
nand U123902 ( n23905, n24208, n4237 );
nor U123903 ( n24208, n24203, n22736 );
nor U123904 ( n23904, n74203, n23905 );
nor U123905 ( n57028, n74204, n57029 );
nand U123906 ( n23889, n23901, n23902 );
nor U123907 ( n23901, n23907, n23908 );
nor U123908 ( n23902, n23903, n23904 );
nor U123909 ( n23907, n74209, n23910 );
nand U123910 ( n57013, n57025, n57026 );
nor U123911 ( n57025, n57031, n57032 );
nor U123912 ( n57026, n57027, n57028 );
nor U123913 ( n57031, n74210, n57034 );
nand U123914 ( n57033, n57335, n6869 );
nor U123915 ( n57335, n57325, n55853 );
nand U123916 ( n23909, n24213, n4237 );
nor U123917 ( n24213, n24203, n22737 );
nor U123918 ( n23908, n74193, n23909 );
nor U123919 ( n57032, n74194, n57033 );
nand U123920 ( n27869, n27806, n27871 );
nand U123921 ( n27871, n27793, n27219 );
nand U123922 ( n61016, n60954, n61018 );
nand U123923 ( n61018, n60941, n60364 );
nand U123924 ( n27547, n27481, n27549 );
nand U123925 ( n27549, n27219, n4282 );
nand U123926 ( n34791, n34726, n34793 );
nand U123927 ( n34793, n34464, n3444 );
nand U123928 ( n69535, n69470, n69537 );
nand U123929 ( n69537, n69214, n6059 );
nand U123930 ( n60699, n60630, n60701 );
nand U123931 ( n60701, n60364, n6914 );
nand U123932 ( n35108, n35047, n35110 );
nand U123933 ( n35110, n35034, n34464 );
nand U123934 ( n69844, n69785, n69846 );
nand U123935 ( n69846, n69772, n69214 );
nand U123936 ( n14688, n4809, n14675 );
nand U123937 ( n57030, n57331, n6869 );
nor U123938 ( n57331, n57325, n57332 );
nand U123939 ( n23906, n24209, n4237 );
nor U123940 ( n24209, n24203, n24210 );
nor U123941 ( n23903, n74215, n23906 );
nor U123942 ( n57027, n74216, n57030 );
nor U123943 ( n24002, n73934, n23905 );
nor U123944 ( n24043, n73865, n23905 );
nor U123945 ( n24083, n73783, n23905 );
nor U123946 ( n57084, n74095, n57029 );
nor U123947 ( n57124, n73935, n57029 );
nor U123948 ( n57165, n73866, n57029 );
nor U123949 ( n57205, n73784, n57029 );
nor U123950 ( n23962, n74096, n23905 );
nor U123951 ( n57246, n73738, n57029 );
nor U123952 ( n57286, n73626, n57029 );
nor U123953 ( n57329, n73690, n57029 );
nor U123954 ( n24124, n73739, n23905 );
nor U123955 ( n24164, n73627, n23905 );
nor U123956 ( n24207, n73691, n23905 );
nand U123957 ( n23991, n23999, n24000 );
nor U123958 ( n23999, n24003, n24004 );
nor U123959 ( n24000, n24001, n24002 );
nor U123960 ( n24003, n73940, n23910 );
nand U123961 ( n24032, n24040, n24041 );
nor U123962 ( n24040, n24044, n24045 );
nor U123963 ( n24041, n24042, n24043 );
nor U123964 ( n24044, n73872, n23910 );
nand U123965 ( n24072, n24080, n24081 );
nor U123966 ( n24080, n24084, n24085 );
nor U123967 ( n24081, n24082, n24083 );
nor U123968 ( n24084, n73789, n23910 );
nand U123969 ( n57073, n57081, n57082 );
nor U123970 ( n57081, n57085, n57086 );
nor U123971 ( n57082, n57083, n57084 );
nor U123972 ( n57085, n74113, n57034 );
nand U123973 ( n57113, n57121, n57122 );
nor U123974 ( n57121, n57125, n57126 );
nor U123975 ( n57122, n57123, n57124 );
nor U123976 ( n57125, n73941, n57034 );
nand U123977 ( n57154, n57162, n57163 );
nor U123978 ( n57162, n57166, n57167 );
nor U123979 ( n57163, n57164, n57165 );
nor U123980 ( n57166, n73873, n57034 );
nand U123981 ( n57194, n57202, n57203 );
nor U123982 ( n57202, n57206, n57207 );
nor U123983 ( n57203, n57204, n57205 );
nor U123984 ( n57206, n73790, n57034 );
nand U123985 ( n23951, n23959, n23960 );
nor U123986 ( n23959, n23963, n23964 );
nor U123987 ( n23960, n23961, n23962 );
nor U123988 ( n23963, n74114, n23910 );
nand U123989 ( n57235, n57243, n57244 );
nor U123990 ( n57243, n57247, n57248 );
nor U123991 ( n57244, n57245, n57246 );
nor U123992 ( n57247, n73732, n57034 );
nand U123993 ( n57275, n57283, n57284 );
nor U123994 ( n57283, n57287, n57288 );
nor U123995 ( n57284, n57285, n57286 );
nor U123996 ( n57287, n73622, n57034 );
nand U123997 ( n57316, n57326, n57327 );
nor U123998 ( n57326, n57333, n57334 );
nor U123999 ( n57327, n57328, n57329 );
nor U124000 ( n57333, n73696, n57034 );
nand U124001 ( n24113, n24121, n24122 );
nor U124002 ( n24121, n24125, n24126 );
nor U124003 ( n24122, n24123, n24124 );
nor U124004 ( n24125, n73733, n23910 );
nand U124005 ( n24153, n24161, n24162 );
nor U124006 ( n24161, n24165, n24166 );
nor U124007 ( n24162, n24163, n24164 );
nor U124008 ( n24165, n73623, n23910 );
nand U124009 ( n24194, n24204, n24205 );
nor U124010 ( n24204, n24211, n24212 );
nor U124011 ( n24205, n24206, n24207 );
nor U124012 ( n24211, n73697, n23910 );
nand U124013 ( n23910, n24214, n4237 );
nor U124014 ( n24214, n24203, n24215 );
nand U124015 ( n57034, n57336, n6869 );
nor U124016 ( n57336, n57325, n57337 );
nor U124017 ( n24004, n73922, n23909 );
nor U124018 ( n24045, n73853, n23909 );
nor U124019 ( n24085, n73771, n23909 );
nor U124020 ( n57086, n74077, n57033 );
nor U124021 ( n57126, n73923, n57033 );
nor U124022 ( n57167, n73854, n57033 );
nor U124023 ( n57207, n73772, n57033 );
nor U124024 ( n23964, n74078, n23909 );
nor U124025 ( n57248, n73720, n57033 );
nor U124026 ( n57288, n73613, n57033 );
nor U124027 ( n57334, n73679, n57033 );
nor U124028 ( n24126, n73721, n23909 );
nor U124029 ( n24166, n73614, n23909 );
nor U124030 ( n24212, n73680, n23909 );
nor U124031 ( n24001, n73946, n23906 );
nor U124032 ( n24042, n73878, n23906 );
nor U124033 ( n24082, n73795, n23906 );
nor U124034 ( n57083, n74119, n57030 );
nor U124035 ( n57123, n73947, n57030 );
nor U124036 ( n57164, n73879, n57030 );
nor U124037 ( n57204, n73796, n57030 );
nor U124038 ( n23961, n74120, n23906 );
nor U124039 ( n57245, n73744, n57030 );
nor U124040 ( n57285, n73631, n57030 );
nor U124041 ( n57328, n73703, n57030 );
nor U124042 ( n24123, n73745, n23906 );
nor U124043 ( n24163, n73632, n23906 );
nor U124044 ( n24206, n73704, n23906 );
nand U124045 ( n14679, n76187, n14675 );
nand U124046 ( n47904, n76177, n47901 );
not U124047 ( n6429, n31914 );
or U124048 ( n30467, n75896, n75897 );
nor U124049 ( n75896, n30471, n74344 );
nor U124050 ( n75897, n30470, n74352 );
or U124051 ( n9877, n75898, n75899 );
nor U124052 ( n75898, n9882, n74363 );
nor U124053 ( n75899, n9880, n74365 );
or U124054 ( n64626, n75900, n75901 );
nor U124055 ( n75900, n64630, n74181 );
nor U124056 ( n75901, n64629, n74205 );
or U124057 ( n43783, n75902, n75903 );
nor U124058 ( n75902, n43787, n74138 );
nor U124059 ( n75903, n43786, n74151 );
nand U124060 ( n10824, n11193, n11169 );
nor U124061 ( n11193, n9380, n11194 );
nand U124062 ( n44592, n44901, n44882 );
nor U124063 ( n44901, n43330, n44902 );
nand U124064 ( n31212, n31516, n31497 );
nor U124065 ( n31516, n30059, n31517 );
nand U124066 ( n65466, n65766, n65747 );
nor U124067 ( n65766, n64076, n65767 );
nor U124068 ( n31211, n74339, n31212 );
nor U124069 ( n31260, n74303, n31212 );
nor U124070 ( n31304, n74261, n31212 );
nor U124071 ( n31345, n74223, n31212 );
nor U124072 ( n31385, n74104, n31212 );
nor U124073 ( n10882, n74323, n10824 );
nor U124074 ( n10932, n74286, n10824 );
nor U124075 ( n10983, n74241, n10824 );
nor U124076 ( n11032, n74140, n10824 );
nor U124077 ( n11082, n74084, n10824 );
nor U124078 ( n11133, n73981, n10824 );
nor U124079 ( n11192, n74017, n10824 );
nor U124080 ( n65514, n74053, n65466 );
nor U124081 ( n65554, n73904, n65466 );
nor U124082 ( n65595, n73837, n65466 );
nor U124083 ( n65635, n73755, n65466 );
nor U124084 ( n44678, n73881, n44592 );
nor U124085 ( n44719, n73807, n44592 );
nor U124086 ( n44758, n73639, n44592 );
nor U124087 ( n44798, n73577, n44592 );
nor U124088 ( n44900, n73555, n44592 );
nor U124089 ( n44839, n73539, n44592 );
nor U124090 ( n44638, n73967, n44592 );
nor U124091 ( n10823, n74359, n10824 );
nor U124092 ( n65465, n74171, n65466 );
nor U124093 ( n44591, n74130, n44592 );
nor U124094 ( n31426, n74024, n31212 );
nor U124095 ( n31466, n73954, n31212 );
nor U124096 ( n31515, n74001, n31212 );
nor U124097 ( n65676, n73714, n65466 );
nor U124098 ( n65716, n73589, n65466 );
nor U124099 ( n65765, n73655, n65466 );
nand U124100 ( n31207, n31208, n31209 );
nor U124101 ( n31208, n31214, n31215 );
nor U124102 ( n31209, n31210, n31211 );
nor U124103 ( n31214, n74343, n31217 );
nand U124104 ( n31256, n31257, n31258 );
nor U124105 ( n31257, n31261, n31262 );
nor U124106 ( n31258, n31259, n31260 );
nor U124107 ( n31261, n74305, n31217 );
nand U124108 ( n31300, n31301, n31302 );
nor U124109 ( n31301, n31305, n31306 );
nor U124110 ( n31302, n31303, n31304 );
nor U124111 ( n31305, n74264, n31217 );
nand U124112 ( n31341, n31342, n31343 );
nor U124113 ( n31342, n31346, n31347 );
nor U124114 ( n31343, n31344, n31345 );
nor U124115 ( n31346, n74226, n31217 );
nand U124116 ( n31381, n31382, n31383 );
nor U124117 ( n31382, n31386, n31387 );
nor U124118 ( n31383, n31384, n31385 );
nor U124119 ( n31386, n74121, n31217 );
nand U124120 ( n10877, n10878, n10879 );
nor U124121 ( n10878, n10883, n10884 );
nor U124122 ( n10879, n10880, n10882 );
nor U124123 ( n10883, n74321, n10830 );
nand U124124 ( n10927, n10928, n10929 );
nor U124125 ( n10928, n10933, n10934 );
nor U124126 ( n10929, n10930, n10932 );
nor U124127 ( n10933, n74284, n10830 );
nand U124128 ( n10978, n10979, n10980 );
nor U124129 ( n10979, n10984, n10985 );
nor U124130 ( n10980, n10982, n10983 );
nor U124131 ( n10984, n74244, n10830 );
nand U124132 ( n11027, n11028, n11029 );
nor U124133 ( n11028, n11033, n11034 );
nor U124134 ( n11029, n11030, n11032 );
nor U124135 ( n11033, n74149, n10830 );
nand U124136 ( n11077, n11078, n11079 );
nor U124137 ( n11078, n11083, n11084 );
nor U124138 ( n11079, n11080, n11082 );
nor U124139 ( n11083, n74072, n10830 );
nand U124140 ( n11128, n11129, n11130 );
nor U124141 ( n11129, n11134, n11135 );
nor U124142 ( n11130, n11132, n11133 );
nor U124143 ( n11134, n73979, n10830 );
nand U124144 ( n11187, n11188, n11189 );
nor U124145 ( n11188, n11197, n11198 );
nor U124146 ( n11189, n11190, n11192 );
nor U124147 ( n11197, n74026, n10830 );
nand U124148 ( n65510, n65511, n65512 );
nor U124149 ( n65511, n65515, n65516 );
nor U124150 ( n65512, n65513, n65514 );
nor U124151 ( n65515, n74065, n65471 );
nand U124152 ( n65550, n65551, n65552 );
nor U124153 ( n65551, n65555, n65556 );
nor U124154 ( n65552, n65553, n65554 );
nor U124155 ( n65555, n73912, n65471 );
nand U124156 ( n65591, n65592, n65593 );
nor U124157 ( n65592, n65596, n65597 );
nor U124158 ( n65593, n65594, n65595 );
nor U124159 ( n65596, n73843, n65471 );
nand U124160 ( n65631, n65632, n65633 );
nor U124161 ( n65632, n65636, n65637 );
nor U124162 ( n65633, n65634, n65635 );
nor U124163 ( n65636, n73761, n65471 );
nand U124164 ( n44674, n44675, n44676 );
nor U124165 ( n44675, n44679, n44680 );
nor U124166 ( n44676, n44677, n44678 );
nor U124167 ( n44679, n73883, n44597 );
nand U124168 ( n44715, n44716, n44717 );
nor U124169 ( n44716, n44720, n44721 );
nor U124170 ( n44717, n44718, n44719 );
nor U124171 ( n44720, n73809, n44597 );
nand U124172 ( n44754, n44755, n44756 );
nor U124173 ( n44755, n44759, n44760 );
nor U124174 ( n44756, n44757, n44758 );
nor U124175 ( n44759, n73644, n44597 );
nand U124176 ( n44794, n44795, n44796 );
nor U124177 ( n44795, n44799, n44800 );
nor U124178 ( n44796, n44797, n44798 );
nor U124179 ( n44799, n73575, n44597 );
nand U124180 ( n44896, n44897, n44898 );
nor U124181 ( n44897, n44904, n44905 );
nor U124182 ( n44898, n44899, n44900 );
nor U124183 ( n44904, n73557, n44597 );
nand U124184 ( n44835, n44836, n44837 );
nor U124185 ( n44836, n44840, n44841 );
nor U124186 ( n44837, n44838, n44839 );
nor U124187 ( n44840, n73537, n44597 );
nand U124188 ( n44634, n44635, n44636 );
nor U124189 ( n44635, n44639, n44640 );
nor U124190 ( n44636, n44637, n44638 );
nor U124191 ( n44639, n73970, n44597 );
nand U124192 ( n10818, n10819, n10820 );
nor U124193 ( n10819, n10827, n10828 );
nor U124194 ( n10820, n10822, n10823 );
nor U124195 ( n10827, n74364, n10830 );
nand U124196 ( n65461, n65462, n65463 );
nor U124197 ( n65462, n65468, n65469 );
nor U124198 ( n65463, n65464, n65465 );
nor U124199 ( n65468, n74180, n65471 );
nand U124200 ( n44587, n44588, n44589 );
nor U124201 ( n44588, n44594, n44595 );
nor U124202 ( n44589, n44590, n44591 );
nor U124203 ( n44594, n74135, n44597 );
nand U124204 ( n31422, n31423, n31424 );
nor U124205 ( n31423, n31427, n31428 );
nor U124206 ( n31424, n31425, n31426 );
nor U124207 ( n31427, n74022, n31217 );
nand U124208 ( n31462, n31463, n31464 );
nor U124209 ( n31463, n31467, n31468 );
nor U124210 ( n31464, n31465, n31466 );
nor U124211 ( n31467, n73952, n31217 );
nand U124212 ( n31511, n31512, n31513 );
nor U124213 ( n31512, n31519, n31520 );
nor U124214 ( n31513, n31514, n31515 );
nor U124215 ( n31519, n74003, n31217 );
nand U124216 ( n65672, n65673, n65674 );
nor U124217 ( n65673, n65677, n65678 );
nor U124218 ( n65674, n65675, n65676 );
nor U124219 ( n65677, n73707, n65471 );
nand U124220 ( n65712, n65713, n65714 );
nor U124221 ( n65713, n65717, n65718 );
nor U124222 ( n65714, n65715, n65716 );
nor U124223 ( n65717, n73585, n65471 );
nand U124224 ( n65761, n65762, n65763 );
nor U124225 ( n65762, n65769, n65770 );
nor U124226 ( n65763, n65764, n65765 );
nor U124227 ( n65769, n73665, n65471 );
or U124228 ( n30473, n30474, n74354 );
or U124229 ( n9884, n9885, n74374 );
or U124230 ( n64632, n64633, n74211 );
or U124231 ( n43789, n43790, n74159 );
nand U124232 ( n10837, n11207, n11169 );
nor U124233 ( n11207, n5147, n9380 );
nand U124234 ( n44602, n44912, n44882 );
nor U124235 ( n44912, n7802, n43330 );
nand U124236 ( n31222, n31527, n31497 );
nor U124237 ( n31527, n3399, n30059 );
nand U124238 ( n65476, n65777, n65747 );
nor U124239 ( n65777, n6014, n64076 );
nor U124240 ( n15810, n16227, n15389 );
nor U124241 ( n16227, n4809, n14947 );
or U124242 ( n23136, n75904, n75905 );
nor U124243 ( n75904, n23140, n74184 );
nor U124244 ( n75905, n23139, n74206 );
or U124245 ( n56257, n75906, n75907 );
nor U124246 ( n75906, n56261, n74185 );
nor U124247 ( n75907, n56260, n74207 );
nor U124248 ( n31219, n31220, n31221 );
nor U124249 ( n31220, n74354, n31223 );
nor U124250 ( n31221, n74349, n31222 );
nor U124251 ( n31264, n31265, n31266 );
nor U124252 ( n31265, n74316, n31223 );
nor U124253 ( n31266, n74310, n31222 );
nor U124254 ( n31308, n31309, n31310 );
nor U124255 ( n31309, n74277, n31223 );
nor U124256 ( n31310, n74270, n31222 );
nor U124257 ( n31349, n31350, n31351 );
nor U124258 ( n31350, n74239, n31223 );
nor U124259 ( n31351, n74231, n31222 );
nor U124260 ( n31389, n31390, n31391 );
nor U124261 ( n31390, n74137, n31223 );
nor U124262 ( n31391, n74127, n31222 );
nor U124263 ( n10887, n10888, n10889 );
nor U124264 ( n10888, n74330, n10838 );
nor U124265 ( n10889, n74326, n10837 );
nor U124266 ( n10937, n10938, n10939 );
nor U124267 ( n10938, n74293, n10838 );
nor U124268 ( n10939, n74289, n10837 );
nor U124269 ( n10988, n10989, n10990 );
nor U124270 ( n10989, n74254, n10838 );
nor U124271 ( n10990, n74249, n10837 );
nor U124272 ( n11037, n11038, n11039 );
nor U124273 ( n11038, n74163, n10838 );
nor U124274 ( n11039, n74155, n10837 );
nor U124275 ( n11087, n11088, n11089 );
nor U124276 ( n11088, n74099, n10838 );
nor U124277 ( n11089, n74089, n10837 );
nor U124278 ( n11138, n11139, n11140 );
nor U124279 ( n11139, n73989, n10838 );
nor U124280 ( n11140, n73984, n10837 );
nor U124281 ( n11203, n11204, n11205 );
nor U124282 ( n11204, n74060, n10838 );
nor U124283 ( n11205, n74039, n10837 );
nor U124284 ( n65518, n65519, n65520 );
nor U124285 ( n65519, n74115, n65477 );
nor U124286 ( n65520, n74083, n65476 );
nor U124287 ( n65558, n65559, n65560 );
nor U124288 ( n65559, n73942, n65477 );
nor U124289 ( n65560, n73927, n65476 );
nor U124290 ( n65599, n65600, n65601 );
nor U124291 ( n65600, n73874, n65477 );
nor U124292 ( n65601, n73858, n65476 );
nor U124293 ( n65639, n65640, n65641 );
nor U124294 ( n65640, n73791, n65477 );
nor U124295 ( n65641, n73776, n65476 );
nor U124296 ( n44682, n44683, n44684 );
nor U124297 ( n44683, n73893, n44603 );
nor U124298 ( n44684, n73888, n44602 );
nor U124299 ( n44723, n44724, n44725 );
nor U124300 ( n44724, n73819, n44603 );
nor U124301 ( n44725, n73814, n44602 );
nor U124302 ( n44762, n44763, n44764 );
nor U124303 ( n44763, n73663, n44603 );
nor U124304 ( n44764, n73649, n44602 );
nor U124305 ( n44802, n44803, n44804 );
nor U124306 ( n44803, n73587, n44603 );
nor U124307 ( n44804, n73581, n44602 );
nor U124308 ( n44909, n44910, n44911 );
nor U124309 ( n44910, n73572, n44603 );
nor U124310 ( n44911, n73563, n44602 );
nor U124311 ( n44843, n44844, n44845 );
nor U124312 ( n44844, n73547, n44603 );
nor U124313 ( n44845, n73542, n44602 );
nor U124314 ( n44642, n44643, n44644 );
nor U124315 ( n44643, n73994, n44603 );
nor U124316 ( n44644, n73975, n44602 );
nor U124317 ( n10833, n10834, n10835 );
nor U124318 ( n10834, n74374, n10838 );
nor U124319 ( n10835, n74369, n10837 );
nor U124320 ( n65473, n65474, n65475 );
nor U124321 ( n65474, n74211, n65477 );
nor U124322 ( n65475, n74195, n65476 );
nor U124323 ( n44599, n44600, n44601 );
nor U124324 ( n44600, n74159, n44603 );
nor U124325 ( n44601, n74146, n44602 );
nor U124326 ( n31430, n31431, n31432 );
nor U124327 ( n31431, n74040, n31223 );
nor U124328 ( n31432, n74032, n31222 );
nor U124329 ( n31470, n31471, n31472 );
nor U124330 ( n31471, n73961, n31223 );
nor U124331 ( n31472, n73957, n31222 );
nor U124332 ( n31524, n31525, n31526 );
nor U124333 ( n31525, n74015, n31223 );
nor U124334 ( n31526, n74009, n31222 );
nor U124335 ( n65680, n65681, n65682 );
nor U124336 ( n65681, n73734, n65477 );
nor U124337 ( n65682, n73722, n65476 );
nor U124338 ( n65720, n65721, n65722 );
nor U124339 ( n65721, n73603, n65477 );
nor U124340 ( n65722, n73594, n65476 );
nor U124341 ( n65774, n65775, n65776 );
nor U124342 ( n65775, n73698, n65477 );
nor U124343 ( n65776, n73681, n65476 );
nand U124344 ( n10825, n11195, n11169 );
nor U124345 ( n11195, n11178, n11194 );
nand U124346 ( n44593, n44903, n44882 );
nor U124347 ( n44903, n44889, n44902 );
nand U124348 ( n31213, n31518, n31497 );
nor U124349 ( n31518, n31504, n31517 );
nand U124350 ( n65467, n65768, n65747 );
nor U124351 ( n65768, n65754, n65767 );
nor U124352 ( n31210, n74345, n31213 );
nor U124353 ( n31259, n74309, n31213 );
nor U124354 ( n31303, n74269, n31213 );
nor U124355 ( n31344, n74230, n31213 );
nor U124356 ( n31384, n74126, n31213 );
nor U124357 ( n10880, n74328, n10825 );
nor U124358 ( n10930, n74291, n10825 );
nor U124359 ( n10982, n74248, n10825 );
nor U124360 ( n11030, n74154, n10825 );
nor U124361 ( n11080, n74097, n10825 );
nor U124362 ( n11132, n73986, n10825 );
nor U124363 ( n11190, n74038, n10825 );
nor U124364 ( n65513, n74079, n65467 );
nor U124365 ( n65553, n73924, n65467 );
nor U124366 ( n65594, n73855, n65467 );
nor U124367 ( n65634, n73773, n65467 );
nor U124368 ( n44677, n73887, n44593 );
nor U124369 ( n44718, n73813, n44593 );
nor U124370 ( n44757, n73648, n44593 );
nor U124371 ( n44797, n73584, n44593 );
nor U124372 ( n44899, n73562, n44593 );
nor U124373 ( n44838, n73545, n44593 );
nor U124374 ( n44637, n73974, n44593 );
nor U124375 ( n10822, n74367, n10825 );
nor U124376 ( n65464, n74186, n65467 );
nor U124377 ( n44590, n74141, n44593 );
nor U124378 ( n31425, n74034, n31213 );
nor U124379 ( n31465, n73959, n31213 );
nor U124380 ( n31514, n74008, n31213 );
nor U124381 ( n65675, n73728, n65467 );
nor U124382 ( n65715, n73596, n65467 );
nor U124383 ( n65764, n73676, n65467 );
or U124384 ( n23142, n23143, n74212 );
or U124385 ( n56263, n56264, n74213 );
nand U124386 ( n10838, n11208, n11169 );
nor U124387 ( n11208, n5147, n11178 );
nand U124388 ( n44603, n44913, n44882 );
nor U124389 ( n44913, n7802, n44889 );
nand U124390 ( n31223, n31528, n31497 );
nor U124391 ( n31528, n3399, n31504 );
nand U124392 ( n65477, n65778, n65747 );
nor U124393 ( n65778, n6014, n65754 );
nand U124394 ( n10829, n11199, n11169 );
nor U124395 ( n11199, n9382, n11194 );
nand U124396 ( n44596, n44906, n44882 );
nor U124397 ( n44906, n43331, n44902 );
nand U124398 ( n31216, n31521, n31497 );
nor U124399 ( n31521, n30060, n31517 );
nand U124400 ( n65470, n65771, n65747 );
nor U124401 ( n65771, n64077, n65767 );
nor U124402 ( n31215, n74338, n31216 );
nor U124403 ( n31262, n74299, n31216 );
nor U124404 ( n31306, n74258, n31216 );
nor U124405 ( n31347, n74221, n31216 );
nor U124406 ( n31387, n74063, n31216 );
nor U124407 ( n10884, n74319, n10829 );
nor U124408 ( n10934, n74280, n10829 );
nor U124409 ( n10985, n74232, n10829 );
nor U124410 ( n11034, n74128, n10829 );
nor U124411 ( n11084, n74046, n10829 );
nor U124412 ( n11135, n73964, n10829 );
nor U124413 ( n11198, n74005, n10829 );
nor U124414 ( n65516, n74027, n65470 );
nor U124415 ( n65556, n73898, n65470 );
nor U124416 ( n65597, n73830, n65470 );
nor U124417 ( n65637, n73749, n65470 );
nor U124418 ( n44680, n73867, n44596 );
nor U124419 ( n44721, n73805, n44596 );
nor U124420 ( n44760, n73636, n44596 );
nor U124421 ( n44800, n73558, n44596 );
nor U124422 ( n44905, n73553, n44596 );
nor U124423 ( n44841, n73534, n44596 );
nor U124424 ( n44640, n73950, n44596 );
nor U124425 ( n10828, n74357, n10829 );
nor U124426 ( n65469, n74167, n65470 );
nor U124427 ( n44595, n74106, n44596 );
nor U124428 ( n31428, n74012, n31216 );
nor U124429 ( n31468, n73949, n31216 );
nor U124430 ( n31520, n73987, n31216 );
nor U124431 ( n65678, n73666, n65470 );
nor U124432 ( n65718, n73564, n65470 );
nor U124433 ( n65770, n73643, n65470 );
or U124434 ( n30472, n30475, n74349 );
or U124435 ( n9883, n9887, n74369 );
or U124436 ( n64631, n64634, n74195 );
or U124437 ( n43788, n43791, n74146 );
nand U124438 ( n10842, n11212, n11169 );
nor U124439 ( n11212, n5147, n9382 );
nand U124440 ( n44606, n44916, n44882 );
nor U124441 ( n44916, n7802, n43331 );
nand U124442 ( n31226, n31531, n31497 );
nor U124443 ( n31531, n3399, n30060 );
nand U124444 ( n65480, n65781, n65747 );
nor U124445 ( n65781, n6014, n64077 );
nor U124446 ( n31218, n31224, n31225 );
nor U124447 ( n31224, n74352, n31227 );
nor U124448 ( n31225, n74344, n31226 );
nor U124449 ( n31263, n31267, n31268 );
nor U124450 ( n31267, n74313, n31227 );
nor U124451 ( n31268, n74306, n31226 );
nor U124452 ( n31307, n31311, n31312 );
nor U124453 ( n31311, n74275, n31227 );
nor U124454 ( n31312, n74265, n31226 );
nor U124455 ( n31348, n31352, n31353 );
nor U124456 ( n31352, n74237, n31227 );
nor U124457 ( n31353, n74227, n31226 );
nor U124458 ( n31388, n31392, n31393 );
nor U124459 ( n31392, n74134, n31227 );
nor U124460 ( n31393, n74122, n31226 );
nor U124461 ( n10885, n10890, n10892 );
nor U124462 ( n10890, n74324, n10843 );
nor U124463 ( n10892, n74320, n10842 );
nor U124464 ( n10987, n10992, n10993 );
nor U124465 ( n10992, n74252, n10843 );
nor U124466 ( n10993, n74245, n10842 );
nor U124467 ( n11035, n11040, n11042 );
nor U124468 ( n11040, n74161, n10843 );
nor U124469 ( n11042, n74150, n10842 );
nor U124470 ( n11137, n11142, n11143 );
nor U124471 ( n11142, n73982, n10843 );
nor U124472 ( n11143, n73978, n10842 );
nor U124473 ( n11202, n11209, n11210 );
nor U124474 ( n11209, n74052, n10843 );
nor U124475 ( n11210, n74031, n10842 );
nor U124476 ( n65517, n65521, n65522 );
nor U124477 ( n65521, n74108, n65481 );
nor U124478 ( n65522, n74066, n65480 );
nor U124479 ( n65557, n65561, n65562 );
nor U124480 ( n65561, n73936, n65481 );
nor U124481 ( n65562, n73913, n65480 );
nor U124482 ( n65598, n65602, n65603 );
nor U124483 ( n65602, n73868, n65481 );
nor U124484 ( n65603, n73844, n65480 );
nor U124485 ( n65638, n65642, n65643 );
nor U124486 ( n65642, n73785, n65481 );
nor U124487 ( n65643, n73762, n65480 );
nor U124488 ( n44681, n44685, n44686 );
nor U124489 ( n44685, n73891, n44607 );
nor U124490 ( n44686, n73884, n44606 );
nor U124491 ( n44722, n44726, n44727 );
nor U124492 ( n44726, n73817, n44607 );
nor U124493 ( n44727, n73810, n44606 );
nor U124494 ( n44761, n44765, n44766 );
nor U124495 ( n44765, n73656, n44607 );
nor U124496 ( n44766, n73645, n44606 );
nor U124497 ( n44801, n44805, n44806 );
nor U124498 ( n44805, n73578, n44607 );
nor U124499 ( n44806, n73573, n44606 );
nor U124500 ( n44908, n44914, n44915 );
nor U124501 ( n44914, n73570, n44607 );
nor U124502 ( n44915, n73559, n44606 );
nor U124503 ( n44842, n44846, n44847 );
nor U124504 ( n44846, n73540, n44607 );
nor U124505 ( n44847, n73536, n44606 );
nor U124506 ( n44641, n44645, n44646 );
nor U124507 ( n44645, n73990, n44607 );
nor U124508 ( n44646, n73971, n44606 );
nor U124509 ( n10832, n10839, n10840 );
nor U124510 ( n10839, n74365, n10843 );
nor U124511 ( n10840, n74363, n10842 );
nor U124512 ( n65472, n65478, n65479 );
nor U124513 ( n65478, n74205, n65481 );
nor U124514 ( n65479, n74181, n65480 );
nor U124515 ( n44598, n44604, n44605 );
nor U124516 ( n44604, n74151, n44607 );
nor U124517 ( n44605, n74138, n44606 );
nor U124518 ( n31429, n31433, n31434 );
nor U124519 ( n31433, n74025, n31227 );
nor U124520 ( n31434, n74021, n31226 );
nor U124521 ( n31469, n31473, n31474 );
nor U124522 ( n31473, n73955, n31227 );
nor U124523 ( n31474, n73951, n31226 );
nor U124524 ( n31523, n31529, n31530 );
nor U124525 ( n31529, n74013, n31227 );
nor U124526 ( n31530, n74004, n31226 );
nor U124527 ( n65679, n65683, n65684 );
nor U124528 ( n65683, n73711, n65481 );
nor U124529 ( n65684, n73701, n65480 );
nor U124530 ( n65719, n65723, n65724 );
nor U124531 ( n65723, n73590, n65481 );
nor U124532 ( n65724, n73583, n65480 );
nor U124533 ( n65773, n65779, n65780 );
nor U124534 ( n65779, n73692, n65481 );
nor U124535 ( n65780, n73667, n65480 );
nor U124536 ( n10935, n10940, n10942 );
nor U124537 ( n10940, n74287, n10843 );
nor U124538 ( n10942, n74283, n10842 );
nor U124539 ( n11085, n11090, n11092 );
nor U124540 ( n11090, n74085, n10843 );
nor U124541 ( n11092, n74071, n10842 );
nand U124542 ( n10830, n11200, n11169 );
nor U124543 ( n11200, n11184, n11194 );
nand U124544 ( n44597, n44907, n44882 );
nor U124545 ( n44907, n44894, n44902 );
nand U124546 ( n31217, n31522, n31497 );
nor U124547 ( n31522, n31509, n31517 );
nand U124548 ( n65471, n65772, n65747 );
nor U124549 ( n65772, n65759, n65767 );
or U124550 ( n23141, n23144, n74196 );
or U124551 ( n56262, n56265, n74197 );
nand U124552 ( n10843, n11213, n11169 );
nor U124553 ( n11213, n5147, n11184 );
nand U124554 ( n44607, n44917, n44882 );
nor U124555 ( n44917, n7802, n44894 );
nand U124556 ( n31227, n31532, n31497 );
nor U124557 ( n31532, n3399, n31509 );
nand U124558 ( n65481, n65782, n65747 );
nor U124559 ( n65782, n6014, n65759 );
nor U124560 ( n14684, n4772, n14693 );
nand U124561 ( n14693, n5207, n14675 );
not U124562 ( n2908, n38361 );
not U124563 ( n1790, n48794 );
nor U124564 ( n34367, n34628, n34629 );
nor U124565 ( n69119, n69374, n69375 );
nand U124566 ( n34455, n34393, n34463 );
nand U124567 ( n34463, n34464, n34367 );
nand U124568 ( n69205, n69145, n69213 );
nand U124569 ( n69213, n69214, n69119 );
nor U124570 ( n27122, n27383, n27384 );
nor U124571 ( n60266, n60531, n60532 );
nand U124572 ( n34539, n34477, n34545 );
nand U124573 ( n34545, n34546, n34367 );
nand U124574 ( n69287, n69227, n69293 );
nand U124575 ( n69293, n69294, n69119 );
nand U124576 ( n27210, n27150, n27218 );
nand U124577 ( n27218, n27219, n27122 );
nand U124578 ( n60355, n60292, n60363 );
nand U124579 ( n60363, n60364, n60266 );
nand U124580 ( n27294, n27232, n27300 );
nand U124581 ( n27300, n27301, n27122 );
nand U124582 ( n60437, n60377, n60443 );
nand U124583 ( n60443, n60444, n60266 );
not U124584 ( n3640, n31178 );
not U124585 ( n6268, n65432 );
not U124586 ( n7160, n57059 );
not U124587 ( n4528, n23935 );
nor U124588 ( n14738, n74538, n14675 );
nor U124589 ( n34703, n34704, n34705 );
nor U124590 ( n27458, n27459, n27460 );
nor U124591 ( n69447, n69448, n69449 );
nor U124592 ( n60607, n60608, n60609 );
nand U124593 ( n57041, n57344, n57325 );
nor U124594 ( n57344, n55852, n57345 );
nand U124595 ( n23917, n24222, n24203 );
nor U124596 ( n24222, n22736, n24223 );
nor U124597 ( n24010, n73905, n23917 );
nor U124598 ( n24051, n73838, n23917 );
nor U124599 ( n24091, n73756, n23917 );
nor U124600 ( n57092, n74054, n57041 );
nor U124601 ( n57132, n73906, n57041 );
nor U124602 ( n57173, n73839, n57041 );
nor U124603 ( n23970, n74055, n23917 );
nor U124604 ( n57254, n73715, n57041 );
nor U124605 ( n57294, n73606, n57041 );
nor U124606 ( n57343, n73657, n57041 );
nor U124607 ( n24132, n73716, n23917 );
nor U124608 ( n24172, n73607, n23917 );
nor U124609 ( n24221, n73658, n23917 );
nor U124610 ( n23916, n74172, n23917 );
nor U124611 ( n57040, n74173, n57041 );
nand U124612 ( n24006, n24007, n24008 );
nor U124613 ( n24007, n24011, n24012 );
nor U124614 ( n24008, n24009, n24010 );
nor U124615 ( n24011, n73914, n23922 );
nand U124616 ( n24047, n24048, n24049 );
nor U124617 ( n24048, n24052, n24053 );
nor U124618 ( n24049, n24050, n24051 );
nor U124619 ( n24052, n73845, n23922 );
nand U124620 ( n24087, n24088, n24089 );
nor U124621 ( n24088, n24092, n24093 );
nor U124622 ( n24089, n24090, n24091 );
nor U124623 ( n24092, n73763, n23922 );
nand U124624 ( n57088, n57089, n57090 );
nor U124625 ( n57089, n57093, n57094 );
nor U124626 ( n57090, n57091, n57092 );
nor U124627 ( n57093, n74067, n57046 );
nand U124628 ( n57128, n57129, n57130 );
nor U124629 ( n57129, n57133, n57134 );
nor U124630 ( n57130, n57131, n57132 );
nor U124631 ( n57133, n73915, n57046 );
nand U124632 ( n57169, n57170, n57171 );
nor U124633 ( n57170, n57174, n57175 );
nor U124634 ( n57171, n57172, n57173 );
nor U124635 ( n57174, n73846, n57046 );
nand U124636 ( n23966, n23967, n23968 );
nor U124637 ( n23967, n23971, n23972 );
nor U124638 ( n23968, n23969, n23970 );
nor U124639 ( n23971, n74068, n23922 );
nand U124640 ( n57250, n57251, n57252 );
nor U124641 ( n57251, n57255, n57256 );
nor U124642 ( n57252, n57253, n57254 );
nor U124643 ( n57255, n73708, n57046 );
nand U124644 ( n57339, n57340, n57341 );
nor U124645 ( n57340, n57347, n57348 );
nor U124646 ( n57341, n57342, n57343 );
nor U124647 ( n57347, n73668, n57046 );
nand U124648 ( n24128, n24129, n24130 );
nor U124649 ( n24129, n24133, n24134 );
nor U124650 ( n24130, n24131, n24132 );
nor U124651 ( n24133, n73709, n23922 );
nand U124652 ( n24217, n24218, n24219 );
nor U124653 ( n24218, n24225, n24226 );
nor U124654 ( n24219, n24220, n24221 );
nor U124655 ( n24225, n73669, n23922 );
nand U124656 ( n23912, n23913, n23914 );
nor U124657 ( n23913, n23919, n23920 );
nor U124658 ( n23914, n23915, n23916 );
nor U124659 ( n23919, n74182, n23922 );
nand U124660 ( n57036, n57037, n57038 );
nor U124661 ( n57037, n57043, n57044 );
nor U124662 ( n57038, n57039, n57040 );
nor U124663 ( n57043, n74183, n57046 );
nor U124664 ( n57213, n73757, n57041 );
and U124665 ( n28115, n27384, n27383 );
and U124666 ( n35350, n34629, n34628 );
and U124667 ( n70082, n69375, n69374 );
and U124668 ( n61270, n60532, n60531 );
nand U124669 ( n57209, n57210, n57211 );
nor U124670 ( n57210, n57214, n57215 );
nor U124671 ( n57211, n57212, n57213 );
nor U124672 ( n57214, n73764, n57046 );
nand U124673 ( n57290, n57291, n57292 );
nor U124674 ( n57291, n57295, n57296 );
nor U124675 ( n57292, n57293, n57294 );
nor U124676 ( n57295, n73600, n57046 );
nand U124677 ( n24168, n24169, n24170 );
nor U124678 ( n24169, n24173, n24174 );
nor U124679 ( n24170, n24171, n24172 );
nor U124680 ( n24173, n73601, n23922 );
nand U124681 ( n23927, n24233, n24203 );
nor U124682 ( n24233, n4237, n22736 );
nand U124683 ( n57051, n57355, n57325 );
nor U124684 ( n57355, n6869, n55852 );
nor U124685 ( n24014, n24015, n24016 );
nor U124686 ( n24015, n73943, n23928 );
nor U124687 ( n24016, n73928, n23927 );
nor U124688 ( n24055, n24056, n24057 );
nor U124689 ( n24056, n73875, n23928 );
nor U124690 ( n24057, n73859, n23927 );
nor U124691 ( n24095, n24096, n24097 );
nor U124692 ( n24096, n73792, n23928 );
nor U124693 ( n24097, n73777, n23927 );
nor U124694 ( n57096, n57097, n57098 );
nor U124695 ( n57097, n74116, n57052 );
nor U124696 ( n57098, n74086, n57051 );
nor U124697 ( n57136, n57137, n57138 );
nor U124698 ( n57137, n73944, n57052 );
nor U124699 ( n57138, n73929, n57051 );
nor U124700 ( n57177, n57178, n57179 );
nor U124701 ( n57178, n73876, n57052 );
nor U124702 ( n57179, n73860, n57051 );
nor U124703 ( n57217, n57218, n57219 );
nor U124704 ( n57218, n73793, n57052 );
nor U124705 ( n57219, n73778, n57051 );
nor U124706 ( n23974, n23975, n23976 );
nor U124707 ( n23975, n74117, n23928 );
nor U124708 ( n23976, n74087, n23927 );
nor U124709 ( n57258, n57259, n57260 );
nor U124710 ( n57259, n73735, n57052 );
nor U124711 ( n57260, n73723, n57051 );
nor U124712 ( n57298, n57299, n57300 );
nor U124713 ( n57299, n73624, n57052 );
nor U124714 ( n57300, n73615, n57051 );
nor U124715 ( n57352, n57353, n57354 );
nor U124716 ( n57353, n73699, n57052 );
nor U124717 ( n57354, n73684, n57051 );
nor U124718 ( n24136, n24137, n24138 );
nor U124719 ( n24137, n73736, n23928 );
nor U124720 ( n24138, n73724, n23927 );
nor U124721 ( n24176, n24177, n24178 );
nor U124722 ( n24177, n73625, n23928 );
nor U124723 ( n24178, n73616, n23927 );
nor U124724 ( n24230, n24231, n24232 );
nor U124725 ( n24231, n73700, n23928 );
nor U124726 ( n24232, n73685, n23927 );
nor U124727 ( n23924, n23925, n23926 );
nor U124728 ( n23925, n74212, n23928 );
nor U124729 ( n23926, n74196, n23927 );
nor U124730 ( n57048, n57049, n57050 );
nor U124731 ( n57049, n74213, n57052 );
nor U124732 ( n57050, n74197, n57051 );
nand U124733 ( n57042, n57346, n57325 );
nor U124734 ( n57346, n57332, n57345 );
nand U124735 ( n23918, n24224, n24203 );
nor U124736 ( n24224, n24210, n24223 );
nor U124737 ( n24009, n73925, n23918 );
nor U124738 ( n24050, n73856, n23918 );
nor U124739 ( n24090, n73774, n23918 );
nor U124740 ( n57091, n74080, n57042 );
nor U124741 ( n57131, n73926, n57042 );
nor U124742 ( n57172, n73857, n57042 );
nor U124743 ( n57212, n73775, n57042 );
nor U124744 ( n23969, n74081, n23918 );
nor U124745 ( n57253, n73729, n57042 );
nor U124746 ( n57293, n73619, n57042 );
nor U124747 ( n57342, n73682, n57042 );
nor U124748 ( n24131, n73730, n23918 );
nor U124749 ( n24171, n73620, n23918 );
nor U124750 ( n24220, n73683, n23918 );
nor U124751 ( n23915, n74187, n23918 );
nor U124752 ( n57039, n74188, n57042 );
nand U124753 ( n23928, n24234, n24203 );
nor U124754 ( n24234, n4237, n24210 );
nand U124755 ( n57052, n57356, n57325 );
nor U124756 ( n57356, n6869, n57332 );
nand U124757 ( n28191, n28128, n28193 );
nand U124758 ( n28193, n28115, n27219 );
nand U124759 ( n61355, n61283, n61357 );
nand U124760 ( n61357, n61270, n60364 );
nand U124761 ( n35424, n35363, n35426 );
nand U124762 ( n35426, n35350, n34464 );
nand U124763 ( n70154, n70095, n70156 );
nand U124764 ( n70156, n70082, n69214 );
nand U124765 ( n57045, n57349, n57325 );
nor U124766 ( n57349, n55853, n57345 );
nand U124767 ( n23921, n24227, n24203 );
nor U124768 ( n24227, n22737, n24223 );
nor U124769 ( n24012, n73899, n23921 );
nor U124770 ( n24053, n73831, n23921 );
nor U124771 ( n24093, n73750, n23921 );
nor U124772 ( n57094, n74028, n57045 );
nor U124773 ( n57134, n73900, n57045 );
nor U124774 ( n57175, n73832, n57045 );
nor U124775 ( n57215, n73751, n57045 );
nor U124776 ( n23972, n74029, n23921 );
nor U124777 ( n57256, n73670, n57045 );
nor U124778 ( n57296, n73568, n57045 );
nor U124779 ( n57348, n73642, n57045 );
nor U124780 ( n24134, n73671, n23921 );
nor U124781 ( n24174, n73569, n23921 );
nor U124782 ( n24226, n73641, n23921 );
nor U124783 ( n23920, n74168, n23921 );
nor U124784 ( n57044, n74169, n57045 );
nand U124785 ( n23931, n24237, n24203 );
nor U124786 ( n24237, n4237, n22737 );
nand U124787 ( n57055, n57359, n57325 );
nor U124788 ( n57359, n6869, n55853 );
nor U124789 ( n24013, n24017, n24018 );
nor U124790 ( n24017, n73937, n23932 );
nor U124791 ( n24018, n73916, n23931 );
nor U124792 ( n24054, n24058, n24059 );
nor U124793 ( n24058, n73869, n23932 );
nor U124794 ( n24059, n73847, n23931 );
nor U124795 ( n24094, n24098, n24099 );
nor U124796 ( n24098, n73786, n23932 );
nor U124797 ( n24099, n73765, n23931 );
nor U124798 ( n57095, n57099, n57100 );
nor U124799 ( n57099, n74109, n57056 );
nor U124800 ( n57100, n74069, n57055 );
nor U124801 ( n57135, n57139, n57140 );
nor U124802 ( n57139, n73938, n57056 );
nor U124803 ( n57140, n73917, n57055 );
nor U124804 ( n57176, n57180, n57181 );
nor U124805 ( n57180, n73870, n57056 );
nor U124806 ( n57181, n73848, n57055 );
nor U124807 ( n57216, n57220, n57221 );
nor U124808 ( n57220, n73787, n57056 );
nor U124809 ( n57221, n73766, n57055 );
nor U124810 ( n23973, n23977, n23978 );
nor U124811 ( n23977, n74110, n23932 );
nor U124812 ( n23978, n74070, n23931 );
nor U124813 ( n57257, n57261, n57262 );
nor U124814 ( n57261, n73717, n57056 );
nor U124815 ( n57262, n73705, n57055 );
nor U124816 ( n57297, n57301, n57302 );
nor U124817 ( n57301, n73608, n57056 );
nor U124818 ( n57302, n73597, n57055 );
nor U124819 ( n57351, n57357, n57358 );
nor U124820 ( n57357, n73693, n57056 );
nor U124821 ( n57358, n73672, n57055 );
nor U124822 ( n24135, n24139, n24140 );
nor U124823 ( n24139, n73718, n23932 );
nor U124824 ( n24140, n73706, n23931 );
nor U124825 ( n24175, n24179, n24180 );
nor U124826 ( n24179, n73609, n23932 );
nor U124827 ( n24180, n73598, n23931 );
nor U124828 ( n24229, n24235, n24236 );
nor U124829 ( n24235, n73694, n23932 );
nor U124830 ( n24236, n73673, n23931 );
nor U124831 ( n23923, n23929, n23930 );
nor U124832 ( n23929, n74206, n23932 );
nor U124833 ( n23930, n74184, n23931 );
nor U124834 ( n57047, n57053, n57054 );
nor U124835 ( n57053, n74207, n57056 );
nor U124836 ( n57054, n74185, n57055 );
nand U124837 ( n23922, n24228, n24203 );
nor U124838 ( n24228, n24215, n24223 );
nand U124839 ( n57046, n57350, n57325 );
nor U124840 ( n57350, n57337, n57345 );
nor U124841 ( n47950, n74525, n47901 );
nand U124842 ( n23932, n24238, n24203 );
nor U124843 ( n24238, n4237, n24215 );
nand U124844 ( n57056, n57360, n57325 );
nor U124845 ( n57360, n6869, n57337 );
not U124846 ( n7453, n47918 );
nand U124847 ( n76045, n76647, n72927 );
nand U124848 ( n76046, n76647, n72927 );
nand U124849 ( n76115, n76501, n72928 );
nand U124850 ( n76116, n76501, n72928 );
not U124851 ( n4809, n14715 );
nor U124852 ( n16217, n74538, n73134 );
nor U124853 ( n49244, n74525, n73133 );
nand U124854 ( n70861, n76647, n72927 );
nand U124855 ( n36141, n76501, n72928 );
not U124856 ( n6124, n67562 );
not U124857 ( n4347, n25557 );
not U124858 ( n6979, n58694 );
not U124859 ( n3509, n32797 );
buf U124860 ( n76922, n76923 );
not U124861 ( n3922, n27028 );
not U124862 ( n6554, n60169 );
not U124863 ( n5679, n69025 );
not U124864 ( n5210, n14697 );
nand U124865 ( n16212, n15384, n16217 );
nand U124866 ( n49240, n48514, n49244 );
not U124867 ( n7464, n48017 );
not U124868 ( n4820, n14812 );
nor U124869 ( n49077, n73140, n74525 );
nor U124870 ( n8771, n75031, n14675 );
nor U124871 ( n46366, n46369, n74986 );
not U124872 ( n7853, n48871 );
nor U124873 ( n16023, n73141, n74538 );
not U124874 ( n5198, n15795 );
not U124875 ( n3639, n31280 );
not U124876 ( n4527, n23986 );
not U124877 ( n6267, n65530 );
not U124878 ( n7159, n57108 );
nor U124879 ( n15506, n75030, n47901 );
not U124880 ( n1799, n49029 );
not U124881 ( n2917, n38395 );
not U124882 ( n249, n57659 );
not U124883 ( n4, n24531 );
not U124884 ( n274, n57675 );
not U124885 ( n268, n57671 );
not U124886 ( n262, n57667 );
not U124887 ( n255, n57663 );
not U124888 ( n292, n57690 );
not U124889 ( n287, n57686 );
not U124890 ( n280, n57682 );
not U124891 ( n24, n24547 );
not U124892 ( n19, n24543 );
not U124893 ( n14, n24539 );
not U124894 ( n9, n24535 );
nor U124895 ( n12697, n74989, n73279 );
not U124896 ( n38, n24559 );
not U124897 ( n34, n24555 );
not U124898 ( n29, n24551 );
not U124899 ( n3458, n34184 );
not U124900 ( n6073, n68938 );
not U124901 ( n4295, n26939 );
not U124902 ( n6928, n60079 );
nor U124903 ( n61267, n73137, n74517 );
nor U124904 ( n28112, n73136, n74516 );
nor U124905 ( n70079, n73139, n74514 );
nor U124906 ( n35347, n73138, n74513 );
nand U124907 ( n15292, n15384, n15385 );
nand U124908 ( n48429, n48514, n48515 );
nor U124909 ( n25425, n25428, n75007 );
nor U124910 ( n58562, n58565, n75008 );
nor U124911 ( n32665, n32668, n75010 );
nor U124912 ( n67430, n67433, n75009 );
not U124913 ( n7917, n46369 );
nand U124914 ( n47968, n74626, n54113 );
nand U124915 ( n54113, n7794, n44889 );
nor U124916 ( n27953, n74555, n73136 );
nor U124917 ( n61106, n74556, n73137 );
nor U124918 ( n35192, n74561, n73138 );
nor U124919 ( n69928, n74562, n73139 );
not U124920 ( n4352, n25428 );
not U124921 ( n3514, n32668 );
not U124922 ( n6129, n67433 );
not U124923 ( n6984, n58565 );
nand U124924 ( n14744, n74646, n21130 );
nand U124925 ( n21130, n5139, n11178 );
nand U124926 ( n60117, n74614, n61741 );
nand U124927 ( n61741, n6862, n57332 );
nand U124928 ( n26977, n74612, n28436 );
nand U124929 ( n28436, n4229, n24210 );
nand U124930 ( n34222, n74611, n35613 );
nand U124931 ( n35613, n3392, n31504 );
nand U124932 ( n68976, n74613, n70341 );
nand U124933 ( n70341, n6007, n65754 );
nor U124934 ( n35641, n73182, n29171 );
nor U124935 ( n70367, n73183, n62893 );
not U124936 ( n7158, n57189 );
not U124937 ( n4525, n24067 );
not U124938 ( n3638, n31361 );
not U124939 ( n6265, n65611 );
not U124940 ( n3078, n34273 );
not U124941 ( n2914, n38424 );
not U124942 ( n1797, n49259 );
nand U124943 ( n12708, n73279, n74989 );
not U124944 ( n7157, n57270 );
not U124945 ( n4524, n24148 );
not U124946 ( n3637, n31442 );
not U124947 ( n6264, n65692 );
nor U124948 ( n21156, n74685, n8297 );
nor U124949 ( n54139, n74686, n42384 );
nor U124950 ( n28462, n73181, n21858 );
nor U124951 ( n61767, n73180, n54949 );
nand U124952 ( n29170, n3078, n29171 );
not U124953 ( n2912, n38456 );
not U124954 ( n1794, n49568 );
nand U124955 ( n62892, n5679, n62893 );
nor U124956 ( n68754, n73076, n68598 );
nor U124957 ( n33998, n73077, n33842 );
nor U124958 ( n14465, n73079, n14262 );
nor U124959 ( n47733, n73071, n47577 );
nor U124960 ( n26753, n73075, n26597 );
nor U124961 ( n59895, n73074, n59739 );
nor U124962 ( n21947, n75064, n73317 );
nor U124963 ( n55059, n75063, n73316 );
nor U124964 ( n63031, n75070, n73319 );
nor U124965 ( n29264, n75069, n73318 );
nand U124966 ( n63004, n63005, n63006 );
nor U124967 ( n63006, n63007, n63008 );
nor U124968 ( n63005, n63009, n63010 );
nand U124969 ( n63007, n75116, n73346 );
nand U124970 ( n29237, n29238, n29239 );
nor U124971 ( n29239, n29240, n29241 );
nor U124972 ( n29238, n29242, n29243 );
nand U124973 ( n29240, n75117, n73347 );
nand U124974 ( n42469, n42470, n42471 );
nor U124975 ( n42471, n42472, n42473 );
nor U124976 ( n42470, n42474, n42475 );
nand U124977 ( n42472, n75118, n72983 );
nand U124978 ( n21920, n21921, n21922 );
nor U124979 ( n21922, n21923, n21924 );
nor U124980 ( n21921, n21925, n21926 );
nand U124981 ( n21923, n75119, n72984 );
nand U124982 ( n55032, n55033, n55034 );
nor U124983 ( n55034, n55035, n55036 );
nor U124984 ( n55033, n55037, n55038 );
nand U124985 ( n55035, n75120, n72985 );
nand U124986 ( n8374, n8375, n8377 );
nor U124987 ( n8377, n8378, n8379 );
nor U124988 ( n8375, n8380, n8382 );
nand U124989 ( n8378, n75121, n72986 );
nand U124990 ( n62994, n75078, n73322 );
nand U124991 ( n29227, n75079, n73323 );
nand U124992 ( n42459, n75080, n73324 );
nand U124993 ( n21910, n75081, n73325 );
nand U124994 ( n55022, n75082, n73326 );
nand U124995 ( n8362, n75083, n73327 );
nand U124996 ( n62990, n62991, n62992 );
nor U124997 ( n62991, n62995, n62996 );
nor U124998 ( n62992, n62993, n62994 );
nand U124999 ( n62995, n75122, n73348 );
nand U125000 ( n29223, n29224, n29225 );
nor U125001 ( n29224, n29228, n29229 );
nor U125002 ( n29225, n29226, n29227 );
nand U125003 ( n29228, n75123, n73349 );
nand U125004 ( n42455, n42456, n42457 );
nor U125005 ( n42456, n42460, n42461 );
nor U125006 ( n42457, n42458, n42459 );
nand U125007 ( n42460, n75124, n73350 );
nand U125008 ( n21906, n21907, n21908 );
nor U125009 ( n21907, n21911, n21912 );
nor U125010 ( n21908, n21909, n21910 );
nand U125011 ( n21911, n75125, n73351 );
nand U125012 ( n55018, n55019, n55020 );
nor U125013 ( n55019, n55023, n55024 );
nor U125014 ( n55020, n55021, n55022 );
nand U125015 ( n55023, n75126, n73352 );
nand U125016 ( n8357, n8358, n8359 );
nor U125017 ( n8358, n8363, n8364 );
nor U125018 ( n8359, n8360, n8362 );
nand U125019 ( n8363, n75127, n73353 );
nand U125020 ( n63008, n75086, n73328 );
nand U125021 ( n62996, n75087, n73329 );
nand U125022 ( n29241, n75088, n73330 );
nand U125023 ( n29229, n75089, n73331 );
nand U125024 ( n42473, n75090, n72971 );
nand U125025 ( n42461, n75091, n72972 );
nand U125026 ( n21924, n75092, n72973 );
nand U125027 ( n21912, n75093, n72974 );
nand U125028 ( n55036, n75094, n72975 );
nand U125029 ( n55024, n75095, n72976 );
nand U125030 ( n8379, n75096, n72977 );
nand U125031 ( n8364, n75097, n72978 );
nand U125032 ( n63010, n75098, n73332 );
nand U125033 ( n29243, n75099, n73333 );
nand U125034 ( n55038, n75100, n72979 );
nand U125035 ( n42475, n75101, n72980 );
nand U125036 ( n21926, n75102, n72981 );
nand U125037 ( n8382, n75103, n72982 );
nor U125038 ( n62919, n73163, n62918 );
nor U125039 ( n29201, n73164, n29200 );
nor U125040 ( n42410, n72962, n42409 );
nor U125041 ( n21884, n72958, n21883 );
nor U125042 ( n54975, n72959, n54974 );
nor U125043 ( n8329, n72963, n8328 );
nand U125044 ( n62993, n75104, n73334 );
nand U125045 ( n29226, n75105, n73335 );
nand U125046 ( n42458, n75106, n73336 );
nand U125047 ( n21909, n75107, n73337 );
nand U125048 ( n55021, n75108, n73338 );
nand U125049 ( n8360, n75109, n73339 );
nor U125050 ( n62998, n62999, n63000 );
nand U125051 ( n62999, n75146, n73368 );
nand U125052 ( n63000, n75110, n73340 );
nor U125053 ( n29231, n29232, n29233 );
nand U125054 ( n29232, n75147, n73369 );
nand U125055 ( n29233, n75111, n73341 );
nor U125056 ( n42463, n42464, n42465 );
nand U125057 ( n42464, n75148, n72991 );
nand U125058 ( n42465, n75112, n73342 );
nor U125059 ( n21914, n21915, n21916 );
nand U125060 ( n21915, n75149, n72992 );
nand U125061 ( n21916, n75113, n73343 );
nor U125062 ( n55026, n55027, n55028 );
nand U125063 ( n55027, n75150, n72993 );
nand U125064 ( n55028, n75114, n73344 );
nor U125065 ( n8367, n8368, n8369 );
nand U125066 ( n8368, n75151, n72994 );
nand U125067 ( n8369, n75115, n73345 );
nand U125068 ( n63003, n63011, n63012 );
nor U125069 ( n63011, n63015, n63016 );
nor U125070 ( n63012, n63013, n63014 );
nand U125071 ( n63015, n75164, n73382 );
nand U125072 ( n29236, n29244, n29245 );
nor U125073 ( n29244, n29248, n29249 );
nor U125074 ( n29245, n29246, n29247 );
nand U125075 ( n29248, n75165, n73383 );
nand U125076 ( n42468, n42476, n42477 );
nor U125077 ( n42476, n42480, n42481 );
nor U125078 ( n42477, n42478, n42479 );
nand U125079 ( n42480, n75166, n72995 );
nand U125080 ( n21919, n21927, n21928 );
nor U125081 ( n21927, n21931, n21932 );
nor U125082 ( n21928, n21929, n21930 );
nand U125083 ( n21931, n75167, n72996 );
nand U125084 ( n55031, n55039, n55040 );
nor U125085 ( n55039, n55043, n55044 );
nor U125086 ( n55040, n55041, n55042 );
nand U125087 ( n55043, n75168, n72997 );
nand U125088 ( n8373, n8383, n8384 );
nor U125089 ( n8383, n8388, n8389 );
nor U125090 ( n8384, n8385, n8387 );
nand U125091 ( n8388, n75169, n72998 );
nand U125092 ( n63014, n75128, n73354 );
nand U125093 ( n29247, n75129, n73355 );
nand U125094 ( n42479, n75130, n73356 );
nand U125095 ( n21930, n75131, n73357 );
nand U125096 ( n55042, n75132, n73358 );
nand U125097 ( n8387, n75133, n73359 );
nor U125098 ( n62997, n63001, n63002 );
nand U125099 ( n63001, n75152, n73370 );
nand U125100 ( n63002, n75134, n73360 );
nor U125101 ( n29230, n29234, n29235 );
nand U125102 ( n29234, n75153, n73371 );
nand U125103 ( n29235, n75135, n73361 );
nor U125104 ( n42462, n42466, n42467 );
nand U125105 ( n42466, n75154, n73372 );
nand U125106 ( n42467, n75136, n73362 );
nor U125107 ( n21913, n21917, n21918 );
nand U125108 ( n21917, n75155, n73373 );
nand U125109 ( n21918, n75137, n73363 );
nor U125110 ( n55025, n55029, n55030 );
nand U125111 ( n55029, n75156, n73374 );
nand U125112 ( n55030, n75138, n73364 );
nor U125113 ( n8365, n8370, n8372 );
nand U125114 ( n8370, n75157, n73375 );
nand U125115 ( n8372, n75139, n73365 );
nand U125116 ( n8295, n4820, n8297 );
nand U125117 ( n42383, n7464, n42384 );
nand U125118 ( n63016, n75140, n73366 );
nand U125119 ( n29249, n75141, n73367 );
nand U125120 ( n42481, n75142, n72987 );
nand U125121 ( n21932, n75143, n72988 );
nand U125122 ( n55044, n75144, n72989 );
nand U125123 ( n8389, n75145, n72990 );
nand U125124 ( n21857, n3922, n21858 );
nand U125125 ( n54948, n6554, n54949 );
nand U125126 ( n63013, n75158, n73376 );
nand U125127 ( n29246, n75159, n73377 );
nand U125128 ( n42478, n75160, n73378 );
nand U125129 ( n21929, n75161, n73379 );
nand U125130 ( n55041, n75162, n73380 );
nand U125131 ( n8385, n75163, n73381 );
not U125132 ( n7155, n57371 );
not U125133 ( n4523, n24246 );
not U125134 ( n3635, n31540 );
not U125135 ( n6263, n65790 );
nor U125136 ( n46586, n74881, n73159 );
not U125137 ( n2909, n38495 );
not U125138 ( n1792, n54632 );
nor U125139 ( n9352, n9353, n5312 );
nor U125140 ( n43307, n43308, n7967 );
nor U125141 ( n64053, n64054, n6178 );
nor U125142 ( n30036, n30037, n3563 );
nor U125143 ( n22713, n22714, n4400 );
nor U125144 ( n55829, n55830, n7033 );
not U125145 ( n7154, n57392 );
not U125146 ( n4522, n24267 );
not U125147 ( n3634, n31561 );
not U125148 ( n6262, n65851 );
nand U125149 ( n14718, n76188, n73134 );
nand U125150 ( n47936, n76178, n73133 );
not U125151 ( n2929, n38527 );
not U125152 ( n1812, n54672 );
nor U125153 ( n21647, n73185, n74713 );
nand U125154 ( n14704, n76189, n14705 );
nand U125155 ( n29186, n72928, n74654 );
nand U125156 ( n47925, n76179, n47926 );
nand U125157 ( n21869, n74651, n73179 );
nand U125158 ( n8310, n74670, n73185 );
nor U125159 ( n36147, n72928, n36122 );
nand U125160 ( n42395, n74650, n73177 );
nor U125161 ( n28974, n74651, n28949 );
nor U125162 ( n54702, n74650, n54661 );
nand U125163 ( n54960, n74636, n73184 );
nand U125164 ( n62904, n72927, n74657 );
nor U125165 ( n21663, n74670, n21639 );
nand U125166 ( n40470, n73051, n73519 );
nand U125167 ( n40469, n73058, n75299 );
nand U125168 ( n49940, DIN_0_, n76930 );
and U125169 ( n48116, n49666, n49451 );
nor U125170 ( n49666, n49667, n49668 );
nor U125171 ( n49668, P2_BUF1_REG_31_, n31928 );
nor U125172 ( n49667, n49669, n49670 );
nand U125173 ( n50537, n50535, n50538 );
nand U125174 ( n50538, P3_DATAO_REG_29_, n50539 );
nand U125175 ( n50539, n76323, n50540 );
nand U125176 ( n50540, n76651, n73405 );
nand U125177 ( n43796, n49658, n49659 );
nand U125178 ( n49658, P2_BUF1_REG_30_, n76478 );
nand U125179 ( n49659, n49660, n76476 );
xnor U125180 ( n49660, n49661, n49662 );
nand U125181 ( n48498, n48499, n48500 );
nand U125182 ( n48500, P2_P1_INSTQUEUE_REG_4__6_, n48426 );
nand U125183 ( n48394, n48395, n48396 );
nand U125184 ( n48396, P2_P1_INSTQUEUE_REG_3__6_, n48344 );
nand U125185 ( n48214, n48215, n48216 );
nand U125186 ( n48216, P2_P1_INSTQUEUE_REG_1__6_, n48149 );
nand U125187 ( n48297, n48298, n48299 );
nand U125188 ( n48299, P2_P1_INSTQUEUE_REG_2__6_, n48247 );
nand U125189 ( n48106, n48107, n48108 );
nand U125190 ( n48108, P2_P1_INSTQUEUE_REG_0__6_, n48024 );
and U125191 ( n50788, n50793, n50794 );
nand U125192 ( n50794, P3_DATAO_REG_28_, n50795 );
nand U125193 ( n50795, n76323, n50796 );
nand U125194 ( n50796, n76651, n73010 );
nand U125195 ( n16983, DIN_0_, n76927 );
nand U125196 ( n17578, n17575, n17579 );
nand U125197 ( n17579, P4_DATAO_REG_29_, n17580 );
nand U125198 ( n17580, n76589, n17581 );
nand U125199 ( n17581, n76656, n73004 );
nand U125200 ( n9893, n16689, n16690 );
nand U125201 ( n16689, P1_BUF1_REG_30_, n76611 );
nand U125202 ( n16690, n16692, n76613 );
xnor U125203 ( n16692, n16693, n16694 );
nand U125204 ( n15364, n15365, n15367 );
nand U125205 ( n15367, P1_P1_INSTQUEUE_REG_4__6_, n15288 );
nand U125206 ( n15365, n15289, n82 );
nand U125207 ( n15249, n15250, n15252 );
nand U125208 ( n15252, P1_P1_INSTQUEUE_REG_3__6_, n15178 );
nand U125209 ( n15250, n15179, n82 );
nand U125210 ( n15139, n15140, n15142 );
nand U125211 ( n15142, P1_P1_INSTQUEUE_REG_2__6_, n15070 );
nand U125212 ( n15140, n15072, n82 );
nand U125213 ( n15029, n15030, n15032 );
nand U125214 ( n15032, P1_P1_INSTQUEUE_REG_1__6_, n14967 );
nand U125215 ( n15030, n14968, n82 );
nand U125216 ( n14905, n14907, n14908 );
nand U125217 ( n14908, P1_P1_INSTQUEUE_REG_0__6_, n14820 );
nand U125218 ( n14907, n82, n14822 );
and U125219 ( n14927, n16708, n16450 );
nor U125220 ( n16708, n16709, n16710 );
nor U125221 ( n16710, P1_BUF1_REG_31_, n76612 );
nor U125222 ( n16709, n16712, n16713 );
nand U125223 ( n51053, n51051, n51054 );
nand U125224 ( n51054, P3_DATAO_REG_27_, n51055 );
nand U125225 ( n51055, n76323, n51056 );
nand U125226 ( n51056, n76651, n73014 );
nand U125227 ( n49923, n8229, P3_DATAO_REG_28_ );
nand U125228 ( n54061, DIN_1_, n76930 );
and U125229 ( n17843, n17848, n17849 );
nand U125230 ( n17849, P4_DATAO_REG_28_, n17850 );
nand U125231 ( n17850, n76589, n17851 );
nand U125232 ( n17851, n76656, n73409 );
nand U125233 ( n20788, n20789, n20790 );
nand U125234 ( n20790, P4_DATAO_REG_15_, n20791 );
nand U125235 ( n20789, P4_DATAO_REG_16_, n20793 );
nand U125236 ( n20791, n16488, n20792 );
nand U125237 ( n20900, n20901, n20902 );
nand U125238 ( n20902, P4_DATAO_REG_14_, n20903 );
nand U125239 ( n20901, P4_DATAO_REG_15_, n20905 );
nand U125240 ( n20903, n16488, n20904 );
nand U125241 ( n53725, n53728, n53729 );
nand U125242 ( n53729, P3_DATAO_REG_14_, n53730 );
nand U125243 ( n53728, P3_DATAO_REG_15_, n53732 );
nand U125244 ( n53730, n49482, n53731 );
nand U125245 ( n53767, n53769, n53770 );
nand U125246 ( n53770, P3_DATAO_REG_15_, n53771 );
nand U125247 ( n53769, P3_DATAO_REG_16_, n53773 );
nand U125248 ( n53771, n49482, n53772 );
nand U125249 ( n18099, n18096, n18100 );
nand U125250 ( n18100, P4_DATAO_REG_27_, n18101 );
nand U125251 ( n18101, n76589, n18102 );
nand U125252 ( n18102, n76656, n73013 );
and U125253 ( n53865, n53861, n53867 );
nand U125254 ( n53867, P3_DATAO_REG_18_, n53868 );
nand U125255 ( n53868, n76323, n53869 );
nand U125256 ( n53869, n76652, n73002 );
nor U125257 ( n16720, n75908, n75909 );
nor U125258 ( n75908, n16726, P4_DATAO_REG_0_ );
and U125259 ( n75909, n2355, n16724 );
nand U125260 ( n53666, n53668, n53669 );
nand U125261 ( n53669, P3_DATAO_REG_13_, n53670 );
nand U125262 ( n53668, P3_DATAO_REG_14_, n53672 );
nand U125263 ( n53670, n49482, n53671 );
nand U125264 ( n50313, n76651, P3_DATAO_REG_30_ );
nand U125265 ( n49922, n50316, n50317 );
nand U125266 ( n50317, n76324, P3_DATAO_REG_30_ );
nor U125267 ( n50316, n1767, n50318 );
nor U125268 ( n50318, P3_DATAO_REG_29_, n50313 );
nand U125269 ( n50311, n50319, n76648 );
and U125270 ( n50319, n50313, P3_DATAO_REG_29_ );
nand U125271 ( n20676, n20741, n20742 );
nand U125272 ( n20742, P4_DATAO_REG_16_, n20743 );
nand U125273 ( n20741, P4_DATAO_REG_17_, n20745 );
nand U125274 ( n20743, n16488, n20744 );
nand U125275 ( n20921, n20922, n20923 );
nand U125276 ( n20923, P4_DATAO_REG_13_, n20924 );
nand U125277 ( n20922, P4_DATAO_REG_14_, n20926 );
nand U125278 ( n20924, n16488, n20925 );
nand U125279 ( n20860, n20862, n20863 );
nand U125280 ( n20863, P4_DATAO_REG_11_, n20864 );
nand U125281 ( n20862, P4_DATAO_REG_12_, n20866 );
nand U125282 ( n20864, n16488, n20865 );
and U125283 ( n53786, n53852, n8233 );
and U125284 ( n53852, n53790, P3_DATAO_REG_15_ );
nand U125285 ( n53780, n53845, n53846 );
nand U125286 ( n53846, P3_DATAO_REG_16_, n53847 );
nand U125287 ( n53845, P3_DATAO_REG_17_, n53849 );
nand U125288 ( n53847, n49482, n53848 );
nand U125289 ( n53522, n53524, n53525 );
nand U125290 ( n53525, P3_DATAO_REG_11_, n53526 );
nand U125291 ( n53524, P3_DATAO_REG_12_, n53528 );
nand U125292 ( n53526, n49482, n53527 );
nand U125293 ( n53597, n53600, n53601 );
nand U125294 ( n53601, P3_DATAO_REG_12_, n53602 );
nand U125295 ( n53600, P3_DATAO_REG_13_, n53604 );
nand U125296 ( n53602, n49482, n53603 );
nand U125297 ( n20910, n20913, n20914 );
nand U125298 ( n20914, P4_DATAO_REG_12_, n20915 );
nand U125299 ( n20913, P4_DATAO_REG_13_, n20917 );
nand U125300 ( n20915, n16488, n20916 );
nand U125301 ( n53471, n53474, n53475 );
nand U125302 ( n53475, P3_DATAO_REG_10_, n53476 );
nand U125303 ( n53474, P3_DATAO_REG_11_, n53478 );
nand U125304 ( n53476, n49482, n53477 );
nand U125305 ( n9954, n16652, n16653 );
nand U125306 ( n16652, P1_BUF1_REG_29_, n76611 );
nand U125307 ( n16653, n16654, n76613 );
xnor U125308 ( n16654, n16655, n16657 );
nand U125309 ( n15353, n15354, n15355 );
nand U125310 ( n15355, P1_P1_INSTQUEUE_REG_4__5_, n15288 );
nand U125311 ( n15354, n15289, n79 );
nand U125312 ( n15239, n15240, n15242 );
nand U125313 ( n15242, P1_P1_INSTQUEUE_REG_3__5_, n15178 );
nand U125314 ( n15240, n15179, n79 );
nand U125315 ( n15129, n15130, n15132 );
nand U125316 ( n15132, P1_P1_INSTQUEUE_REG_2__5_, n15070 );
nand U125317 ( n15130, n15072, n79 );
nand U125318 ( n15019, n15020, n15022 );
nand U125319 ( n15022, P1_P1_INSTQUEUE_REG_1__5_, n14967 );
nand U125320 ( n15020, n14968, n79 );
nand U125321 ( n20829, n20832, n20833 );
nand U125322 ( n20833, P4_DATAO_REG_10_, n20834 );
nand U125323 ( n20832, P4_DATAO_REG_11_, n20836 );
nand U125324 ( n20834, n16488, n20835 );
nand U125325 ( n14892, n14893, n14894 );
nand U125326 ( n14894, P1_P1_INSTQUEUE_REG_0__5_, n14820 );
nand U125327 ( n14893, n79, n14822 );
and U125328 ( n20662, n20667, n20668 );
nand U125329 ( n20668, P4_DATAO_REG_18_, n20669 );
nand U125330 ( n20669, n76589, n20670 );
nand U125331 ( n20670, n76655, n73408 );
nand U125332 ( n43845, n49628, n49629 );
nand U125333 ( n49628, P2_BUF1_REG_29_, n76478 );
nand U125334 ( n49629, n49630, n76476 );
nand U125335 ( n48489, n48490, n48491 );
nand U125336 ( n48491, P2_P1_INSTQUEUE_REG_4__5_, n48426 );
nand U125337 ( n48490, n48427, n342 );
nand U125338 ( n48386, n48387, n48388 );
nand U125339 ( n48388, P2_P1_INSTQUEUE_REG_3__5_, n48344 );
nand U125340 ( n48387, n48345, n342 );
nand U125341 ( n48289, n48290, n48291 );
nand U125342 ( n48291, P2_P1_INSTQUEUE_REG_2__5_, n48247 );
nand U125343 ( n48290, n48248, n342 );
nand U125344 ( n48191, n48192, n48193 );
nand U125345 ( n48193, P2_P1_INSTQUEUE_REG_1__5_, n48149 );
nand U125346 ( n48192, n48150, n342 );
nand U125347 ( n48095, n48096, n48097 );
nand U125348 ( n48097, P2_P1_INSTQUEUE_REG_0__5_, n48024 );
nand U125349 ( n48096, n342, n48025 );
nand U125350 ( n17369, n17370, n17371 );
nor U125351 ( n17370, n2882, n17372 );
nand U125352 ( n17371, P4_DATAO_REG_30_, n76590 );
and U125353 ( n17372, n73399, n17367 );
nand U125354 ( n53341, n53344, n53345 );
nand U125355 ( n53344, P3_DATAO_REG_9_, n53348 );
nand U125356 ( n53345, P3_DATAO_REG_10_, n53346 );
nand U125357 ( n53348, n49482, n53349 );
nor U125358 ( n20586, n75910, n75911 );
nand U125359 ( n75910, n20584, n8225 );
xor U125360 ( n49751, n49757, n49758 );
xor U125361 ( n49757, n50002, n50003 );
xor U125362 ( n49758, n49759, n49760 );
nand U125363 ( n50002, n8239, P3_DATAO_REG_8_ );
and U125364 ( n53640, n53703, n8234 );
and U125365 ( n53703, n53644, P3_DATAO_REG_12_ );
nand U125366 ( n20483, n20486, n20487 );
nand U125367 ( n20486, P4_DATAO_REG_9_, n20490 );
nand U125368 ( n20487, P4_DATAO_REG_10_, n20488 );
nand U125369 ( n20490, n16488, n20491 );
nand U125370 ( n51476, n51474, n51477 );
nand U125371 ( n51477, P3_DATAO_REG_25_, n51478 );
nand U125372 ( n51478, n76323, n51479 );
nand U125373 ( n51479, n76651, n73016 );
nand U125374 ( n52886, n52884, n52887 );
nand U125375 ( n52887, P3_DATAO_REG_21_, n52888 );
nand U125376 ( n52888, n76323, n52889 );
nand U125377 ( n52889, n76651, n73401 );
nand U125378 ( n53878, n53876, n53879 );
nand U125379 ( n53879, P3_DATAO_REG_19_, n53880 );
nand U125380 ( n53880, n76323, n53881 );
nand U125381 ( n53881, n76652, n73403 );
and U125382 ( n53826, n53831, n53832 );
nand U125383 ( n53832, P3_DATAO_REG_20_, n53833 );
nand U125384 ( n53833, n76323, n53834 );
nand U125385 ( n53834, n76652, n73005 );
nand U125386 ( n16988, P4_DATAO_REG_28_, n8220 );
nand U125387 ( n48480, n48481, n48482 );
nand U125388 ( n48482, P2_P1_INSTQUEUE_REG_4__4_, n48426 );
nand U125389 ( n48481, n48427, n339 );
nand U125390 ( n43893, n49600, n49601 );
nand U125391 ( n49600, P2_BUF1_REG_28_, n76478 );
nand U125392 ( n49601, n49602, n76476 );
xor U125393 ( n49602, n49603, n49604 );
nand U125394 ( n48378, n48379, n48380 );
nand U125395 ( n48380, P2_P1_INSTQUEUE_REG_3__4_, n48344 );
nand U125396 ( n48379, n48345, n339 );
nand U125397 ( n48281, n48282, n48283 );
nand U125398 ( n48283, P2_P1_INSTQUEUE_REG_2__4_, n48247 );
nand U125399 ( n48282, n48248, n339 );
nand U125400 ( n48183, n48184, n48185 );
nand U125401 ( n48185, P2_P1_INSTQUEUE_REG_1__4_, n48149 );
nand U125402 ( n48184, n48150, n339 );
nand U125403 ( n53141, n53235, n53236 );
nand U125404 ( n53236, P3_DATAO_REG_8_, n53237 );
nand U125405 ( n53235, P3_DATAO_REG_9_, n53239 );
nand U125406 ( n53237, n49482, n53238 );
and U125407 ( n50529, n50799, P3_DATAO_REG_27_ );
nand U125408 ( n48084, n48085, n48086 );
nand U125409 ( n48086, P2_P1_INSTQUEUE_REG_0__4_, n48024 );
nand U125410 ( n48085, n339, n48025 );
nand U125411 ( n17374, DIN_1_, n76927 );
nand U125412 ( n9970, n16615, n16617 );
nand U125413 ( n16615, P1_BUF1_REG_28_, n76611 );
nand U125414 ( n16617, n16618, n76613 );
xor U125415 ( n16618, n16619, n16620 );
nand U125416 ( n15335, n15337, n15338 );
nand U125417 ( n15338, P1_P1_INSTQUEUE_REG_4__4_, n15288 );
nand U125418 ( n15337, n15289, n76 );
nand U125419 ( n15229, n15230, n15232 );
nand U125420 ( n15232, P1_P1_INSTQUEUE_REG_3__4_, n15178 );
nand U125421 ( n15230, n15179, n76 );
nand U125422 ( n15119, n15120, n15122 );
nand U125423 ( n15122, P1_P1_INSTQUEUE_REG_2__4_, n15070 );
nand U125424 ( n15120, n15072, n76 );
nand U125425 ( n15009, n15010, n15012 );
nand U125426 ( n15012, P1_P1_INSTQUEUE_REG_1__4_, n14967 );
nand U125427 ( n15010, n14968, n76 );
nand U125428 ( n14878, n14879, n14880 );
nand U125429 ( n14880, P1_P1_INSTQUEUE_REG_0__4_, n14820 );
nand U125430 ( n14879, n76, n14822 );
nor U125431 ( n20264, n75912, n75913 );
nand U125432 ( n75912, n20262, n8219 );
or U125433 ( n52025, n52478, n75914 );
and U125434 ( n75914, n8237, P3_DATAO_REG_12_ );
and U125435 ( n49931, DIN_2_, n76929 );
nand U125436 ( n50312, n76319, P3_DATAO_REG_28_ );
nand U125437 ( n52997, n53135, n53136 );
nand U125438 ( n53136, P3_DATAO_REG_7_, n53137 );
nand U125439 ( n53135, P3_DATAO_REG_8_, n53139 );
nand U125440 ( n53137, n49482, n53138 );
and U125441 ( n50802, n50799, P3_DATAO_REG_25_ );
nand U125442 ( n43974, n49555, n49556 );
nand U125443 ( n49555, P2_BUF1_REG_27_, n76478 );
nand U125444 ( n49556, n49557, n76476 );
xor U125445 ( n49557, n49558, n49559 );
nand U125446 ( n48471, n48472, n48473 );
nand U125447 ( n48473, P2_P1_INSTQUEUE_REG_4__3_, n48426 );
nand U125448 ( n48472, n48427, n335 );
nand U125449 ( n48370, n48371, n48372 );
nand U125450 ( n48372, P2_P1_INSTQUEUE_REG_3__3_, n48344 );
nand U125451 ( n48371, n48345, n335 );
nand U125452 ( n48273, n48274, n48275 );
nand U125453 ( n48275, P2_P1_INSTQUEUE_REG_2__3_, n48247 );
nand U125454 ( n48274, n48248, n335 );
nand U125455 ( n48175, n48176, n48177 );
nand U125456 ( n48177, P2_P1_INSTQUEUE_REG_1__3_, n48149 );
nand U125457 ( n48176, n48150, n335 );
nand U125458 ( n48059, n48060, n48061 );
nand U125459 ( n48061, P2_P1_INSTQUEUE_REG_0__3_, n48024 );
nand U125460 ( n48060, n335, n48025 );
nand U125461 ( n20595, n20592, n20596 );
nand U125462 ( n20596, P4_DATAO_REG_19_, n20597 );
nand U125463 ( n20597, n76589, n20598 );
nand U125464 ( n20598, n76655, n73007 );
and U125465 ( n19911, n20270, P4_DATAO_REG_15_ );
nor U125466 ( n20270, n2767, n76587 );
and U125467 ( n20295, n20300, n20301 );
nand U125468 ( n20301, P4_DATAO_REG_20_, n20302 );
nand U125469 ( n20302, n76589, n20303 );
nand U125470 ( n20303, n76655, n73011 );
nand U125471 ( n52995, n53976, n53977 );
nand U125472 ( n53977, P3_DATAO_REG_6_, n53978 );
nand U125473 ( n53976, P3_DATAO_REG_7_, n53980 );
nand U125474 ( n53978, n49482, n53979 );
nand U125475 ( n19933, n19930, n19934 );
nand U125476 ( n19934, P4_DATAO_REG_21_, n19935 );
nand U125477 ( n19935, n76589, n19936 );
nand U125478 ( n19936, n76655, n73407 );
nand U125479 ( n20186, n20381, n20382 );
nand U125480 ( n20382, P4_DATAO_REG_8_, n20383 );
nand U125481 ( n20381, P4_DATAO_REG_9_, n20385 );
nand U125482 ( n20383, n16488, n20384 );
xor U125483 ( n16796, n16802, n16803 );
xor U125484 ( n16802, n17048, n17049 );
xor U125485 ( n16803, n16804, n16805 );
nand U125486 ( n17048, n8213, P4_DATAO_REG_8_ );
xor U125487 ( n49766, n49771, n49772 );
xor U125488 ( n49771, n49987, n49988 );
xor U125489 ( n49772, n49773, n49774 );
nand U125490 ( n49987, n49990, P3_DATAO_REG_13_ );
nand U125491 ( n18512, n18509, n18513 );
nand U125492 ( n18513, P4_DATAO_REG_25_, n18514 );
nand U125493 ( n18514, n76589, n18515 );
nand U125494 ( n18515, n76656, n73417 );
nand U125495 ( n10058, n16579, n16580 );
nand U125496 ( n16579, P1_BUF1_REG_27_, n76611 );
nand U125497 ( n16580, n16582, n76613 );
xnor U125498 ( n16582, n16583, n16584 );
nand U125499 ( n15324, n15325, n15327 );
nand U125500 ( n15327, P1_P1_INSTQUEUE_REG_4__3_, n15288 );
nand U125501 ( n15325, n15289, n73 );
nand U125502 ( n15219, n15220, n15222 );
nand U125503 ( n15222, P1_P1_INSTQUEUE_REG_3__3_, n15178 );
nand U125504 ( n15220, n15179, n73 );
nand U125505 ( n15109, n15110, n15112 );
nand U125506 ( n15112, P1_P1_INSTQUEUE_REG_2__3_, n15070 );
nand U125507 ( n15110, n15072, n73 );
nand U125508 ( n14999, n15000, n15002 );
nand U125509 ( n15002, P1_P1_INSTQUEUE_REG_1__3_, n14967 );
nand U125510 ( n15000, n14968, n73 );
nand U125511 ( n14864, n14865, n14867 );
nand U125512 ( n14867, P1_P1_INSTQUEUE_REG_0__3_, n14820 );
nand U125513 ( n14865, n73, n14822 );
nand U125514 ( n51615, n51613, n51616 );
nand U125515 ( n51616, P3_DATAO_REG_24_, n51617 );
nand U125516 ( n51617, n76323, n51618 );
nand U125517 ( n51618, n76651, n73416 );
and U125518 ( n50534, n76319, P3_DATAO_REG_27_ );
and U125519 ( n53675, n53727, P3_DATAO_REG_13_ );
nand U125520 ( n20042, n20179, n20180 );
nand U125521 ( n20180, P4_DATAO_REG_7_, n20181 );
nand U125522 ( n20179, P4_DATAO_REG_8_, n20183 );
nand U125523 ( n20181, n16488, n20182 );
and U125524 ( n53735, n53727, P3_DATAO_REG_15_ );
nand U125525 ( n19069, n19295, n19296 );
nand U125526 ( n19296, P4_DATAO_REG_12_, n8215 );
nand U125527 ( n20039, n21080, n21081 );
nand U125528 ( n21081, P4_DATAO_REG_6_, n21082 );
nand U125529 ( n21080, P4_DATAO_REG_7_, n21084 );
nand U125530 ( n21082, n16488, n21083 );
and U125531 ( n53857, n53866, P3_DATAO_REG_16_ );
nand U125532 ( n53972, n54057, n54058 );
nand U125533 ( n54058, P3_DATAO_REG_5_, n54059 );
nand U125534 ( n54057, P3_DATAO_REG_6_, n54062 );
nand U125535 ( n54059, n49482, n54060 );
and U125536 ( n53607, n53599, P3_DATAO_REG_13_ );
nand U125537 ( n20747, n20748, P4_DATAO_REG_16_ );
nor U125538 ( n20748, n18105, n75911 );
and U125539 ( n53531, n53599, P3_DATAO_REG_11_ );
and U125540 ( n53481, n53473, P3_DATAO_REG_11_ );
nand U125541 ( n44019, n49525, n49526 );
nand U125542 ( n49525, P2_BUF1_REG_26_, n76478 );
nand U125543 ( n49526, n49527, n31928 );
xor U125544 ( n49527, n49528, n49529 );
nand U125545 ( n48462, n48463, n48464 );
nand U125546 ( n48464, P2_P1_INSTQUEUE_REG_4__2_, n48426 );
nand U125547 ( n48463, n48427, n330 );
nand U125548 ( n48362, n48363, n48364 );
nand U125549 ( n48364, P2_P1_INSTQUEUE_REG_3__2_, n48344 );
nand U125550 ( n48363, n48345, n330 );
nand U125551 ( n48265, n48266, n48267 );
nand U125552 ( n48267, P2_P1_INSTQUEUE_REG_2__2_, n48247 );
nand U125553 ( n48266, n48248, n330 );
nand U125554 ( n48167, n48168, n48169 );
nand U125555 ( n48169, P2_P1_INSTQUEUE_REG_1__2_, n48149 );
nand U125556 ( n48168, n48150, n330 );
and U125557 ( n17585, P4_DATAO_REG_27_, n17854 );
and U125558 ( n53351, n53473, P3_DATAO_REG_9_ );
nand U125559 ( n48048, n48049, n48050 );
nand U125560 ( n48050, P2_P1_INSTQUEUE_REG_0__2_, n48024 );
nand U125561 ( n48049, n330, n48025 );
and U125562 ( n20734, P4_DATAO_REG_15_, n20786 );
xor U125563 ( n16811, n16816, n16817 );
xor U125564 ( n16816, n17033, n17034 );
xor U125565 ( n16817, n16818, n16819 );
nand U125566 ( n17033, n17036, P4_DATAO_REG_13_ );
nand U125567 ( n51287, n76651, P3_DATAO_REG_26_ );
nand U125568 ( n51288, n51295, n76648 );
and U125569 ( n51295, n51287, P3_DATAO_REG_25_ );
nand U125570 ( n51291, n51292, n51293 );
nand U125571 ( n51293, n76324, P3_DATAO_REG_26_ );
nor U125572 ( n51292, n1752, n51294 );
nor U125573 ( n51294, P3_DATAO_REG_25_, n51287 );
buf U125574 ( n76320, n49911 );
nand U125575 ( n49911, DIN_4_, n76930 );
nand U125576 ( n52001, n8229, P3_DATAO_REG_21_ );
nand U125577 ( n21077, n21100, n21101 );
nand U125578 ( n21101, P4_DATAO_REG_5_, n21102 );
nand U125579 ( n21100, P4_DATAO_REG_6_, n21104 );
nand U125580 ( n21102, n16488, n21103 );
nand U125581 ( n18655, n18652, n18656 );
nand U125582 ( n18656, P4_DATAO_REG_24_, n18657 );
nand U125583 ( n18657, n76589, n18658 );
nand U125584 ( n18658, n76655, n73000 );
nand U125585 ( n50789, n76319, P3_DATAO_REG_26_ );
nand U125586 ( n54033, n54049, n54050 );
nand U125587 ( n54050, P3_DATAO_REG_4_, n54051 );
nand U125588 ( n54049, P3_DATAO_REG_5_, n54053 );
nand U125589 ( n54051, n49482, n54052 );
and U125590 ( n20783, n20786, P4_DATAO_REG_13_ );
and U125591 ( n17838, n17854, P4_DATAO_REG_25_ );
and U125592 ( n20839, P4_DATAO_REG_11_, n20831 );
nand U125593 ( n16974, DIN_2_, n76928 );
buf U125594 ( n76928, SEL );
and U125595 ( n51050, n76319, P3_DATAO_REG_25_ );
and U125596 ( n20896, P4_DATAO_REG_13_, n20912 );
nand U125597 ( n10114, n16542, n16543 );
nand U125598 ( n16542, P1_BUF1_REG_26_, n76610 );
nand U125599 ( n16543, n16544, n76613 );
xor U125600 ( n16544, n16545, n16547 );
nand U125601 ( n15313, n15314, n15315 );
nand U125602 ( n15315, P1_P1_INSTQUEUE_REG_4__2_, n15288 );
nand U125603 ( n15314, n15289, n70 );
nand U125604 ( n15200, n15202, n15203 );
nand U125605 ( n15203, P1_P1_INSTQUEUE_REG_3__2_, n15178 );
nand U125606 ( n15202, n15179, n70 );
nand U125607 ( n15099, n15100, n15102 );
nand U125608 ( n15102, P1_P1_INSTQUEUE_REG_2__2_, n15070 );
nand U125609 ( n15100, n15072, n70 );
nand U125610 ( n14989, n14990, n14992 );
nand U125611 ( n14992, P1_P1_INSTQUEUE_REG_1__2_, n14967 );
nand U125612 ( n14990, n14968, n70 );
nand U125613 ( n14850, n14852, n14853 );
nand U125614 ( n14853, P1_P1_INSTQUEUE_REG_0__2_, n14820 );
nand U125615 ( n14852, n70, n14822 );
nor U125616 ( n50953, n51181, n49989 );
nand U125617 ( n51181, n50951, P3_DATAO_REG_7_ );
nand U125618 ( n44065, n49496, n49497 );
nand U125619 ( n49496, P2_BUF1_REG_25_, n76478 );
nand U125620 ( n49497, n49498, n31928 );
xor U125621 ( n49498, n49499, n49500 );
nand U125622 ( n48437, n48438, n48439 );
nand U125623 ( n48439, P2_P1_INSTQUEUE_REG_4__1_, n48426 );
nand U125624 ( n48438, n48427, n327 );
nand U125625 ( n51998, n76651, P3_DATAO_REG_23_ );
nand U125626 ( n52000, n52002, n52003 );
nand U125627 ( n52003, n76324, P3_DATAO_REG_23_ );
nor U125628 ( n52002, n1724, n52004 );
nor U125629 ( n52004, P3_DATAO_REG_22_, n51998 );
nand U125630 ( n51996, n52005, n76648 );
and U125631 ( n52005, n51998, P3_DATAO_REG_22_ );
nand U125632 ( n48354, n48355, n48356 );
nand U125633 ( n48356, P2_P1_INSTQUEUE_REG_3__1_, n48344 );
nand U125634 ( n48355, n48345, n327 );
nand U125635 ( n48257, n48258, n48259 );
nand U125636 ( n48259, P2_P1_INSTQUEUE_REG_2__1_, n48247 );
nand U125637 ( n48258, n48248, n327 );
nand U125638 ( n48159, n48160, n48161 );
nand U125639 ( n48161, P2_P1_INSTQUEUE_REG_1__1_, n48149 );
nand U125640 ( n48160, n48150, n327 );
nand U125641 ( n52453, n76651, P3_DATAO_REG_22_ );
nand U125642 ( n52455, n52456, n52457 );
nand U125643 ( n52457, n76324, P3_DATAO_REG_22_ );
nor U125644 ( n52456, n1710, n52458 );
nor U125645 ( n52458, P3_DATAO_REG_21_, n52453 );
nand U125646 ( n52451, n52459, n76649 );
and U125647 ( n52459, n52453, P3_DATAO_REG_21_ );
nand U125648 ( n48037, n48038, n48039 );
nand U125649 ( n48039, P2_P1_INSTQUEUE_REG_0__1_, n48024 );
nand U125650 ( n48038, n327, n48025 );
nand U125651 ( n18335, n18336, n18337 );
nor U125652 ( n18336, n18333, n18338 );
nand U125653 ( n18337, P4_DATAO_REG_26_, n76590 );
nor U125654 ( n18338, P4_DATAO_REG_25_, n18332 );
and U125655 ( n20493, n20831, P4_DATAO_REG_9_ );
and U125656 ( n52462, n52892, P3_DATAO_REG_20_ );
and U125657 ( n20869, n20912, P4_DATAO_REG_11_ );
nand U125658 ( n21049, n21093, n21094 );
nand U125659 ( n21094, P4_DATAO_REG_4_, n21095 );
nand U125660 ( n21093, P4_DATAO_REG_5_, n21097 );
nand U125661 ( n21095, n16488, n21096 );
and U125662 ( n53839, n53866, P3_DATAO_REG_18_ );
and U125663 ( n51299, n51482, P3_DATAO_REG_24_ );
and U125664 ( n52878, n52892, P3_DATAO_REG_18_ );
nand U125665 ( n54025, n54027, n54028 );
nand U125666 ( n54028, P3_DATAO_REG_3_, n54029 );
nand U125667 ( n54027, P3_DATAO_REG_4_, n54031 );
nand U125668 ( n54029, n49482, n54030 );
and U125669 ( n53768, n76318, P3_DATAO_REG_14_ );
and U125670 ( n20603, n20601, P4_DATAO_REG_16_ );
and U125671 ( n53726, n76318, P3_DATAO_REG_13_ );
nand U125672 ( n17366, n17373, P4_DATAO_REG_29_ );
nor U125673 ( n17373, n17367, n17374 );
and U125674 ( n53667, n76318, P3_DATAO_REG_12_ );
nand U125675 ( n53862, n76319, P3_DATAO_REG_16_ );
nand U125676 ( n53778, n76319, P3_DATAO_REG_15_ );
nor U125677 ( n17995, n18225, n17035 );
nand U125678 ( n18225, n17993, P4_DATAO_REG_7_ );
nand U125679 ( n19370, n19371, n19372 );
nor U125680 ( n19371, n2827, n19373 );
nand U125681 ( n19372, n76590, P4_DATAO_REG_22_ );
and U125682 ( n19373, n73006, n19368 );
and U125683 ( n20388, n20485, P4_DATAO_REG_9_ );
nor U125684 ( n20485, n18105, n73418 );
and U125685 ( n53598, n76318, P3_DATAO_REG_11_ );
nand U125686 ( n49887, n8227, P3_DATAO_REG_25_ );
nand U125687 ( n18332, P4_DATAO_REG_26_, n76654 );
nor U125688 ( n18333, n75915, n75916 );
nand U125689 ( n75915, n18332, n8222 );
nand U125690 ( n51289, n76319, P3_DATAO_REG_24_ );
nand U125691 ( n44112, n49463, n49464 );
nand U125692 ( n49463, P2_BUF1_REG_24_, n76477 );
nand U125693 ( n49464, n49465, n31928 );
xnor U125694 ( n49465, n49466, n49467 );
nand U125695 ( n48423, n48424, n48425 );
nand U125696 ( n48425, P2_P1_INSTQUEUE_REG_4__0_, n48426 );
nand U125697 ( n48424, n48427, n324 );
nand U125698 ( n48341, n48342, n48343 );
nand U125699 ( n48343, P2_P1_INSTQUEUE_REG_3__0_, n48344 );
nand U125700 ( n48342, n48345, n324 );
nand U125701 ( n48244, n48245, n48246 );
nand U125702 ( n48246, P2_P1_INSTQUEUE_REG_2__0_, n48247 );
nand U125703 ( n48245, n48248, n324 );
nand U125704 ( n48146, n48147, n48148 );
nand U125705 ( n48148, P2_P1_INSTQUEUE_REG_1__0_, n48149 );
nand U125706 ( n48147, n48150, n324 );
nand U125707 ( n21040, n21042, n21043 );
nand U125708 ( n21043, P4_DATAO_REG_3_, n21044 );
nand U125709 ( n21042, P4_DATAO_REG_4_, n21046 );
nand U125710 ( n21044, n16488, n21045 );
nand U125711 ( n48021, n48022, n48023 );
nand U125712 ( n48023, P2_P1_INSTQUEUE_REG_0__0_, n48024 );
nand U125713 ( n48022, n324, n48025 );
nand U125714 ( n19048, n19050, n19051 );
nor U125715 ( n19050, n2839, n19052 );
nand U125716 ( n19051, P4_DATAO_REG_23_, n76590 );
and U125717 ( n19052, n73398, n19046 );
and U125718 ( n53523, n76318, P3_DATAO_REG_10_ );
and U125719 ( n53472, n76318, P3_DATAO_REG_9_ );
nand U125720 ( n19049, P4_DATAO_REG_21_, n8220 );
nand U125721 ( n10177, n16505, n16507 );
nand U125722 ( n16505, P1_BUF1_REG_25_, n76610 );
nand U125723 ( n16507, n16508, n76613 );
xor U125724 ( n16508, n16509, n16510 );
nand U125725 ( n15302, n15303, n15304 );
nand U125726 ( n15304, P1_P1_INSTQUEUE_REG_4__1_, n15288 );
nand U125727 ( n15303, n15289, n67 );
nand U125728 ( n15190, n15192, n15193 );
nand U125729 ( n15193, P1_P1_INSTQUEUE_REG_3__1_, n15178 );
nand U125730 ( n15192, n15179, n67 );
nand U125731 ( n15089, n15090, n15092 );
nand U125732 ( n15092, P1_P1_INSTQUEUE_REG_2__1_, n15070 );
nand U125733 ( n15090, n15072, n67 );
nand U125734 ( n14979, n14980, n14982 );
nand U125735 ( n14982, P1_P1_INSTQUEUE_REG_1__1_, n14967 );
nand U125736 ( n14980, n14968, n67 );
nand U125737 ( n14837, n14838, n14839 );
nand U125738 ( n14839, P1_P1_INSTQUEUE_REG_0__1_, n14820 );
nand U125739 ( n14838, n67, n14822 );
and U125740 ( n18108, n18340, P4_DATAO_REG_25_ );
nor U125741 ( n18340, n18105, n73417 );
nand U125742 ( n53689, n8233, P3_DATAO_REG_13_ );
and U125743 ( n51468, n51482, P3_DATAO_REG_22_ );
nand U125744 ( n53545, n8233, P3_DATAO_REG_11_ );
and U125745 ( n53342, n76318, P3_DATAO_REG_8_ );
and U125746 ( n20290, P4_DATAO_REG_18_, n20601 );
nand U125747 ( n53621, n8233, P3_DATAO_REG_12_ );
nand U125748 ( n17575, n17582, P4_DATAO_REG_28_ );
nor U125749 ( n17582, n17583, n17374 );
and U125750 ( n19377, P4_DATAO_REG_20_, n19939 );
nand U125751 ( n51997, n76319, P3_DATAO_REG_21_ );
nand U125752 ( n44210, n51672, n51673 );
nand U125753 ( n51672, P2_BUF1_REG_23_, n76477 );
nand U125754 ( n51673, n51674, n76476 );
xnor U125755 ( n51674, n50620, n51675 );
nand U125756 ( n54008, n54011, n54012 );
nand U125757 ( n54012, P3_DATAO_REG_2_, n54013 );
nand U125758 ( n54011, P3_DATAO_REG_3_, n54015 );
nand U125759 ( n54013, n49482, n54014 );
nand U125760 ( n52452, n76319, P3_DATAO_REG_20_ );
nand U125761 ( n48697, n48698, n48699 );
nor U125762 ( n48699, n48700, n48701 );
nor U125763 ( n48698, n48709, n48710 );
and U125764 ( n48700, n48624, P2_P1_INSTQUEUE_REG_6__7_ );
nand U125765 ( n48603, n48604, n48605 );
nor U125766 ( n48605, n48606, n48607 );
nor U125767 ( n48604, n48615, n48616 );
and U125768 ( n48606, n48530, P2_P1_INSTQUEUE_REG_5__7_ );
nand U125769 ( n49063, n49064, n49065 );
nor U125770 ( n49065, n49066, n49067 );
nor U125771 ( n49064, n49075, n49076 );
and U125772 ( n49066, n48990, P2_P1_INSTQUEUE_REG_10__7_ );
nand U125773 ( n48968, n48969, n48970 );
nor U125774 ( n48970, n48971, n48972 );
nor U125775 ( n48969, n48980, n48981 );
and U125776 ( n48971, n48891, P2_P1_INSTQUEUE_REG_9__7_ );
nand U125777 ( n49332, n49333, n49334 );
nor U125778 ( n49334, n49335, n49336 );
nor U125779 ( n49333, n49344, n49345 );
and U125780 ( n49335, n49275, P2_P1_INSTQUEUE_REG_13__7_ );
nand U125781 ( n49425, n49426, n49427 );
nor U125782 ( n49427, n49428, n49429 );
nor U125783 ( n49426, n49437, n49438 );
and U125784 ( n49428, n49353, P2_P1_INSTQUEUE_REG_14__7_ );
and U125785 ( n20188, n20380, P4_DATAO_REG_8_ );
nor U125786 ( n20380, n18105, n73018 );
and U125787 ( n53875, n76318, P3_DATAO_REG_17_ );
and U125788 ( n19941, n19939, P4_DATAO_REG_18_ );
and U125789 ( n51473, n76319, P3_DATAO_REG_23_ );
and U125790 ( n18343, P4_DATAO_REG_24_, n18518 );
nand U125791 ( n53334, n8233, P3_DATAO_REG_9_ );
and U125792 ( n53144, n76318, P3_DATAO_REG_7_ );
and U125793 ( n52883, n76319, P3_DATAO_REG_19_ );
nand U125794 ( n17340, P4_DATAO_REG_26_, n76583 );
and U125795 ( n16957, DIN_4_, n76927 );
nand U125796 ( n53827, n76319, P3_DATAO_REG_18_ );
and U125797 ( n20044, n20178, P4_DATAO_REG_7_ );
nor U125798 ( n20178, n73420, n18105 );
nand U125799 ( n10235, n16464, n16465 );
nand U125800 ( n16464, P1_BUF1_REG_24_, n76610 );
nand U125801 ( n16465, n16467, n76612 );
xnor U125802 ( n16467, n16468, n16469 );
nand U125803 ( n15284, n15285, n15287 );
nand U125804 ( n15287, P1_P1_INSTQUEUE_REG_4__0_, n15288 );
nand U125805 ( n15285, n15289, n64 );
nand U125806 ( n15174, n15175, n15177 );
nand U125807 ( n15177, P1_P1_INSTQUEUE_REG_3__0_, n15178 );
nand U125808 ( n15175, n15179, n64 );
nand U125809 ( n15067, n15068, n15069 );
nand U125810 ( n15069, P1_P1_INSTQUEUE_REG_2__0_, n15070 );
nand U125811 ( n15068, n15072, n64 );
nand U125812 ( n14963, n14964, n14965 );
nand U125813 ( n14965, P1_P1_INSTQUEUE_REG_1__0_, n14967 );
nand U125814 ( n14964, n14968, n64 );
nand U125815 ( n53225, n8233, P3_DATAO_REG_8_ );
nand U125816 ( n14817, n14818, n14819 );
nand U125817 ( n14819, P1_P1_INSTQUEUE_REG_0__0_, n14820 );
nand U125818 ( n14818, n64, n14822 );
and U125819 ( n53000, n76319, P3_DATAO_REG_6_ );
buf U125820 ( n76315, n49943 );
nand U125821 ( n49943, DIN_6_, n76930 );
nand U125822 ( n17848, n17852, P4_DATAO_REG_27_ );
nor U125823 ( n17852, n17853, n17374 );
nand U125824 ( n21009, n21012, n21013 );
nand U125825 ( n21013, P4_DATAO_REG_2_, n21014 );
nand U125826 ( n21012, P4_DATAO_REG_3_, n21016 );
nand U125827 ( n21014, n16488, n21015 );
and U125828 ( n52996, n76318, P3_DATAO_REG_5_ );
and U125829 ( n54018, n54010, P3_DATAO_REG_3_ );
nand U125830 ( n18096, n18103, P4_DATAO_REG_26_ );
nor U125831 ( n18103, n18104, n17374 );
nand U125832 ( n53125, n8233, P3_DATAO_REG_7_ );
nand U125833 ( n10358, n18716, n18717 );
nand U125834 ( n18716, P1_BUF1_REG_23_, n76611 );
nand U125835 ( n18717, n18718, n76613 );
xnor U125836 ( n18718, n17664, n18719 );
nor U125837 ( n21075, n75917, n75919 );
or U125838 ( n75917, n73020, n18105 );
nand U125839 ( n16104, n16105, n16107 );
nor U125840 ( n16107, n16108, n16109 );
nor U125841 ( n16105, n16119, n16120 );
and U125842 ( n16108, n16033, P1_P1_INSTQUEUE_REG_11__7_ );
nand U125843 ( n16005, n16007, n16008 );
nor U125844 ( n16008, n16009, n16010 );
nor U125845 ( n16007, n16020, n16022 );
and U125846 ( n16009, n15925, P1_P1_INSTQUEUE_REG_10__7_ );
nand U125847 ( n15898, n15899, n15900 );
nor U125848 ( n15900, n15902, n15903 );
nor U125849 ( n15899, n15913, n15914 );
and U125850 ( n15902, n15820, P1_P1_INSTQUEUE_REG_9__7_ );
nand U125851 ( n15583, n15584, n15585 );
nor U125852 ( n15585, n15587, n15588 );
nor U125853 ( n15584, n15598, n15599 );
and U125854 ( n15587, n15512, P1_P1_INSTQUEUE_REG_6__7_ );
nand U125855 ( n15485, n15487, n15488 );
nor U125856 ( n15488, n15489, n15490 );
nor U125857 ( n15487, n15500, n15502 );
and U125858 ( n15489, n15405, P1_P1_INSTQUEUE_REG_5__7_ );
nand U125859 ( n16315, n16317, n16318 );
nor U125860 ( n16318, n16319, n16320 );
nor U125861 ( n16317, n16329, n16330 );
and U125862 ( n16319, n16235, P1_P1_INSTQUEUE_REG_13__7_ );
nand U125863 ( n16418, n16419, n16420 );
nor U125864 ( n16420, n16422, n16423 );
nor U125865 ( n16419, n16433, n16434 );
and U125866 ( n16422, n16340, P1_P1_INSTQUEUE_REG_14__7_ );
and U125867 ( n51612, n76319, P3_DATAO_REG_22_ );
and U125868 ( n18521, n18518, P4_DATAO_REG_22_ );
nand U125869 ( n16956, DIN_5_, n76928 );
nand U125870 ( n17562, P4_DATAO_REG_25_, n76583 );
nand U125871 ( n53010, n8233, P3_DATAO_REG_6_ );
and U125872 ( n53973, n76318, P3_DATAO_REG_4_ );
nand U125873 ( n20779, P4_DATAO_REG_13_, n8225 );
nand U125874 ( n20892, P4_DATAO_REG_12_, n8225 );
nand U125875 ( n52752, n8233, P3_DATAO_REG_5_ );
nand U125876 ( n44253, n49649, n49650 );
nand U125877 ( n49649, P2_BUF1_REG_22_, n76478 );
nand U125878 ( n49650, n49651, n76476 );
xor U125879 ( n49651, n49652, n49653 );
nand U125880 ( n20667, n20671, P4_DATAO_REG_17_ );
nor U125881 ( n20671, n20672, n17374 );
nand U125882 ( n20822, P4_DATAO_REG_10_, n8225 );
nand U125883 ( n20883, P4_DATAO_REG_11_, n8225 );
nor U125884 ( n21051, n75918, n75919 );
or U125885 ( n75918, n73022, n18105 );
xor U125886 ( n16884, n16892, n16893 );
xor U125887 ( n16892, n17012, n17013 );
xor U125888 ( n16893, n16894, n16895 );
nand U125889 ( n17012, P4_DATAO_REG_19_, n76170 );
nand U125890 ( n20685, P4_DATAO_REG_13_, n76581 );
nand U125891 ( n20769, P4_DATAO_REG_11_, n76581 );
and U125892 ( n54036, n76318, P3_DATAO_REG_3_ );
nand U125893 ( n53962, n8233, P3_DATAO_REG_4_ );
nand U125894 ( n20476, P4_DATAO_REG_9_, n8225 );
and U125895 ( n53913, n54010, P3_DATAO_REG_1_ );
nand U125896 ( n53499, n8227, P3_DATAO_REG_10_ );
nand U125897 ( n53559, n8227, P3_DATAO_REG_11_ );
nand U125898 ( n53633, n8227, P3_DATAO_REG_12_ );
nand U125899 ( n44297, n49619, n49620 );
nand U125900 ( n49619, P2_BUF1_REG_21_, n76478 );
nand U125901 ( n49620, n49621, n76476 );
xor U125902 ( n49621, n49622, n49623 );
nand U125903 ( n10412, n16678, n16679 );
nand U125904 ( n16678, P1_BUF1_REG_22_, n76611 );
nand U125905 ( n16679, n16680, n76613 );
xor U125906 ( n16680, n16682, n16683 );
nand U125907 ( n19367, n19374, P4_DATAO_REG_21_ );
nor U125908 ( n19374, n19368, n17374 );
nand U125909 ( n20499, P4_DATAO_REG_9_, n76582 );
and U125910 ( n17592, P4_DATAO_REG_24_, n76581 );
and U125911 ( n21019, n21011, P4_DATAO_REG_3_ );
nand U125912 ( n19045, n19053, P4_DATAO_REG_22_ );
nor U125913 ( n19053, n19046, n17374 );
nand U125914 ( n53209, n8227, P3_DATAO_REG_8_ );
and U125915 ( n54026, n76318, P3_DATAO_REG_2_ );
nand U125916 ( n20371, P4_DATAO_REG_8_, n8225 );
nand U125917 ( n20721, P4_DATAO_REG_12_, n76581 );
nand U125918 ( n20844, P4_DATAO_REG_10_, n76581 );
nand U125919 ( n50250, n8234, P3_DATAO_REG_23_ );
nand U125920 ( n20592, n20599, P4_DATAO_REG_18_ );
nor U125921 ( n20599, n20600, n17374 );
nand U125922 ( n54039, n8233, P3_DATAO_REG_3_ );
nand U125923 ( n20300, n20304, P4_DATAO_REG_19_ );
nor U125924 ( n20304, n20305, n17374 );
nand U125925 ( n19930, n19937, P4_DATAO_REG_20_ );
nor U125926 ( n19937, n19938, n17374 );
nand U125927 ( n18509, n18516, P4_DATAO_REG_24_ );
nor U125928 ( n18516, n18517, n17374 );
nand U125929 ( n20394, P4_DATAO_REG_8_, n76582 );
nand U125930 ( n18083, P4_DATAO_REG_23_, n76582 );
nand U125931 ( n10467, n16640, n16642 );
nand U125932 ( n16640, P1_BUF1_REG_21_, n76611 );
nand U125933 ( n16642, n16643, n76613 );
xor U125934 ( n16643, n16644, n16645 );
nand U125935 ( n53109, n8227, P3_DATAO_REG_7_ );
nand U125936 ( n52981, n8227, P3_DATAO_REG_6_ );
buf U125937 ( n76578, n16967 );
nand U125938 ( n16967, DIN_6_, n76927 );
nand U125939 ( n54002, n8233, P3_DATAO_REG_2_ );
nand U125940 ( n20169, P4_DATAO_REG_7_, n8225 );
nand U125941 ( n44305, n49591, n49592 );
nand U125942 ( n49591, P2_BUF1_REG_20_, n76478 );
nand U125943 ( n49592, n49593, n76476 );
xor U125944 ( n49593, n49594, n49595 );
nand U125945 ( n20278, P4_DATAO_REG_16_, n76582 );
nand U125946 ( n20575, P4_DATAO_REG_14_, n76582 );
buf U125947 ( n76312, n49946 );
nand U125948 ( n49946, DIN_8_, n76930 );
nand U125949 ( n20579, P4_DATAO_REG_15_, n76581 );
and U125950 ( n20192, P4_DATAO_REG_7_, n76581 );
nand U125951 ( n19917, P4_DATAO_REG_17_, n76582 );
nand U125952 ( n19350, P4_DATAO_REG_18_, n76582 );
and U125953 ( n54009, n76318, P3_DATAO_REG_1_ );
nand U125954 ( n52729, n8227, P3_DATAO_REG_5_ );
nand U125955 ( n20054, P4_DATAO_REG_6_, n8225 );
and U125956 ( n20957, n21011, P4_DATAO_REG_1_ );
nand U125957 ( n19796, P4_DATAO_REG_5_, n8225 );
nand U125958 ( n19028, P4_DATAO_REG_19_, n76582 );
nand U125959 ( n18652, n18659, P4_DATAO_REG_23_ );
nor U125960 ( n18659, n18660, n17374 );
nand U125961 ( n18316, P4_DATAO_REG_22_, n76582 );
nand U125962 ( n52613, n8227, P3_DATAO_REG_4_ );
nand U125963 ( n10477, n16604, n16605 );
nand U125964 ( n16604, P1_BUF1_REG_20_, n76611 );
nand U125965 ( n16605, n16607, n76613 );
xor U125966 ( n16607, n16608, n16609 );
nand U125967 ( n20060, P4_DATAO_REG_6_, n76582 );
buf U125968 ( n76309, n49947 );
nand U125969 ( n49947, DIN_9_, n76930 );
nand U125970 ( n21067, P4_DATAO_REG_4_, n8225 );
nand U125971 ( n53924, n8233, P3_DATAO_REG_1_ );
nand U125972 ( n49512, n53906, n53907 );
nand U125973 ( n53907, P3_DATAO_REG_1_, n53908 );
nand U125974 ( n53906, P3_DATAO_REG_2_, n53910 );
nand U125975 ( n53908, n49482, n53909 );
nand U125976 ( n18496, P4_DATAO_REG_21_, n76582 );
nand U125977 ( n52293, n8227, P3_DATAO_REG_3_ );
and U125978 ( n19801, P4_DATAO_REG_5_, n76581 );
nand U125979 ( n53262, n8234, P3_DATAO_REG_8_ );
and U125980 ( n19646, P4_DATAO_REG_4_, n76581 );
nand U125981 ( n53441, n8234, P3_DATAO_REG_10_ );
nand U125982 ( n53383, n8234, P3_DATAO_REG_9_ );
nand U125983 ( n44382, n49546, n49547 );
nand U125984 ( n49546, P2_BUF1_REG_19_, n76478 );
nand U125985 ( n49547, n49548, n31928 );
xor U125986 ( n49548, n49549, n49550 );
nand U125987 ( n17304, P4_DATAO_REG_23_, n8219 );
nand U125988 ( n21061, n8225, P4_DATAO_REG_3_ );
nand U125989 ( n18639, P4_DATAO_REG_20_, n76582 );
nand U125990 ( n52414, n8234, P3_DATAO_REG_15_ );
nand U125991 ( n53569, n8234, P3_DATAO_REG_11_ );
nand U125992 ( n53947, n8227, P3_DATAO_REG_2_ );
nand U125993 ( n52904, n8234, P3_DATAO_REG_13_ );
nand U125994 ( n52964, n8234, P3_DATAO_REG_6_ );
and U125995 ( n19640, P4_DATAO_REG_3_, n76581 );
nand U125996 ( n16527, n20950, n20951 );
nand U125997 ( n20951, P4_DATAO_REG_1_, n20952 );
nand U125998 ( n20950, P4_DATAO_REG_2_, n20954 );
nand U125999 ( n20952, n16488, n20953 );
nand U126000 ( n21003, P4_DATAO_REG_2_, n8225 );
nand U126001 ( n10573, n16568, n16569 );
nand U126002 ( n16568, P1_BUF1_REG_19_, n76610 );
nand U126003 ( n16569, n16570, n76613 );
xor U126004 ( n16570, n16572, n16573 );
nand U126005 ( n52712, n8234, P3_DATAO_REG_5_ );
buf U126006 ( n76571, n16991 );
nand U126007 ( n16991, DIN_8_, n76928 );
nand U126008 ( n20693, P4_DATAO_REG_10_, n8219 );
and U126009 ( n21024, P4_DATAO_REG_2_, n76581 );
nand U126010 ( n52584, n8234, P3_DATAO_REG_4_ );
nand U126011 ( n44440, n49516, n49517 );
nand U126012 ( n49516, P2_BUF1_REG_18_, n76478 );
nand U126013 ( n49517, n49518, n31928 );
xor U126014 ( n49518, n49519, n49520 );
nand U126015 ( n53941, n8227, P3_DATAO_REG_1_ );
nand U126016 ( n20525, P4_DATAO_REG_9_, n8219 );
nand U126017 ( n20408, n8219, P4_DATAO_REG_8_ );
nand U126018 ( n52272, n8234, P3_DATAO_REG_3_ );
buf U126019 ( n76568, n16992 );
nand U126020 ( n16992, DIN_9_, n76928 );
nand U126021 ( n20548, P4_DATAO_REG_11_, n8219 );
nand U126022 ( n52118, n8234, P3_DATAO_REG_2_ );
nand U126023 ( n20968, n8225, P4_DATAO_REG_1_ );
nand U126024 ( n19892, P4_DATAO_REG_13_, n8219 );
nand U126025 ( n49932, n49934, n49935 );
nor U126026 ( n49934, n49936, n49937 );
nand U126027 ( n49935, n8229, P3_DATAO_REG_30_ );
nor U126028 ( n49937, P3_DATAO_REG_31_, n49938 );
nand U126029 ( n10628, n16530, n16532 );
nand U126030 ( n16530, P1_BUF1_REG_18_, n76610 );
nand U126031 ( n16532, n16533, n76613 );
xor U126032 ( n16533, n16534, n16535 );
nand U126033 ( n44482, n49487, n49488 );
nand U126034 ( n49487, P2_BUF1_REG_17_, n76478 );
nand U126035 ( n49488, n49489, n31928 );
xor U126036 ( n49489, n49490, n49491 );
nand U126037 ( n50217, n8237, P3_DATAO_REG_20_ );
nand U126038 ( n19325, P4_DATAO_REG_15_, n8219 );
nand U126039 ( n20974, n76583, P4_DATAO_REG_1_ );
nand U126040 ( n49938, n76649, P3_DATAO_REG_30_ );
nand U126041 ( n52835, n8237, P3_DATAO_REG_11_ );
nand U126042 ( n44493, n49452, n49453 );
nand U126043 ( n49452, P2_BUF1_REG_16_, n76477 );
nand U126044 ( n49453, n49454, n31928 );
xor U126045 ( n49454, n49455, n49456 );
nand U126046 ( n53503, n8237, P3_DATAO_REG_10_ );
nand U126047 ( n13174, n70986, n848 );
nor U126048 ( n70986, P3_IR_REG_18_, P3_IR_REG_17_ );
nand U126049 ( n11399, n70980, n70976 );
nor U126050 ( n70980, P3_IR_REG_26_, P3_IR_REG_25_ );
nand U126051 ( n16703, n70994, n73024 );
nor U126052 ( n70994, P3_IR_REG_2_, P3_IR_REG_1_ );
nor U126053 ( n12652, n13174, P3_IR_REG_19_ );
nand U126054 ( n15214, n70989, n869 );
nor U126055 ( n70989, P3_IR_REG_12_, P3_IR_REG_11_ );
nand U126056 ( n14375, n70987, n855 );
nor U126057 ( n70987, P3_IR_REG_16_, P3_IR_REG_15_ );
nand U126058 ( n16270, n70993, n909 );
nor U126059 ( n70993, P3_IR_REG_4_, P3_IR_REG_3_ );
nand U126060 ( n15745, n70991, n889 );
nor U126061 ( n70991, P3_IR_REG_8_, P3_IR_REG_7_ );
nand U126062 ( n15482, n70990, n883 );
nor U126063 ( n70990, P3_IR_REG_9_, P3_IR_REG_10_ );
nand U126064 ( n16002, n70992, n899 );
nor U126065 ( n70992, P3_IR_REG_6_, P3_IR_REG_5_ );
nand U126066 ( n14923, n70988, n860 );
nor U126067 ( n70988, P3_IR_REG_14_, P3_IR_REG_13_ );
nor U126068 ( n70976, n11633, P3_IR_REG_24_ );
nand U126069 ( n41382, n42282, n42283 );
nand U126070 ( n42283, P3_IR_REG_0_, n604 );
nor U126071 ( n42282, n42284, n42285 );
nor U126072 ( n42284, n624, n40830 );
nand U126073 ( n67242, n67256, n815 );
nor U126074 ( n67256, P3_IR_REG_28_, P3_IR_REG_27_ );
nand U126075 ( n67314, n70985, n67316 );
nor U126076 ( n70985, P3_IR_REG_22_, P3_IR_REG_21_ );
nand U126077 ( n11340, n67241, n67242 );
nand U126078 ( n67241, P3_IR_REG_28_, n67243 );
nand U126079 ( n67243, n815, n73506 );
nor U126080 ( n67316, n844, P3_IR_REG_20_ );
or U126081 ( n11633, n67314, P3_IR_REG_23_ );
nand U126082 ( n41769, n67228, n67229 );
nand U126083 ( n67229, n76390, P3_IR_REG_0_ );
nand U126084 ( n67228, P1_P3_DATAO_REG_0_, n76389 );
nand U126085 ( n41449, n67239, n67240 );
nand U126086 ( n67239, P3_IR_REG_28_, n76841 );
or U126087 ( n67240, n11340, n76840 );
nand U126088 ( n1971, n40807, n40808 );
nor U126089 ( n40807, n40848, n40849 );
nor U126090 ( n40808, n40809, n40810 );
and U126091 ( n40848, n76042, P3_REG3_REG_28_ );
nand U126092 ( n20008, n8219, P4_DATAO_REG_6_ );
and U126093 ( n49515, n76318, P3_DATAO_REG_0_ );
nand U126094 ( n1871, n41204, n41205 );
nor U126095 ( n41204, n41304, n41305 );
nor U126096 ( n41205, n41206, n41207 );
and U126097 ( n41304, n76042, P3_REG3_REG_26_ );
xor U126098 ( n49901, n49909, n49910 );
nand U126099 ( n49909, n8227, P3_DATAO_REG_26_ );
nor U126100 ( n49910, n73010, n76322 );
nand U126101 ( n37080, n40340, n40341 );
nand U126102 ( n40340, P4_IR_REG_28_, n76795 );
nand U126103 ( n40341, n40342, P4_IR_REG_31_ );
nand U126104 ( n39626, n40570, n2202 );
nor U126105 ( n40570, P4_IR_REG_16_, P4_IR_REG_15_ );
nand U126106 ( n37764, n40338, n40339 );
nand U126107 ( n40339, P4_IR_REG_0_, n76459 );
nand U126108 ( n40338, P2_P3_DATAO_REG_0_, n76457 );
nor U126109 ( n39501, n39626, P4_IR_REG_17_ );
nor U126110 ( n40450, n40530, P4_IR_REG_22_ );
nor U126111 ( n40479, n40489, P4_IR_REG_28_ );
nand U126112 ( n40289, n40651, n73023 );
nor U126113 ( n40651, P4_IR_REG_2_, P4_IR_REG_1_ );
nand U126114 ( n39856, n40592, n2204 );
nor U126115 ( n40592, P4_IR_REG_12_, P4_IR_REG_11_ );
nand U126116 ( n40035, n40614, n2207 );
nor U126117 ( n40614, P4_IR_REG_8_, P4_IR_REG_7_ );
nand U126118 ( n40205, n40640, n2209 );
nor U126119 ( n40640, P4_IR_REG_4_, P4_IR_REG_3_ );
nand U126120 ( n39755, n40581, n2203 );
nor U126121 ( n40581, P4_IR_REG_14_, P4_IR_REG_13_ );
nand U126122 ( n39955, n40603, n2205 );
nor U126123 ( n40603, P4_IR_REG_9_, P4_IR_REG_10_ );
nand U126124 ( n40128, n40629, n2208 );
nor U126125 ( n40629, P4_IR_REG_6_, P4_IR_REG_5_ );
nand U126126 ( n40530, n40540, n40541 );
nor U126127 ( n40540, P4_IR_REG_21_, P4_IR_REG_20_ );
nor U126128 ( n40541, n40547, P4_IR_REG_19_ );
nor U126129 ( n40496, n40524, P4_IR_REG_24_ );
nand U126130 ( n37016, n37767, n37768 );
nand U126131 ( n37768, P4_IR_REG_0_, n2088 );
nor U126132 ( n37767, n37769, n37770 );
nor U126133 ( n37769, n2155, n37766 );
and U126134 ( n40346, n40495, n40496 );
nor U126135 ( n40495, P4_IR_REG_26_, P4_IR_REG_25_ );
nand U126136 ( n3196, n36404, n36405 );
nor U126137 ( n36404, n36447, n36448 );
nor U126138 ( n36405, n36406, n36407 );
and U126139 ( n36447, n76922, P4_REG3_REG_28_ );
nand U126140 ( n51933, n8237, P3_DATAO_REG_13_ );
nand U126141 ( n51771, n8234, P3_DATAO_REG_1_ );
nand U126142 ( n19756, n8219, P4_DATAO_REG_5_ );
nand U126143 ( n10680, n16494, n16495 );
nand U126144 ( n16494, P1_BUF1_REG_17_, n76610 );
nand U126145 ( n16495, n16497, n76613 );
xor U126146 ( n16497, n16498, n16499 );
nand U126147 ( n3096, n36823, n36824 );
nor U126148 ( n36823, n36936, n36937 );
nor U126149 ( n36824, n36825, n36826 );
and U126150 ( n36936, n76922, P4_REG3_REG_26_ );
nor U126151 ( n11394, P3_IR_REG_27_, n815 );
nand U126152 ( n41972, n67230, n67231 );
nand U126153 ( n67231, P3_IR_REG_27_, n67232 );
nand U126154 ( n67230, n11394, P3_IR_REG_31_ );
nand U126155 ( n67232, P3_IR_REG_31_, n11399 );
nand U126156 ( n16985, n16986, P4_DATAO_REG_29_ );
nor U126157 ( n16986, n16987, n16988 );
nand U126158 ( n53407, n8237, P3_DATAO_REG_9_ );
nand U126159 ( n37022, n40311, n40312 );
nand U126160 ( n40312, n76459, n37706 );
nand U126161 ( n40311, P2_P3_DATAO_REG_1_, n76458 );
nand U126162 ( n53172, n8237, P3_DATAO_REG_7_ );
nand U126163 ( n37300, n40413, n40414 );
nand U126164 ( n40413, P4_IR_REG_20_, n76796 );
or U126165 ( n40414, n40415, n76793 );
xor U126166 ( n40415, n40541, P4_IR_REG_20_ );
nand U126167 ( n19628, n8219, P4_DATAO_REG_4_ );
nand U126168 ( n37102, n40419, n40420 );
nand U126169 ( n40419, P4_IR_REG_22_, n76796 );
or U126170 ( n40420, n40421, n76793 );
nand U126171 ( n50742, n8237, P3_DATAO_REG_18_ );
nand U126172 ( n37609, n40343, n40344 );
nand U126173 ( n40343, P4_IR_REG_27_, n40348 );
nand U126174 ( n40344, n40345, P4_IR_REG_31_ );
nand U126175 ( n40348, n40347, P4_IR_REG_31_ );
nand U126176 ( n10694, n16452, n16453 );
nand U126177 ( n16452, P1_BUF1_REG_16_, n76610 );
nand U126178 ( n16453, n16454, n76612 );
xor U126179 ( n16454, n16455, n16457 );
nand U126180 ( n1926, n41012, n41013 );
nor U126181 ( n41012, n41020, n41021 );
nor U126182 ( n41013, n41014, n41015 );
and U126183 ( n41020, n76042, P3_REG3_REG_24_ );
nand U126184 ( n16975, n16977, n16978 );
nor U126185 ( n16977, n16979, n16980 );
nand U126186 ( n16978, P4_DATAO_REG_30_, n8220 );
nor U126187 ( n16980, P4_DATAO_REG_31_, n16981 );
nand U126188 ( n19479, n8219, P4_DATAO_REG_3_ );
nand U126189 ( n3086, n37115, n37116 );
nand U126190 ( n37115, P4_B_REG, n37601 );
nand U126191 ( n37116, n37117, n37118 );
nand U126192 ( n37601, n37602, n37603 );
nand U126193 ( n50201, n8238, P3_DATAO_REG_18_ );
nand U126194 ( n41378, n67011, n67012 );
nand U126195 ( n67012, n76391, n45201 );
nand U126196 ( n67011, P1_P3_DATAO_REG_1_, n76389 );
nand U126197 ( n2481, n38888, n38889 );
nand U126198 ( n38888, P4_REG0_REG_27_, n76422 );
nand U126199 ( n38889, n76012, n38633 );
nand U126200 ( n2641, n38631, n38632 );
nand U126201 ( n38631, P4_REG1_REG_27_, n76425 );
nand U126202 ( n38632, n76015, n38633 );
nand U126203 ( n53072, n8238, P3_DATAO_REG_7_ );
nand U126204 ( n19162, n8219, P4_DATAO_REG_2_ );
nand U126205 ( n41369, n66754, n66755 );
nand U126206 ( n66755, n76391, n42229 );
nand U126207 ( n66754, P1_P3_DATAO_REG_2_, n76389 );
nand U126208 ( n2651, n38625, n38626 );
nand U126209 ( n38625, P4_REG1_REG_29_, n76425 );
nand U126210 ( n38626, n76015, n38627 );
nand U126211 ( n2491, n38758, n38759 );
nand U126212 ( n38758, P4_REG0_REG_29_, n76421 );
nand U126213 ( n38759, n76012, n38627 );
nand U126214 ( n51005, n8237, P3_DATAO_REG_17_ );
nand U126215 ( n53040, n8238, P3_DATAO_REG_6_ );
nand U126216 ( n37007, n40284, n40285 );
nand U126217 ( n40285, n76460, n37721 );
nand U126218 ( n40284, P2_P3_DATAO_REG_2_, n76458 );
nand U126219 ( n17271, P4_DATAO_REG_20_, n8215 );
nand U126220 ( n3151, n36619, n36620 );
nor U126221 ( n36619, n36634, n36635 );
nor U126222 ( n36620, n36621, n36622 );
and U126223 ( n36634, n76922, P4_REG3_REG_24_ );
nand U126224 ( n52780, n8238, P3_DATAO_REG_5_ );
nand U126225 ( n2486, n38824, n38825 );
nand U126226 ( n38824, P4_REG0_REG_28_, n76422 );
nand U126227 ( n38825, n76012, n38630 );
nand U126228 ( n2646, n38628, n38629 );
nand U126229 ( n38628, P4_REG1_REG_28_, n38617 );
nand U126230 ( n38629, n76015, n38630 );
nand U126231 ( n49933, n76319, P3_DATAO_REG_29_ );
nand U126232 ( n40789, n66443, n66444 );
nand U126233 ( n66444, n76391, n42251 );
nand U126234 ( n66443, P1_P3_DATAO_REG_3_, n76389 );
nand U126235 ( n51409, n8237, P3_DATAO_REG_15_ );
nand U126236 ( n36386, n40238, n40239 );
nand U126237 ( n40239, n76460, n37740 );
nand U126238 ( n40238, P2_P3_DATAO_REG_3_, n76458 );
nand U126239 ( n51498, n8238, P3_DATAO_REG_13_ );
nand U126240 ( n19873, P4_DATAO_REG_11_, n8215 );
nand U126241 ( n20238, P4_DATAO_REG_10_, n8215 );
nand U126242 ( n1426, n55788, n55789 );
nand U126243 ( n55788, P3_REG1_REG_29_, n76288 );
nand U126244 ( n55789, n76002, n55790 );
nand U126245 ( n1266, n61390, n61391 );
nand U126246 ( n61390, P3_REG0_REG_29_, n76255 );
nand U126247 ( n61391, n75994, n55790 );
nand U126248 ( n1261, n61579, n61580 );
nand U126249 ( n61579, P3_REG0_REG_28_, n76255 );
nand U126250 ( n61580, n75994, n55954 );
nand U126251 ( n1421, n55952, n55953 );
nand U126252 ( n55952, P3_REG1_REG_28_, n76288 );
nand U126253 ( n55953, n76002, n55954 );
nand U126254 ( n20533, P4_DATAO_REG_9_, n8215 );
nand U126255 ( n49969, DIN_12_, n76930 );
nand U126256 ( n52550, n8238, P3_DATAO_REG_4_ );
nand U126257 ( n51225, n8237, P3_DATAO_REG_16_ );
nand U126258 ( n20216, P4_DATAO_REG_7_, n8215 );
nand U126259 ( n49941, n8234, P3_DATAO_REG_24_ );
nand U126260 ( n36655, n40200, n40201 );
nand U126261 ( n40201, n76460, n37783 );
nand U126262 ( n40200, P2_P3_DATAO_REG_4_, n76458 );
nand U126263 ( n36822, n40123, n40124 );
nand U126264 ( n40124, n76460, n37816 );
nand U126265 ( n40123, P2_P3_DATAO_REG_6_, n76458 );
nand U126266 ( n18977, P4_DATAO_REG_13_, n8215 );
nand U126267 ( n2636, n38634, n38635 );
nand U126268 ( n38634, P4_REG1_REG_26_, n38617 );
nand U126269 ( n38635, n76015, n38636 );
nand U126270 ( n2476, n38957, n38958 );
nand U126271 ( n38957, P4_REG0_REG_26_, n76421 );
nand U126272 ( n38958, n76012, n38636 );
nand U126273 ( n36594, n40163, n40164 );
nand U126274 ( n40164, n76460, n37799 );
nand U126275 ( n40163, P2_P3_DATAO_REG_5_, n76458 );
nand U126276 ( n37097, n40416, n40417 );
nand U126277 ( n40416, P4_IR_REG_21_, n76796 );
or U126278 ( n40417, n40418, n76793 );
nand U126279 ( n40418, n40539, n40530 );
nand U126280 ( n40539, P4_IR_REG_21_, n40542 );
nand U126281 ( n40542, n40541, n73042 );
nor U126282 ( n67262, n75920, n75921 );
and U126283 ( n75920, P3_IR_REG_26_, n76842 );
nor U126284 ( n75921, n11455, n76839 );
nand U126285 ( n11455, n70979, n11399 );
nand U126286 ( n70979, P3_IR_REG_26_, n70981 );
or U126287 ( n70981, n622, P3_IR_REG_25_ );
nand U126288 ( n1896, n41120, n41121 );
nor U126289 ( n41120, n41130, n41131 );
nor U126290 ( n41121, n41122, n41123 );
and U126291 ( n41130, n76042, P3_REG3_REG_22_ );
nand U126292 ( n18815, n8219, P4_DATAO_REG_1_ );
and U126293 ( n44560, n45510, n45511 );
nand U126294 ( n45510, P2_BUF1_REG_15_, n76478 );
nand U126295 ( n45511, n45512, n31928 );
xor U126296 ( n45512, n45513, n45514 );
nand U126297 ( n15851, n45505, n45506 );
nand U126298 ( n45506, P2_P1_LWORD_REG_15_, n76352 );
nor U126299 ( n45505, n45507, n45508 );
nor U126300 ( n45507, n74865, n76349 );
nand U126301 ( n1906, n41076, n41077 );
nor U126302 ( n41076, n41086, n41087 );
nor U126303 ( n41077, n41078, n41079 );
and U126304 ( n41086, n76042, P3_REG3_REG_20_ );
nand U126305 ( n3121, n36736, n36737 );
nor U126306 ( n36736, n36748, n36749 );
nor U126307 ( n36737, n36738, n36739 );
and U126308 ( n36748, n76922, P4_REG3_REG_22_ );
nand U126309 ( n49970, DIN_13_, n76929 );
nand U126310 ( n52094, n8238, P3_DATAO_REG_2_ );
xor U126311 ( n16946, n16954, n16955 );
nand U126312 ( n16954, P4_DATAO_REG_27_, n76581 );
nor U126313 ( n16955, n76586, n73013 );
nand U126314 ( n16981, P4_DATAO_REG_30_, n8222 );
nand U126315 ( n1256, n62236, n62237 );
nand U126316 ( n62236, P3_REG0_REG_27_, n76255 );
nand U126317 ( n62237, n75994, n56052 );
nand U126318 ( n1416, n56050, n56051 );
nand U126319 ( n56050, P3_REG1_REG_27_, n76288 );
nand U126320 ( n56051, n76002, n56052 );
nand U126321 ( n46000, n46001, n46002 );
nand U126322 ( n46001, P3_REG2_REG_27_, n45363 );
nand U126323 ( n46002, n76858, n46003 );
nand U126324 ( n70965, n70982, n70983 );
nand U126325 ( n70982, P3_IR_REG_24_, n76840 );
nand U126326 ( n70983, n70984, P3_IR_REG_31_ );
and U126327 ( n70984, n622, n11574 );
xnor U126328 ( n10769, n10120, P3_IR_REG_30_ );
nand U126329 ( n67249, n67254, n67255 );
nand U126330 ( n67254, P3_IR_REG_30_, n76842 );
or U126331 ( n67255, n10769, n76839 );
or U126332 ( n10120, n67242, P3_IR_REG_29_ );
nand U126333 ( n20116, n8217, P4_DATAO_REG_7_ );
nand U126334 ( n2471, n39022, n39023 );
nand U126335 ( n39022, P4_REG0_REG_25_, n76422 );
nand U126336 ( n39023, n76012, n38639 );
nand U126337 ( n2631, n38637, n38638 );
nand U126338 ( n38637, P4_REG1_REG_25_, n38617 );
nand U126339 ( n38638, n76015, n38639 );
nand U126340 ( n41042, n66372, n66373 );
nand U126341 ( n66373, n76391, n42299 );
nand U126342 ( n66372, P1_P3_DATAO_REG_4_, n76389 );
buf U126343 ( n76792, n2250 );
not U126344 ( n2250, P4_IR_REG_31_ );
nand U126345 ( n17783, P4_DATAO_REG_18_, n8215 );
nand U126346 ( n2461, n39138, n39139 );
nand U126347 ( n39138, P4_REG0_REG_23_, n76422 );
nand U126348 ( n39139, n76012, n38645 );
nand U126349 ( n2621, n38643, n38644 );
nand U126350 ( n38643, P4_REG1_REG_23_, n76425 );
nand U126351 ( n38644, n76015, n38645 );
nand U126352 ( n41466, n67309, n67310 );
nand U126353 ( n67309, P3_IR_REG_21_, n76842 );
or U126354 ( n67310, n12109, n76839 );
xnor U126355 ( n12109, n843, P3_IR_REG_21_ );
nand U126356 ( n3131, n36685, n36686 );
nor U126357 ( n36685, n36703, n36704 );
nor U126358 ( n36686, n36687, n36688 );
and U126359 ( n36703, n76922, P4_REG3_REG_20_ );
nand U126360 ( n11574, P3_IR_REG_24_, n11633 );
xor U126361 ( n11518, P3_IR_REG_25_, n70976 );
nand U126362 ( n70968, n70974, n70975 );
nand U126363 ( n70974, P3_IR_REG_25_, n76842 );
or U126364 ( n70975, n11518, n76839 );
nand U126365 ( n71021, n72897, n73430 );
nand U126366 ( n72897, n73396, n72898 );
nand U126367 ( n72898, P4_DATAO_REG_29_, n72899 );
nand U126368 ( n72899, n72900, n72901 );
nor U126369 ( n72890, n2362, P3_WR_REG );
nand U126370 ( n71259, n72758, n72759 );
nor U126371 ( n72758, n72762, n72763 );
nor U126372 ( n72759, n72760, n72761 );
and U126373 ( n72763, P3_ADDR_REG_2_, P3_WR_REG );
nor U126374 ( n72761, n73439, n71104 );
nand U126375 ( n20084, n8217, P4_DATAO_REG_6_ );
and U126376 ( n67238, n76254, P3_REG0_REG_0_ );
nor U126377 ( n72901, n72902, n72903 );
nand U126378 ( n72903, n72904, n72905 );
nand U126379 ( n72902, n72909, n72910 );
nor U126380 ( n72904, P4_DATAO_REG_22_, n72908 );
and U126381 ( n43798, n45498, n45499 );
nand U126382 ( n45498, P2_BUF1_REG_14_, n76477 );
nand U126383 ( n45499, n45500, n31928 );
xnor U126384 ( n45500, n45501, n45502 );
nand U126385 ( n15931, n45384, n45385 );
nand U126386 ( n45385, P2_P1_UWORD_REG_14_, n76352 );
nor U126387 ( n45384, n45386, n45387 );
nor U126388 ( n45387, n75404, n76350 );
nand U126389 ( n15856, n45495, n45496 );
nand U126390 ( n45496, P2_P1_LWORD_REG_14_, n76352 );
nor U126391 ( n45495, n45386, n45497 );
nor U126392 ( n45497, n73251, n76349 );
nand U126393 ( n71012, n72852, n73431 );
nand U126394 ( n72852, n72853, n72854 );
nor U126395 ( n72853, P3_DATAO_REG_30_, P3_DATAO_REG_29_ );
nand U126396 ( n72854, P3_DATAO_REG_28_, n72855 );
nor U126397 ( n72830, n1244, P4_WR_REG );
nor U126398 ( n72779, n73447, n71283 );
nand U126399 ( n72870, n72877, n72878 );
nor U126400 ( n72877, P3_DATAO_REG_16_, n72881 );
nor U126401 ( n72878, n72879, n72880 );
nand U126402 ( n72881, n73002, n73403 );
nor U126403 ( n72768, n73443, n71283 );
nand U126404 ( n41493, n67306, n67307 );
nand U126405 ( n67306, P3_IR_REG_20_, n76842 );
nand U126406 ( n67307, n67308, P3_IR_REG_31_ );
and U126407 ( n67308, n843, n12409 );
nand U126408 ( n72859, n72860, n72861 );
nor U126409 ( n72860, P3_DATAO_REG_22_, n72864 );
nor U126410 ( n72861, n72862, n72863 );
nand U126411 ( n72864, n73416, n73016 );
nand U126412 ( n17255, P4_DATAO_REG_18_, n8217 );
nand U126413 ( n16236, n44608, n44609 );
nor U126414 ( n44609, n44610, n44611 );
nor U126415 ( n44608, n44615, n44616 );
nor U126416 ( n44610, P2_P1_EAX_REG_14_, n44556 );
nand U126417 ( n72795, P3_WR_REG, P3_ADDR_REG_0_ );
nand U126418 ( n72796, n71001, n73026 );
nand U126419 ( n71001, n72797, n72798 );
nand U126420 ( n72798, n2362, P2_P1_ADDRESS_REG_0_ );
nor U126421 ( n72797, n72799, n72800 );
nor U126422 ( n72799, n73435, n71017 );
nor U126423 ( n72800, n73434, n71022 );
nand U126424 ( n40989, n66300, n66301 );
nand U126425 ( n66301, n76391, n42344 );
nand U126426 ( n66300, P1_P3_DATAO_REG_5_, n76389 );
xnor U126427 ( n40362, n40478, P4_IR_REG_30_ );
nand U126428 ( n40478, n40479, n73058 );
nand U126429 ( n40354, n40360, n40361 );
nand U126430 ( n40360, P4_IR_REG_30_, n76795 );
or U126431 ( n40361, n40362, n76793 );
nor U126432 ( n72865, P3_DATAO_REG_3_, n72869 );
nand U126433 ( n72869, n73021, n73421 );
nor U126434 ( n72748, n73441, n71283 );
nor U126435 ( n72786, n73449, n71283 );
nand U126436 ( n37303, n40410, n40411 );
nand U126437 ( n40410, P4_IR_REG_19_, n76796 );
or U126438 ( n40411, n40412, n76793 );
and U126439 ( n16602, n76583, P4_DATAO_REG_0_ );
nand U126440 ( n1251, n62292, n62293 );
nand U126441 ( n62292, P3_REG0_REG_26_, n76255 );
nand U126442 ( n62293, n75994, n56148 );
nand U126443 ( n1411, n56146, n56147 );
nand U126444 ( n56146, P3_REG1_REG_26_, n76288 );
nand U126445 ( n56147, n76002, n56148 );
nand U126446 ( n46222, n46223, n46224 );
nand U126447 ( n46223, P3_REG2_REG_26_, n45363 );
nand U126448 ( n46224, n76858, n46225 );
nand U126449 ( n67248, n67252, n67253 );
nand U126450 ( n67252, P3_IR_REG_29_, n76841 );
nand U126451 ( n67253, P3_IR_REG_31_, n11245 );
nand U126452 ( n11245, P3_IR_REG_29_, n67242 );
nand U126453 ( n40442, n40459, n40460 );
nand U126454 ( n40459, P4_IR_REG_24_, n76796 );
nand U126455 ( n40460, n40461, P4_IR_REG_31_ );
nand U126456 ( n2626, n38640, n38641 );
nand U126457 ( n38640, P4_REG1_REG_24_, n38617 );
nand U126458 ( n38641, n76015, n38642 );
nand U126459 ( n2466, n39074, n39075 );
nand U126460 ( n39074, P4_REG0_REG_24_, n76421 );
nand U126461 ( n39075, n76012, n38642 );
nand U126462 ( n12409, P3_IR_REG_20_, n844 );
nor U126463 ( n72917, P4_DATAO_REG_0_, n72921 );
nand U126464 ( n72921, n73414, n73012 );
nand U126465 ( n40353, n40357, n40358 );
nand U126466 ( n40357, P4_IR_REG_29_, n76795 );
or U126467 ( n40358, n40359, n76794 );
and U126468 ( n10784, n11734, n11735 );
nand U126469 ( n11734, P1_BUF1_REG_15_, n76610 );
nand U126470 ( n11735, n11737, n76612 );
xor U126471 ( n11737, n11738, n11739 );
nand U126472 ( n9116, n11728, n11729 );
nand U126473 ( n11729, P1_P1_LWORD_REG_15_, n11504 );
nor U126474 ( n11728, n11730, n11732 );
nor U126475 ( n11730, n74864, n76615 );
nand U126476 ( n72871, n72872, n72873 );
nor U126477 ( n72873, n72874, n72875 );
nor U126478 ( n72872, P3_DATAO_REG_0_, n72876 );
nand U126479 ( n72874, n73400, n72999 );
nand U126480 ( n1236, n62535, n62536 );
nand U126481 ( n62535, P3_REG0_REG_23_, n76255 );
nand U126482 ( n62536, n75994, n57363 );
nand U126483 ( n1396, n57361, n57362 );
nand U126484 ( n57361, P3_REG1_REG_23_, n76288 );
nand U126485 ( n57362, n76002, n57363 );
nand U126486 ( n51790, n8238, P3_DATAO_REG_1_ );
nand U126487 ( n47417, n47418, n47419 );
nand U126488 ( n47418, P3_REG2_REG_23_, n45363 );
nand U126489 ( n47419, n76858, n47420 );
nand U126490 ( n18047, P4_DATAO_REG_17_, n8215 );
nor U126491 ( n72552, n73457, n71283 );
nand U126492 ( n41203, n66220, n66221 );
nand U126493 ( n66221, n76391, n45184 );
nand U126494 ( n66220, P1_P3_DATAO_REG_6_, n76389 );
nor U126495 ( n72922, P4_DATAO_REG_16_, n72926 );
nand U126496 ( n72926, n73408, n73007 );
and U126497 ( n40356, n76420, P4_REG0_REG_0_ );
nand U126498 ( n18453, P4_DATAO_REG_15_, n8215 );
nor U126499 ( n72794, n73438, n71022 );
nand U126500 ( n71024, n72791, n72792 );
nand U126501 ( n72792, n2362, P2_P1_ADDRESS_REG_1_ );
nor U126502 ( n72791, n72793, n72794 );
nor U126503 ( n72793, n73437, n71017 );
nor U126504 ( n72724, n73453, n71283 );
nand U126505 ( n19824, n8217, P4_DATAO_REG_5_ );
nand U126506 ( n41908, n67303, n67304 );
nand U126507 ( n67303, P3_IR_REG_19_, n76842 );
nand U126508 ( n67304, n67305, P3_IR_REG_31_ );
nor U126509 ( n67305, n12652, n12650 );
buf U126510 ( n76838, n934 );
not U126511 ( n934, P3_IR_REG_31_ );
and U126512 ( n40335, n76420, P4_REG0_REG_1_ );
nand U126513 ( n1246, n62352, n62353 );
nand U126514 ( n62352, P3_REG0_REG_25_, n76255 );
nand U126515 ( n62353, n75994, n56372 );
nand U126516 ( n1406, n56370, n56371 );
nand U126517 ( n56370, P3_REG1_REG_25_, n76288 );
nand U126518 ( n56371, n76002, n56372 );
nor U126519 ( n72474, n73469, n71283 );
and U126520 ( n12650, P3_IR_REG_19_, n13174 );
nand U126521 ( n18542, P4_DATAO_REG_13_, n8217 );
and U126522 ( n49834, DIN_14_, n76929 );
and U126523 ( n52035, n49834, P3_DATAO_REG_8_ );
and U126524 ( n43846, n45478, n45479 );
nand U126525 ( n45478, P2_BUF1_REG_13_, n76477 );
nand U126526 ( n45479, n45480, n31928 );
xor U126527 ( n45480, n45481, n45482 );
nand U126528 ( n15936, n45380, n45381 );
nand U126529 ( n45381, P2_P1_UWORD_REG_13_, n76352 );
nor U126530 ( n45380, n45382, n45383 );
nor U126531 ( n45383, n75218, n76350 );
nand U126532 ( n15861, n45475, n45476 );
nand U126533 ( n45476, P2_P1_LWORD_REG_13_, n76352 );
nor U126534 ( n45475, n45382, n45477 );
nor U126535 ( n45477, n74842, n76349 );
nor U126536 ( n72829, n73461, n71283 );
nand U126537 ( n36293, n40074, n40075 );
nand U126538 ( n40075, n76460, n37827 );
nand U126539 ( n40074, P2_P3_DATAO_REG_7_, n76458 );
nand U126540 ( n41471, n67311, n67312 );
nand U126541 ( n67311, P3_IR_REG_22_, n76842 );
or U126542 ( n67312, n11785, n76839 );
nand U126543 ( n11785, n67313, n67314 );
nand U126544 ( n67313, P3_IR_REG_22_, n67315 );
or U126545 ( n67315, n843, P3_IR_REG_21_ );
nand U126546 ( n2456, n39199, n39200 );
nand U126547 ( n39199, P4_REG0_REG_22_, n76422 );
nand U126548 ( n39200, n76012, n38648 );
nand U126549 ( n2616, n38646, n38647 );
nand U126550 ( n38646, P4_REG1_REG_22_, n76425 );
nand U126551 ( n38647, n76015, n38648 );
nand U126552 ( n66120, n76391, n42678 );
nand U126553 ( n66119, P1_P3_DATAO_REG_7_, n76389 );
nor U126554 ( n40262, n76414, n73999 );
and U126555 ( n67251, n76254, P3_REG0_REG_1_ );
nor U126556 ( n72386, n73471, n71283 );
nor U126557 ( n72811, n73462, n71283 );
nor U126558 ( n72689, n73465, n71283 );
and U126559 ( n9895, n11719, n11720 );
nand U126560 ( n11719, P1_BUF1_REG_14_, n76610 );
nand U126561 ( n11720, n11722, n76612 );
xnor U126562 ( n11722, n11723, n11724 );
nand U126563 ( n9196, n11585, n11587 );
nand U126564 ( n11587, P1_P1_UWORD_REG_14_, n76618 );
nor U126565 ( n11585, n11588, n11589 );
nor U126566 ( n11589, n75405, n76616 );
nand U126567 ( n9121, n11715, n11717 );
nand U126568 ( n11717, P1_P1_LWORD_REG_14_, n76618 );
nor U126569 ( n11715, n11588, n11718 );
nor U126570 ( n11718, n73252, n76615 );
and U126571 ( n67004, n76254, P3_REG0_REG_2_ );
nor U126572 ( n40261, P4_REG3_REG_3_, n76403 );
nand U126573 ( n19594, n8217, P4_DATAO_REG_4_ );
nand U126574 ( n9501, n10844, n10845 );
nor U126575 ( n10845, n10847, n10848 );
nor U126576 ( n10844, n10853, n10854 );
nor U126577 ( n10847, P1_P1_EAX_REG_14_, n10779 );
nand U126578 ( n18273, P4_DATAO_REG_16_, n8215 );
nand U126579 ( n51907, n49834, P3_DATAO_REG_9_ );
nor U126580 ( n66731, P3_REG3_REG_3_, n76241 );
nand U126581 ( n17247, P4_DATAO_REG_18_, n76166 );
and U126582 ( n17015, DIN_12_, n76927 );
nand U126583 ( n36467, n40030, n40031 );
nand U126584 ( n40031, n76460, n37841 );
nand U126585 ( n40030, P2_P3_DATAO_REG_8_, n76458 );
nand U126586 ( n36360, n39950, n39951 );
nand U126587 ( n39951, n76459, n37872 );
nand U126588 ( n39950, P2_P3_DATAO_REG_10_, n76458 );
nand U126589 ( n1241, n62419, n62420 );
nand U126590 ( n62419, P3_REG0_REG_24_, n76255 );
nand U126591 ( n62420, n75994, n56888 );
nand U126592 ( n1401, n56886, n56887 );
nand U126593 ( n56886, P3_REG1_REG_24_, n76288 );
nand U126594 ( n56887, n76002, n56888 );
and U126595 ( n51504, n49834, P3_DATAO_REG_10_ );
nand U126596 ( n46939, n46940, n46941 );
nand U126597 ( n46940, P3_REG2_REG_24_, n45363 );
nand U126598 ( n46941, n76858, n46942 );
nand U126599 ( n36672, n39986, n39987 );
nand U126600 ( n39987, n76460, n37855 );
nand U126601 ( n39986, P2_P3_DATAO_REG_9_, n76458 );
nand U126602 ( n1231, n62627, n62628 );
nand U126603 ( n62627, P3_REG0_REG_22_, n76255 );
nand U126604 ( n62628, n75994, n57455 );
nand U126605 ( n1391, n57453, n57454 );
nand U126606 ( n57453, P3_REG1_REG_22_, n76288 );
nand U126607 ( n57454, n76002, n57455 );
and U126608 ( n40263, n76420, P4_REG0_REG_3_ );
nor U126609 ( n72754, n73474, n71104 );
nand U126610 ( n50169, n49834, P3_DATAO_REG_16_ );
nand U126611 ( n40765, n65827, n65828 );
nand U126612 ( n65828, n76390, n45243 );
nand U126613 ( n65827, P1_P3_DATAO_REG_10_, n76389 );
nand U126614 ( n2451, n39261, n39262 );
nand U126615 ( n39261, P4_REG0_REG_21_, n76422 );
nand U126616 ( n39262, n76012, n38651 );
nand U126617 ( n2611, n38649, n38650 );
nand U126618 ( n38649, P4_REG1_REG_21_, n76425 );
nand U126619 ( n38650, n76015, n38651 );
and U126620 ( n66733, n76254, P3_REG0_REG_3_ );
nand U126621 ( n41059, n65950, n65951 );
nand U126622 ( n65951, n76390, n43230 );
nand U126623 ( n65950, P1_P3_DATAO_REG_9_, n76389 );
and U126624 ( n40304, n76420, P4_REG0_REG_2_ );
nand U126625 ( n18964, P4_DATAO_REG_11_, n76169 );
nand U126626 ( n51388, n49834, P3_DATAO_REG_11_ );
nand U126627 ( n71143, n72285, n72286 );
nor U126628 ( n72285, n72289, n72290 );
nor U126629 ( n72286, n72287, n72288 );
and U126630 ( n72290, P4_ADDR_REG_4_, P4_WR_REG );
nor U126631 ( n72288, n73478, n71283 );
buf U126632 ( n76384, n41511 );
nand U126633 ( n41511, LOGIC0, n76389 );
nand U126634 ( n52808, n49834, P3_DATAO_REG_7_ );
and U126635 ( n9955, n11707, n11708 );
nand U126636 ( n11707, P1_BUF1_REG_13_, n76610 );
nand U126637 ( n11708, n11709, n76612 );
xor U126638 ( n11709, n11710, n11712 );
nand U126639 ( n9201, n11580, n11582 );
nand U126640 ( n11582, P1_P1_UWORD_REG_13_, n76618 );
nor U126641 ( n11580, n11583, n11584 );
nor U126642 ( n11584, n75219, n76616 );
nand U126643 ( n9126, n11703, n11704 );
nand U126644 ( n11704, P1_P1_LWORD_REG_13_, n76618 );
nor U126645 ( n11703, n11583, n11705 );
nor U126646 ( n11705, n74843, n76615 );
nand U126647 ( n20220, P4_DATAO_REG_7_, n76171 );
nand U126648 ( n41150, n65355, n65356 );
nand U126649 ( n65356, n76390, n43559 );
nand U126650 ( n65355, P1_P3_DATAO_REG_11_, n76389 );
nor U126651 ( n40184, n76414, n74166 );
and U126652 ( n43896, n45468, n45469 );
nand U126653 ( n45468, P2_BUF1_REG_12_, n76477 );
nand U126654 ( n45469, n45470, n31928 );
xnor U126655 ( n45470, n45471, n45472 );
nand U126656 ( n15941, n45376, n45377 );
nand U126657 ( n45377, P2_P1_UWORD_REG_12_, n76352 );
nor U126658 ( n45376, n45378, n45379 );
nor U126659 ( n45379, n75324, n76350 );
nand U126660 ( n15866, n45465, n45466 );
nand U126661 ( n45466, P2_P1_LWORD_REG_12_, n76352 );
nor U126662 ( n45465, n45378, n45467 );
nor U126663 ( n45467, n74803, n76349 );
nand U126664 ( n1226, n62728, n62729 );
nand U126665 ( n62728, P3_REG0_REG_21_, n76255 );
nand U126666 ( n62729, n75994, n57498 );
nand U126667 ( n1386, n57496, n57497 );
nand U126668 ( n57496, P3_REG1_REG_21_, n76288 );
nand U126669 ( n57497, n76002, n57498 );
nand U126670 ( n48076, n48077, n48078 );
nand U126671 ( n48077, P3_REG2_REG_21_, n45363 );
nand U126672 ( n48078, n76858, n48079 );
nand U126673 ( n40869, n66036, n66037 );
nand U126674 ( n66037, n76391, n42957 );
nand U126675 ( n66036, P1_P3_DATAO_REG_8_, n76389 );
nand U126676 ( n19138, n8217, P4_DATAO_REG_2_ );
nand U126677 ( n19292, P4_DATAO_REG_10_, n76169 );
nand U126678 ( n52922, n49834, P3_DATAO_REG_6_ );
nand U126679 ( n19392, P4_DATAO_REG_9_, n76167 );
nand U126680 ( n20088, P4_DATAO_REG_6_, n76166 );
nand U126681 ( n36767, n39909, n39910 );
nand U126682 ( n39910, n76459, n37883 );
nand U126683 ( n39909, P2_P3_DATAO_REG_11_, n76458 );
nand U126684 ( n19960, P4_DATAO_REG_8_, n76165 );
nand U126685 ( n40457, n40510, n40511 );
nor U126686 ( n40510, P4_IR_REG_25_, n39626 );
nor U126687 ( n40437, n75922, n75923 );
and U126688 ( n75922, P4_IR_REG_26_, n76796 );
nor U126689 ( n75923, n40464, n76793 );
nand U126690 ( n17016, n76928, DIN_13_ );
nor U126691 ( n40143, n76414, n74236 );
nor U126692 ( n41483, n41484, n41485 );
nand U126693 ( n41485, n41471, n41460 );
nor U126694 ( n41484, n41486, P3_B_REG );
nor U126695 ( n41486, n41487, n41488 );
and U126696 ( n40185, n76420, P4_REG0_REG_5_ );
nor U126697 ( n72180, n73485, n71283 );
nand U126698 ( n17504, P4_DATAO_REG_17_, n76165 );
nand U126699 ( n72801, n72891, n72892 );
nand U126700 ( n72892, P2_P3_DATAO_REG_30_, n73429 );
nor U126701 ( n72891, n72893, n72894 );
nor U126702 ( n72893, P2_P1_DATAO_REG_31_, n73428 );
nor U126703 ( n72894, P2_P2_DATAO_REG_31_, n73427 );
and U126704 ( n18447, P4_DATAO_REG_12_, n76167 );
nand U126705 ( n50446, n49834, P3_DATAO_REG_15_ );
nand U126706 ( n52790, n49834, P3_DATAO_REG_5_ );
and U126707 ( n40220, n76420, P4_REG0_REG_4_ );
and U126708 ( n40144, n76419, P4_REG0_REG_6_ );
nand U126709 ( n1376, n57587, n57588 );
nand U126710 ( n57587, P3_REG1_REG_19_, n76288 );
nand U126711 ( n57588, n76003, n57589 );
nand U126712 ( n1216, n62933, n62934 );
nand U126713 ( n62933, P3_REG0_REG_19_, n76255 );
nand U126714 ( n62934, n75995, n57589 );
and U126715 ( n18267, P4_DATAO_REG_13_, n76168 );
nand U126716 ( n36537, n39851, n39852 );
nand U126717 ( n39852, n76459, n37897 );
nand U126718 ( n39851, P2_P3_DATAO_REG_12_, n76458 );
nand U126719 ( n2601, n38659, n38660 );
nand U126720 ( n38659, P4_REG1_REG_19_, n76425 );
nand U126721 ( n38660, n76016, n38661 );
nand U126722 ( n2441, n39379, n39380 );
nand U126723 ( n39379, P4_REG0_REG_19_, n76422 );
nand U126724 ( n39380, n76013, n38661 );
nand U126725 ( n2606, n38656, n38657 );
nand U126726 ( n38656, P4_REG1_REG_20_, n76425 );
nand U126727 ( n38657, n76015, n38658 );
nand U126728 ( n2446, n39324, n39325 );
nand U126729 ( n39324, P4_REG0_REG_20_, n76422 );
nand U126730 ( n39325, n76012, n38658 );
nand U126731 ( n46482, n46578, n46579 );
nand U126732 ( n46578, n46581, n76341 );
nand U126733 ( n46579, P2_P1_INSTADDRPOINTER_REG_24_, n46580 );
or U126734 ( n46580, n46581, n76342 );
nand U126735 ( n44548, P2_P1_INSTQUEUERD_ADDR_REG_2_, n73497 );
nand U126736 ( n47204, n47234, n47235 );
nand U126737 ( n47234, n47237, n76341 );
nand U126738 ( n47235, P2_P1_INSTADDRPOINTER_REG_7_, n47236 );
or U126739 ( n47236, n47237, n76342 );
nand U126740 ( n46311, n46371, n46372 );
nand U126741 ( n46371, P2_P1_INSTADDRPOINTER_REG_29_, n46373 );
nand U126742 ( n46372, n46313, n76342 );
nand U126743 ( n45627, n46478, n46479 );
nand U126744 ( n46479, P2_P1_INSTADDRPOINTER_REG_26_, n46480 );
nand U126745 ( n46480, n76345, n46481 );
nand U126746 ( n46481, P2_P1_INSTADDRPOINTER_REG_25_, n46482 );
nand U126747 ( n46617, n46649, n46650 );
nor U126748 ( n46649, n7534, n46651 );
nor U126749 ( n46651, P2_P1_INSTADDRPOINTER_REG_22_, n76341 );
nor U126750 ( n46440, n45627, P2_P1_INSTADDRPOINTER_REG_27_ );
nor U126751 ( n47021, n47121, n47122 );
and U126752 ( n47122, P2_P1_INSTADDRPOINTER_REG_10_, n47123 );
nand U126753 ( n47123, n76345, n47124 );
nand U126754 ( n46320, P2_P1_INSTADDRPOINTER_REG_30_, n46311 );
nand U126755 ( n46373, n46396, n46397 );
nand U126756 ( n46397, P2_P1_INSTADDRPOINTER_REG_28_, n76341 );
nor U126757 ( n46396, n45630, n46398 );
nor U126758 ( n46398, n7533, n46369 );
nand U126759 ( n46692, n46837, n46838 );
nand U126760 ( n46838, P2_P1_INSTADDRPOINTER_REG_17_, n76341 );
nor U126761 ( n46837, n7537, n46839 );
nor U126762 ( n46839, n7538, n46818 );
nor U126763 ( n46315, n46317, n46318 );
nor U126764 ( n46318, P2_P1_INSTADDRPOINTER_REG_30_, n46311 );
nor U126765 ( n46317, n46319, n76341 );
nor U126766 ( n46319, n75052, n46320 );
nand U126767 ( n47124, n47160, P2_P1_INSTADDRPOINTER_REG_8_ );
nor U126768 ( n47160, n7544, n73078 );
or U126769 ( n46313, n46373, P2_P1_INSTADDRPOINTER_REG_29_ );
and U126770 ( n45546, n46305, n46306 );
nand U126771 ( n46306, n46307, n46308 );
nand U126772 ( n46305, n46315, n46316 );
nand U126773 ( n46308, n76006, P2_P1_INSTADDRPOINTER_REG_31_ );
nand U126774 ( n15686, n46294, n46295 );
nand U126775 ( n46295, n76859, P2_P1_INSTADDRPOINTER_REG_31_ );
nor U126776 ( n46294, n46296, n46297 );
nor U126777 ( n46297, n75328, n76334 );
nand U126778 ( n46875, n46911, n46912 );
nand U126779 ( n46911, n46914, n76341 );
nand U126780 ( n46912, P2_P1_INSTADDRPOINTER_REG_15_, n46913 );
or U126781 ( n46913, n46914, n76342 );
nand U126782 ( n36735, n39804, n39805 );
nand U126783 ( n39805, n76459, n37913 );
nand U126784 ( n39804, P2_P3_DATAO_REG_13_, n76458 );
nand U126785 ( n72831, n72882, n72883 );
nand U126786 ( n72883, P1_P3_DATAO_REG_30_, n73436 );
nor U126787 ( n72882, n72884, n72885 );
nor U126788 ( n72884, P1_P1_DATAO_REG_31_, n73433 );
nor U126789 ( n72885, P1_P2_DATAO_REG_31_, n73432 );
and U126790 ( n9974, n11694, n11695 );
nand U126791 ( n11694, P1_BUF1_REG_12_, n76610 );
nand U126792 ( n11695, n11697, n76612 );
xnor U126793 ( n11697, n11698, n11699 );
nand U126794 ( n9206, n11575, n11577 );
nand U126795 ( n11577, P1_P1_UWORD_REG_12_, n76618 );
nor U126796 ( n11575, n11578, n11579 );
nor U126797 ( n11579, n75325, n76616 );
nand U126798 ( n9131, n11690, n11692 );
nand U126799 ( n11692, P1_P1_LWORD_REG_12_, n76618 );
nor U126800 ( n11690, n11578, n11693 );
nor U126801 ( n11693, n74802, n76615 );
nor U126802 ( n72702, n73487, n71104 );
nand U126803 ( n71243, n72699, n72700 );
nor U126804 ( n72699, n72703, n72704 );
nor U126805 ( n72700, n72701, n72702 );
and U126806 ( n72704, P3_ADDR_REG_4_, P3_WR_REG );
nand U126807 ( n1221, n62818, n62819 );
nand U126808 ( n62818, P3_REG0_REG_20_, n76255 );
nand U126809 ( n62819, n75994, n57542 );
nand U126810 ( n1381, n57540, n57541 );
nand U126811 ( n57540, P3_REG1_REG_20_, n76288 );
nand U126812 ( n57541, n76002, n57542 );
nand U126813 ( n44894, P2_P1_INSTQUEUERD_ADDR_REG_1_, P2_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U126814 ( n40458, P4_IR_REG_25_, n40512 );
nand U126815 ( n40512, n40511, n2200 );
not U126816 ( n2200, n39626 );
nand U126817 ( n40445, n40454, n40455 );
nand U126818 ( n40454, P4_IR_REG_25_, n76796 );
nand U126819 ( n40455, n40456, P4_IR_REG_31_ );
and U126820 ( n40456, n40457, n40458 );
and U126821 ( n66429, n76254, P3_REG0_REG_4_ );
nand U126822 ( n36955, n39679, n39680 );
nand U126823 ( n39680, n76459, n37941 );
nand U126824 ( n39679, P2_P3_DATAO_REG_15_, n76458 );
nand U126825 ( n65423, P2_P3_INSTQUEUERD_ADDR_REG_2_, n73502 );
nand U126826 ( n67376, n67435, n67436 );
nand U126827 ( n67435, P2_P3_INSTADDRPOINTER_REG_29_, n67437 );
nand U126828 ( n67436, n67378, n76198 );
nor U126829 ( n67380, n67382, n67383 );
nor U126830 ( n67383, P2_P3_INSTADDRPOINTER_REG_30_, n67376 );
nor U126831 ( n67382, n67384, n76197 );
nor U126832 ( n67384, n75068, n67385 );
nand U126833 ( n71327, n72058, n72059 );
nor U126834 ( n72058, n72062, n72063 );
nor U126835 ( n72059, n72060, n72061 );
and U126836 ( n72063, P4_ADDR_REG_2_, P4_WR_REG );
nand U126837 ( n23877, P1_P2_INSTQUEUERD_ADDR_REG_2_, n73503 );
nand U126838 ( n57001, P2_P2_INSTQUEUERD_ADDR_REG_2_, n73504 );
nand U126839 ( n68235, n68265, n68266 );
nand U126840 ( n68265, n68268, n76197 );
nand U126841 ( n68266, P2_P3_INSTADDRPOINTER_REG_7_, n68267 );
or U126842 ( n68267, n68268, n76198 );
nand U126843 ( n26234, n26264, n26265 );
nand U126844 ( n26264, n26267, n76521 );
nand U126845 ( n26265, P1_P2_INSTADDRPOINTER_REG_7_, n26266 );
or U126846 ( n26266, n26267, n76522 );
nand U126847 ( n59373, n59403, n59404 );
nand U126848 ( n59403, n59406, n76263 );
nand U126849 ( n59404, P2_P2_INSTADDRPOINTER_REG_7_, n59405 );
or U126850 ( n59405, n59406, n76264 );
nand U126851 ( n25371, n25430, n25431 );
nand U126852 ( n25430, P1_P2_INSTADDRPOINTER_REG_29_, n25432 );
nand U126853 ( n25431, n25373, n76522 );
nand U126854 ( n58508, n58567, n58568 );
nand U126855 ( n58567, P2_P2_INSTADDRPOINTER_REG_29_, n58569 );
nand U126856 ( n58568, n58510, n76264 );
nand U126857 ( n24717, n25536, n25537 );
nand U126858 ( n25537, P1_P2_INSTADDRPOINTER_REG_26_, n25538 );
nand U126859 ( n25538, n76525, n25539 );
nand U126860 ( n25539, P1_P2_INSTADDRPOINTER_REG_25_, n25540 );
nand U126861 ( n66552, n67541, n67542 );
nand U126862 ( n67542, P2_P3_INSTADDRPOINTER_REG_26_, n67543 );
nand U126863 ( n67543, n76201, n67544 );
nand U126864 ( n67544, P2_P3_INSTADDRPOINTER_REG_25_, n67545 );
nand U126865 ( n57851, n58673, n58674 );
nand U126866 ( n58674, P2_P2_INSTADDRPOINTER_REG_26_, n58675 );
nand U126867 ( n58675, n76267, n58676 );
nand U126868 ( n58676, P2_P2_INSTADDRPOINTER_REG_25_, n58677 );
nand U126869 ( n67664, n67696, n67697 );
nor U126870 ( n67696, n5748, n67698 );
nor U126871 ( n67698, P2_P3_INSTADDRPOINTER_REG_22_, n76197 );
nand U126872 ( n25659, n25691, n25692 );
nor U126873 ( n25691, n3990, n25693 );
nor U126874 ( n25693, P1_P2_INSTADDRPOINTER_REG_22_, n76521 );
nand U126875 ( n58799, n58831, n58832 );
nor U126876 ( n58831, n6623, n58833 );
nor U126877 ( n58833, P2_P2_INSTADDRPOINTER_REG_22_, n76263 );
nor U126878 ( n25499, n24717, P1_P2_INSTADDRPOINTER_REG_27_ );
nor U126879 ( n67504, n66552, P2_P3_INSTADDRPOINTER_REG_27_ );
nor U126880 ( n58636, n57851, P2_P2_INSTADDRPOINTER_REG_27_ );
nor U126881 ( n68056, n68152, n68153 );
and U126882 ( n68153, P2_P3_INSTADDRPOINTER_REG_10_, n68154 );
nand U126883 ( n68154, n76201, n68155 );
nor U126884 ( n26053, n26151, n26152 );
and U126885 ( n26152, P1_P2_INSTADDRPOINTER_REG_10_, n26153 );
nand U126886 ( n26153, n76525, n26154 );
nor U126887 ( n59194, n59290, n59291 );
and U126888 ( n59291, P2_P2_INSTADDRPOINTER_REG_10_, n59292 );
nand U126889 ( n59292, n76267, n59293 );
nand U126890 ( n25380, P1_P2_INSTADDRPOINTER_REG_30_, n25371 );
nand U126891 ( n67385, P2_P3_INSTADDRPOINTER_REG_30_, n67376 );
nand U126892 ( n58517, P2_P2_INSTADDRPOINTER_REG_30_, n58508 );
nand U126893 ( n25432, n25455, n25456 );
nand U126894 ( n25456, P1_P2_INSTADDRPOINTER_REG_28_, n76521 );
nor U126895 ( n25455, n24719, n25457 );
nor U126896 ( n25457, n3989, n25428 );
nand U126897 ( n67437, n67460, n67461 );
nand U126898 ( n67461, P2_P3_INSTADDRPOINTER_REG_28_, n76197 );
nor U126899 ( n67460, n66554, n67462 );
nor U126900 ( n67462, n5747, n67433 );
nand U126901 ( n58569, n58592, n58593 );
nand U126902 ( n58593, P2_P2_INSTADDRPOINTER_REG_28_, n76263 );
nor U126903 ( n58592, n57853, n58594 );
nor U126904 ( n58594, n6622, n58565 );
nand U126905 ( n67739, n67884, n67885 );
nand U126906 ( n67885, P2_P3_INSTADDRPOINTER_REG_17_, n76197 );
nor U126907 ( n67884, n5750, n67886 );
nor U126908 ( n67886, n5752, n67865 );
nand U126909 ( n58874, n59019, n59020 );
nand U126910 ( n59020, P2_P2_INSTADDRPOINTER_REG_17_, n76263 );
nor U126911 ( n59019, n6625, n59021 );
nor U126912 ( n59021, n6627, n59000 );
nand U126913 ( n66470, n67370, n67371 );
nand U126914 ( n67371, n67372, n67373 );
nand U126915 ( n67370, n67380, n67381 );
nand U126916 ( n67373, n75990, P2_P3_INSTADDRPOINTER_REG_31_ );
nor U126917 ( n25375, n25377, n25378 );
nor U126918 ( n25378, P1_P2_INSTADDRPOINTER_REG_30_, n25371 );
nor U126919 ( n25377, n25379, n76521 );
nor U126920 ( n25379, n75066, n25380 );
nor U126921 ( n58512, n58514, n58515 );
nor U126922 ( n58515, P2_P2_INSTADDRPOINTER_REG_30_, n58508 );
nor U126923 ( n58514, n58516, n76263 );
nor U126924 ( n58516, n75067, n58517 );
nand U126925 ( n68155, n68191, P2_P3_INSTADDRPOINTER_REG_8_ );
nor U126926 ( n68191, n5758, n73084 );
nand U126927 ( n26154, n26190, P1_P2_INSTADDRPOINTER_REG_8_ );
nor U126928 ( n26190, n4000, n73085 );
nand U126929 ( n59293, n59329, P2_P2_INSTADDRPOINTER_REG_8_ );
nor U126930 ( n59329, n6633, n73086 );
nand U126931 ( n25734, n25881, n25882 );
nand U126932 ( n25882, P1_P2_INSTADDRPOINTER_REG_17_, n76521 );
nor U126933 ( n25881, n3993, n25883 );
nor U126934 ( n25883, n3994, n25862 );
nor U126935 ( n72061, n73491, n71283 );
nand U126936 ( n24633, n25365, n25366 );
nand U126937 ( n25366, n25367, n25368 );
nand U126938 ( n25365, n25375, n25376 );
nand U126939 ( n25368, n76027, P1_P2_INSTADDRPOINTER_REG_31_ );
nand U126940 ( n57765, n58502, n58503 );
nand U126941 ( n58503, n58504, n58505 );
nand U126942 ( n58502, n58512, n58513 );
nand U126943 ( n58505, n75998, P2_P2_INSTADDRPOINTER_REG_31_ );
or U126944 ( n25373, n25432, P1_P2_INSTADDRPOINTER_REG_29_ );
or U126945 ( n67378, n67437, P2_P3_INSTADDRPOINTER_REG_29_ );
or U126946 ( n58510, n58569, P2_P2_INSTADDRPOINTER_REG_29_ );
nand U126947 ( n67922, n67958, n67959 );
nand U126948 ( n67958, n67961, n76197 );
nand U126949 ( n67959, P2_P3_INSTADDRPOINTER_REG_15_, n67960 );
or U126950 ( n67960, n67961, n76198 );
nand U126951 ( n25919, n25955, n25956 );
nand U126952 ( n25955, n25958, n76521 );
nand U126953 ( n25956, P1_P2_INSTADDRPOINTER_REG_15_, n25957 );
or U126954 ( n25957, n25958, n76522 );
nand U126955 ( n59057, n59093, n59094 );
nand U126956 ( n59093, n59096, n76263 );
nand U126957 ( n59094, P2_P2_INSTADDRPOINTER_REG_15_, n59095 );
or U126958 ( n59095, n59096, n76264 );
nand U126959 ( n67545, n67625, n67626 );
nand U126960 ( n67625, n67628, n76197 );
nand U126961 ( n67626, P2_P3_INSTADDRPOINTER_REG_24_, n67627 );
or U126962 ( n67627, n67628, n76198 );
nand U126963 ( n25540, n25620, n25621 );
nand U126964 ( n25620, n25623, n76521 );
nand U126965 ( n25621, P1_P2_INSTADDRPOINTER_REG_24_, n25622 );
or U126966 ( n25622, n25623, n76522 );
nand U126967 ( n58677, n58757, n58758 );
nand U126968 ( n58757, n58760, n76263 );
nand U126969 ( n58758, P2_P2_INSTADDRPOINTER_REG_24_, n58759 );
or U126970 ( n58759, n58760, n76264 );
and U126971 ( n51092, n49834, P3_DATAO_REG_12_ );
nor U126972 ( n71611, n73481, n71283 );
nand U126973 ( n18834, n8217, P4_DATAO_REG_1_ );
and U126974 ( n49809, DIN_16_, n76929 );
nand U126975 ( n51538, n49809, P3_DATAO_REG_8_ );
nand U126976 ( n24215, P1_P2_INSTQUEUERD_ADDR_REG_1_, P1_P2_INSTQUEUERD_ADDR_REG_0_ );
nand U126977 ( n57337, P2_P2_INSTQUEUERD_ADDR_REG_1_, P2_P2_INSTQUEUERD_ADDR_REG_0_ );
nand U126978 ( n65759, P2_P3_INSTQUEUERD_ADDR_REG_1_, P2_P3_INSTQUEUERD_ADDR_REG_0_ );
nor U126979 ( n71610, n73482, n71284 );
and U126980 ( n52317, n49834, P3_DATAO_REG_3_ );
nand U126981 ( n41119, n64526, n64527 );
nand U126982 ( n64527, n76390, n43866 );
nand U126983 ( n64526, P1_P3_DATAO_REG_13_, n76389 );
nand U126984 ( n40935, n64815, n64816 );
nand U126985 ( n64816, n76390, n43666 );
nand U126986 ( n64815, P1_P3_DATAO_REG_12_, n76389 );
nor U126987 ( n71612, n73483, n71287 );
nand U126988 ( n2586, n38668, n38669 );
nand U126989 ( n38668, P4_REG1_REG_16_, n76425 );
nand U126990 ( n38669, n76016, n38670 );
nand U126991 ( n2426, n39562, n39563 );
nand U126992 ( n39562, P4_REG0_REG_16_, n76422 );
nand U126993 ( n39563, n76013, n38670 );
and U126994 ( n19829, P4_DATAO_REG_5_, n76170 );
nand U126995 ( n51894, n49809, P3_DATAO_REG_7_ );
nor U126996 ( n46307, n46309, n46310 );
nor U126997 ( n46309, n76005, n46312 );
and U126998 ( n46310, n46311, P2_P1_INSTADDRPOINTER_REG_30_ );
nor U126999 ( n46312, n46313, n46314 );
and U127000 ( n16879, DIN_14_, n76927 );
nand U127001 ( n19079, n16879, P4_DATAO_REG_8_ );
nand U127002 ( n17770, P4_DATAO_REG_16_, n76171 );
nor U127003 ( n25367, n25369, n25370 );
nor U127004 ( n25369, n76026, n25372 );
and U127005 ( n25370, n25371, P1_P2_INSTADDRPOINTER_REG_30_ );
nor U127006 ( n25372, n25373, n25374 );
nor U127007 ( n67372, n67374, n67375 );
nor U127008 ( n67374, n75989, n67377 );
and U127009 ( n67375, n67376, P2_P3_INSTADDRPOINTER_REG_30_ );
nor U127010 ( n67377, n67378, n67379 );
nor U127011 ( n58504, n58506, n58507 );
nor U127012 ( n58506, n75997, n58509 );
and U127013 ( n58507, n58508, P2_P2_INSTADDRPOINTER_REG_30_ );
nor U127014 ( n58509, n58510, n58511 );
nand U127015 ( n52663, n49834, P3_DATAO_REG_4_ );
and U127016 ( n19674, P4_DATAO_REG_4_, n76165 );
nand U127017 ( n44515, n7809, P2_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U127018 ( n2596, n38662, n38663 );
nand U127019 ( n38662, P4_REG1_REG_18_, n76425 );
nand U127020 ( n38663, n76016, n38664 );
nand U127021 ( n2436, n39433, n39434 );
nand U127022 ( n39433, P4_REG0_REG_18_, n76422 );
nand U127023 ( n39434, n76013, n38664 );
nand U127024 ( n36327, n39750, n39751 );
nand U127025 ( n39751, n76459, n37930 );
nand U127026 ( n39750, P2_P3_DATAO_REG_14_, n76458 );
nor U127027 ( n44132, n44894, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nor U127028 ( n71453, n73493, n71283 );
and U127029 ( n66280, n76253, P3_REG0_REG_6_ );
nand U127030 ( n52169, n49834, P3_DATAO_REG_2_ );
nand U127031 ( n50716, n49834, P3_DATAO_REG_14_ );
nand U127032 ( n18951, n16879, P4_DATAO_REG_9_ );
nand U127033 ( n65390, n6022, P2_P3_INSTQUEUERD_ADDR_REG_0_ );
nand U127034 ( n23844, n4244, P1_P2_INSTQUEUERD_ADDR_REG_0_ );
nand U127035 ( n56968, n6877, P2_P2_INSTQUEUERD_ADDR_REG_0_ );
nor U127036 ( n56587, n57337, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nor U127037 ( n23465, n24215, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nor U127038 ( n64974, n65759, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U127039 ( n19519, P4_DATAO_REG_3_, n76168 );
nand U127040 ( n51375, n49809, P3_DATAO_REG_9_ );
and U127041 ( n46344, n75924, n75925 );
nand U127042 ( n75924, n45563, n76657 );
nand U127043 ( n75925, n46329, P2_P1_INSTADDRPOINTER_REG_30_ );
nand U127044 ( n15681, n46335, n46336 );
nand U127045 ( n46336, n76859, P2_P1_INSTADDRPOINTER_REG_30_ );
nor U127046 ( n46335, n46337, n46338 );
nor U127047 ( n46338, n75237, n76334 );
nand U127048 ( n36577, n39621, n39622 );
nand U127049 ( n39622, n76459, n37955 );
nand U127050 ( n39621, P2_P3_DATAO_REG_16_, n76457 );
and U127051 ( n25403, n75926, n75927 );
nand U127052 ( n75926, n24651, n76751 );
nand U127053 ( n75927, n25388, P1_P2_INSTADDRPOINTER_REG_30_ );
and U127054 ( n58540, n75928, n75929 );
nand U127055 ( n75928, n57787, n76684 );
nand U127056 ( n75929, n58525, P2_P2_INSTADDRPOINTER_REG_30_ );
and U127057 ( n67408, n75930, n75931 );
nand U127058 ( n75930, n66488, n76705 );
nand U127059 ( n75931, n67393, P2_P3_INSTADDRPOINTER_REG_30_ );
nand U127060 ( n6701, n25394, n25395 );
nand U127061 ( n25395, n76520, P1_P2_INSTADDRPOINTER_REG_30_ );
nor U127062 ( n25394, n25396, n25397 );
nor U127063 ( n25397, n75064, n76908 );
nand U127064 ( n13436, n58531, n58532 );
nand U127065 ( n58532, n76262, P2_P2_INSTADDRPOINTER_REG_30_ );
nor U127066 ( n58531, n58533, n58534 );
nor U127067 ( n58534, n75063, n76882 );
nand U127068 ( n11191, n67399, n67400 );
nand U127069 ( n67400, n76196, P2_P3_INSTADDRPOINTER_REG_30_ );
nor U127070 ( n67399, n67401, n67402 );
nor U127071 ( n67402, n75070, n76873 );
buf U127072 ( n76787, n2358 );
not U127073 ( n2358, P4_DATAO_REG_0_ );
and U127074 ( n66356, n76254, P3_REG0_REG_5_ );
nor U127075 ( n72695, n73500, n71104 );
and U127076 ( n52513, n49809, P3_DATAO_REG_5_ );
nand U127077 ( n46425, P2_P1_INSTADDRPOINTER_REG_28_, n46426 );
nand U127078 ( n46426, n46427, n46428 );
nor U127079 ( n46427, n46388, n46435 );
nor U127080 ( n46428, n46429, n46430 );
nand U127081 ( n15671, n46417, n46418 );
nand U127082 ( n46418, n76859, P2_P1_INSTADDRPOINTER_REG_28_ );
nor U127083 ( n46417, n46419, n46420 );
nor U127084 ( n46420, n75302, n76334 );
nand U127085 ( n67489, P2_P3_INSTADDRPOINTER_REG_28_, n67490 );
nand U127086 ( n67490, n67491, n67492 );
nor U127087 ( n67491, n67452, n67499 );
nor U127088 ( n67492, n67493, n67494 );
nand U127089 ( n25484, P1_P2_INSTADDRPOINTER_REG_28_, n25485 );
nand U127090 ( n25485, n25486, n25487 );
nor U127091 ( n25486, n25447, n25494 );
nor U127092 ( n25487, n25488, n25489 );
nand U127093 ( n58621, P2_P2_INSTADDRPOINTER_REG_28_, n58622 );
nand U127094 ( n58622, n58623, n58624 );
nor U127095 ( n58623, n58584, n58631 );
nor U127096 ( n58624, n58625, n58626 );
nand U127097 ( n11181, n67481, n67482 );
nand U127098 ( n67482, n76196, P2_P3_INSTADDRPOINTER_REG_28_ );
nor U127099 ( n67481, n67483, n67484 );
nor U127100 ( n67484, n75361, n76873 );
nand U127101 ( n6691, n25476, n25477 );
nand U127102 ( n25477, n76520, P1_P2_INSTADDRPOINTER_REG_28_ );
nor U127103 ( n25476, n25478, n25479 );
nor U127104 ( n25479, n75301, n76908 );
nand U127105 ( n13426, n58613, n58614 );
nand U127106 ( n58614, n76262, P2_P2_INSTADDRPOINTER_REG_28_ );
nor U127107 ( n58613, n58615, n58616 );
nor U127108 ( n58616, n75300, n76882 );
nand U127109 ( n19966, n16879, P4_DATAO_REG_6_ );
nand U127110 ( n44511, P2_P1_INSTQUEUERD_ADDR_REG_0_, n47864 );
nor U127111 ( n40096, n76414, n74318 );
nand U127112 ( n40732, n64388, n64389 );
nand U127113 ( n64389, n76390, n44395 );
nand U127114 ( n64388, P1_P3_DATAO_REG_14_, n76389 );
nand U127115 ( n1361, n57726, n57727 );
nand U127116 ( n57726, P3_REG1_REG_16_, n76288 );
nand U127117 ( n57727, n76003, n57728 );
nand U127118 ( n1201, n63978, n63979 );
nand U127119 ( n63978, P3_REG0_REG_16_, n76255 );
nand U127120 ( n63979, n75995, n57728 );
nand U127121 ( n51889, n49809, P3_DATAO_REG_6_ );
nand U127122 ( n41323, n64234, n64235 );
nand U127123 ( n64235, n76390, n44857 );
nand U127124 ( n64234, P1_P3_DATAO_REG_15_, n76389 );
and U127125 ( n18548, n16879, P4_DATAO_REG_10_ );
nand U127126 ( n1211, n63253, n63254 );
nand U127127 ( n63253, P3_REG0_REG_18_, n76255 );
nand U127128 ( n63254, n75995, n57634 );
nand U127129 ( n1371, n57632, n57633 );
nand U127130 ( n57632, P3_REG1_REG_18_, n76288 );
nand U127131 ( n57633, n76003, n57634 );
nand U127132 ( n65386, P2_P3_INSTQUEUERD_ADDR_REG_0_, n68884 );
nand U127133 ( n23840, P1_P2_INSTQUEUERD_ADDR_REG_0_, n26885 );
nand U127134 ( n56964, P2_P2_INSTQUEUERD_ADDR_REG_0_, n60025 );
and U127135 ( n19197, P4_DATAO_REG_2_, n76166 );
nand U127136 ( n71096, n72834, n72835 );
nand U127137 ( n72834, P4_WR_REG, P4_ADDR_REG_1_ );
nand U127138 ( n72835, n71000, n73025 );
nand U127139 ( n71000, n72836, n72837 );
nand U127140 ( n72837, n1244, P1_P1_ADDRESS_REG_1_ );
nor U127141 ( n72836, n72838, n72839 );
nor U127142 ( n72838, n73488, n71009 );
nor U127143 ( n72839, n73486, n71013 );
nand U127144 ( n19852, n16879, P4_DATAO_REG_7_ );
and U127145 ( n43975, n45458, n45459 );
nand U127146 ( n45458, P2_BUF1_REG_11_, n76477 );
nand U127147 ( n45459, n45460, n31928 );
xor U127148 ( n45460, n45461, n45462 );
nand U127149 ( n15946, n45372, n45373 );
nand U127150 ( n45373, P2_P1_UWORD_REG_11_, n76352 );
nor U127151 ( n45372, n45374, n45375 );
nor U127152 ( n45375, n73320, n76350 );
nand U127153 ( n15871, n45455, n45456 );
nand U127154 ( n45456, P2_P1_LWORD_REG_11_, n76352 );
nor U127155 ( n45455, n45374, n45457 );
nor U127156 ( n45457, n73237, n76349 );
nand U127157 ( n16221, n44728, n44729 );
nor U127158 ( n44729, n44730, n44731 );
nor U127159 ( n44728, n44735, n44736 );
nor U127160 ( n44730, P2_P1_EAX_REG_11_, n44694 );
nand U127161 ( n40972, n64033, n64034 );
nand U127162 ( n64034, n76390, n45007 );
nand U127163 ( n64033, P1_P3_DATAO_REG_16_, n76389 );
buf U127164 ( n76833, n1217 );
not U127165 ( n1217, P3_DATAO_REG_0_ );
nand U127166 ( n18432, n16879, P4_DATAO_REG_11_ );
and U127167 ( n40097, n76419, P4_REG0_REG_7_ );
nand U127168 ( n2591, n38665, n38666 );
nand U127169 ( n38665, P4_REG1_REG_17_, n76425 );
nand U127170 ( n38666, n76016, n38667 );
nand U127171 ( n2431, n39504, n39505 );
nand U127172 ( n39504, P4_REG0_REG_17_, n76422 );
nand U127173 ( n39505, n76013, n38667 );
nand U127174 ( n17223, P4_DATAO_REG_16_, n16879 );
nand U127175 ( n18034, P4_DATAO_REG_15_, n76170 );
nor U127176 ( n39971, n76414, n74358 );
nand U127177 ( n36618, n39557, n39558 );
nand U127178 ( n39558, n76459, n37969 );
nand U127179 ( n39557, P2_P3_DATAO_REG_17_, n76457 );
nor U127180 ( n40005, n76414, n74366 );
and U127181 ( n50834, n49834, P3_DATAO_REG_13_ );
nand U127182 ( n2581, n38671, n38672 );
nand U127183 ( n38671, P4_REG1_REG_15_, n76425 );
nand U127184 ( n38672, n76016, n38673 );
nand U127185 ( n2421, n39628, n39629 );
nand U127186 ( n39628, P4_REG0_REG_15_, n76422 );
nand U127187 ( n39629, n76013, n38673 );
and U127188 ( n66187, n76253, P3_REG0_REG_7_ );
nand U127189 ( n50145, n49809, P3_DATAO_REG_14_ );
nand U127190 ( n1366, n57676, n57677 );
nand U127191 ( n57676, P3_REG1_REG_17_, n76288 );
nand U127192 ( n57677, n76003, n57678 );
nand U127193 ( n1206, n63653, n63654 );
nand U127194 ( n63653, P3_REG0_REG_17_, n76255 );
nand U127195 ( n63654, n75995, n57678 );
and U127196 ( n51800, n49834, P3_DATAO_REG_1_ );
nand U127197 ( n51202, n49809, P3_DATAO_REG_10_ );
nand U127198 ( n49967, n8238, P3_DATAO_REG_20_ );
and U127199 ( n39972, n76419, P4_REG0_REG_10_ );
nand U127200 ( n47157, P2_P1_INSTADDRPOINTER_REG_8_, n76341 );
nand U127201 ( n19834, n16879, P4_DATAO_REG_5_ );
and U127202 ( n40006, n76419, P4_REG0_REG_9_ );
xor U127203 ( n45605, n46395, n46373 );
xor U127204 ( n46395, n76342, P2_P1_INSTADDRPOINTER_REG_29_ );
nand U127205 ( n15676, n46374, n46375 );
nand U127206 ( n46375, n76859, P2_P1_INSTADDRPOINTER_REG_29_ );
nor U127207 ( n46374, n46376, n46377 );
nor U127208 ( n46377, n73391, n76334 );
xor U127209 ( n66530, n67459, n67437 );
xor U127210 ( n67459, n76198, P2_P3_INSTADDRPOINTER_REG_29_ );
xor U127211 ( n24695, n25454, n25432 );
xor U127212 ( n25454, n76522, P1_P2_INSTADDRPOINTER_REG_29_ );
xor U127213 ( n57829, n58591, n58569 );
xor U127214 ( n58591, n76264, P2_P2_INSTADDRPOINTER_REG_29_ );
nand U127215 ( n11186, n67438, n67439 );
nand U127216 ( n67439, n76196, P2_P3_INSTADDRPOINTER_REG_29_ );
nor U127217 ( n67438, n67440, n67441 );
nor U127218 ( n67441, n73319, n76873 );
nand U127219 ( n6696, n25433, n25434 );
nand U127220 ( n25434, n76520, P1_P2_INSTADDRPOINTER_REG_29_ );
nor U127221 ( n25433, n25435, n25436 );
nor U127222 ( n25436, n73317, n76908 );
nand U127223 ( n13431, n58570, n58571 );
nand U127224 ( n58571, n76262, P2_P2_INSTADDRPOINTER_REG_29_ );
nor U127225 ( n58570, n58572, n58573 );
nor U127226 ( n58573, n73316, n76882 );
nand U127227 ( n49849, n8237, P3_DATAO_REG_21_ );
and U127228 ( n44020, n45448, n45449 );
nand U127229 ( n45448, P2_BUF1_REG_10_, n76477 );
nand U127230 ( n45449, n45450, n31928 );
xnor U127231 ( n45450, n45451, n45452 );
nand U127232 ( n15876, n45445, n45446 );
nand U127233 ( n45446, P2_P1_LWORD_REG_10_, n76352 );
nor U127234 ( n45445, n45370, n45447 );
nor U127235 ( n45447, n74786, n76349 );
nand U127236 ( n15951, n45368, n45369 );
nand U127237 ( n45369, P2_P1_UWORD_REG_10_, n76352 );
nor U127238 ( n45368, n45370, n45371 );
nor U127239 ( n45371, n75084, n76350 );
nand U127240 ( n68188, P2_P3_INSTADDRPOINTER_REG_8_, n76197 );
nand U127241 ( n26187, P1_P2_INSTADDRPOINTER_REG_8_, n76521 );
nand U127242 ( n59326, P2_P2_INSTADDRPOINTER_REG_8_, n76263 );
and U127243 ( n40051, n76419, P4_REG0_REG_8_ );
and U127244 ( n65808, n76253, P3_REG0_REG_11_ );
and U127245 ( n10059, n11682, n11683 );
nand U127246 ( n11682, P1_BUF1_REG_11_, n76610 );
nand U127247 ( n11683, n11684, n76612 );
xor U127248 ( n11684, n11685, n11687 );
nand U127249 ( n9211, n11564, n11565 );
nand U127250 ( n11565, P1_P1_UWORD_REG_11_, n76618 );
nor U127251 ( n11564, n11567, n11568 );
nor U127252 ( n11568, n73321, n76616 );
nand U127253 ( n9136, n11678, n11679 );
nand U127254 ( n11679, P1_P1_LWORD_REG_11_, n76618 );
nor U127255 ( n11678, n11567, n11680 );
nor U127256 ( n11680, n73238, n76615 );
and U127257 ( n18027, P4_DATAO_REG_14_, n76169 );
nand U127258 ( n9486, n10994, n10995 );
nor U127259 ( n10995, n10997, n10998 );
nor U127260 ( n10994, n11003, n11004 );
nor U127261 ( n10997, P1_P1_EAX_REG_11_, n10952 );
nand U127262 ( n1196, n64185, n64186 );
nand U127263 ( n64185, P3_REG0_REG_15_, n76255 );
nand U127264 ( n64186, n75995, n57998 );
nand U127265 ( n1356, n57996, n57997 );
nand U127266 ( n57996, P3_REG1_REG_15_, n76288 );
nand U127267 ( n57997, n76003, n57998 );
and U127268 ( n65932, n76253, P3_REG0_REG_10_ );
nor U127269 ( n66097, n76248, n74383 );
nand U127270 ( n18839, P4_DATAO_REG_1_, n76167 );
nand U127271 ( n41011, n63710, n63711 );
nand U127272 ( n63711, n76390, n45077 );
nand U127273 ( n63710, P1_P3_DATAO_REG_17_, n76389 );
nand U127274 ( n2416, n39684, n39685 );
nand U127275 ( n39684, P4_REG0_REG_14_, n76422 );
nand U127276 ( n39685, n76013, n38676 );
nand U127277 ( n2576, n38674, n38675 );
nand U127278 ( n38674, P4_REG1_REG_14_, n76425 );
nand U127279 ( n38675, n76016, n38676 );
nand U127280 ( n31169, P1_P3_INSTQUEUERD_ADDR_REG_2_, n73524 );
nand U127281 ( n32867, n33128, n33129 );
nand U127282 ( n33129, P1_P3_INSTADDRPOINTER_REG_17_, n76472 );
nor U127283 ( n33128, n32229, n33130 );
nor U127284 ( n33130, n3152, n33109 );
nand U127285 ( n32611, n32670, n32671 );
nand U127286 ( n32670, P1_P3_INSTADDRPOINTER_REG_29_, n32672 );
nand U127287 ( n32671, n32613, n76472 );
nand U127288 ( n31949, n32776, n32777 );
nand U127289 ( n32777, P1_P3_INSTADDRPOINTER_REG_26_, n32778 );
nand U127290 ( n32778, n76475, n32779 );
nand U127291 ( n32779, P1_P3_INSTADDRPOINTER_REG_25_, n32780 );
nor U127292 ( n32739, n31949, P1_P3_INSTADDRPOINTER_REG_27_ );
nor U127293 ( n33165, n32227, P1_P3_INSTADDRPOINTER_REG_16_ );
nand U127294 ( n32227, n33203, n33204 );
nand U127295 ( n33203, n33206, n76472 );
nand U127296 ( n33204, P1_P3_INSTADDRPOINTER_REG_15_, n33205 );
or U127297 ( n33205, n33206, n76471 );
nand U127298 ( n32620, P1_P3_INSTADDRPOINTER_REG_30_, n32611 );
nand U127299 ( n33484, n33510, n33511 );
nand U127300 ( n33510, n33513, n76472 );
nand U127301 ( n33511, P1_P3_INSTADDRPOINTER_REG_7_, n33512 );
or U127302 ( n33512, n33513, n76472 );
nand U127303 ( n32672, n32695, n32696 );
nand U127304 ( n32696, P1_P3_INSTADDRPOINTER_REG_28_, n76472 );
nor U127305 ( n32695, n31951, n32697 );
nor U127306 ( n32697, n3150, n32668 );
nand U127307 ( n33206, n33242, n33243 );
nand U127308 ( n33242, n33245, n76472 );
nand U127309 ( n33243, P1_P3_INSTADDRPOINTER_REG_14_, n33244 );
or U127310 ( n33244, n33245, n76472 );
nand U127311 ( n31847, n32605, n32606 );
nand U127312 ( n32606, n32607, n32608 );
nand U127313 ( n32605, n32615, n32616 );
nand U127314 ( n32608, n76475, P1_P3_INSTADDRPOINTER_REG_31_ );
nor U127315 ( n32615, n32617, n32618 );
nor U127316 ( n32618, P1_P3_INSTADDRPOINTER_REG_30_, n32611 );
nor U127317 ( n32617, n32619, n76470 );
nor U127318 ( n32619, n75065, n32620 );
or U127319 ( n32613, n32672, P1_P3_INSTADDRPOINTER_REG_29_ );
nand U127320 ( n33370, n33481, n33482 );
nand U127321 ( n33481, n33484, n76472 );
nand U127322 ( n33482, P1_P3_INSTADDRPOINTER_REG_8_, n33483 );
or U127323 ( n33483, n33484, n76471 );
nand U127324 ( n31509, P1_P3_INSTQUEUERD_ADDR_REG_1_, P1_P3_INSTQUEUERD_ADDR_REG_0_ );
nand U127325 ( n52655, n49809, P3_DATAO_REG_4_ );
nand U127326 ( n17491, P4_DATAO_REG_15_, n16879 );
nand U127327 ( n72789, P3_WR_REG, P3_ADDR_REG_1_ );
and U127328 ( n66098, n76253, P3_REG0_REG_8_ );
and U127329 ( n49990, DIN_18_, n76929 );
nand U127330 ( n51514, n49990, P3_DATAO_REG_6_ );
and U127331 ( n50704, n49809, P3_DATAO_REG_11_ );
and U127332 ( n66012, n76253, P3_REG0_REG_9_ );
and U127333 ( n16854, DIN_16_, n76927 );
nand U127334 ( n50433, n49809, P3_DATAO_REG_13_ );
nand U127335 ( n18582, n16854, P4_DATAO_REG_8_ );
nand U127336 ( n1191, n64333, n64334 );
nand U127337 ( n64333, P3_REG0_REG_14_, n76255 );
nand U127338 ( n64334, n75995, n58227 );
nand U127339 ( n1351, n58225, n58226 );
nand U127340 ( n58225, P3_REG1_REG_14_, n76288 );
nand U127341 ( n58226, n76003, n58227 );
nor U127342 ( n32607, n32609, n32610 );
nor U127343 ( n32609, n76021, n32612 );
and U127344 ( n32610, n32611, P1_P3_INSTADDRPOINTER_REG_30_ );
nor U127345 ( n32612, n32613, n32614 );
nor U127346 ( n30772, n31509, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nor U127347 ( n39928, n76414, n74394 );
nand U127348 ( n45609, n45619, n45620 );
nand U127349 ( n45619, n45631, P2_P1_PHYADDRPOINTER_REG_27_ );
nand U127350 ( n45620, n45621, n45622 );
and U127351 ( n45631, n74891, n45632 );
nand U127352 ( n24699, n24709, n24710 );
nand U127353 ( n24709, n24720, P1_P2_PHYADDRPOINTER_REG_27_ );
nand U127354 ( n24710, n24711, n24712 );
and U127355 ( n24720, n75243, n24721 );
nand U127356 ( n66534, n66544, n66545 );
nand U127357 ( n66544, n66555, P2_P3_PHYADDRPOINTER_REG_27_ );
nand U127358 ( n66545, n66546, n66547 );
and U127359 ( n66555, n75244, n66556 );
nand U127360 ( n57833, n57843, n57844 );
nand U127361 ( n57843, n57854, P2_P2_PHYADDRPOINTER_REG_27_ );
nand U127362 ( n57844, n57845, n57846 );
and U127363 ( n57854, n75245, n57855 );
nand U127364 ( n18938, n16854, P4_DATAO_REG_7_ );
nand U127365 ( n36802, n39496, n39497 );
nand U127366 ( n39497, n76459, n38038 );
nand U127367 ( n39496, P2_P3_DATAO_REG_18_, n76457 );
and U127368 ( n10115, n11669, n11670 );
nand U127369 ( n11669, P1_BUF1_REG_10_, n76610 );
nand U127370 ( n11670, n11672, n76612 );
xnor U127371 ( n11672, n11673, n11674 );
nand U127372 ( n9141, n11665, n11667 );
nand U127373 ( n11667, P1_P1_LWORD_REG_10_, n76618 );
nor U127374 ( n11665, n11562, n11668 );
nor U127375 ( n11668, n74787, n76615 );
nand U127376 ( n9216, n11559, n11560 );
nand U127377 ( n11560, P1_P1_UWORD_REG_10_, n76618 );
nor U127378 ( n11559, n11562, n11563 );
nor U127379 ( n11563, n75085, n76616 );
and U127380 ( n18129, n16879, P4_DATAO_REG_12_ );
nand U127381 ( n51362, n49990, P3_DATAO_REG_7_ );
nand U127382 ( n1346, n58433, n58434 );
nand U127383 ( n58433, P3_REG1_REG_13_, n76288 );
nand U127384 ( n58434, n76003, n58435 );
nand U127385 ( n1186, n64486, n64487 );
nand U127386 ( n64486, P3_REG0_REG_13_, n76255 );
nand U127387 ( n64487, n75995, n58435 );
nand U127388 ( n31136, n3407, P1_P3_INSTQUEUERD_ADDR_REG_0_ );
nand U127389 ( n41183, n63313, n63314 );
nand U127390 ( n63314, n76390, n45270 );
nand U127391 ( n63313, P1_P3_DATAO_REG_18_, n76389 );
nand U127392 ( n51875, n49990, P3_DATAO_REG_5_ );
and U127393 ( n32643, n75932, n75933 );
nand U127394 ( n75932, n31865, n76772 );
nand U127395 ( n75933, n32628, P1_P3_INSTADDRPOINTER_REG_30_ );
nand U127396 ( n4456, n32634, n32635 );
nand U127397 ( n32635, n76469, P1_P3_INSTADDRPOINTER_REG_30_ );
nor U127398 ( n32634, n32636, n32637 );
nor U127399 ( n32637, n75069, n76899 );
nand U127400 ( n19707, n16879, P4_DATAO_REG_4_ );
nand U127401 ( n2571, n38677, n38678 );
nand U127402 ( n38677, P4_REG1_REG_13_, n76425 );
nand U127403 ( n38678, n76016, n38679 );
nand U127404 ( n2411, n39757, n39758 );
nand U127405 ( n39757, P4_REG0_REG_13_, n76422 );
nand U127406 ( n39758, n76013, n38679 );
nand U127407 ( n2501, n38730, n38731 );
nand U127408 ( n38730, P4_REG0_REG_31_, n76422 );
nand U127409 ( n38731, n76012, n38616 );
nand U127410 ( n2661, n38614, n38615 );
nand U127411 ( n38614, P4_REG1_REG_31_, n38617 );
nand U127412 ( n38615, n76015, n38616 );
nand U127413 ( n19524, n16879, P4_DATAO_REG_3_ );
nand U127414 ( n40806, n62980, n62981 );
nand U127415 ( n62981, n76390, n41908 );
nand U127416 ( n62980, P1_P3_DATAO_REG_19_, n76389 );
nand U127417 ( n18933, n16854, P4_DATAO_REG_6_ );
nor U127418 ( n72805, n73522, n71104 );
xor U127419 ( n45653, n7533, n46476 );
nor U127420 ( n46476, n46477, n46434 );
nor U127421 ( n46477, P2_P1_INSTADDRPOINTER_REG_27_, n76005 );
nand U127422 ( n15666, n46465, n46466 );
nand U127423 ( n46466, n76859, P2_P1_INSTADDRPOINTER_REG_27_ );
nor U127424 ( n46465, n46467, n46468 );
nor U127425 ( n46468, n75014, n76334 );
nand U127426 ( n32724, P1_P3_INSTADDRPOINTER_REG_28_, n32725 );
nand U127427 ( n32725, n32726, n32727 );
nor U127428 ( n32726, n32687, n32734 );
nor U127429 ( n32727, n32728, n32729 );
nand U127430 ( n4446, n32716, n32717 );
nand U127431 ( n32717, n76469, P1_P3_INSTADDRPOINTER_REG_28_ );
nor U127432 ( n32716, n32718, n32719 );
nor U127433 ( n32719, n75362, n76899 );
xor U127434 ( n24742, n3989, n25534 );
nor U127435 ( n25534, n25535, n25493 );
nor U127436 ( n25535, P1_P2_INSTADDRPOINTER_REG_27_, n76026 );
xor U127437 ( n66577, n5747, n67539 );
nor U127438 ( n67539, n67540, n67498 );
nor U127439 ( n67540, P2_P3_INSTADDRPOINTER_REG_27_, n75989 );
xor U127440 ( n57876, n6622, n58671 );
nor U127441 ( n58671, n58672, n58630 );
nor U127442 ( n58672, P2_P2_INSTADDRPOINTER_REG_27_, n75997 );
nand U127443 ( n6686, n25523, n25524 );
nand U127444 ( n25524, n76520, P1_P2_INSTADDRPOINTER_REG_27_ );
nor U127445 ( n25523, n25525, n25526 );
nor U127446 ( n25526, n74999, n76908 );
nand U127447 ( n11176, n67528, n67529 );
nand U127448 ( n67529, n76196, P2_P3_INSTADDRPOINTER_REG_27_ );
nor U127449 ( n67528, n67530, n67531 );
nor U127450 ( n67531, n75003, n76873 );
nand U127451 ( n13421, n58660, n58661 );
nand U127452 ( n58661, n76262, P2_P2_INSTADDRPOINTER_REG_27_ );
nor U127453 ( n58660, n58662, n58663 );
nor U127454 ( n58663, n75000, n76882 );
and U127455 ( n52173, n49809, P3_DATAO_REG_2_ );
and U127456 ( n39929, n76419, P4_REG0_REG_11_ );
nand U127457 ( n31132, P1_P3_INSTQUEUERD_ADDR_REG_0_, n34130 );
nor U127458 ( n71282, n73510, n71283 );
and U127459 ( n19398, n16854, P4_DATAO_REG_5_ );
nand U127460 ( n2656, n38622, n38623 );
nand U127461 ( n38622, P4_REG1_REG_30_, n38617 );
nand U127462 ( n38623, n76015, n38624 );
nand U127463 ( n2496, n38739, n38740 );
nand U127464 ( n38739, P4_REG0_REG_30_, n76421 );
nand U127465 ( n38740, n76012, n38624 );
nand U127466 ( n36915, P2_P3_DATAO_REG_20_, n76457 );
nand U127467 ( n51871, n49990, P3_DATAO_REG_4_ );
nand U127468 ( n52330, n49809, P3_DATAO_REG_3_ );
nand U127469 ( n19213, n16879, P4_DATAO_REG_2_ );
nand U127470 ( n18419, n16854, P4_DATAO_REG_9_ );
and U127471 ( n39873, n76419, P4_REG0_REG_12_ );
nand U127472 ( n17757, n16879, P4_DATAO_REG_14_ );
nand U127473 ( n36403, n39431, n39432 );
nand U127474 ( n39432, n76459, n37303 );
nand U127475 ( n39431, P2_P3_DATAO_REG_19_, n76457 );
and U127476 ( n50560, n49809, P3_DATAO_REG_12_ );
and U127477 ( n39828, n76419, P4_REG0_REG_13_ );
nand U127478 ( n39260, P2_P3_DATAO_REG_22_, n76457 );
nand U127479 ( n2566, n38680, n38681 );
nand U127480 ( n38680, P4_REG1_REG_12_, n76425 );
nand U127481 ( n38681, n76016, n38682 );
nand U127482 ( n2406, n39813, n39814 );
nand U127483 ( n39813, P4_REG0_REG_12_, n76422 );
nand U127484 ( n39814, n76013, n38682 );
nor U127485 ( n39827, n76415, n74404 );
nor U127486 ( n46575, P2_P1_INSTADDRPOINTER_REG_25_, n46577 );
xor U127487 ( n46577, n46482, n76006 );
nand U127488 ( n15656, n46556, n46557 );
nand U127489 ( n46557, n76859, P2_P1_INSTADDRPOINTER_REG_25_ );
nor U127490 ( n46556, n46558, n46559 );
nor U127491 ( n46559, n73304, n76334 );
nor U127492 ( n67622, P2_P3_INSTADDRPOINTER_REG_25_, n67624 );
xor U127493 ( n67624, n67545, n75990 );
nor U127494 ( n25617, P1_P2_INSTADDRPOINTER_REG_25_, n25619 );
xor U127495 ( n25619, n25540, n76027 );
nor U127496 ( n58754, P2_P2_INSTADDRPOINTER_REG_25_, n58756 );
xor U127497 ( n58756, n58677, n75998 );
nand U127498 ( n11166, n67603, n67604 );
nand U127499 ( n67604, n76196, P2_P3_INSTADDRPOINTER_REG_25_ );
nor U127500 ( n67603, n67605, n67606 );
nor U127501 ( n67606, n73292, n76873 );
nand U127502 ( n6676, n25598, n25599 );
nand U127503 ( n25599, n76520, P1_P2_INSTADDRPOINTER_REG_25_ );
nor U127504 ( n25598, n25600, n25601 );
nor U127505 ( n25601, n73291, n76908 );
nand U127506 ( n13411, n58735, n58736 );
nand U127507 ( n58736, n76262, P2_P2_INSTADDRPOINTER_REG_25_ );
nor U127508 ( n58735, n58737, n58738 );
nor U127509 ( n58738, n73290, n76882 );
nand U127510 ( n1341, n58780, n58781 );
nand U127511 ( n58780, P3_REG1_REG_12_, n76288 );
nand U127512 ( n58781, n76003, n58782 );
nand U127513 ( n1181, n64774, n64775 );
nand U127514 ( n64774, P3_REG0_REG_12_, n76255 );
nand U127515 ( n64775, n75995, n58782 );
and U127516 ( n65325, n76253, P3_REG0_REG_12_ );
nand U127517 ( n51803, n49809, P3_DATAO_REG_1_ );
and U127518 ( n44066, n45438, n45439 );
nand U127519 ( n45438, P2_BUF1_REG_9_, n76477 );
nand U127520 ( n45439, n45440, n31928 );
xor U127521 ( n45440, n45441, n45442 );
nand U127522 ( n15956, n45364, n45365 );
nand U127523 ( n45365, P2_P1_UWORD_REG_9_, n76352 );
nor U127524 ( n45364, n45366, n45367 );
nor U127525 ( n45367, n75061, n76350 );
nand U127526 ( n15881, n45435, n45436 );
nand U127527 ( n45436, P2_P1_LWORD_REG_9_, n76352 );
nor U127528 ( n45435, n45366, n45437 );
nor U127529 ( n45437, n74757, n76349 );
nand U127530 ( n15661, n46503, n46504 );
nand U127531 ( n46504, n76859, P2_P1_INSTADDRPOINTER_REG_26_ );
nor U127532 ( n46503, n46505, n46506 );
nor U127533 ( n46506, n73308, n76334 );
nand U127534 ( n11171, n67564, n67565 );
nand U127535 ( n67565, n76196, P2_P3_INSTADDRPOINTER_REG_26_ );
nor U127536 ( n67564, n67566, n67567 );
nor U127537 ( n67567, n73296, n76873 );
nand U127538 ( n6681, n25559, n25560 );
nand U127539 ( n25560, n76520, P1_P2_INSTADDRPOINTER_REG_26_ );
nor U127540 ( n25559, n25561, n25562 );
nor U127541 ( n25562, n73294, n76908 );
nand U127542 ( n13416, n58696, n58697 );
nand U127543 ( n58697, n76262, P2_P2_INSTADDRPOINTER_REG_26_ );
nor U127544 ( n58696, n58698, n58699 );
nor U127545 ( n58699, n73295, n76882 );
nor U127546 ( n39771, n76415, n74414 );
nand U127547 ( n51189, n49990, P3_DATAO_REG_8_ );
nor U127548 ( n46525, n46527, n46528 );
and U127549 ( n46527, n46529, P2_P1_INSTADDRPOINTER_REG_26_ );
nor U127550 ( n46528, n46521, n46482 );
nor U127551 ( n67586, n67588, n67589 );
and U127552 ( n67588, n67590, P2_P3_INSTADDRPOINTER_REG_26_ );
nor U127553 ( n67589, n67582, n67545 );
nor U127554 ( n25581, n25583, n25584 );
and U127555 ( n25583, n25585, P1_P2_INSTADDRPOINTER_REG_26_ );
nor U127556 ( n25584, n25577, n25540 );
nor U127557 ( n58718, n58720, n58721 );
and U127558 ( n58720, n58722, P2_P2_INSTADDRPOINTER_REG_26_ );
nor U127559 ( n58721, n58714, n58677 );
nor U127560 ( n46520, n46523, n46524 );
xor U127561 ( n46524, n76342, P2_P1_INSTADDRPOINTER_REG_26_ );
and U127562 ( n46523, n46482, P2_P1_INSTADDRPOINTER_REG_25_ );
nor U127563 ( n67581, n67584, n67585 );
xor U127564 ( n67585, n76198, P2_P3_INSTADDRPOINTER_REG_26_ );
and U127565 ( n67584, n67545, P2_P3_INSTADDRPOINTER_REG_25_ );
nor U127566 ( n25576, n25579, n25580 );
xor U127567 ( n25580, n76522, P1_P2_INSTADDRPOINTER_REG_26_ );
and U127568 ( n25579, n25540, P1_P2_INSTADDRPOINTER_REG_25_ );
nor U127569 ( n58713, n58716, n58717 );
xor U127570 ( n58717, n76264, P2_P2_INSTADDRPOINTER_REG_26_ );
and U127571 ( n58716, n58677, P2_P2_INSTADDRPOINTER_REG_25_ );
nor U127572 ( n39701, n76415, n74422 );
nand U127573 ( n46968, n76006, n47052 );
nand U127574 ( n47052, P2_P1_INSTADDRPOINTER_REG_12_, P2_P1_INSTADDRPOINTER_REG_13_ );
and U127575 ( n64791, n76253, P3_REG0_REG_13_ );
nand U127576 ( n36907, P2_P3_DATAO_REG_21_, n76457 );
and U127577 ( n64351, n76253, P3_REG0_REG_15_ );
nand U127578 ( n1331, n59659, n59660 );
nand U127579 ( n59659, P3_REG1_REG_10_, n55262 );
nand U127580 ( n59660, n76003, n59661 );
nand U127581 ( n1171, n65793, n65794 );
nand U127582 ( n65793, P3_REG0_REG_10_, n61177 );
nand U127583 ( n65794, n75995, n59661 );
nand U127584 ( n2561, n38683, n38684 );
nand U127585 ( n38683, P4_REG1_REG_11_, n38617 );
nand U127586 ( n38684, n76016, n38685 );
nand U127587 ( n2401, n39858, n39859 );
nand U127588 ( n39858, P4_REG0_REG_11_, n76421 );
nand U127589 ( n39859, n76013, n38685 );
nand U127590 ( n50959, n49990, P3_DATAO_REG_9_ );
nand U127591 ( n26000, n76027, n26080 );
nand U127592 ( n26080, P1_P2_INSTADDRPOINTER_REG_12_, P1_P2_INSTADDRPOINTER_REG_13_ );
nand U127593 ( n59138, n75998, n59221 );
nand U127594 ( n59221, P2_P2_INSTADDRPOINTER_REG_12_, P2_P2_INSTADDRPOINTER_REG_13_ );
nand U127595 ( n68003, n75990, n68083 );
nand U127596 ( n68083, P2_P3_INSTADDRPOINTER_REG_12_, P2_P3_INSTADDRPOINTER_REG_13_ );
xor U127597 ( n31907, n32694, n32672 );
xor U127598 ( n32694, n76471, P1_P3_INSTADDRPOINTER_REG_29_ );
nand U127599 ( n4451, n32673, n32674 );
nand U127600 ( n32674, n76469, P1_P3_INSTADDRPOINTER_REG_29_ );
nor U127601 ( n32673, n32675, n32676 );
nor U127602 ( n32676, n73318, n76899 );
and U127603 ( n45503, n49834, P3_DATAO_REG_0_ );
nand U127604 ( n2556, n38690, n38691 );
nand U127605 ( n38690, P4_REG1_REG_10_, n38617 );
nand U127606 ( n38691, n76016, n38692 );
nand U127607 ( n2396, n39914, n39915 );
nand U127608 ( n39914, P4_REG0_REG_10_, n76421 );
nand U127609 ( n39915, n76013, n38692 );
nor U127610 ( n47516, P2_P1_INSTADDRPOINTER_REG_3_, n47517 );
nand U127611 ( n47285, n47326, n47327 );
or U127612 ( n47326, n47330, n47329 );
nand U127613 ( n47327, P2_P1_INSTADDRPOINTER_REG_5_, n47328 );
nand U127614 ( n47328, n47329, n47330 );
nand U127615 ( n47436, n47510, n47511 );
nand U127616 ( n47510, n47517, P2_P1_INSTADDRPOINTER_REG_3_ );
nand U127617 ( n47511, n47512, n47513 );
nand U127618 ( n47513, n7623, n47514 );
nand U127619 ( n1336, n59152, n59153 );
nand U127620 ( n59152, P3_REG1_REG_11_, n55262 );
nand U127621 ( n59153, n76003, n59154 );
nand U127622 ( n1176, n65307, n65308 );
nand U127623 ( n65307, P3_REG0_REG_11_, n61177 );
nand U127624 ( n65308, n75995, n59154 );
and U127625 ( n39642, n76419, P4_REG0_REG_16_ );
and U127626 ( n39772, n76419, P4_REG0_REG_14_ );
nand U127627 ( n33296, n76472, n33372 );
nand U127628 ( n33372, n33373, n73115 );
nor U127629 ( n33373, P1_P3_INSTADDRPOINTER_REG_9_, P1_P3_INSTADDRPOINTER_REG_11_ );
and U127630 ( n39702, n76419, P4_REG0_REG_15_ );
nor U127631 ( n26536, P1_P2_INSTADDRPOINTER_REG_3_, n26537 );
nor U127632 ( n59678, P2_P2_INSTADDRPOINTER_REG_3_, n59679 );
nand U127633 ( n26315, n26357, n26358 );
or U127634 ( n26357, n26361, n26360 );
nand U127635 ( n26358, P1_P2_INSTADDRPOINTER_REG_5_, n26359 );
nand U127636 ( n26359, n26360, n26361 );
nand U127637 ( n59454, n59496, n59497 );
or U127638 ( n59496, n59500, n59499 );
nand U127639 ( n59497, P2_P2_INSTADDRPOINTER_REG_5_, n59498 );
nand U127640 ( n59498, n59499, n59500 );
nand U127641 ( n26456, n26530, n26531 );
nand U127642 ( n26530, n26537, P1_P2_INSTADDRPOINTER_REG_3_ );
nand U127643 ( n26531, n26532, n26533 );
nand U127644 ( n26533, n4064, n26534 );
nand U127645 ( n59595, n59672, n59673 );
nand U127646 ( n59672, n59679, P2_P2_INSTADDRPOINTER_REG_3_ );
nand U127647 ( n59673, n59674, n59675 );
nand U127648 ( n59675, n6697, n59676 );
nor U127649 ( n68537, P2_P3_INSTADDRPOINTER_REG_3_, n68538 );
nand U127650 ( n68316, n68358, n68359 );
or U127651 ( n68358, n68362, n68361 );
nand U127652 ( n68359, P2_P3_INSTADDRPOINTER_REG_5_, n68360 );
nand U127653 ( n68360, n68361, n68362 );
nand U127654 ( n68457, n68531, n68532 );
nand U127655 ( n68531, n68538, P2_P3_INSTADDRPOINTER_REG_3_ );
nand U127656 ( n68532, n68533, n68534 );
nand U127657 ( n68534, n5835, n68535 );
and U127658 ( n17875, n16879, P4_DATAO_REG_13_ );
nor U127659 ( n72817, n73530, n71104 );
and U127660 ( n18844, n16879, P4_DATAO_REG_1_ );
and U127661 ( n64201, n76253, P3_REG0_REG_16_ );
nand U127662 ( n17199, n16854, P4_DATAO_REG_14_ );
nand U127663 ( n18250, n16854, P4_DATAO_REG_10_ );
nand U127664 ( n1326, n60120, n60121 );
nand U127665 ( n60120, P3_REG1_REG_9_, n55262 );
nand U127666 ( n60121, n76003, n60122 );
nand U127667 ( n1166, n65916, n65917 );
nand U127668 ( n65916, P3_REG0_REG_9_, n61177 );
nand U127669 ( n65917, n75995, n60122 );
nor U127670 ( n48776, n48777, n48778 );
and U127671 ( n48777, n48718, P2_P1_INSTQUEUE_REG_7__7_ );
nor U127672 ( n48778, n48139, n48769 );
nand U127673 ( n45424, n53886, n53887 );
nand U127674 ( n53886, P2_BUF1_REG_7_, n76477 );
nand U127675 ( n53887, n53888, n31928 );
xor U127676 ( n53888, n51762, n53889 );
nor U127677 ( n49160, n49161, n49162 );
and U127678 ( n49161, n49085, P2_P1_INSTQUEUE_REG_11__7_ );
nor U127679 ( n49162, n48139, n49152 );
nor U127680 ( n48306, n48307, n48308 );
and U127681 ( n48307, n48247, P2_P1_INSTQUEUE_REG_2__7_ );
nor U127682 ( n48308, n48139, n48249 );
nor U127683 ( n48223, n48224, n48225 );
and U127684 ( n48224, n48149, P2_P1_INSTQUEUE_REG_1__7_ );
nor U127685 ( n48225, n48139, n48151 );
nor U127686 ( n48403, n48404, n48405 );
and U127687 ( n48404, n48344, P2_P1_INSTQUEUE_REG_3__7_ );
nor U127688 ( n48405, n48139, n48346 );
nand U127689 ( n10763, P1_P1_INSTQUEUERD_ADDR_REG_2_, n73525 );
nand U127690 ( n13039, n13374, n13375 );
nand U127691 ( n13375, P1_P1_INSTADDRPOINTER_REG_17_, n76035 );
nor U127692 ( n13374, n12224, n13377 );
nor U127693 ( n13377, n4892, n13350 );
nor U127694 ( n13420, n12220, P1_P1_INSTADDRPOINTER_REG_16_ );
nand U127695 ( n12220, n13468, n13469 );
nand U127696 ( n13468, n13472, n76606 );
nand U127697 ( n13469, P1_P1_INSTADDRPOINTER_REG_15_, n13470 );
or U127698 ( n13470, n13472, n76035 );
nor U127699 ( n12710, n12809, P1_P1_INSTADDRPOINTER_REG_28_ );
nand U127700 ( n13525, n13717, n13718 );
nand U127701 ( n13718, P1_P1_INSTADDRPOINTER_REG_10_, n13719 );
nand U127702 ( n13719, n76602, n13720 );
nand U127703 ( n13720, n13762, P1_P1_INSTADDRPOINTER_REG_8_ );
nor U127704 ( n13762, n13763, n73109 );
nand U127705 ( n11879, n12925, n12927 );
nand U127706 ( n12927, P1_P1_INSTADDRPOINTER_REG_26_, n12928 );
nand U127707 ( n12928, n76603, n12929 );
nand U127708 ( n12929, P1_P1_INSTADDRPOINTER_REG_25_, n12930 );
and U127709 ( n13763, n13849, n13850 );
nand U127710 ( n13849, n13853, n76606 );
nand U127711 ( n13850, P1_P1_INSTADDRPOINTER_REG_7_, n13852 );
or U127712 ( n13852, n13853, n76035 );
nand U127713 ( n12719, n12805, n12807 );
nand U127714 ( n12807, n12808, P1_P1_INSTADDRPOINTER_REG_28_ );
or U127715 ( n12805, n12710, n76603 );
nor U127716 ( n12712, n12714, n12715 );
nor U127717 ( n12714, n12717, n76034 );
nor U127718 ( n12715, P1_P1_INSTADDRPOINTER_REG_30_, n12705 );
nor U127719 ( n12717, n75051, n12718 );
and U127720 ( n11779, n12698, n12699 );
nand U127721 ( n12699, n12700, n12702 );
nand U127722 ( n12698, n12712, n12713 );
nand U127723 ( n12702, n76603, P1_P1_INSTADDRPOINTER_REG_31_ );
nand U127724 ( n8951, n12682, n12683 );
nand U127725 ( n12683, n76886, P1_P1_INSTADDRPOINTER_REG_31_ );
nor U127726 ( n12682, n12684, n12685 );
nor U127727 ( n12685, n75329, n76600 );
nand U127728 ( n12705, n12784, n12785 );
nand U127729 ( n12784, n12719, n76606 );
nand U127730 ( n12785, P1_P1_INSTADDRPOINTER_REG_29_, n12787 );
or U127731 ( n12787, n12719, n76035 );
nand U127732 ( n19699, n16854, P4_DATAO_REG_4_ );
nand U127733 ( n47729, P2_P1_INSTADDRPOINTER_REG_0_, n47682 );
nand U127734 ( n47650, n47726, n47727 );
or U127735 ( n47726, n47729, n44985 );
nand U127736 ( n47727, P2_P1_INSTADDRPOINTER_REG_1_, n47728 );
nand U127737 ( n47728, n47729, n44985 );
and U127738 ( n10178, n11657, n11658 );
nand U127739 ( n11657, P1_BUF1_REG_9_, n76610 );
nand U127740 ( n11658, n11659, n76612 );
xor U127741 ( n11659, n11660, n11662 );
nand U127742 ( n9221, n11554, n11555 );
nand U127743 ( n11555, P1_P1_UWORD_REG_9_, n76618 );
nor U127744 ( n11554, n11557, n11558 );
nor U127745 ( n11558, n75062, n76616 );
nand U127746 ( n9146, n11653, n11654 );
nand U127747 ( n11654, P1_P1_LWORD_REG_9_, n76618 );
nor U127748 ( n11653, n11557, n11655 );
nor U127749 ( n11655, n74756, n76615 );
and U127750 ( n50427, n49990, P3_DATAO_REG_10_ );
nand U127751 ( n49833, n49834, P3_DATAO_REG_17_ );
nand U127752 ( n50121, n49990, P3_DATAO_REG_12_ );
and U127753 ( n64500, n76253, P3_REG0_REG_14_ );
nand U127754 ( n16894, P4_DATAO_REG_21_, n8215 );
nand U127755 ( n2391, n39957, n39958 );
nand U127756 ( n39957, P4_REG0_REG_9_, n76421 );
nand U127757 ( n39958, n76013, n38695 );
nand U127758 ( n2551, n38693, n38694 );
nand U127759 ( n38693, P4_REG1_REG_9_, n38617 );
nand U127760 ( n38694, n76016, n38695 );
nor U127761 ( n12862, n12865, n12867 );
nor U127762 ( n12867, n12868, n74946 );
nor U127763 ( n12865, P1_P1_INSTADDRPOINTER_REG_28_, n12882 );
nor U127764 ( n12868, n12869, n12870 );
and U127765 ( n11870, n12888, n12889 );
nand U127766 ( n12889, n76603, P1_P1_INSTADDRPOINTER_REG_28_ );
nor U127767 ( n12888, n12890, n12808 );
nor U127768 ( n12890, n76602, n12892 );
nand U127769 ( n8936, n12842, n12843 );
nand U127770 ( n12843, n76886, P1_P1_INSTADDRPOINTER_REG_28_ );
nor U127771 ( n12842, n12844, n12845 );
nor U127772 ( n12845, n75303, n76600 );
nand U127773 ( n26749, P1_P2_INSTADDRPOINTER_REG_0_, n26702 );
nand U127774 ( n59891, P2_P2_INSTADDRPOINTER_REG_0_, n59844 );
nand U127775 ( n68750, P2_P3_INSTADDRPOINTER_REG_0_, n68703 );
nand U127776 ( n68671, n68747, n68748 );
or U127777 ( n68747, n68750, n65893 );
nand U127778 ( n68748, P2_P3_INSTADDRPOINTER_REG_1_, n68749 );
nand U127779 ( n68749, n68750, n65893 );
nand U127780 ( n26670, n26746, n26747 );
or U127781 ( n26746, n26749, n24311 );
nand U127782 ( n26747, P1_P2_INSTADDRPOINTER_REG_1_, n26748 );
nand U127783 ( n26748, n26749, n24311 );
nand U127784 ( n59812, n59888, n59889 );
or U127785 ( n59888, n59891, n57434 );
nand U127786 ( n59889, P2_P2_INSTADDRPOINTER_REG_1_, n59890 );
nand U127787 ( n59890, n59891, n57434 );
nor U127788 ( n47515, n47690, P2_P1_INSTADDRPOINTER_REG_2_ );
nor U127789 ( n12700, n12703, n12704 );
nor U127790 ( n12703, n76602, n12707 );
and U127791 ( n12704, n12705, P1_P1_INSTADDRPOINTER_REG_30_ );
nor U127792 ( n12707, n12708, n12709 );
nand U127793 ( n33302, n76022, n33326 );
nand U127794 ( n33326, P1_P3_INSTADDRPOINTER_REG_12_, P1_P3_INSTADDRPOINTER_REG_13_ );
nand U127795 ( n71098, n72846, n72847 );
nand U127796 ( n72846, P4_WR_REG, P4_ADDR_REG_0_ );
nand U127797 ( n72847, n71018, n73025 );
nor U127798 ( n72851, n73513, n71013 );
nand U127799 ( n71018, n72848, n72849 );
nand U127800 ( n72849, n1244, P1_P1_ADDRESS_REG_0_ );
nor U127801 ( n72848, n72850, n72851 );
nor U127802 ( n72850, n73514, n71009 );
nand U127803 ( n47514, P2_P1_INSTADDRPOINTER_REG_2_, n47690 );
nand U127804 ( n52349, n49990, P3_DATAO_REG_3_ );
nor U127805 ( n68536, n68711, P2_P3_INSTADDRPOINTER_REG_2_ );
nor U127806 ( n26535, n26710, P1_P2_INSTADDRPOINTER_REG_2_ );
nor U127807 ( n59677, n59852, P2_P2_INSTADDRPOINTER_REG_2_ );
nand U127808 ( n11184, P1_P1_INSTQUEUERD_ADDR_REG_1_, P1_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U127809 ( n31931, n31941, n31942 );
nand U127810 ( n31941, n31952, P1_P3_PHYADDRPOINTER_REG_27_ );
nand U127811 ( n31942, n31943, n31944 );
and U127812 ( n31952, n75246, n31953 );
and U127813 ( n44113, n45428, n45429 );
nand U127814 ( n45428, P2_BUF1_REG_8_, n76478 );
nand U127815 ( n45429, n45430, n31928 );
xor U127816 ( n45430, n45431, n45432 );
nand U127817 ( n15886, n45425, n45426 );
nand U127818 ( n45426, P2_P1_LWORD_REG_8_, n76352 );
nor U127819 ( n45425, n45359, n45427 );
nor U127820 ( n45427, n73218, n76349 );
nand U127821 ( n15961, n45357, n45358 );
nand U127822 ( n45358, P2_P1_UWORD_REG_8_, n76352 );
nor U127823 ( n45357, n45359, n45360 );
nor U127824 ( n45360, n73306, n76350 );
nand U127825 ( n68535, P2_P3_INSTADDRPOINTER_REG_2_, n68711 );
nand U127826 ( n26534, P1_P2_INSTADDRPOINTER_REG_2_, n26710 );
nand U127827 ( n59676, P2_P2_INSTADDRPOINTER_REG_2_, n59852 );
and U127828 ( n17036, DIN_18_, n76927 );
nand U127829 ( n18558, n17036, P4_DATAO_REG_6_ );
nand U127830 ( n16206, n44862, n44863 );
nor U127831 ( n44863, n44864, n44865 );
nor U127832 ( n44862, n44869, n44870 );
nor U127833 ( n44864, P2_P1_EAX_REG_8_, n44814 );
nor U127834 ( n10260, n11184, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
or U127835 ( n47433, n75934, n47483 );
and U127836 ( n12750, n75935, n75936 );
nand U127837 ( n75935, n11805, n76724 );
nand U127838 ( n75936, n12729, P1_P1_INSTADDRPOINTER_REG_30_ );
nand U127839 ( n8946, n12737, n12738 );
nand U127840 ( n12738, n76886, P1_P1_INSTADDRPOINTER_REG_30_ );
nor U127841 ( n12737, n12739, n12740 );
nor U127842 ( n12740, n75238, n76600 );
and U127843 ( n50117, n49990, P3_DATAO_REG_11_ );
nand U127844 ( n39085, P2_P3_DATAO_REG_23_, n76457 );
nand U127845 ( n1591, n45361, n45405 );
nand U127846 ( n45405, P3_REG2_REG_30_, n45363 );
nand U127847 ( n1596, n45361, n45362 );
nand U127848 ( n45362, P3_REG2_REG_31_, n45363 );
or U127849 ( n68454, n75937, n68504 );
or U127850 ( n26453, n75938, n26503 );
or U127851 ( n59592, n75939, n59642 );
nand U127852 ( n13717, n13764, n76606 );
nand U127853 ( n13764, n13765, n13763 );
nor U127854 ( n13765, P1_P1_INSTADDRPOINTER_REG_9_, P1_P1_INSTADDRPOINTER_REG_8_ );
and U127855 ( n17745, n16854, P4_DATAO_REG_11_ );
nand U127856 ( n18919, n17036, P4_DATAO_REG_5_ );
xor U127857 ( n31974, n3150, n32774 );
nor U127858 ( n32774, n32775, n32733 );
nor U127859 ( n32775, P1_P3_INSTADDRPOINTER_REG_27_, n76021 );
nand U127860 ( n4441, n32763, n32764 );
nand U127861 ( n32764, n76469, P1_P3_INSTADDRPOINTER_REG_27_ );
nor U127862 ( n32763, n32765, n32766 );
nor U127863 ( n32766, n75004, n76899 );
nand U127864 ( n2386, n39991, n39992 );
nand U127865 ( n39991, P4_REG0_REG_8_, n76421 );
nand U127866 ( n39992, n76013, n38698 );
nand U127867 ( n2546, n38696, n38697 );
nand U127868 ( n38696, P4_REG1_REG_8_, n38617 );
nand U127869 ( n38697, n76016, n38698 );
nand U127870 ( n15631, n46750, n46751 );
nand U127871 ( n46751, n76859, P2_P1_INSTADDRPOINTER_REG_20_ );
nor U127872 ( n46750, n46752, n46753 );
nor U127873 ( n46753, n74951, n76333 );
nand U127874 ( n11141, n67797, n67798 );
nand U127875 ( n67798, n76196, P2_P3_INSTADDRPOINTER_REG_20_ );
nor U127876 ( n67797, n67799, n67800 );
nor U127877 ( n67800, n74928, n76872 );
nand U127878 ( n6651, n25794, n25795 );
nand U127879 ( n25795, n76520, P1_P2_INSTADDRPOINTER_REG_20_ );
nor U127880 ( n25794, n25796, n25797 );
nor U127881 ( n25797, n74926, n76907 );
nand U127882 ( n13386, n58932, n58933 );
nand U127883 ( n58933, n76262, P2_P2_INSTADDRPOINTER_REG_20_ );
nor U127884 ( n58932, n58934, n58935 );
nor U127885 ( n58935, n74925, n76881 );
nand U127886 ( n47282, P2_P1_INSTADDRPOINTER_REG_6_, n7562 );
nand U127887 ( n17478, n16854, P4_DATAO_REG_13_ );
nand U127888 ( n10717, P1_P1_INSTQUEUERD_ADDR_REG_0_, n14629 );
nand U127889 ( n18406, n17036, P4_DATAO_REG_7_ );
and U127890 ( n52189, n49990, P3_DATAO_REG_2_ );
nand U127891 ( n68313, P2_P3_INSTADDRPOINTER_REG_6_, n5774 );
nand U127892 ( n26312, P1_P2_INSTADDRPOINTER_REG_6_, n4015 );
nand U127893 ( n59451, P2_P2_INSTADDRPOINTER_REG_6_, n6648 );
nor U127894 ( n15260, n15262, n15263 );
and U127895 ( n15262, n15178, P1_P1_INSTQUEUE_REG_3__7_ );
nor U127896 ( n15263, n14954, n15180 );
nor U127897 ( n15150, n15152, n15153 );
and U127898 ( n15152, n15070, P1_P1_INSTQUEUE_REG_2__7_ );
nor U127899 ( n15153, n14954, n15073 );
nor U127900 ( n15040, n15042, n15043 );
and U127901 ( n15042, n14967, P1_P1_INSTQUEUE_REG_1__7_ );
nor U127902 ( n15043, n14954, n14969 );
nand U127903 ( n11638, n20930, n20931 );
nand U127904 ( n20930, P1_BUF1_REG_7_, n76611 );
nand U127905 ( n20931, n20932, n76612 );
xor U127906 ( n20932, n18806, n20933 );
nand U127907 ( n15651, n46601, n46602 );
nand U127908 ( n46602, n76859, P2_P1_INSTADDRPOINTER_REG_24_ );
nor U127909 ( n46601, n46603, n46604 );
nor U127910 ( n46604, n75005, n76334 );
nand U127911 ( n10722, n5154, P1_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U127912 ( n11161, n67648, n67649 );
nand U127913 ( n67649, n76196, P2_P3_INSTADDRPOINTER_REG_24_ );
nor U127914 ( n67648, n67650, n67651 );
nor U127915 ( n67651, n74993, n76873 );
nand U127916 ( n6671, n25643, n25644 );
nand U127917 ( n25644, n76520, P1_P2_INSTADDRPOINTER_REG_24_ );
nor U127918 ( n25643, n25645, n25646 );
nor U127919 ( n25646, n74991, n76908 );
nand U127920 ( n13406, n58783, n58784 );
nand U127921 ( n58784, n76262, P2_P2_INSTADDRPOINTER_REG_24_ );
nor U127922 ( n58783, n58785, n58786 );
nor U127923 ( n58786, n74990, n76882 );
and U127924 ( n63992, n76253, P3_REG0_REG_17_ );
nand U127925 ( n18915, n17036, P4_DATAO_REG_4_ );
nand U127926 ( n13589, n76603, n13620 );
nand U127927 ( n13620, P1_P1_INSTADDRPOINTER_REG_12_, P1_P1_INSTADDRPOINTER_REG_13_ );
and U127928 ( n39580, n76419, P4_REG0_REG_17_ );
nand U127929 ( n2541, n38699, n38700 );
nand U127930 ( n38699, P4_REG1_REG_7_, n38617 );
nand U127931 ( n38700, n76017, n38701 );
nand U127932 ( n2381, n40037, n40038 );
nand U127933 ( n40037, P4_REG0_REG_7_, n76421 );
nand U127934 ( n40038, n76014, n38701 );
nand U127935 ( n12709, n12710, P1_P1_INSTADDRPOINTER_REG_31_ );
xnor U127936 ( n45815, n46728, n46729 );
xor U127937 ( n46728, n76342, P2_P1_INSTADDRPOINTER_REG_21_ );
nor U127938 ( n46729, n46730, n46731 );
nor U127939 ( n46730, n7535, n46734 );
nand U127940 ( n15636, n46712, n46713 );
nand U127941 ( n46713, n76859, P2_P1_INSTADDRPOINTER_REG_21_ );
nor U127942 ( n46712, n46714, n46715 );
nor U127943 ( n46715, n74958, n76333 );
xnor U127944 ( n66766, n67775, n67776 );
xor U127945 ( n67775, n76198, P2_P3_INSTADDRPOINTER_REG_21_ );
nor U127946 ( n67776, n67777, n67778 );
nor U127947 ( n67777, n5749, n67781 );
xnor U127948 ( n24888, n25772, n25773 );
xor U127949 ( n25772, n76522, P1_P2_INSTADDRPOINTER_REG_21_ );
nor U127950 ( n25773, n25774, n25775 );
nor U127951 ( n25774, n3992, n25778 );
xnor U127952 ( n58025, n58910, n58911 );
xor U127953 ( n58910, n76264, P2_P2_INSTADDRPOINTER_REG_21_ );
nor U127954 ( n58911, n58912, n58913 );
nor U127955 ( n58912, n6624, n58916 );
nand U127956 ( n11146, n67759, n67760 );
nand U127957 ( n67760, n76196, P2_P3_INSTADDRPOINTER_REG_21_ );
nor U127958 ( n67759, n67761, n67762 );
nor U127959 ( n67762, n74944, n76872 );
nand U127960 ( n6656, n25756, n25757 );
nand U127961 ( n25757, n76520, P1_P2_INSTADDRPOINTER_REG_21_ );
nor U127962 ( n25756, n25758, n25759 );
nor U127963 ( n25759, n74939, n76907 );
nand U127964 ( n13391, n58894, n58895 );
nand U127965 ( n58895, n76262, P2_P2_INSTADDRPOINTER_REG_21_ );
nor U127966 ( n58894, n58896, n58897 );
nor U127967 ( n58897, n74938, n76881 );
nand U127968 ( n1431, n55521, n55522 );
nand U127969 ( n55521, P3_REG1_REG_30_, n55262 );
nand U127970 ( n55522, n76002, n55523 );
nand U127971 ( n1271, n61284, n61285 );
nand U127972 ( n61284, P3_REG0_REG_30_, n76255 );
nand U127973 ( n61285, n75994, n55523 );
and U127974 ( n11700, n76168, P4_DATAO_REG_0_ );
nor U127975 ( n32857, P1_P3_INSTADDRPOINTER_REG_25_, n32859 );
xor U127976 ( n32859, n32780, n76022 );
nand U127977 ( n4431, n32838, n32839 );
nand U127978 ( n32839, n76469, P1_P3_INSTADDRPOINTER_REG_25_ );
nor U127979 ( n32838, n32840, n32841 );
nor U127980 ( n32841, n73293, n76899 );
and U127981 ( n19217, n16854, P4_DATAO_REG_2_ );
nor U127982 ( n15688, n15689, n15690 );
and U127983 ( n15689, n15609, P1_P1_INSTQUEUE_REG_7__7_ );
nor U127984 ( n15690, n14954, n15678 );
nand U127985 ( n1321, n60230, n60231 );
nand U127986 ( n60230, P3_REG1_REG_8_, n55262 );
nand U127987 ( n60231, n76003, n60232 );
nand U127988 ( n1161, n65994, n65995 );
nand U127989 ( n65994, P3_REG0_REG_8_, n61177 );
nand U127990 ( n65995, n75995, n60232 );
nand U127991 ( n1276, n61168, n61169 );
nand U127992 ( n61168, P3_REG0_REG_31_, n61177 );
nand U127993 ( n61169, n75994, n55261 );
nand U127994 ( n1436, n55259, n55260 );
nand U127995 ( n55259, P3_REG1_REG_31_, n76288 );
nand U127996 ( n55260, n76002, n55261 );
nand U127997 ( n4436, n32799, n32800 );
nand U127998 ( n32800, n76469, P1_P3_INSTADDRPOINTER_REG_26_ );
nor U127999 ( n32799, n32801, n32802 );
nor U128000 ( n32802, n73297, n76899 );
nor U128001 ( n72823, n73544, n71104 );
xnor U128002 ( n32120, n33019, n33020 );
xor U128003 ( n33019, n76471, P1_P3_INSTADDRPOINTER_REG_21_ );
nor U128004 ( n33020, n3147, n33021 );
nand U128005 ( n33021, n33022, n33023 );
nand U128006 ( n4411, n33003, n33004 );
nand U128007 ( n33004, n76469, P1_P3_INSTADDRPOINTER_REG_21_ );
nor U128008 ( n33003, n33005, n33006 );
nor U128009 ( n33006, n74945, n76898 );
nand U128010 ( n36848, P2_P3_DATAO_REG_24_, n76457 );
nand U128011 ( n49457, n49809, P3_DATAO_REG_0_ );
nand U128012 ( n19538, n16854, P4_DATAO_REG_3_ );
nor U128013 ( n32821, n32823, n32824 );
and U128014 ( n32823, n32825, P1_P3_INSTADDRPOINTER_REG_26_ );
nor U128015 ( n32824, n32817, n32780 );
and U128016 ( n10237, n11643, n11644 );
nand U128017 ( n11643, P1_BUF1_REG_8_, n76610 );
nand U128018 ( n11644, n11645, n76613 );
xor U128019 ( n11645, n11648, n11649 );
nand U128020 ( n9151, n11639, n11640 );
nand U128021 ( n11640, P1_P1_LWORD_REG_8_, n76618 );
nor U128022 ( n11639, n11552, n11642 );
nor U128023 ( n11642, n73219, n76615 );
nand U128024 ( n9226, n11549, n11550 );
nand U128025 ( n11550, P1_P1_UWORD_REG_8_, n76618 );
nor U128026 ( n11549, n11552, n11553 );
nor U128027 ( n11553, n73307, n76616 );
nand U128028 ( n33301, n76475, n33369 );
nand U128029 ( n33369, P1_P3_INSTADDRPOINTER_REG_10_, P1_P3_INSTADDRPOINTER_REG_11_ );
nand U128030 ( n9471, n11144, n11145 );
nor U128031 ( n11145, n11147, n11148 );
nor U128032 ( n11144, n11153, n11154 );
nor U128033 ( n11147, P1_P1_EAX_REG_8_, n11102 );
nor U128034 ( n32816, n32819, n32820 );
xor U128035 ( n32820, n76471, P1_P3_INSTADDRPOINTER_REG_26_ );
and U128036 ( n32819, n32780, P1_P3_INSTADDRPOINTER_REG_25_ );
nand U128037 ( n37706, n40313, n40314 );
nand U128038 ( n40314, P4_IR_REG_31_, n40315 );
nand U128039 ( n40313, P4_IR_REG_1_, n76795 );
and U128040 ( n51820, n49990, P3_DATAO_REG_1_ );
nand U128041 ( n2536, n38702, n38703 );
nand U128042 ( n38702, P4_REG1_REG_6_, n38617 );
nand U128043 ( n38703, n76017, n38704 );
nand U128044 ( n2376, n40079, n40080 );
nand U128045 ( n40079, P4_REG0_REG_6_, n76421 );
nand U128046 ( n40080, n76014, n38704 );
and U128047 ( n17603, n16854, P4_DATAO_REG_12_ );
nand U128048 ( n15891, n45421, n45422 );
nand U128049 ( n45422, P2_P1_LWORD_REG_7_, n76352 );
nor U128050 ( n45421, n45423, n45356 );
nor U128051 ( n45423, n74738, n76349 );
nand U128052 ( n15966, n45353, n45354 );
nand U128053 ( n45354, P2_P1_UWORD_REG_7_, n45325 );
nor U128054 ( n45353, n45355, n45356 );
nor U128055 ( n45355, n75012, n76350 );
nor U128056 ( n33781, P1_P3_INSTADDRPOINTER_REG_3_, n33782 );
nand U128057 ( n33560, n33602, n33603 );
or U128058 ( n33602, n33606, n33605 );
nand U128059 ( n33603, P1_P3_INSTADDRPOINTER_REG_5_, n33604 );
nand U128060 ( n33604, n33605, n33606 );
nand U128061 ( n33701, n33775, n33776 );
nand U128062 ( n33775, n33782, P1_P3_INSTADDRPOINTER_REG_3_ );
nand U128063 ( n33776, n33777, n33778 );
nand U128064 ( n33778, n3236, n33779 );
nand U128065 ( n49808, n49809, P3_DATAO_REG_15_ );
nand U128066 ( n18847, n16854, P4_DATAO_REG_1_ );
nand U128067 ( n1316, n60342, n60343 );
nand U128068 ( n60342, P3_REG1_REG_7_, n55262 );
nand U128069 ( n60343, n76004, n60344 );
nand U128070 ( n1156, n66083, n66084 );
nand U128071 ( n66083, P3_REG0_REG_7_, n61177 );
nand U128072 ( n66084, n75996, n60344 );
nand U128073 ( n32940, n32903, n32944 );
nand U128074 ( n32944, n3149, P1_P3_INSTADDRPOINTER_REG_22_ );
nand U128075 ( n4421, n32918, n32919 );
nand U128076 ( n32919, n76469, P1_P3_INSTADDRPOINTER_REG_23_ );
nor U128077 ( n32918, n32920, n32921 );
nor U128078 ( n32921, n74988, n76898 );
nand U128079 ( n4406, n33043, n33044 );
nand U128080 ( n33044, n76469, P1_P3_INSTADDRPOINTER_REG_20_ );
nor U128081 ( n33043, n33045, n33046 );
nor U128082 ( n33046, n74929, n76898 );
nand U128083 ( n8941, n12788, n12789 );
nand U128084 ( n12789, n76886, P1_P1_INSTADDRPOINTER_REG_29_ );
nor U128085 ( n12788, n12790, n12792 );
nor U128086 ( n12792, n73392, n76600 );
nand U128087 ( n50089, DIN_21_, n76930 );
nand U128088 ( n51172, n8235, P3_DATAO_REG_4_ );
and U128089 ( n63677, n76253, P3_REG0_REG_18_ );
and U128090 ( n39518, n76419, P4_REG0_REG_18_ );
nor U128091 ( n62946, n76249, n74501 );
nand U128092 ( n39021, P2_P3_DATAO_REG_25_, n76457 );
nor U128093 ( n33054, n33057, n33058 );
xor U128094 ( n33058, n76471, P1_P3_INSTADDRPOINTER_REG_20_ );
nor U128095 ( n33057, n33025, n74610 );
nor U128096 ( n63268, n76249, n74498 );
and U128097 ( n63269, n76252, P3_REG0_REG_19_ );
and U128098 ( n62947, n76252, P3_REG0_REG_20_ );
nand U128099 ( n18233, n17036, P4_DATAO_REG_8_ );
nor U128100 ( n39274, n76415, n74530 );
nand U128101 ( n15646, n46632, n46633 );
nand U128102 ( n46633, n76859, P2_P1_INSTADDRPOINTER_REG_23_ );
nor U128103 ( n46632, n46634, n46635 );
nor U128104 ( n46635, n74995, n76333 );
nand U128105 ( n11156, n67679, n67680 );
nand U128106 ( n67680, n76196, P2_P3_INSTADDRPOINTER_REG_23_ );
nor U128107 ( n67679, n67681, n67682 );
nor U128108 ( n67682, n74987, n76872 );
nand U128109 ( n6666, n25674, n25675 );
nand U128110 ( n25675, n76520, P1_P2_INSTADDRPOINTER_REG_23_ );
nor U128111 ( n25674, n25676, n25677 );
nor U128112 ( n25677, n74970, n76907 );
nand U128113 ( n13401, n58814, n58815 );
nand U128114 ( n58815, n76262, P2_P2_INSTADDRPOINTER_REG_23_ );
nor U128115 ( n58814, n58816, n58817 );
nor U128116 ( n58817, n74969, n76881 );
nand U128117 ( n45420, n49641, n49642 );
nand U128118 ( n49641, P2_BUF1_REG_6_, n76478 );
nand U128119 ( n49642, n49643, n76476 );
xor U128120 ( n49643, n49644, n49645 );
nand U128121 ( n48766, n48767, n48768 );
nand U128122 ( n48768, P2_P1_INSTQUEUE_REG_7__6_, n48718 );
nand U128123 ( n48767, n7447, n283 );
nand U128124 ( n49417, n49418, n49419 );
nand U128125 ( n49419, P2_P1_INSTQUEUE_REG_14__6_, n49353 );
nand U128126 ( n49418, n7440, n283 );
nand U128127 ( n49324, n49325, n49326 );
nand U128128 ( n49326, P2_P1_INSTQUEUE_REG_13__6_, n49275 );
nand U128129 ( n49325, n7442, n283 );
nand U128130 ( n49149, n49150, n49151 );
nand U128131 ( n49151, P2_P1_INSTQUEUE_REG_11__6_, n49085 );
nand U128132 ( n49150, n7443, n283 );
nand U128133 ( n49055, n49056, n49057 );
nand U128134 ( n49057, P2_P1_INSTQUEUE_REG_10__6_, n48990 );
nand U128135 ( n49056, n7444, n283 );
nand U128136 ( n48960, n48961, n48962 );
nand U128137 ( n48962, P2_P1_INSTQUEUE_REG_9__6_, n48891 );
nand U128138 ( n48961, n7445, n283 );
nand U128139 ( n48689, n48690, n48691 );
nand U128140 ( n48691, P2_P1_INSTQUEUE_REG_6__6_, n48624 );
nand U128141 ( n48690, n7448, n283 );
nand U128142 ( n48595, n48596, n48597 );
nand U128143 ( n48597, P2_P1_INSTQUEUE_REG_5__6_, n48530 );
nand U128144 ( n48596, n7449, n283 );
nand U128145 ( n50939, n8235, P3_DATAO_REG_5_ );
nand U128146 ( n2531, n38705, n38706 );
nand U128147 ( n38705, P4_REG1_REG_5_, n38617 );
nand U128148 ( n38706, n76017, n38707 );
nand U128149 ( n2371, n40130, n40131 );
nand U128150 ( n40130, P4_REG0_REG_5_, n76421 );
nand U128151 ( n40131, n76014, n38707 );
nand U128152 ( n33994, P1_P3_INSTADDRPOINTER_REG_0_, n33947 );
nand U128153 ( n33915, n33991, n33992 );
or U128154 ( n33991, n33994, n31607 );
nand U128155 ( n33992, P1_P3_INSTADDRPOINTER_REG_1_, n33993 );
nand U128156 ( n33993, n31607, n33994 );
nand U128157 ( n42229, n66756, n66757 );
nand U128158 ( n66757, n66758, P3_IR_REG_31_ );
nand U128159 ( n66756, P3_IR_REG_2_, n76841 );
and U128160 ( n66758, n16703, n16702 );
nor U128161 ( n39450, n76415, n74511 );
nand U128162 ( n45201, n67013, n67014 );
nand U128163 ( n67014, P3_IR_REG_31_, n21629 );
nand U128164 ( n67013, P3_IR_REG_1_, n76841 );
nand U128165 ( n36935, P2_P3_DATAO_REG_26_, n76457 );
nand U128166 ( n15626, n46790, n46791 );
nand U128167 ( n46791, n76860, P2_P1_INSTADDRPOINTER_REG_19_ );
nor U128168 ( n46790, n46792, n46793 );
nor U128169 ( n46793, n73267, n76333 );
nand U128170 ( n11136, n67837, n67838 );
nand U128171 ( n67838, n76196, P2_P3_INSTADDRPOINTER_REG_19_ );
nor U128172 ( n67837, n67839, n67840 );
nor U128173 ( n67840, n73263, n76872 );
nand U128174 ( n6646, n25834, n25835 );
nand U128175 ( n25835, n76520, P1_P2_INSTADDRPOINTER_REG_19_ );
nor U128176 ( n25834, n25836, n25837 );
nor U128177 ( n25837, n73262, n76907 );
nand U128178 ( n13381, n58972, n58973 );
nand U128179 ( n58973, n76262, P2_P2_INSTADDRPOINTER_REG_19_ );
nor U128180 ( n58972, n58974, n58975 );
nor U128181 ( n58975, n73261, n76881 );
nor U128182 ( n11869, n11870, n11872 );
nor U128183 ( n11872, n4890, n11873 );
nor U128184 ( n11873, n11874, n11875 );
nor U128185 ( n11875, P1_P1_INSTADDRPOINTER_REG_28_, n76602 );
nand U128186 ( n11857, n11867, n11868 );
nand U128187 ( n11867, n11880, P1_P1_PHYADDRPOINTER_REG_27_ );
nand U128188 ( n11868, n11869, n76729 );
and U128189 ( n11880, n74880, n11882 );
nand U128190 ( n18001, n17036, P4_DATAO_REG_9_ );
nor U128191 ( n14185, P1_P1_INSTADDRPOINTER_REG_3_, n14187 );
nand U128192 ( n13912, n13979, n13980 );
or U128193 ( n13979, n13984, n13983 );
nand U128194 ( n13980, P1_P1_INSTADDRPOINTER_REG_5_, n13982 );
nand U128195 ( n13982, n13983, n13984 );
nand U128196 ( n14085, n14178, n14179 );
nand U128197 ( n14178, n14187, P1_P1_INSTADDRPOINTER_REG_3_ );
nand U128198 ( n14179, n14180, n14182 );
nand U128199 ( n14182, n4969, n14183 );
nor U128200 ( n33780, n33955, P1_P3_INSTADDRPOINTER_REG_2_ );
nand U128201 ( n54865, n54866, n54867 );
or U128202 ( n54866, n54868, n573 );
nand U128203 ( n54867, n76335, P3_REG3_REG_2_ );
nand U128204 ( n54992, n54993, n54994 );
nand U128205 ( n54993, n76858, n54995 );
nand U128206 ( n54994, n76335, P3_REG3_REG_0_ );
nand U128207 ( n54910, n54916, n54917 );
nand U128208 ( n54917, n76338, n40784 );
nand U128209 ( n54916, n76335, P3_REG3_REG_1_ );
xnor U128210 ( n45795, n46686, n46687 );
xor U128211 ( n46686, n76342, P2_P1_INSTADDRPOINTER_REG_22_ );
nor U128212 ( n46687, n46688, n46689 );
nand U128213 ( n46688, n46655, n46654 );
nand U128214 ( n15641, n46675, n46676 );
nand U128215 ( n46676, n76859, P2_P1_INSTADDRPOINTER_REG_22_ );
nor U128216 ( n46675, n46677, n46678 );
nor U128217 ( n46678, n73280, n76333 );
xnor U128218 ( n66703, n67733, n67734 );
xor U128219 ( n67733, n76198, P2_P3_INSTADDRPOINTER_REG_22_ );
nor U128220 ( n67734, n67735, n67736 );
nand U128221 ( n67735, n67702, n67701 );
xnor U128222 ( n24868, n25728, n25729 );
xor U128223 ( n25728, n76522, P1_P2_INSTADDRPOINTER_REG_22_ );
nor U128224 ( n25729, n25730, n25731 );
nand U128225 ( n25730, n25697, n25696 );
xnor U128226 ( n58005, n58868, n58869 );
xor U128227 ( n58868, n76264, P2_P2_INSTADDRPOINTER_REG_22_ );
nor U128228 ( n58869, n58870, n58871 );
nand U128229 ( n58870, n58837, n58836 );
nand U128230 ( n11151, n67722, n67723 );
nand U128231 ( n67723, n76196, P2_P3_INSTADDRPOINTER_REG_22_ );
nor U128232 ( n67722, n67724, n67725 );
nor U128233 ( n67725, n73277, n76872 );
nand U128234 ( n6661, n25717, n25718 );
nand U128235 ( n25718, n76520, P1_P2_INSTADDRPOINTER_REG_22_ );
nor U128236 ( n25717, n25719, n25720 );
nor U128237 ( n25720, n73276, n76907 );
nand U128238 ( n13396, n58857, n58858 );
nand U128239 ( n58858, n76262, P2_P2_INSTADDRPOINTER_REG_22_ );
nor U128240 ( n58857, n58859, n58860 );
nor U128241 ( n58860, n73275, n76881 );
nand U128242 ( n37354, P2_P3_DATAO_REG_31_, n76457 );
nand U128243 ( n1306, n60562, n60563 );
nand U128244 ( n60562, P3_REG1_REG_5_, n55262 );
nand U128245 ( n60563, n76004, n60564 );
nand U128246 ( n1146, n66266, n66267 );
nand U128247 ( n66266, P3_REG0_REG_5_, n61177 );
nand U128248 ( n66267, n75996, n60564 );
nand U128249 ( n33779, P1_P3_INSTADDRPOINTER_REG_2_, n33955 );
nor U128250 ( n62872, n76249, n74521 );
nand U128251 ( n42251, n66445, n66446 );
nand U128252 ( n66445, P3_IR_REG_3_, n76841 );
or U128253 ( n66446, n16393, n76839 );
nand U128254 ( n36425, P2_P3_DATAO_REG_28_, n76457 );
nor U128255 ( n39392, n76415, n74519 );
nand U128256 ( n4416, n32968, n32969 );
nand U128257 ( n32969, n76469, P1_P3_INSTADDRPOINTER_REG_22_ );
nor U128258 ( n32968, n32970, n32971 );
nor U128259 ( n32971, n73278, n76898 );
nor U128260 ( n72480, n73824, n71104 );
and U128261 ( n62873, n76252, P3_REG0_REG_21_ );
and U128262 ( n39393, n76418, P4_REG0_REG_20_ );
and U128263 ( n39275, n76418, P4_REG0_REG_22_ );
nand U128264 ( n37721, n40286, n40287 );
nand U128265 ( n40287, n40288, P4_IR_REG_31_ );
nand U128266 ( n40286, P4_IR_REG_2_, n76795 );
and U128267 ( n40288, n40289, n40290 );
nand U128268 ( n37600, P2_P3_DATAO_REG_29_, n76457 );
nand U128269 ( n37740, n40240, n40241 );
nand U128270 ( n40240, P4_IR_REG_3_, n76795 );
or U128271 ( n40241, n40242, n76793 );
nand U128272 ( n33152, P1_P3_INSTADDRPOINTER_REG_17_, n33153 );
nand U128273 ( n33153, n33154, n33155 );
nor U128274 ( n33154, n33163, n33137 );
nor U128275 ( n33155, n33156, n33157 );
nand U128276 ( n4391, n33144, n33145 );
nand U128277 ( n33145, n76468, P1_P3_INSTADDRPOINTER_REG_17_ );
nor U128278 ( n33144, n33146, n33147 );
nor U128279 ( n33147, n74885, n76898 );
nand U128280 ( n36446, P2_P3_DATAO_REG_27_, n76457 );
and U128281 ( n11725, n16879, P4_DATAO_REG_0_ );
and U128282 ( n39451, n76418, P4_REG0_REG_19_ );
nand U128283 ( n4401, n33081, n33082 );
nand U128284 ( n33082, n76469, P1_P3_INSTADDRPOINTER_REG_19_ );
nor U128285 ( n33081, n33083, n33084 );
nor U128286 ( n33084, n73264, n76898 );
or U128287 ( n33698, n75940, n33748 );
nand U128288 ( n9231, n11544, n11545 );
nand U128289 ( n11545, P1_P1_UWORD_REG_7_, n76618 );
nor U128290 ( n11544, n11547, n11548 );
nor U128291 ( n11547, n75013, n76616 );
nand U128292 ( n9156, n11634, n11635 );
nand U128293 ( n11635, P1_P1_LWORD_REG_7_, n11504 );
nor U128294 ( n11634, n11637, n11548 );
nor U128295 ( n11637, n74739, n76615 );
nor U128296 ( n39341, n76415, n74545 );
nand U128297 ( n1151, n66169, n66170 );
nand U128298 ( n66169, P3_REG0_REG_6_, n61177 );
nand U128299 ( n66170, n75996, n60461 );
nand U128300 ( n1311, n60459, n60460 );
nand U128301 ( n60459, P3_REG1_REG_6_, n55262 );
nand U128302 ( n60460, n76004, n60461 );
nor U128303 ( n11874, n11877, n11878 );
nand U128304 ( n11878, P1_P1_INSTADDRPOINTER_REG_28_, n11879 );
nor U128305 ( n62739, n76249, n74551 );
nand U128306 ( n1141, n66339, n66340 );
nand U128307 ( n66339, P3_REG0_REG_4_, n61177 );
nand U128308 ( n66340, n75996, n60669 );
nand U128309 ( n1301, n60667, n60668 );
nand U128310 ( n60667, P3_REG1_REG_4_, n55262 );
nand U128311 ( n60668, n76004, n60669 );
nand U128312 ( n14460, P1_P1_INSTADDRPOINTER_REG_0_, n14410 );
nand U128313 ( n14353, n14457, n14458 );
or U128314 ( n14457, n14460, n11304 );
nand U128315 ( n14458, P1_P1_INSTADDRPOINTER_REG_1_, n14459 );
nand U128316 ( n14459, n11304, n14460 );
nand U128317 ( n15621, n46825, n46826 );
nand U128318 ( n46826, n76860, P2_P1_INSTADDRPOINTER_REG_18_ );
nor U128319 ( n46825, n46827, n46828 );
nor U128320 ( n46828, n74914, n76333 );
nand U128321 ( n11131, n67872, n67873 );
nand U128322 ( n67873, n76195, P2_P3_INSTADDRPOINTER_REG_18_ );
nor U128323 ( n67872, n67874, n67875 );
nor U128324 ( n67875, n74900, n76872 );
nand U128325 ( n6641, n25869, n25870 );
nand U128326 ( n25870, n76519, P1_P2_INSTADDRPOINTER_REG_18_ );
nor U128327 ( n25869, n25871, n25872 );
nor U128328 ( n25872, n74899, n76907 );
nand U128329 ( n13376, n59007, n59008 );
nand U128330 ( n59008, n76261, P2_P2_INSTADDRPOINTER_REG_18_ );
nor U128331 ( n59007, n59009, n59010 );
nor U128332 ( n59010, n74898, n76881 );
nand U128333 ( n16878, P4_DATAO_REG_17_, n16879 );
and U128334 ( n39342, n76418, P4_REG0_REG_21_ );
and U128335 ( n17472, n17036, P4_DATAO_REG_10_ );
nand U128336 ( n17175, n17036, P4_DATAO_REG_12_ );
nand U128337 ( n33557, P1_P3_INSTADDRPOINTER_REG_6_, n3175 );
nor U128338 ( n14184, n14392, P1_P1_INSTADDRPOINTER_REG_2_ );
nand U128339 ( n46655, P2_P1_INSTADDRPOINTER_REG_20_, n76341 );
nand U128340 ( n19556, n17036, P4_DATAO_REG_3_ );
nand U128341 ( n15971, n45349, n45350 );
nand U128342 ( n45350, P2_P1_UWORD_REG_6_, n76352 );
nor U128343 ( n45349, n45351, n45352 );
nor U128344 ( n45351, n75001, n76351 );
nand U128345 ( n15896, n45417, n45418 );
nand U128346 ( n45418, P2_P1_LWORD_REG_6_, n76352 );
nor U128347 ( n45417, n45419, n45352 );
nor U128348 ( n45419, n74704, n76349 );
xnor U128349 ( n11905, n11879, n12923 );
nor U128350 ( n12923, n12924, n4896 );
nor U128351 ( n12924, P1_P1_INSTADDRPOINTER_REG_27_, n76602 );
nand U128352 ( n8931, n12899, n12900 );
nand U128353 ( n12900, n76886, P1_P1_INSTADDRPOINTER_REG_27_ );
nor U128354 ( n12899, n12902, n12903 );
nor U128355 ( n12903, n75015, n76600 );
nand U128356 ( n46654, P2_P1_INSTADDRPOINTER_REG_18_, n76341 );
nor U128357 ( n62639, n76249, n74553 );
nand U128358 ( n14183, P1_P1_INSTADDRPOINTER_REG_2_, n14392 );
nand U128359 ( n11625, n16668, n16669 );
nand U128360 ( n16668, P1_BUF1_REG_6_, n76611 );
nand U128361 ( n16669, n16670, n76613 );
xnor U128362 ( n16670, n16672, n16673 );
nand U128363 ( n67702, P2_P3_INSTADDRPOINTER_REG_20_, n76197 );
nand U128364 ( n25697, P1_P2_INSTADDRPOINTER_REG_20_, n76521 );
nand U128365 ( n58837, P2_P2_INSTADDRPOINTER_REG_20_, n76263 );
nand U128366 ( n4426, n32887, n32888 );
nand U128367 ( n32888, n76469, P1_P3_INSTADDRPOINTER_REG_24_ );
nor U128368 ( n32887, n32889, n32890 );
nor U128369 ( n32890, n74994, n76899 );
nand U128370 ( n16408, n16409, n16410 );
nand U128371 ( n16410, P1_P1_INSTQUEUE_REG_14__6_, n16340 );
nand U128372 ( n16409, n4797, n31 );
nand U128373 ( n16305, n16307, n16308 );
nand U128374 ( n16308, P1_P1_INSTQUEUE_REG_13__6_, n16235 );
nand U128375 ( n16307, n4798, n31 );
nand U128376 ( n16094, n16095, n16097 );
nand U128377 ( n16097, P1_P1_INSTQUEUE_REG_11__6_, n16033 );
nand U128378 ( n16095, n4799, n31 );
nand U128379 ( n15987, n15988, n15989 );
nand U128380 ( n15989, P1_P1_INSTQUEUE_REG_10__6_, n15925 );
nand U128381 ( n15988, n4800, n31 );
nand U128382 ( n15888, n15889, n15890 );
nand U128383 ( n15890, P1_P1_INSTQUEUE_REG_9__6_, n15820 );
nand U128384 ( n15889, n4802, n31 );
nand U128385 ( n15674, n15675, n15677 );
nand U128386 ( n15677, P1_P1_INSTQUEUE_REG_7__6_, n15609 );
nand U128387 ( n15675, n4803, n31 );
nand U128388 ( n15573, n15574, n15575 );
nand U128389 ( n15575, P1_P1_INSTQUEUE_REG_6__6_, n15512 );
nand U128390 ( n15574, n4804, n31 );
nand U128391 ( n15467, n15468, n15469 );
nand U128392 ( n15469, P1_P1_INSTQUEUE_REG_5__6_, n15405 );
nand U128393 ( n15468, n4805, n31 );
nand U128394 ( n2366, n40168, n40169 );
nand U128395 ( n40168, P4_REG0_REG_4_, n76421 );
nand U128396 ( n40169, n76014, n38710 );
nand U128397 ( n2526, n38708, n38709 );
nand U128398 ( n38708, P4_REG1_REG_4_, n38617 );
nand U128399 ( n38709, n76017, n38710 );
nor U128400 ( n46872, n46876, n46877 );
xor U128401 ( n46876, n76342, P2_P1_INSTADDRPOINTER_REG_17_ );
nand U128402 ( n46877, n46878, n46871 );
nand U128403 ( n46878, P2_P1_INSTADDRPOINTER_REG_16_, n46875 );
nand U128404 ( n15616, n46853, n46854 );
nand U128405 ( n46854, n76860, P2_P1_INSTADDRPOINTER_REG_17_ );
nor U128406 ( n46853, n46855, n46856 );
nor U128407 ( n46856, n74904, n76333 );
and U128408 ( n62740, n76252, P3_REG0_REG_22_ );
nor U128409 ( n67919, n67923, n67924 );
xor U128410 ( n67923, n76198, P2_P3_INSTADDRPOINTER_REG_17_ );
nand U128411 ( n67924, n67925, n67918 );
nand U128412 ( n67925, P2_P3_INSTADDRPOINTER_REG_16_, n67922 );
nor U128413 ( n25916, n25920, n25921 );
xor U128414 ( n25920, n76522, P1_P2_INSTADDRPOINTER_REG_17_ );
nand U128415 ( n25921, n25922, n25915 );
nand U128416 ( n25922, P1_P2_INSTADDRPOINTER_REG_16_, n25919 );
nor U128417 ( n59054, n59058, n59059 );
xor U128418 ( n59058, n76264, P2_P2_INSTADDRPOINTER_REG_17_ );
nand U128419 ( n59059, n59060, n59053 );
nand U128420 ( n59060, P2_P2_INSTADDRPOINTER_REG_16_, n59057 );
nand U128421 ( n11126, n67900, n67901 );
nand U128422 ( n67901, n76195, P2_P3_INSTADDRPOINTER_REG_17_ );
nor U128423 ( n67900, n67902, n67903 );
nor U128424 ( n67903, n74884, n76872 );
nand U128425 ( n6636, n25897, n25898 );
nand U128426 ( n25898, n76519, P1_P2_INSTADDRPOINTER_REG_17_ );
nor U128427 ( n25897, n25899, n25900 );
nor U128428 ( n25900, n74883, n76907 );
nand U128429 ( n13371, n59035, n59036 );
nand U128430 ( n59036, n76261, P2_P2_INSTADDRPOINTER_REG_17_ );
nor U128431 ( n59035, n59037, n59038 );
nor U128432 ( n59038, n74882, n76881 );
nand U128433 ( n67701, P2_P3_INSTADDRPOINTER_REG_18_, n76197 );
nand U128434 ( n25696, P1_P2_INSTADDRPOINTER_REG_18_, n76521 );
nand U128435 ( n58836, P2_P2_INSTADDRPOINTER_REG_18_, n76263 );
nand U128436 ( n51131, n8235, P3_DATAO_REG_2_ );
or U128437 ( n14082, n75941, n14144 );
nand U128438 ( n33023, P1_P3_INSTADDRPOINTER_REG_20_, n76472 );
and U128439 ( n17171, n17036, P4_DATAO_REG_11_ );
nand U128440 ( n45416, n49612, n49613 );
nand U128441 ( n49612, P2_BUF1_REG_5_, n76478 );
nand U128442 ( n49613, n49614, n76476 );
xor U128443 ( n49614, n49615, n49616 );
nand U128444 ( n49316, n49317, n49318 );
nand U128445 ( n49318, P2_P1_INSTQUEUE_REG_13__5_, n49275 );
nand U128446 ( n49317, n7442, n277 );
nand U128447 ( n49125, n49126, n49127 );
nand U128448 ( n49127, P2_P1_INSTQUEUE_REG_11__5_, n49085 );
nand U128449 ( n49126, n7443, n277 );
nand U128450 ( n49047, n49048, n49049 );
nand U128451 ( n49049, P2_P1_INSTQUEUE_REG_10__5_, n48990 );
nand U128452 ( n49048, n7444, n277 );
nand U128453 ( n48952, n48953, n48954 );
nand U128454 ( n48954, P2_P1_INSTQUEUE_REG_9__5_, n48891 );
nand U128455 ( n48953, n7445, n277 );
nand U128456 ( n48758, n48759, n48760 );
nand U128457 ( n48760, P2_P1_INSTQUEUE_REG_7__5_, n48718 );
nand U128458 ( n48759, n7447, n277 );
nand U128459 ( n48665, n48666, n48667 );
nand U128460 ( n48667, P2_P1_INSTQUEUE_REG_6__5_, n48624 );
nand U128461 ( n48666, n7448, n277 );
nand U128462 ( n48587, n48588, n48589 );
nand U128463 ( n48589, P2_P1_INSTQUEUE_REG_5__5_, n48530 );
nand U128464 ( n48588, n7449, n277 );
nand U128465 ( n49409, n49410, n49411 );
nand U128466 ( n49411, P2_P1_INSTQUEUE_REG_14__5_, n49353 );
nand U128467 ( n49410, n7440, n277 );
and U128468 ( n49522, n49990, P3_DATAO_REG_0_ );
and U128469 ( n50006, DIN_22_, n76929 );
nand U128470 ( n51121, n50006, P3_DATAO_REG_3_ );
nand U128471 ( n37783, n40202, n40203 );
nand U128472 ( n40203, n40204, P4_IR_REG_31_ );
nand U128473 ( n40202, P4_IR_REG_4_, n76795 );
and U128474 ( n40204, n40205, n40206 );
nor U128475 ( n13027, P1_P1_INSTADDRPOINTER_REG_25_, n13029 );
xor U128476 ( n13029, n12930, n76603 );
nand U128477 ( n8921, n13004, n13005 );
nand U128478 ( n13005, n76886, P1_P1_INSTADDRPOINTER_REG_25_ );
nor U128479 ( n13004, n13007, n13008 );
nor U128480 ( n13008, n73305, n76600 );
nand U128481 ( n37799, n40165, n40166 );
nand U128482 ( n40165, P4_IR_REG_5_, n76795 );
or U128483 ( n40166, n40167, n76794 );
nand U128484 ( n36771, n36772, n36773 );
nand U128485 ( n36772, P4_REG3_REG_2_, n36488 );
nand U128486 ( n36773, n76830, n36774 );
nand U128487 ( n36774, n36775, n36776 );
nand U128488 ( n37298, P2_P3_DATAO_REG_30_, n76457 );
and U128489 ( n62640, n76252, P3_REG0_REG_23_ );
and U128490 ( n51105, n50006, P3_DATAO_REG_4_ );
nand U128491 ( n41154, n41155, n41156 );
nand U128492 ( n41155, P3_REG3_REG_2_, n40881 );
nand U128493 ( n41156, n76850, n41157 );
nand U128494 ( n41157, n41158, n41159 );
nand U128495 ( n37816, n40125, n40126 );
nand U128496 ( n40126, n40127, P4_IR_REG_31_ );
nand U128497 ( n40125, P4_IR_REG_6_, n76795 );
and U128498 ( n40127, n40128, n40129 );
nor U128499 ( n12974, n12977, n12978 );
and U128500 ( n12977, n12979, P1_P1_INSTADDRPOINTER_REG_26_ );
nor U128501 ( n12978, n12969, n12930 );
nand U128502 ( n8926, n12954, n12955 );
nand U128503 ( n12955, n76886, P1_P1_INSTADDRPOINTER_REG_26_ );
nor U128504 ( n12954, n12957, n12958 );
nor U128505 ( n12958, n73309, n76600 );
nand U128506 ( n4396, n33116, n33117 );
nand U128507 ( n33117, n76468, P1_P3_INSTADDRPOINTER_REG_18_ );
nor U128508 ( n33116, n33118, n33119 );
nor U128509 ( n33119, n74901, n76898 );
nand U128510 ( n51848, n8235, P3_DATAO_REG_1_ );
nand U128511 ( n13908, P1_P1_INSTADDRPOINTER_REG_6_, n4912 );
nand U128512 ( n2521, n38711, n38712 );
nand U128513 ( n38711, P4_REG1_REG_3_, n38617 );
nand U128514 ( n38712, n76017, n38713 );
nand U128515 ( n2361, n40207, n40208 );
nand U128516 ( n40207, P4_REG0_REG_3_, n76421 );
nand U128517 ( n40208, n76014, n38713 );
and U128518 ( n19233, n17036, P4_DATAO_REG_2_ );
nand U128519 ( n1136, n66416, n66417 );
nand U128520 ( n66416, P3_REG0_REG_3_, n61177 );
nand U128521 ( n66417, n75996, n60768 );
nand U128522 ( n1296, n60766, n60767 );
nand U128523 ( n60766, P3_REG1_REG_3_, n55262 );
nand U128524 ( n60767, n76004, n60768 );
nand U128525 ( n50927, n50006, P3_DATAO_REG_5_ );
nor U128526 ( n39216, n76415, n74600 );
and U128527 ( n12972, n12930, P1_P1_INSTADDRPOINTER_REG_25_ );
nor U128528 ( n72301, n74020, n71104 );
nand U128529 ( n40873, n40874, n40875 );
nand U128530 ( n40874, P3_REG3_REG_1_, n40881 );
nand U128531 ( n40875, n76851, n40876 );
xor U128532 ( n40876, n40877, n40878 );
nand U128533 ( n1291, n60873, n60874 );
nand U128534 ( n60873, P3_REG1_REG_2_, n55262 );
nand U128535 ( n60874, n76004, n60875 );
nand U128536 ( n1131, n66717, n66718 );
nand U128537 ( n66717, P3_REG0_REG_2_, n61177 );
nand U128538 ( n66718, n75996, n60875 );
xnor U128539 ( n12080, n13240, n13242 );
xor U128540 ( n13240, n76035, P1_P1_INSTADDRPOINTER_REG_21_ );
nor U128541 ( n13242, n4887, n13243 );
nand U128542 ( n13243, n13244, n13245 );
nand U128543 ( n8901, n13220, n13222 );
nand U128544 ( n13222, n76886, P1_P1_INSTADDRPOINTER_REG_21_ );
nor U128545 ( n13220, n13223, n13224 );
nor U128546 ( n13224, n74959, n76599 );
nand U128547 ( n2356, n40247, n40248 );
nand U128548 ( n40247, P4_REG0_REG_2_, n76421 );
nand U128549 ( n40248, n76014, n38716 );
nand U128550 ( n2516, n38714, n38715 );
nand U128551 ( n38714, P4_REG1_REG_2_, n38617 );
nand U128552 ( n38715, n76017, n38716 );
nand U128553 ( n13132, n13085, n13137 );
nand U128554 ( n13137, n4889, P1_P1_INSTADDRPOINTER_REG_22_ );
nand U128555 ( n8911, n13104, n13105 );
nand U128556 ( n13105, n76886, P1_P1_INSTADDRPOINTER_REG_23_ );
nor U128557 ( n13104, n13107, n13108 );
nor U128558 ( n13108, n74996, n76599 );
nand U128559 ( n50395, DIN_23_, n76929 );
nand U128560 ( n51145, n8239, P3_DATAO_REG_3_ );
nand U128561 ( n50670, n50006, P3_DATAO_REG_6_ );
nand U128562 ( n9236, n11539, n11540 );
nand U128563 ( n11540, P1_P1_UWORD_REG_6_, n76618 );
nor U128564 ( n11539, n11542, n11543 );
nor U128565 ( n11542, n75002, n76617 );
nand U128566 ( n9161, n11622, n11623 );
nand U128567 ( n11623, P1_P1_LWORD_REG_6_, n11504 );
nor U128568 ( n11622, n11624, n11543 );
nor U128569 ( n11624, n74705, n76615 );
nand U128570 ( n8896, n13269, n13270 );
nand U128571 ( n13270, n76886, P1_P1_INSTADDRPOINTER_REG_20_ );
nor U128572 ( n13269, n13272, n13273 );
nor U128573 ( n13273, n74952, n76599 );
nand U128574 ( n42299, n66374, n66375 );
nand U128575 ( n66375, n66376, P3_IR_REG_31_ );
nand U128576 ( n66374, P3_IR_REG_4_, n76841 );
and U128577 ( n66376, n16270, n16269 );
nand U128578 ( n36471, n36472, n36473 );
nand U128579 ( n36472, P4_REG3_REG_1_, n36488 );
nand U128580 ( n36473, n76831, n36474 );
nand U128581 ( n36474, n36475, n36476 );
and U128582 ( n18863, n17036, P4_DATAO_REG_1_ );
nand U128583 ( n15976, n45345, n45346 );
nand U128584 ( n45346, P2_P1_UWORD_REG_5_, n76352 );
nor U128585 ( n45345, n45347, n45348 );
nor U128586 ( n45347, n73288, n76351 );
nand U128587 ( n15901, n45413, n45414 );
nand U128588 ( n45414, P2_P1_LWORD_REG_5_, n76352 );
nor U128589 ( n45413, n45415, n45348 );
nor U128590 ( n45415, n73195, n76349 );
and U128591 ( n39217, n76418, P4_REG0_REG_23_ );
nor U128592 ( n62546, n76250, n74647 );
nand U128593 ( n32904, P1_P3_INSTADDRPOINTER_REG_23_, n76472 );
nand U128594 ( n32210, n32220, n32221 );
nand U128595 ( n32220, n32230, n32231 );
nand U128596 ( n32221, n32222, n32223 );
nor U128597 ( n32231, P1_P3_PHYADDRPOINTER_REG_17_, n32201 );
nand U128598 ( n16191, n44939, n44940 );
nor U128599 ( n44940, n44941, n44942 );
nor U128600 ( n44939, n44946, n44947 );
nor U128601 ( n44941, P2_P1_EAX_REG_5_, n44935 );
nor U128602 ( n42188, n42189, n73024 );
nor U128603 ( n42189, n42190, n42191 );
nor U128604 ( n42190, P3_REG1_REG_0_, n42194 );
nand U128605 ( n42191, n42192, n42193 );
nand U128606 ( n11620, n16632, n16633 );
nand U128607 ( n16632, P1_BUF1_REG_5_, n76611 );
nand U128608 ( n16633, n16634, n76613 );
xor U128609 ( n16634, n16635, n16637 );
nand U128610 ( n16458, n16854, P4_DATAO_REG_0_ );
nand U128611 ( n16398, n16399, n16400 );
nand U128612 ( n16400, P1_P1_INSTQUEUE_REG_14__5_, n16340 );
nand U128613 ( n16399, n4797, n26 );
nand U128614 ( n16295, n16297, n16298 );
nand U128615 ( n16298, P1_P1_INSTQUEUE_REG_13__5_, n16235 );
nand U128616 ( n16297, n4798, n26 );
nand U128617 ( n16084, n16085, n16087 );
nand U128618 ( n16087, P1_P1_INSTQUEUE_REG_11__5_, n16033 );
nand U128619 ( n16085, n4799, n26 );
nand U128620 ( n15977, n15978, n15979 );
nand U128621 ( n15979, P1_P1_INSTQUEUE_REG_10__5_, n15925 );
nand U128622 ( n15978, n4800, n26 );
nand U128623 ( n15878, n15879, n15880 );
nand U128624 ( n15880, P1_P1_INSTQUEUE_REG_9__5_, n15820 );
nand U128625 ( n15879, n4802, n26 );
nand U128626 ( n15664, n15665, n15667 );
nand U128627 ( n15667, P1_P1_INSTQUEUE_REG_7__5_, n15609 );
nand U128628 ( n15665, n4803, n26 );
nand U128629 ( n15563, n15564, n15565 );
nand U128630 ( n15565, P1_P1_INSTQUEUE_REG_6__5_, n15512 );
nand U128631 ( n15564, n4804, n26 );
nand U128632 ( n15457, n15458, n15459 );
nand U128633 ( n15459, P1_P1_INSTQUEUE_REG_5__5_, n15405 );
nand U128634 ( n15458, n4805, n26 );
nand U128635 ( n15611, n46899, n46900 );
nand U128636 ( n46900, n76860, P2_P1_INSTADDRPOINTER_REG_16_ );
nor U128637 ( n46899, n46901, n46902 );
nor U128638 ( n46902, n73253, n76333 );
nand U128639 ( n11121, n67946, n67947 );
nand U128640 ( n67947, n76195, P2_P3_INSTADDRPOINTER_REG_16_ );
nor U128641 ( n67946, n67948, n67949 );
nor U128642 ( n67949, n73249, n76872 );
nand U128643 ( n6631, n25943, n25944 );
nand U128644 ( n25944, n76519, P1_P2_INSTADDRPOINTER_REG_16_ );
nor U128645 ( n25943, n25945, n25946 );
nor U128646 ( n25946, n73248, n76907 );
nand U128647 ( n13366, n59081, n59082 );
nand U128648 ( n59082, n76261, P2_P2_INSTADDRPOINTER_REG_16_ );
nor U128649 ( n59081, n59083, n59084 );
nor U128650 ( n59084, n73247, n76881 );
nand U128651 ( n50399, n50006, P3_DATAO_REG_7_ );
nand U128652 ( n50897, n50006, P3_DATAO_REG_2_ );
nand U128653 ( n17052, DIN_21_, n76928 );
nand U128654 ( n18216, n8218, P4_DATAO_REG_4_ );
nand U128655 ( n42344, n66302, n66303 );
nand U128656 ( n66302, P3_IR_REG_5_, n76841 );
or U128657 ( n66303, n16142, n76839 );
nand U128658 ( n42234, n42235, n42236 );
nand U128659 ( n42235, P3_ADDR_REG_2_, n42201 );
nand U128660 ( n42236, n574, n42229 );
nor U128661 ( n39151, n76416, n74707 );
and U128662 ( n62547, n76252, P3_REG0_REG_24_ );
nand U128663 ( n45412, n49584, n49585 );
nand U128664 ( n49584, P2_BUF1_REG_4_, n76478 );
nand U128665 ( n49585, n49586, n76476 );
xor U128666 ( n49586, n49587, n49588 );
xor U128667 ( n32247, n3152, n33201 );
nor U128668 ( n33201, n33202, n33162 );
nor U128669 ( n33202, P1_P3_INSTADDRPOINTER_REG_16_, n76021 );
nand U128670 ( n4386, n33190, n33191 );
nand U128671 ( n33191, n76468, P1_P3_INSTADDRPOINTER_REG_16_ );
nor U128672 ( n33190, n33192, n33193 );
nor U128673 ( n33193, n73250, n76898 );
nor U128674 ( n37684, n37685, n73023 );
nor U128675 ( n37685, n37686, n37687 );
nor U128676 ( n37686, P4_REG2_REG_0_, n37690 );
nand U128677 ( n37687, n37688, n37689 );
nand U128678 ( n49308, n49309, n49310 );
nand U128679 ( n49310, P2_P1_INSTQUEUE_REG_13__4_, n49275 );
nand U128680 ( n49309, n7442, n270 );
nand U128681 ( n49117, n49118, n49119 );
nand U128682 ( n49119, P2_P1_INSTQUEUE_REG_11__4_, n49085 );
nand U128683 ( n49118, n7443, n270 );
nand U128684 ( n49039, n49040, n49041 );
nand U128685 ( n49041, P2_P1_INSTQUEUE_REG_10__4_, n48990 );
nand U128686 ( n49040, n7444, n270 );
nand U128687 ( n48944, n48945, n48946 );
nand U128688 ( n48946, P2_P1_INSTQUEUE_REG_9__4_, n48891 );
nand U128689 ( n48945, n7445, n270 );
nand U128690 ( n48657, n48658, n48659 );
nand U128691 ( n48659, P2_P1_INSTQUEUE_REG_6__4_, n48624 );
nand U128692 ( n48658, n7448, n270 );
nand U128693 ( n48579, n48580, n48581 );
nand U128694 ( n48581, P2_P1_INSTQUEUE_REG_5__4_, n48530 );
nand U128695 ( n48580, n7449, n270 );
nand U128696 ( n49401, n49402, n49403 );
nand U128697 ( n49403, P2_P1_INSTQUEUE_REG_14__4_, n49353 );
nand U128698 ( n49402, n7440, n270 );
nand U128699 ( n48750, n48751, n48752 );
nand U128700 ( n48752, P2_P1_INSTQUEUE_REG_7__4_, n48718 );
nand U128701 ( n48751, n7447, n270 );
nand U128702 ( n16853, P4_DATAO_REG_15_, n16854 );
nand U128703 ( n1286, n60971, n60972 );
nand U128704 ( n60971, P3_REG1_REG_1_, n55262 );
nand U128705 ( n60972, n76004, n60973 );
nand U128706 ( n1126, n66991, n66992 );
nand U128707 ( n66991, P3_REG0_REG_1_, n61177 );
nand U128708 ( n66992, n75996, n60973 );
nand U128709 ( n2511, n38717, n38718 );
nand U128710 ( n38717, P4_REG1_REG_1_, n38617 );
nand U128711 ( n38718, n76017, n38719 );
nand U128712 ( n2351, n40291, n40292 );
nand U128713 ( n40291, P4_REG0_REG_1_, n76421 );
nand U128714 ( n40292, n76014, n38719 );
nand U128715 ( n8906, n13175, n13177 );
nand U128716 ( n13177, n76886, P1_P1_INSTADDRPOINTER_REG_22_ );
nor U128717 ( n13175, n13178, n13179 );
nor U128718 ( n13179, n73281, n76599 );
nand U128719 ( n17981, n8218, P4_DATAO_REG_5_ );
nand U128720 ( n40393, n2093, n40394 );
nand U128721 ( n40394, n40395, n74741 );
nor U128722 ( n40395, P4_D_REG_24_, P4_D_REG_23_ );
nand U128723 ( n47046, n47093, n47094 );
nand U128724 ( n47093, P2_P1_INSTADDRPOINTER_REG_11_, n76342 );
nand U128725 ( n47094, n47020, n7539 );
and U128726 ( n46024, n47040, n47041 );
nand U128727 ( n47040, n47049, n47050 );
nand U128728 ( n47041, n47042, n47043 );
nand U128729 ( n47050, P2_P1_INSTADDRPOINTER_REG_13_, n76342 );
nand U128730 ( n15596, n47029, n47030 );
nand U128731 ( n47030, n76860, P2_P1_INSTADDRPOINTER_REG_13_ );
nor U128732 ( n47029, n47031, n47032 );
nor U128733 ( n47032, n73239, n76333 );
nand U128734 ( n68077, n68124, n68125 );
nand U128735 ( n68124, P2_P3_INSTADDRPOINTER_REG_11_, n76198 );
nand U128736 ( n68125, n68055, n5753 );
nand U128737 ( n26074, n26121, n26122 );
nand U128738 ( n26121, P1_P2_INSTADDRPOINTER_REG_11_, n76522 );
nand U128739 ( n26122, n26052, n3995 );
nand U128740 ( n59215, n59262, n59263 );
nand U128741 ( n59262, P2_P2_INSTADDRPOINTER_REG_11_, n76264 );
nand U128742 ( n59263, n59193, n6628 );
and U128743 ( n66964, n68071, n68072 );
nand U128744 ( n68071, n68080, n68081 );
nand U128745 ( n68072, n68073, n68074 );
nand U128746 ( n68081, P2_P3_INSTADDRPOINTER_REG_13_, n76198 );
and U128747 ( n25088, n26068, n26069 );
nand U128748 ( n26068, n26077, n26078 );
nand U128749 ( n26069, n26070, n26071 );
nand U128750 ( n26078, P1_P2_INSTADDRPOINTER_REG_13_, n76522 );
and U128751 ( n58223, n59209, n59210 );
nand U128752 ( n59209, n59218, n59219 );
nand U128753 ( n59210, n59211, n59212 );
nand U128754 ( n59219, P2_P2_INSTADDRPOINTER_REG_13_, n76264 );
nand U128755 ( n11106, n68060, n68061 );
nand U128756 ( n68061, n76195, P2_P3_INSTADDRPOINTER_REG_13_ );
nor U128757 ( n68060, n68062, n68063 );
nor U128758 ( n68063, n73236, n76872 );
nand U128759 ( n6616, n26057, n26058 );
nand U128760 ( n26058, n76519, P1_P2_INSTADDRPOINTER_REG_13_ );
nor U128761 ( n26057, n26059, n26060 );
nor U128762 ( n26060, n73234, n76907 );
nand U128763 ( n13351, n59198, n59199 );
nand U128764 ( n59199, n76261, P2_P2_INSTADDRPOINTER_REG_13_ );
nor U128765 ( n59198, n59200, n59201 );
nor U128766 ( n59201, n73233, n76881 );
nand U128767 ( n40392, n2093, n40396 );
nand U128768 ( n40396, n40397, n40398 );
nor U128769 ( n40397, P4_D_REG_19_, P4_D_REG_18_ );
nor U128770 ( n40398, P4_D_REG_21_, P4_D_REG_20_ );
nor U128771 ( n42187, P3_IR_REG_0_, n42195 );
nor U128772 ( n42195, n42196, n42197 );
nor U128773 ( n42196, n73633, n42198 );
nor U128774 ( n42197, n73579, n42194 );
nand U128775 ( n16702, P3_IR_REG_2_, n66759 );
nand U128776 ( n66759, n73024, n73566 );
nand U128777 ( n50011, n8239, P3_DATAO_REG_7_ );
nand U128778 ( n13404, P1_P1_INSTADDRPOINTER_REG_17_, n13405 );
nand U128779 ( n13405, n13407, n13408 );
nor U128780 ( n13407, n13418, n13385 );
nor U128781 ( n13408, n13409, n13410 );
nand U128782 ( n8881, n13394, n13395 );
nand U128783 ( n13395, n76887, P1_P1_INSTADDRPOINTER_REG_17_ );
nor U128784 ( n13394, n13397, n13398 );
nor U128785 ( n13398, n74905, n76599 );
nor U128786 ( n62430, n76250, n74725 );
nand U128787 ( n8891, n13315, n13317 );
nand U128788 ( n13317, n76887, P1_P1_INSTADDRPOINTER_REG_19_ );
nor U128789 ( n13315, n13318, n13319 );
nor U128790 ( n13319, n73268, n76599 );
xnor U128791 ( n40315, n73535, P4_IR_REG_0_ );
and U128792 ( n49743, n50006, P3_DATAO_REG_8_ );
nor U128793 ( n47090, P2_P1_INSTADDRPOINTER_REG_12_, n47091 );
xor U128794 ( n47091, n47046, n76006 );
nand U128795 ( n15591, n47070, n47071 );
nand U128796 ( n47071, n76860, P2_P1_INSTADDRPOINTER_REG_12_ );
nor U128797 ( n47070, n47072, n47073 );
nor U128798 ( n47073, n74815, n76333 );
nor U128799 ( n68121, P2_P3_INSTADDRPOINTER_REG_12_, n68122 );
xor U128800 ( n68122, n68077, n75990 );
nor U128801 ( n26118, P1_P2_INSTADDRPOINTER_REG_12_, n26119 );
xor U128802 ( n26119, n26074, n76027 );
nor U128803 ( n59259, P2_P2_INSTADDRPOINTER_REG_12_, n59260 );
xor U128804 ( n59260, n59215, n75998 );
nand U128805 ( n11101, n68101, n68102 );
nand U128806 ( n68102, n76195, P2_P3_INSTADDRPOINTER_REG_12_ );
nor U128807 ( n68101, n68103, n68104 );
nor U128808 ( n68104, n74800, n76872 );
nand U128809 ( n6611, n26098, n26099 );
nand U128810 ( n26099, n76519, P1_P2_INSTADDRPOINTER_REG_12_ );
nor U128811 ( n26098, n26100, n26101 );
nor U128812 ( n26101, n74799, n76907 );
nand U128813 ( n13346, n59239, n59240 );
nand U128814 ( n59240, n76261, P2_P2_INSTADDRPOINTER_REG_12_ );
nor U128815 ( n59239, n59241, n59242 );
nor U128816 ( n59242, n74798, n76881 );
and U128817 ( n39152, n76418, P4_REG0_REG_24_ );
nand U128818 ( n50624, n8239, P3_DATAO_REG_1_ );
nor U128819 ( n37683, P4_IR_REG_0_, n37691 );
nor U128820 ( n37691, n37692, n37693 );
nor U128821 ( n37692, n73798, n37694 );
nor U128822 ( n37693, n73799, n37690 );
nor U128823 ( n39037, n76416, n74716 );
nand U128824 ( n50884, n50006, P3_DATAO_REG_1_ );
xor U128825 ( n45547, n46321, n75052 );
nand U128826 ( n46321, n45599, P2_P1_INSTADDRPOINTER_REG_30_ );
nand U128827 ( n47611, P2_P1_INSTADDRPOINTER_REG_2_, n47674 );
nand U128828 ( n47175, n47190, n47191 );
or U128829 ( n47190, n47194, n47193 );
nand U128830 ( n47191, P2_P1_INSTADDRPOINTER_REG_8_, n47192 );
nand U128831 ( n47192, n47193, n47194 );
nor U128832 ( n47338, n47341, n47342 );
nor U128833 ( n47341, P2_P1_INSTADDRPOINTER_REG_5_, n47337 );
or U128834 ( n47342, n7594, n47343 );
and U128835 ( n47244, n47289, n47290 );
or U128836 ( n47289, n47293, n47292 );
nand U128837 ( n47290, P2_P1_INSTADDRPOINTER_REG_6_, n47291 );
nand U128838 ( n47291, n47292, n47293 );
and U128839 ( n47193, n47241, n47242 );
or U128840 ( n47241, n47245, n47244 );
nand U128841 ( n47242, P2_P1_INSTADDRPOINTER_REG_7_, n47243 );
nand U128842 ( n47243, n47244, n47245 );
nor U128843 ( n39092, n76416, n74706 );
nor U128844 ( n72294, n74274, n71104 );
nand U128845 ( n9241, n11534, n11535 );
nand U128846 ( n11535, P1_P1_UWORD_REG_5_, n76618 );
nor U128847 ( n11534, n11537, n11538 );
nor U128848 ( n11537, n73289, n76617 );
nand U128849 ( n9166, n11617, n11618 );
nand U128850 ( n11618, P1_P1_LWORD_REG_5_, n11504 );
nor U128851 ( n11617, n11619, n11538 );
nor U128852 ( n11619, n73196, n76615 );
nand U128853 ( n37726, n37727, n37728 );
nand U128854 ( n37727, P4_ADDR_REG_2_, n2080 );
nand U128855 ( n37728, n2077, n37721 );
and U128856 ( n39093, n76418, P4_REG0_REG_25_ );
nand U128857 ( n2506, n38724, n38725 );
nand U128858 ( n38724, P4_REG1_REG_0_, n38617 );
nand U128859 ( n38725, n76017, n38726 );
nand U128860 ( n2346, n40316, n40317 );
nand U128861 ( n40316, P4_REG0_REG_0_, n76421 );
nand U128862 ( n40317, n76014, n38726 );
nand U128863 ( n1281, n61068, n61069 );
nand U128864 ( n61068, P3_REG1_REG_0_, n55262 );
nand U128865 ( n61069, n76004, n61070 );
nand U128866 ( n1121, n67210, n67211 );
nand U128867 ( n67210, P3_REG0_REG_0_, n61177 );
nand U128868 ( n67211, n75996, n61070 );
nor U128869 ( n47608, n47674, P2_P1_INSTADDRPOINTER_REG_2_ );
and U128870 ( n39038, n76418, P4_REG0_REG_26_ );
and U128871 ( n37114, n40404, n40405 );
nand U128872 ( n40405, n40406, n40402 );
nand U128873 ( n40404, P4_D_REG_1_, n2093 );
nand U128874 ( n40129, P4_IR_REG_6_, n40630 );
nand U128875 ( n40630, n2208, n73948 );
nand U128876 ( n9456, n11247, n11248 );
nor U128877 ( n11248, n11249, n11250 );
nor U128878 ( n11247, n11255, n11257 );
nor U128879 ( n11249, P1_P1_EAX_REG_5_, n11235 );
nor U128880 ( n47042, n47047, n47048 );
nor U128881 ( n47048, n73099, n76341 );
and U128882 ( n47047, n47046, P2_P1_INSTADDRPOINTER_REG_12_ );
nor U128883 ( n68073, n68078, n68079 );
nor U128884 ( n68079, n73104, n76197 );
and U128885 ( n68078, n68077, P2_P3_INSTADDRPOINTER_REG_12_ );
nor U128886 ( n26070, n26075, n26076 );
nor U128887 ( n26076, n73105, n76521 );
and U128888 ( n26075, n26074, P1_P2_INSTADDRPOINTER_REG_12_ );
nor U128889 ( n59211, n59216, n59217 );
nor U128890 ( n59217, n73106, n76263 );
and U128891 ( n59216, n59215, P2_P2_INSTADDRPOINTER_REG_12_ );
and U128892 ( n62431, n76252, P3_REG0_REG_25_ );
nand U128893 ( n13245, P1_P1_INSTADDRPOINTER_REG_20_, n76035 );
nand U128894 ( n45184, n66222, n66223 );
nand U128895 ( n66223, n66224, P3_IR_REG_31_ );
nand U128896 ( n66222, P3_IR_REG_6_, n76841 );
and U128897 ( n66224, n16002, n16000 );
nand U128898 ( n40290, P4_IR_REG_2_, n40652 );
nand U128899 ( n40652, n73023, n73535 );
nand U128900 ( n8916, n13065, n13067 );
nand U128901 ( n13067, n76886, P1_P1_INSTADDRPOINTER_REG_24_ );
nor U128902 ( n13065, n13068, n13069 );
nor U128903 ( n13069, n75006, n76600 );
nand U128904 ( n37827, n40076, n40077 );
nand U128905 ( n40076, P4_IR_REG_7_, n76795 );
or U128906 ( n40077, n40078, n76794 );
xor U128907 ( n45575, n45599, P2_P1_INSTADDRPOINTER_REG_30_ );
and U128908 ( n37113, n40399, n40400 );
nand U128909 ( n40400, n40401, n40402 );
nand U128910 ( n40399, P4_D_REG_0_, n2093 );
xor U128911 ( n45960, n46961, n46914 );
xor U128912 ( n46961, n76342, P2_P1_INSTADDRPOINTER_REG_15_ );
nand U128913 ( n15606, n46943, n46944 );
nand U128914 ( n46944, n76860, P2_P1_INSTADDRPOINTER_REG_15_ );
nor U128915 ( n46943, n46945, n46946 );
nor U128916 ( n46946, n74868, n76333 );
xor U128917 ( n66911, n67996, n67961 );
xor U128918 ( n67996, n76198, P2_P3_INSTADDRPOINTER_REG_15_ );
xor U128919 ( n25035, n25993, n25958 );
xor U128920 ( n25993, n76522, P1_P2_INSTADDRPOINTER_REG_15_ );
xor U128921 ( n58170, n59131, n59096 );
xor U128922 ( n59131, n76264, P2_P2_INSTADDRPOINTER_REG_15_ );
nand U128923 ( n11116, n67978, n67979 );
nand U128924 ( n67979, n76195, P2_P3_INSTADDRPOINTER_REG_15_ );
nor U128925 ( n67978, n67980, n67981 );
nor U128926 ( n67981, n74840, n76872 );
nand U128927 ( n6626, n25975, n25976 );
nand U128928 ( n25976, n76519, P1_P2_INSTADDRPOINTER_REG_15_ );
nor U128929 ( n25975, n25977, n25978 );
nor U128930 ( n25978, n74838, n76907 );
nand U128931 ( n13361, n59113, n59114 );
nand U128932 ( n59114, n76261, P2_P2_INSTADDRPOINTER_REG_15_ );
nor U128933 ( n59113, n59115, n59116 );
nor U128934 ( n59116, n74837, n76881 );
nand U128935 ( n47531, n47676, n47677 );
nand U128936 ( n47676, n47680, n47679 );
nand U128937 ( n47677, P2_P1_INSTADDRPOINTER_REG_1_, n47678 );
or U128938 ( n47678, n47679, n47680 );
nand U128939 ( n42678, n66121, n66122 );
nand U128940 ( n66121, P3_IR_REG_7_, n76841 );
or U128941 ( n66122, n15873, n76840 );
nand U128942 ( n38606, n38607, n38608 );
nand U128943 ( n38608, n76446, P4_REG3_REG_0_ );
nand U128944 ( n38607, n38609, n76811 );
nand U128945 ( n17053, DIN_22_, n76928 );
nand U128946 ( n18164, n8214, P4_DATAO_REG_3_ );
nand U128947 ( n37943, n37996, n37997 );
nand U128948 ( n37996, n37928, n37930 );
nand U128949 ( n37997, P4_REG1_REG_14_, n37998 );
or U128950 ( n37998, n37928, n37930 );
nand U128951 ( n37881, n38008, n38009 );
nand U128952 ( n38008, n37870, n37872 );
nand U128953 ( n38009, P4_REG1_REG_10_, n38010 );
or U128954 ( n38010, n37870, n37872 );
nand U128955 ( n37825, n38020, n38021 );
nand U128956 ( n38020, n37811, n37816 );
nand U128957 ( n38021, P4_REG1_REG_6_, n38022 );
or U128958 ( n38022, n37811, n37816 );
nand U128959 ( n37915, n38002, n38003 );
nand U128960 ( n38002, n37895, n37897 );
nand U128961 ( n38003, P4_REG1_REG_12_, n38004 );
or U128962 ( n38004, n37895, n37897 );
nand U128963 ( n37853, n38014, n38015 );
nand U128964 ( n38014, n37843, n37841 );
nand U128965 ( n38015, P4_REG1_REG_8_, n38016 );
or U128966 ( n38016, n37843, n37841 );
nand U128967 ( n37742, n38032, n38033 );
nand U128968 ( n38032, n37719, n37721 );
nand U128969 ( n38033, P4_REG1_REG_2_, n38034 );
or U128970 ( n38034, n37719, n37721 );
nand U128971 ( n37953, n37993, n37994 );
nand U128972 ( n37993, n37943, n37941 );
nand U128973 ( n37994, P4_REG1_REG_15_, n37995 );
or U128974 ( n37995, n37943, n37941 );
nand U128975 ( n37928, n37999, n38000 );
nand U128976 ( n37999, n37915, n37913 );
nand U128977 ( n38000, P4_REG1_REG_13_, n38001 );
or U128978 ( n38001, n37915, n37913 );
nand U128979 ( n37895, n38005, n38006 );
nand U128980 ( n38005, n37881, n37883 );
nand U128981 ( n38006, P4_REG1_REG_11_, n38007 );
or U128982 ( n38007, n37881, n37883 );
nand U128983 ( n37870, n38011, n38012 );
nand U128984 ( n38011, n37853, n37855 );
nand U128985 ( n38012, P4_REG1_REG_9_, n38013 );
or U128986 ( n38013, n37853, n37855 );
nand U128987 ( n37843, n38017, n38018 );
nand U128988 ( n38017, n37825, n37827 );
nand U128989 ( n38018, P4_REG1_REG_7_, n38019 );
or U128990 ( n38019, n37825, n37827 );
nand U128991 ( n37811, n38023, n38024 );
nand U128992 ( n38023, n37801, n37799 );
nand U128993 ( n38024, P4_REG1_REG_5_, n38025 );
or U128994 ( n38025, n37801, n37799 );
nand U128995 ( n37781, n38029, n38030 );
nand U128996 ( n38029, n37742, n37740 );
nand U128997 ( n38030, P4_REG1_REG_3_, n38031 );
or U128998 ( n38031, n37742, n37740 );
nand U128999 ( n37719, n38035, n38036 );
nand U129000 ( n38035, n37704, n37706 );
nand U129001 ( n38036, P4_REG1_REG_1_, n38037 );
or U129002 ( n38037, n37706, n37704 );
nand U129003 ( n15981, n45341, n45342 );
nand U129004 ( n45342, P2_P1_UWORD_REG_4_, n76352 );
nor U129005 ( n45341, n45343, n45344 );
nor U129006 ( n45343, n74965, n76351 );
nand U129007 ( n15906, n45409, n45410 );
nand U129008 ( n45410, P2_P1_LWORD_REG_4_, n76352 );
nor U129009 ( n45409, n45411, n45344 );
nor U129010 ( n45411, n74681, n76349 );
nand U129011 ( n37982, n37983, n37984 );
nand U129012 ( n37984, n37985, n37986 );
nand U129013 ( n37986, P4_REG1_REG_17_, n37987 );
nand U129014 ( n37967, n37990, n37991 );
nand U129015 ( n37990, n37953, n37955 );
nand U129016 ( n37991, P4_REG1_REG_16_, n37992 );
or U129017 ( n37992, n37953, n37955 );
nand U129018 ( n37801, n38026, n38027 );
nand U129019 ( n38026, n37781, n37783 );
nand U129020 ( n38027, P4_REG1_REG_4_, n38028 );
or U129021 ( n38028, n37781, n37783 );
nand U129022 ( n37786, n38089, n38090 );
nand U129023 ( n38089, n37738, n37740 );
nand U129024 ( n38090, P4_REG2_REG_3_, n38091 );
or U129025 ( n38091, n37738, n37740 );
nand U129026 ( n37724, n38095, n38096 );
nand U129027 ( n38095, n37708, n37706 );
nand U129028 ( n38096, P4_REG2_REG_1_, n38097 );
or U129029 ( n38097, n37706, n37708 );
nand U129030 ( n37738, n38092, n38093 );
nand U129031 ( n38092, n37724, n37721 );
nand U129032 ( n38093, P4_REG2_REG_2_, n38094 );
or U129033 ( n38094, n37724, n37721 );
nand U129034 ( n37814, n38083, n38084 );
nand U129035 ( n38083, n37797, n37799 );
nand U129036 ( n38084, P4_REG2_REG_5_, n38085 );
or U129037 ( n38085, n37797, n37799 );
nand U129038 ( n37839, n38077, n38078 );
nand U129039 ( n38077, n37829, n37827 );
nand U129040 ( n38078, P4_REG2_REG_7_, n38079 );
or U129041 ( n38079, n37829, n37827 );
nand U129042 ( n37867, n38071, n38072 );
nand U129043 ( n38071, n37857, n37855 );
nand U129044 ( n38072, P4_REG2_REG_9_, n38073 );
or U129045 ( n38073, n37857, n37855 );
nand U129046 ( n37899, n38065, n38066 );
nand U129047 ( n38065, n37885, n37883 );
nand U129048 ( n38066, P4_REG2_REG_11_, n38067 );
or U129049 ( n38067, n37885, n37883 );
nand U129050 ( n37925, n38059, n38060 );
nand U129051 ( n38059, n37911, n37913 );
nand U129052 ( n38060, P4_REG2_REG_13_, n38061 );
or U129053 ( n38061, n37911, n37913 );
nand U129054 ( n37957, n38053, n38054 );
nand U129055 ( n38053, n37939, n37941 );
nand U129056 ( n38054, P4_REG2_REG_15_, n38055 );
or U129057 ( n38055, n37939, n37941 );
nand U129058 ( n37829, n38080, n38081 );
nand U129059 ( n38080, n37814, n37816 );
nand U129060 ( n38081, P4_REG2_REG_6_, n38082 );
or U129061 ( n38082, n37814, n37816 );
nand U129062 ( n37885, n38068, n38069 );
nand U129063 ( n38068, n37867, n37872 );
nand U129064 ( n38069, P4_REG2_REG_10_, n38070 );
or U129065 ( n38070, n37867, n37872 );
nand U129066 ( n37939, n38056, n38057 );
nand U129067 ( n38056, n37925, n37930 );
nand U129068 ( n38057, P4_REG2_REG_14_, n38058 );
or U129069 ( n38058, n37925, n37930 );
nand U129070 ( n38044, n38045, n38046 );
nand U129071 ( n38046, P4_REG2_REG_17_, n38047 );
nand U129072 ( n37857, n38074, n38075 );
nand U129073 ( n38074, n37839, n37841 );
nand U129074 ( n38075, P4_REG2_REG_8_, n38076 );
or U129075 ( n38076, n37839, n37841 );
nand U129076 ( n37911, n38062, n38063 );
nand U129077 ( n38062, n37899, n37897 );
nand U129078 ( n38063, P4_REG2_REG_12_, n38064 );
or U129079 ( n38064, n37899, n37897 );
nand U129080 ( n37971, n38050, n38051 );
nand U129081 ( n38050, n37957, n37955 );
nand U129082 ( n38051, P4_REG2_REG_16_, n38052 );
or U129083 ( n38052, n37957, n37955 );
nand U129084 ( n37797, n38086, n38087 );
nand U129085 ( n38086, n37786, n37783 );
nand U129086 ( n38087, P4_REG2_REG_4_, n38088 );
or U129087 ( n38088, n37786, n37783 );
nor U129088 ( n62364, n76250, n74768 );
nor U129089 ( n47529, P2_P1_INSTADDRPOINTER_REG_3_, n47525 );
and U129090 ( n62365, n76252, P3_REG0_REG_26_ );
nand U129091 ( n33455, n33470, n33471 );
or U129092 ( n33470, n33474, n33473 );
nand U129093 ( n33471, P1_P3_INSTADDRPOINTER_REG_8_, n33472 );
nand U129094 ( n33472, n33473, n33474 );
nand U129095 ( n33876, P1_P3_INSTADDRPOINTER_REG_2_, n33939 );
nor U129096 ( n33614, n33617, n33618 );
nor U129097 ( n33617, P1_P3_INSTADDRPOINTER_REG_5_, n33613 );
or U129098 ( n33618, n3208, n33619 );
and U129099 ( n33473, n33517, n33518 );
or U129100 ( n33517, n33521, n33520 );
nand U129101 ( n33518, P1_P3_INSTADDRPOINTER_REG_7_, n33519 );
nand U129102 ( n33519, n33520, n33521 );
and U129103 ( n33520, n33564, n33565 );
or U129104 ( n33564, n33568, n33567 );
nand U129105 ( n33565, P1_P3_INSTADDRPOINTER_REG_6_, n33566 );
nand U129106 ( n33566, n33567, n33568 );
nand U129107 ( n11615, n16595, n16597 );
nand U129108 ( n16595, P1_BUF1_REG_4_, n76611 );
nand U129109 ( n16597, n16598, n76613 );
xnor U129110 ( n16598, n16599, n16600 );
nand U129111 ( n68632, P2_P3_INSTADDRPOINTER_REG_2_, n68695 );
nand U129112 ( n26631, P1_P2_INSTADDRPOINTER_REG_2_, n26694 );
nand U129113 ( n59773, P2_P2_INSTADDRPOINTER_REG_2_, n59836 );
nand U129114 ( n26205, n26220, n26221 );
or U129115 ( n26220, n26224, n26223 );
nand U129116 ( n26221, P1_P2_INSTADDRPOINTER_REG_8_, n26222 );
nand U129117 ( n26222, n26223, n26224 );
nand U129118 ( n59344, n59359, n59360 );
or U129119 ( n59359, n59363, n59362 );
nand U129120 ( n59360, P2_P2_INSTADDRPOINTER_REG_8_, n59361 );
nand U129121 ( n59361, n59362, n59363 );
nor U129122 ( n68370, n68373, n68374 );
nor U129123 ( n68373, P2_P3_INSTADDRPOINTER_REG_5_, n68369 );
or U129124 ( n68374, n5807, n68375 );
nor U129125 ( n26369, n26372, n26373 );
nor U129126 ( n26372, P1_P2_INSTADDRPOINTER_REG_5_, n26368 );
or U129127 ( n26373, n4040, n26374 );
nor U129128 ( n59508, n59511, n59512 );
nor U129129 ( n59511, P2_P2_INSTADDRPOINTER_REG_5_, n59507 );
or U129130 ( n59512, n6673, n59513 );
and U129131 ( n68275, n68320, n68321 );
or U129132 ( n68320, n68324, n68323 );
nand U129133 ( n68321, P2_P3_INSTADDRPOINTER_REG_6_, n68322 );
nand U129134 ( n68322, n68323, n68324 );
and U129135 ( n68224, n68272, n68273 );
or U129136 ( n68272, n68276, n68275 );
nand U129137 ( n68273, P2_P3_INSTADDRPOINTER_REG_7_, n68274 );
nand U129138 ( n68274, n68275, n68276 );
and U129139 ( n26223, n26271, n26272 );
or U129140 ( n26271, n26275, n26274 );
nand U129141 ( n26272, P1_P2_INSTADDRPOINTER_REG_7_, n26273 );
nand U129142 ( n26273, n26274, n26275 );
and U129143 ( n59362, n59410, n59411 );
or U129144 ( n59410, n59414, n59413 );
nand U129145 ( n59411, P2_P2_INSTADDRPOINTER_REG_7_, n59412 );
nand U129146 ( n59412, n59413, n59414 );
and U129147 ( n26274, n26319, n26320 );
or U129148 ( n26319, n26323, n26322 );
nand U129149 ( n26320, P1_P2_INSTADDRPOINTER_REG_6_, n26321 );
nand U129150 ( n26321, n26322, n26323 );
and U129151 ( n59413, n59458, n59459 );
or U129152 ( n59458, n59462, n59461 );
nand U129153 ( n59459, P2_P2_INSTADDRPOINTER_REG_6_, n59460 );
nand U129154 ( n59460, n59461, n59462 );
nand U129155 ( n68206, n68221, n68222 );
or U129156 ( n68221, n68225, n68224 );
nand U129157 ( n68222, P2_P3_INSTADDRPOINTER_REG_8_, n68223 );
nand U129158 ( n68223, n68224, n68225 );
nand U129159 ( n45618, n74974, n46462 );
nand U129160 ( n46462, n45688, P2_P1_INSTADDRPOINTER_REG_27_ );
nand U129161 ( n16285, n16287, n16288 );
nand U129162 ( n16288, P1_P1_INSTQUEUE_REG_13__4_, n16235 );
nand U129163 ( n16287, n4798, n21 );
nand U129164 ( n16074, n16075, n16077 );
nand U129165 ( n16077, P1_P1_INSTQUEUE_REG_11__4_, n16033 );
nand U129166 ( n16075, n4799, n21 );
nand U129167 ( n15967, n15968, n15969 );
nand U129168 ( n15969, P1_P1_INSTQUEUE_REG_10__4_, n15925 );
nand U129169 ( n15968, n4800, n21 );
nand U129170 ( n15862, n15863, n15864 );
nand U129171 ( n15864, P1_P1_INSTQUEUE_REG_9__4_, n15820 );
nand U129172 ( n15863, n4802, n21 );
nand U129173 ( n15553, n15554, n15555 );
nand U129174 ( n15555, P1_P1_INSTQUEUE_REG_6__4_, n15512 );
nand U129175 ( n15554, n4804, n21 );
nand U129176 ( n15447, n15448, n15449 );
nand U129177 ( n15449, P1_P1_INSTQUEUE_REG_5__4_, n15405 );
nand U129178 ( n15448, n4805, n21 );
nand U129179 ( n16382, n16383, n16384 );
nand U129180 ( n16384, P1_P1_INSTQUEUE_REG_14__4_, n16340 );
nand U129181 ( n16383, n4797, n21 );
nand U129182 ( n15654, n15655, n15657 );
nand U129183 ( n15657, P1_P1_INSTQUEUE_REG_7__4_, n15609 );
nand U129184 ( n15655, n4803, n21 );
xor U129185 ( n12180, n13373, n13039 );
xor U129186 ( n13373, n76035, P1_P1_INSTADDRPOINTER_REG_18_ );
nand U129187 ( n8886, n13359, n13360 );
nand U129188 ( n13360, n76887, P1_P1_INSTADDRPOINTER_REG_18_ );
nor U129189 ( n13359, n13362, n13363 );
nor U129190 ( n13363, n74915, n76599 );
nor U129191 ( n38845, n76416, n74784 );
nand U129192 ( n40206, P4_IR_REG_4_, n40641 );
nand U129193 ( n40641, n2209, n73803 );
nor U129194 ( n38911, n76416, n74783 );
nor U129195 ( n38970, n76416, n74781 );
nor U129196 ( n33873, n33939, P1_P3_INSTADDRPOINTER_REG_2_ );
nor U129197 ( n62247, n76250, n74813 );
nor U129198 ( n68629, n68695, P2_P3_INSTADDRPOINTER_REG_2_ );
nor U129199 ( n26628, n26694, P1_P2_INSTADDRPOINTER_REG_2_ );
nor U129200 ( n59770, n59836, P2_P2_INSTADDRPOINTER_REG_2_ );
nand U129201 ( n67294, n619, n67295 );
nand U129202 ( n67295, n67296, n74623 );
nor U129203 ( n67296, P3_D_REG_24_, P3_D_REG_23_ );
xnor U129204 ( n31849, n32603, P1_P3_INSTADDRPOINTER_REG_31_ );
nand U129205 ( n32603, n31901, P1_P3_INSTADDRPOINTER_REG_30_ );
nor U129206 ( n33364, P1_P3_INSTADDRPOINTER_REG_12_, n33365 );
xor U129207 ( n33365, n76471, n3153 );
nand U129208 ( n67293, n619, n67297 );
nand U129209 ( n67297, n67298, n67299 );
nor U129210 ( n67298, P3_D_REG_19_, P3_D_REG_18_ );
nor U129211 ( n67299, P3_D_REG_21_, P3_D_REG_20_ );
nand U129212 ( n4366, n33344, n33345 );
nand U129213 ( n33345, n76468, P1_P3_INSTADDRPOINTER_REG_12_ );
nor U129214 ( n33344, n33346, n33347 );
nor U129215 ( n33347, n74801, n76898 );
xnor U129216 ( n66472, n67368, P2_P3_INSTADDRPOINTER_REG_31_ );
nand U129217 ( n67368, n66524, P2_P3_INSTADDRPOINTER_REG_30_ );
xnor U129218 ( n24635, n25363, P1_P2_INSTADDRPOINTER_REG_31_ );
nand U129219 ( n25363, n24689, P1_P2_INSTADDRPOINTER_REG_30_ );
xnor U129220 ( n57767, n58500, P2_P2_INSTADDRPOINTER_REG_31_ );
nand U129221 ( n58500, n57823, P2_P2_INSTADDRPOINTER_REG_30_ );
nor U129222 ( n37748, n37784, n37690 );
xnor U129223 ( n37784, n37785, n37786 );
xor U129224 ( n37785, n37783, P4_REG2_REG_4_ );
nor U129225 ( n37714, n37722, n37690 );
xnor U129226 ( n37722, n37723, n37724 );
xor U129227 ( n37723, n37721, P4_REG2_REG_2_ );
nand U129228 ( n15601, n46982, n46983 );
nand U129229 ( n46983, n76860, P2_P1_INSTADDRPOINTER_REG_14_ );
nor U129230 ( n46982, n46984, n46985 );
nor U129231 ( n46985, n74860, n76333 );
nand U129232 ( n11111, n68017, n68018 );
nand U129233 ( n68018, n76195, P2_P3_INSTADDRPOINTER_REG_14_ );
nor U129234 ( n68017, n68019, n68020 );
nor U129235 ( n68020, n74830, n76872 );
nand U129236 ( n6621, n26014, n26015 );
nand U129237 ( n26015, n76519, P1_P2_INSTADDRPOINTER_REG_14_ );
nor U129238 ( n26014, n26016, n26017 );
nor U129239 ( n26017, n74828, n76907 );
nand U129240 ( n13356, n59155, n59156 );
nand U129241 ( n59156, n76261, P2_P2_INSTADDRPOINTER_REG_14_ );
nor U129242 ( n59155, n59157, n59158 );
nor U129243 ( n59158, n74827, n76881 );
nand U129244 ( n47178, P2_P1_INSTADDRPOINTER_REG_8_, n47189 );
xor U129245 ( n45533, n46324, n75052 );
nand U129246 ( n46324, P2_P1_INSTADDRPOINTER_REG_30_, n45596 );
nand U129247 ( n47299, n47346, n47347 );
or U129248 ( n47346, n47350, n47349 );
nand U129249 ( n47347, P2_P1_INSTADDRPOINTER_REG_5_, n47348 );
nand U129250 ( n47348, n47349, n47350 );
nand U129251 ( n47189, n47249, n47250 );
nand U129252 ( n47249, n7564, n47252 );
nand U129253 ( n47250, P2_P1_INSTADDRPOINTER_REG_7_, n47251 );
or U129254 ( n47251, n47252, n7564 );
nand U129255 ( n37353, n38751, n38752 );
nand U129256 ( n38752, P4_REG0_REG_31_, n76418 );
nor U129257 ( n38751, n38754, n38755 );
nor U129258 ( n38754, n76410, n74773 );
nor U129259 ( n38755, n76416, n74771 );
nand U129260 ( n4381, n33223, n33224 );
nand U129261 ( n33224, n76468, P1_P3_INSTADDRPOINTER_REG_15_ );
nor U129262 ( n33223, n33225, n33226 );
nor U129263 ( n33226, n74839, n76898 );
xor U129264 ( n31877, n31901, P1_P3_INSTADDRPOINTER_REG_30_ );
and U129265 ( n32325, n33314, n33315 );
nand U129266 ( n33314, n33323, n33324 );
nand U129267 ( n33315, n33316, n33317 );
nand U129268 ( n33324, P1_P3_INSTADDRPOINTER_REG_13_, n76472 );
nand U129269 ( n4371, n33303, n33304 );
nand U129270 ( n33304, n76468, P1_P3_INSTADDRPOINTER_REG_13_ );
nor U129271 ( n33303, n33305, n33306 );
nor U129272 ( n33306, n73235, n76898 );
xor U129273 ( n24663, n24689, P1_P2_INSTADDRPOINTER_REG_30_ );
xor U129274 ( n57799, n57823, P2_P2_INSTADDRPOINTER_REG_30_ );
xor U129275 ( n66500, n66524, P2_P3_INSTADDRPOINTER_REG_30_ );
nand U129276 ( n50857, n50007, P3_DATAO_REG_3_ );
nand U129277 ( n18174, n8218, P4_DATAO_REG_2_ );
and U129278 ( n50007, DIN_24_, n76929 );
nand U129279 ( n17969, n8214, P4_DATAO_REG_5_ );
nand U129280 ( n50657, n50007, P3_DATAO_REG_4_ );
nand U129281 ( n33796, n33941, n33942 );
nand U129282 ( n33941, n33945, n33944 );
nand U129283 ( n33942, P1_P3_INSTADDRPOINTER_REG_1_, n33943 );
or U129284 ( n33943, n33944, n33945 );
nand U129285 ( n26551, n26696, n26697 );
nand U129286 ( n26696, n26700, n26699 );
nand U129287 ( n26697, P1_P2_INSTADDRPOINTER_REG_1_, n26698 );
or U129288 ( n26698, n26699, n26700 );
nand U129289 ( n59693, n59838, n59839 );
nand U129290 ( n59838, n59842, n59841 );
nand U129291 ( n59839, P2_P2_INSTADDRPOINTER_REG_1_, n59840 );
or U129292 ( n59840, n59841, n59842 );
nand U129293 ( n68552, n68697, n68698 );
nand U129294 ( n68697, n68701, n68700 );
nand U129295 ( n68698, P2_P3_INSTADDRPOINTER_REG_1_, n68699 );
or U129296 ( n68699, n68700, n68701 );
nand U129297 ( n37855, n39988, n39989 );
nand U129298 ( n39988, P4_IR_REG_9_, n76794 );
or U129299 ( n39989, n39990, n76793 );
nand U129300 ( n50381, n50007, P3_DATAO_REG_5_ );
nand U129301 ( n17715, n8214, P4_DATAO_REG_6_ );
nand U129302 ( n37841, n40032, n40033 );
nand U129303 ( n40033, n40034, P4_IR_REG_31_ );
nand U129304 ( n40032, P4_IR_REG_8_, n76794 );
and U129305 ( n40034, n40035, n40036 );
xor U129306 ( n45574, n45596, P2_P1_INSTADDRPOINTER_REG_30_ );
nor U129307 ( n33794, P1_P3_INSTADDRPOINTER_REG_3_, n33790 );
nor U129308 ( n68550, P2_P3_INSTADDRPOINTER_REG_3_, n68546 );
nor U129309 ( n26549, P1_P2_INSTADDRPOINTER_REG_3_, n26545 );
nor U129310 ( n59691, P2_P2_INSTADDRPOINTER_REG_3_, n59687 );
nand U129311 ( n45404, n49538, n49539 );
nand U129312 ( n49538, P2_BUF1_REG_3_, n76478 );
nand U129313 ( n49539, n49540, n76476 );
xor U129314 ( n49540, n49541, n49542 );
nand U129315 ( n18892, n8218, P4_DATAO_REG_1_ );
nand U129316 ( n49393, n49394, n49395 );
nand U129317 ( n49395, P2_P1_INSTQUEUE_REG_14__3_, n49353 );
nand U129318 ( n49394, n7440, n264 );
nand U129319 ( n49300, n49301, n49302 );
nand U129320 ( n49302, P2_P1_INSTQUEUE_REG_13__3_, n49275 );
nand U129321 ( n49301, n7442, n264 );
nand U129322 ( n49109, n49110, n49111 );
nand U129323 ( n49111, P2_P1_INSTQUEUE_REG_11__3_, n49085 );
nand U129324 ( n49110, n7443, n264 );
nand U129325 ( n49015, n49016, n49017 );
nand U129326 ( n49017, P2_P1_INSTQUEUE_REG_10__3_, n48990 );
nand U129327 ( n49016, n7444, n264 );
nand U129328 ( n48932, n48933, n48934 );
nand U129329 ( n48934, P2_P1_INSTQUEUE_REG_9__3_, n48891 );
nand U129330 ( n48933, n7445, n264 );
nand U129331 ( n48649, n48650, n48651 );
nand U129332 ( n48651, P2_P1_INSTQUEUE_REG_6__3_, n48624 );
nand U129333 ( n48650, n7448, n264 );
nand U129334 ( n48555, n48556, n48557 );
nand U129335 ( n48557, P2_P1_INSTQUEUE_REG_5__3_, n48530 );
nand U129336 ( n48556, n7449, n264 );
nand U129337 ( n48742, n48743, n48744 );
nand U129338 ( n48744, P2_P1_INSTQUEUE_REG_7__3_, n48718 );
nand U129339 ( n48743, n7447, n264 );
and U129340 ( n38971, n76418, P4_REG0_REG_27_ );
nand U129341 ( n37872, n39952, n39953 );
nand U129342 ( n39953, n39954, P4_IR_REG_31_ );
nand U129343 ( n39952, P4_IR_REG_10_, n76794 );
and U129344 ( n39954, n39955, n39956 );
nor U129345 ( n38777, n2193, n38794 );
nor U129346 ( n38794, n38795, n38796 );
nor U129347 ( n38795, P4_B_REG, n38604 );
nor U129348 ( n38796, n76457, n36264 );
nand U129349 ( n31940, n74973, n32760 );
nand U129350 ( n32760, n32009, P1_P3_INSTADDRPOINTER_REG_27_ );
and U129351 ( n38912, n76418, P4_REG0_REG_28_ );
and U129352 ( n62248, n76252, P3_REG0_REG_28_ );
nand U129353 ( n66543, n74976, n67525 );
nand U129354 ( n67525, n66612, P2_P3_INSTADDRPOINTER_REG_27_ );
nand U129355 ( n24708, n74975, n25520 );
nand U129356 ( n25520, n24777, P1_P2_INSTADDRPOINTER_REG_27_ );
nand U129357 ( n57842, n74977, n58657 );
nand U129358 ( n58657, n57911, P2_P2_INSTADDRPOINTER_REG_27_ );
and U129359 ( n16538, n17036, P4_DATAO_REG_0_ );
and U129360 ( n38846, n76418, P4_REG0_REG_29_ );
nand U129361 ( n50873, n50007, P3_DATAO_REG_2_ );
nand U129362 ( n16269, P3_IR_REG_4_, n66377 );
nand U129363 ( n66377, n909, n73797 );
nand U129364 ( n13784, n13802, n13803 );
or U129365 ( n13802, n13807, n13805 );
nand U129366 ( n13803, P1_P1_INSTADDRPOINTER_REG_8_, n13804 );
nand U129367 ( n13804, n13805, n13807 );
nand U129368 ( n14304, P1_P1_INSTADDRPOINTER_REG_2_, n14400 );
nor U129369 ( n13970, n13974, n13975 );
nor U129370 ( n13974, P1_P1_INSTADDRPOINTER_REG_5_, n13969 );
or U129371 ( n13975, n4940, n13977 );
and U129372 ( n13805, n13858, n13859 );
or U129373 ( n13858, n13863, n13862 );
nand U129374 ( n13859, P1_P1_INSTADDRPOINTER_REG_7_, n13860 );
nand U129375 ( n13860, n13862, n13863 );
and U129376 ( n13862, n13917, n13918 );
or U129377 ( n13917, n13922, n13920 );
nand U129378 ( n13918, P1_P1_INSTADDRPOINTER_REG_6_, n13919 );
nand U129379 ( n13919, n13920, n13922 );
xor U129380 ( n11820, n12749, n74989 );
nand U129381 ( n12749, n4882, P1_P1_INSTADDRPOINTER_REG_29_ );
nand U129382 ( n43230, n65952, n65953 );
nand U129383 ( n65952, P3_IR_REG_9_, n76840 );
or U129384 ( n65953, n15619, n76839 );
nand U129385 ( n41510, n61289, n61290 );
nand U129386 ( n61290, P3_REG0_REG_31_, n76252 );
nor U129387 ( n61289, n61292, n61293 );
nor U129388 ( n61292, n76244, n74846 );
nor U129389 ( n61293, n76250, n74844 );
and U129390 ( n55000, n67259, n67260 );
nand U129391 ( n67260, n9650, n67261 );
nand U129392 ( n67259, n619, P3_D_REG_1_ );
nand U129393 ( n50017, n50007, P3_DATAO_REG_6_ );
nand U129394 ( n43559, n65357, n65358 );
nand U129395 ( n65357, P3_IR_REG_11_, n76840 );
or U129396 ( n65358, n15348, n76839 );
xor U129397 ( n37970, n37971, n37972 );
xor U129398 ( n37972, n37969, P4_REG2_REG_17_ );
nand U129399 ( n41948, n61416, n61417 );
nand U129400 ( n61417, P3_REG0_REG_30_, n76252 );
nor U129401 ( n61416, n61418, n61419 );
nor U129402 ( n61418, n76244, n74867 );
nor U129403 ( n61419, n76250, n74866 );
xor U129404 ( n45664, n45688, P2_P1_INSTADDRPOINTER_REG_27_ );
nor U129405 ( n14300, n14400, P1_P1_INSTADDRPOINTER_REG_2_ );
nor U129406 ( n62303, n76250, n74824 );
nand U129407 ( n11919, n12910, n12912 );
nand U129408 ( n12912, P1_P1_INSTADDRPOINTER_REG_27_, n4881 );
nor U129409 ( n12910, n12913, n12914 );
nor U129410 ( n12914, n4881, n12915 );
nand U129411 ( n4376, n33258, n33259 );
nand U129412 ( n33259, n76468, P1_P3_INSTADDRPOINTER_REG_14_ );
nor U129413 ( n33258, n33260, n33261 );
nor U129414 ( n33261, n74829, n76898 );
xor U129415 ( n50003, n50004, n50005 );
nand U129416 ( n50004, n50006, P3_DATAO_REG_9_ );
nand U129417 ( n50005, n8235, P3_DATAO_REG_10_ );
nor U129418 ( n47343, n47521, P2_P1_INSTADDRPOINTER_REG_4_ );
nor U129419 ( n45689, P2_P1_INSTADDRPOINTER_REG_26_, n46540 );
nor U129420 ( n61395, n780, n61413 );
nor U129421 ( n61413, n61414, n61415 );
nor U129422 ( n61414, P3_B_REG, n76062 );
nor U129423 ( n61415, n76389, n40664 );
nand U129424 ( n45615, n74974, n46464 );
nand U129425 ( n46464, n45685, P2_P1_INSTADDRPOINTER_REG_27_ );
nor U129426 ( n61597, n76250, n74863 );
nand U129427 ( n33458, P1_P3_INSTADDRPOINTER_REG_8_, n33469 );
nand U129428 ( n33574, n33622, n33623 );
or U129429 ( n33622, n33626, n33625 );
nand U129430 ( n33623, P1_P3_INSTADDRPOINTER_REG_5_, n33624 );
nand U129431 ( n33624, n33625, n33626 );
nand U129432 ( n33469, n33524, n33525 );
nand U129433 ( n33524, n3178, n33527 );
nand U129434 ( n33525, P1_P3_INSTADDRPOINTER_REG_7_, n33526 );
or U129435 ( n33526, n33527, n3178 );
xor U129436 ( n11853, n4882, P1_P1_INSTADDRPOINTER_REG_29_ );
nand U129437 ( n68209, P2_P3_INSTADDRPOINTER_REG_8_, n68220 );
nand U129438 ( n26208, P1_P2_INSTADDRPOINTER_REG_8_, n26219 );
nand U129439 ( n59347, P2_P2_INSTADDRPOINTER_REG_8_, n59358 );
nand U129440 ( n68330, n68378, n68379 );
or U129441 ( n68378, n68382, n68381 );
nand U129442 ( n68379, P2_P3_INSTADDRPOINTER_REG_5_, n68380 );
nand U129443 ( n68380, n68381, n68382 );
nand U129444 ( n26329, n26377, n26378 );
or U129445 ( n26377, n26381, n26380 );
nand U129446 ( n26378, P1_P2_INSTADDRPOINTER_REG_5_, n26379 );
nand U129447 ( n26379, n26380, n26381 );
nand U129448 ( n59468, n59516, n59517 );
or U129449 ( n59516, n59520, n59519 );
nand U129450 ( n59517, P2_P2_INSTADDRPOINTER_REG_5_, n59518 );
nand U129451 ( n59518, n59519, n59520 );
nand U129452 ( n68220, n68280, n68281 );
nand U129453 ( n68280, n5777, n68283 );
nand U129454 ( n68281, P2_P3_INSTADDRPOINTER_REG_7_, n68282 );
or U129455 ( n68282, n68283, n5777 );
nand U129456 ( n26219, n26279, n26280 );
nand U129457 ( n26279, n4018, n26282 );
nand U129458 ( n26280, P1_P2_INSTADDRPOINTER_REG_7_, n26281 );
or U129459 ( n26281, n26282, n4018 );
nand U129460 ( n59358, n59418, n59419 );
nand U129461 ( n59418, n6650, n59421 );
nand U129462 ( n59419, P2_P2_INSTADDRPOINTER_REG_7_, n59420 );
or U129463 ( n59420, n59421, n6650 );
nand U129464 ( n37788, P4_ADDR_REG_4_, n2080 );
nor U129465 ( n72074, n74342, n71104 );
nand U129466 ( n14204, n14403, n14404 );
nand U129467 ( n14403, n14408, n14407 );
nand U129468 ( n14404, P1_P1_INSTADDRPOINTER_REG_1_, n14405 );
or U129469 ( n14405, n14407, n14408 );
xor U129470 ( n46057, n47120, n7539 );
xor U129471 ( n47120, n76342, P2_P1_INSTADDRPOINTER_REG_11_ );
nand U129472 ( n15586, n47109, n47110 );
nand U129473 ( n47110, n76860, P2_P1_INSTADDRPOINTER_REG_11_ );
nor U129474 ( n47109, n47111, n47112 );
nor U129475 ( n47112, n74811, n76332 );
xor U129476 ( n67021, n68151, n5753 );
xor U129477 ( n68151, n76198, P2_P3_INSTADDRPOINTER_REG_11_ );
xor U129478 ( n25121, n26150, n3995 );
xor U129479 ( n26150, n76522, P1_P2_INSTADDRPOINTER_REG_11_ );
xor U129480 ( n58259, n59289, n6628 );
xor U129481 ( n59289, n76264, P2_P2_INSTADDRPOINTER_REG_11_ );
nand U129482 ( n11096, n68140, n68141 );
nand U129483 ( n68141, n76195, P2_P3_INSTADDRPOINTER_REG_11_ );
nor U129484 ( n68140, n68142, n68143 );
nor U129485 ( n68143, n74790, n76871 );
nand U129486 ( n6606, n26139, n26140 );
nand U129487 ( n26140, n76519, P1_P2_INSTADDRPOINTER_REG_11_ );
nor U129488 ( n26139, n26141, n26142 );
nor U129489 ( n26142, n74789, n76906 );
nand U129490 ( n13341, n59278, n59279 );
nand U129491 ( n59279, n76261, P2_P2_INSTADDRPOINTER_REG_11_ );
nor U129492 ( n59278, n59280, n59281 );
nor U129493 ( n59281, n74788, n76880 );
nand U129494 ( n50331, DIN_25_, n76929 );
nand U129495 ( n37299, n38797, n38798 );
nand U129496 ( n38798, P4_REG0_REG_30_, n76418 );
nor U129497 ( n38797, n38799, n38800 );
nor U129498 ( n38799, n76410, n74826 );
nor U129499 ( n38800, n76416, n74825 );
nand U129500 ( n9246, n11529, n11530 );
nand U129501 ( n11530, P1_P1_UWORD_REG_4_, n76618 );
nor U129502 ( n11529, n11532, n11533 );
nor U129503 ( n11532, n74966, n76617 );
nand U129504 ( n9171, n11612, n11613 );
nand U129505 ( n11613, P1_P1_LWORD_REG_4_, n11504 );
nor U129506 ( n11612, n11614, n11533 );
nor U129507 ( n11614, n74682, n76615 );
nand U129508 ( n45243, n65829, n65830 );
nand U129509 ( n65830, n65831, P3_IR_REG_31_ );
nand U129510 ( n65829, P3_IR_REG_10_, n76840 );
and U129511 ( n65831, n15482, n15480 );
and U129512 ( n62304, n76252, P3_REG0_REG_27_ );
nand U129513 ( n17440, DIN_23_, n76928 );
nand U129514 ( n18189, n8213, P4_DATAO_REG_3_ );
nand U129515 ( n12198, n12210, n12212 );
nand U129516 ( n12210, n12225, n12227 );
nand U129517 ( n12212, n12213, n12214 );
nor U129518 ( n12227, P1_P1_PHYADDRPOINTER_REG_17_, n12187 );
nand U129519 ( n17444, n8214, P4_DATAO_REG_7_ );
nand U129520 ( n42957, n66038, n66039 );
nand U129521 ( n66039, n66040, P3_IR_REG_31_ );
nand U129522 ( n66038, P3_IR_REG_8_, n76841 );
and U129523 ( n66040, n15745, n15744 );
xor U129524 ( n31876, n31898, P1_P3_INSTADDRPOINTER_REG_30_ );
xor U129525 ( n24662, n24686, P1_P2_INSTADDRPOINTER_REG_30_ );
xor U129526 ( n57798, n57820, P2_P2_INSTADDRPOINTER_REG_30_ );
xor U129527 ( n66499, n66521, P2_P3_INSTADDRPOINTER_REG_30_ );
and U129528 ( n49655, n50006, P3_DATAO_REG_0_ );
nor U129529 ( n14202, P1_P1_INSTADDRPOINTER_REG_3_, n14197 );
nand U129530 ( n37883, n39911, n39912 );
nand U129531 ( n39911, P4_IR_REG_11_, n76795 );
or U129532 ( n39912, n39913, n76793 );
and U129533 ( n37710, n2080, P4_ADDR_REG_1_ );
and U129534 ( n37695, n2080, P4_ADDR_REG_0_ );
nand U129535 ( n40142, P4_REG3_REG_4_, P4_REG3_REG_3_ );
nand U129536 ( n61073, n67317, n67318 );
nand U129537 ( n67318, n9768, n67261 );
nand U129538 ( n67317, n619, P3_D_REG_0_ );
nand U129539 ( n17941, n8214, P4_DATAO_REG_2_ );
xnor U129540 ( n32358, n33399, n33400 );
xor U129541 ( n33400, n74755, n76470 );
nand U129542 ( n33399, n33401, n33402 );
nand U129543 ( n33402, P1_P3_INSTADDRPOINTER_REG_10_, n76472 );
nor U129544 ( n33401, n3158, n33403 );
not U129545 ( n3158, n33405 );
nor U129546 ( n33403, n33404, n33299 );
nor U129547 ( n33404, P1_P3_INSTADDRPOINTER_REG_10_, n76470 );
nand U129548 ( n4361, n33388, n33389 );
nand U129549 ( n33389, n76468, P1_P3_INSTADDRPOINTER_REG_11_ );
nor U129550 ( n33388, n33390, n33391 );
nor U129551 ( n33391, n74791, n76897 );
and U129552 ( n61598, n76252, P3_REG0_REG_29_ );
xor U129553 ( n31985, n32009, P1_P3_INSTADDRPOINTER_REG_27_ );
nand U129554 ( n39956, P4_IR_REG_10_, n40604 );
nand U129555 ( n40604, n2205, n74298 );
xor U129556 ( n24753, n24777, P1_P2_INSTADDRPOINTER_REG_27_ );
xor U129557 ( n66588, n66612, P2_P3_INSTADDRPOINTER_REG_27_ );
xor U129558 ( n57887, n57911, P2_P2_INSTADDRPOINTER_REG_27_ );
nand U129559 ( n50652, n8240, P3_DATAO_REG_2_ );
xor U129560 ( n38527, n40142, P4_REG3_REG_5_ );
nand U129561 ( n13788, P1_P1_INSTADDRPOINTER_REG_8_, n13817 );
nand U129562 ( n13817, n13867, n13868 );
nand U129563 ( n13867, n4914, n13870 );
nand U129564 ( n13868, P1_P1_INSTADDRPOINTER_REG_7_, n13869 );
or U129565 ( n13869, n13870, n4914 );
nand U129566 ( n11918, n12919, n12920 );
nand U129567 ( n12920, P1_P1_INSTADDRPOINTER_REG_27_, n4907 );
nor U129568 ( n12919, n12913, n12922 );
nor U129569 ( n12922, n4907, n12915 );
nand U129570 ( n13929, n13988, n13989 );
or U129571 ( n13988, n13993, n13992 );
nand U129572 ( n13989, P1_P1_INSTADDRPOINTER_REG_5_, n13990 );
nand U129573 ( n13990, n13992, n13993 );
xor U129574 ( n31834, n32623, n75065 );
nand U129575 ( n32623, P1_P3_INSTADDRPOINTER_REG_30_, n31898 );
xor U129576 ( n24620, n25383, n75066 );
nand U129577 ( n25383, P1_P2_INSTADDRPOINTER_REG_30_, n24686 );
xor U129578 ( n57752, n58520, n75067 );
nand U129579 ( n58520, P2_P2_INSTADDRPOINTER_REG_30_, n57820 );
xor U129580 ( n66457, n67388, n75068 );
nand U129581 ( n67388, P2_P3_INSTADDRPOINTER_REG_30_, n66521 );
xor U129582 ( n12247, n4892, n13465 );
nor U129583 ( n13465, n13467, n13417 );
nor U129584 ( n13467, P1_P1_INSTADDRPOINTER_REG_16_, n76602 );
nand U129585 ( n8876, n13452, n13453 );
nand U129586 ( n13453, n76887, P1_P1_INSTADDRPOINTER_REG_16_ );
nor U129587 ( n13452, n13454, n13455 );
nor U129588 ( n13455, n73254, n76599 );
nand U129589 ( n16000, P3_IR_REG_6_, n66225 );
nand U129590 ( n66225, n899, n74105 );
nand U129591 ( n37941, n39681, n39682 );
nand U129592 ( n39681, P4_IR_REG_15_, n76795 );
or U129593 ( n39682, n39683, n76793 );
nor U129594 ( n33619, n33786, P1_P3_INSTADDRPOINTER_REG_4_ );
nor U129595 ( n26374, n26541, P1_P2_INSTADDRPOINTER_REG_4_ );
nor U129596 ( n59513, n59683, P2_P2_INSTADDRPOINTER_REG_4_ );
nor U129597 ( n68375, n68542, P2_P3_INSTADDRPOINTER_REG_4_ );
nand U129598 ( n50375, n8240, P3_DATAO_REG_3_ );
nand U129599 ( n15480, P3_IR_REG_10_, n65832 );
nand U129600 ( n65832, n883, n74300 );
xor U129601 ( n11953, n12859, P1_P1_INSTADDRPOINTER_REG_26_ );
xor U129602 ( n11819, n12748, n74989 );
nand U129603 ( n12748, n4908, P1_P1_INSTADDRPOINTER_REG_29_ );
nand U129604 ( n31937, n74973, n32762 );
nand U129605 ( n32762, n32006, P1_P3_INSTADDRPOINTER_REG_27_ );
xor U129606 ( n45663, n45685, P2_P1_INSTADDRPOINTER_REG_27_ );
nand U129607 ( n15986, n45337, n45338 );
nand U129608 ( n45338, P2_P1_UWORD_REG_3_, n76352 );
nor U129609 ( n45337, n45339, n45340 );
nor U129610 ( n45339, n74953, n76351 );
nand U129611 ( n15911, n45401, n45402 );
nand U129612 ( n45402, P2_P1_LWORD_REG_3_, n45325 );
nor U129613 ( n45401, n45403, n45340 );
nor U129614 ( n45403, n74631, n76350 );
nand U129615 ( n24705, n74975, n25522 );
nand U129616 ( n25522, n24774, P1_P2_INSTADDRPOINTER_REG_27_ );
nand U129617 ( n66540, n74976, n67527 );
nand U129618 ( n67527, n66609, P2_P3_INSTADDRPOINTER_REG_27_ );
nand U129619 ( n57839, n74977, n58659 );
nand U129620 ( n58659, n57908, P2_P2_INSTADDRPOINTER_REG_27_ );
nand U129621 ( n32025, n73232, n32883 );
nand U129622 ( n32883, n32882, P1_P3_INSTADDRPOINTER_REG_24_ );
nand U129623 ( n66628, n73223, n67644 );
nand U129624 ( n67644, n67643, P2_P3_INSTADDRPOINTER_REG_24_ );
nand U129625 ( n24793, n73224, n25639 );
nand U129626 ( n25639, n25638, P1_P2_INSTADDRPOINTER_REG_24_ );
nand U129627 ( n57927, n73225, n58776 );
nand U129628 ( n58776, n58775, P2_P2_INSTADDRPOINTER_REG_24_ );
nand U129629 ( n11610, n16558, n16559 );
nand U129630 ( n16558, P1_BUF1_REG_3_, n76610 );
nand U129631 ( n16559, n16560, n76613 );
xor U129632 ( n16560, n16562, n16563 );
nand U129633 ( n16372, n16373, n16374 );
nand U129634 ( n16374, P1_P1_INSTQUEUE_REG_14__3_, n16340 );
nand U129635 ( n16373, n4797, n16 );
nand U129636 ( n16275, n16277, n16278 );
nand U129637 ( n16278, P1_P1_INSTQUEUE_REG_13__3_, n16235 );
nand U129638 ( n16277, n4798, n16 );
nand U129639 ( n16064, n16065, n16067 );
nand U129640 ( n16067, P1_P1_INSTQUEUE_REG_11__3_, n16033 );
nand U129641 ( n16065, n4799, n16 );
nand U129642 ( n15957, n15958, n15959 );
nand U129643 ( n15959, P1_P1_INSTQUEUE_REG_10__3_, n15925 );
nand U129644 ( n15958, n4800, n16 );
nand U129645 ( n15852, n15853, n15854 );
nand U129646 ( n15854, P1_P1_INSTQUEUE_REG_9__3_, n15820 );
nand U129647 ( n15853, n4802, n16 );
nand U129648 ( n15543, n15544, n15545 );
nand U129649 ( n15545, P1_P1_INSTQUEUE_REG_6__3_, n15512 );
nand U129650 ( n15544, n4804, n16 );
nand U129651 ( n15437, n15438, n15439 );
nand U129652 ( n15439, P1_P1_INSTQUEUE_REG_5__3_, n15405 );
nand U129653 ( n15438, n4805, n16 );
nand U129654 ( n15644, n15645, n15647 );
nand U129655 ( n15647, P1_P1_INSTQUEUE_REG_7__3_, n15609 );
nand U129656 ( n15645, n4803, n16 );
nand U129657 ( n45703, n73220, n46596 );
nand U129658 ( n46596, n46597, P2_P1_INSTADDRPOINTER_REG_24_ );
nand U129659 ( n11974, n74774, n13058 );
nand U129660 ( n13058, n13059, P1_P1_INSTADDRPOINTER_REG_24_ );
nand U129661 ( n42313, P3_ADDR_REG_4_, n42201 );
nand U129662 ( n40036, P4_IR_REG_8_, n40615 );
nand U129663 ( n40615, n2207, n74257 );
nand U129664 ( n37913, n39806, n39807 );
nand U129665 ( n39806, P4_IR_REG_13_, n76794 );
or U129666 ( n39807, n39808, n76793 );
and U129667 ( n50628, n50007, P3_DATAO_REG_1_ );
nand U129668 ( n37955, n39623, n39624 );
nand U129669 ( n39623, P4_IR_REG_16_, n76794 );
nand U129670 ( n39624, n39625, P4_IR_REG_31_ );
and U129671 ( n39625, n39626, n39627 );
xor U129672 ( n11852, P1_P1_INSTADDRPOINTER_REG_29_, n4908 );
nand U129673 ( n45400, n49509, n49510 );
nand U129674 ( n49509, P2_BUF1_REG_2_, n76478 );
nand U129675 ( n49510, n49511, n76476 );
xor U129676 ( n49511, n49512, n49513 );
nand U129677 ( n49385, n49386, n49387 );
nand U129678 ( n49387, P2_P1_INSTQUEUE_REG_14__2_, n49353 );
nand U129679 ( n49386, n7440, n258 );
nand U129680 ( n49292, n49293, n49294 );
nand U129681 ( n49294, P2_P1_INSTQUEUE_REG_13__2_, n49275 );
nand U129682 ( n49293, n7442, n258 );
nand U129683 ( n49101, n49102, n49103 );
nand U129684 ( n49103, P2_P1_INSTQUEUE_REG_11__2_, n49085 );
nand U129685 ( n49102, n7443, n258 );
nand U129686 ( n49007, n49008, n49009 );
nand U129687 ( n49009, P2_P1_INSTQUEUE_REG_10__2_, n48990 );
nand U129688 ( n49008, n7444, n258 );
nand U129689 ( n48924, n48925, n48926 );
nand U129690 ( n48926, P2_P1_INSTQUEUE_REG_9__2_, n48891 );
nand U129691 ( n48925, n7445, n258 );
nand U129692 ( n48641, n48642, n48643 );
nand U129693 ( n48643, P2_P1_INSTQUEUE_REG_6__2_, n48624 );
nand U129694 ( n48642, n7448, n258 );
nand U129695 ( n48547, n48548, n48549 );
nand U129696 ( n48549, P2_P1_INSTQUEUE_REG_5__2_, n48530 );
nand U129697 ( n48548, n7449, n258 );
nand U129698 ( n48734, n48735, n48736 );
nand U129699 ( n48736, P2_P1_INSTQUEUE_REG_7__2_, n48718 );
nand U129700 ( n48735, n7447, n258 );
nor U129701 ( n45686, P2_P1_INSTADDRPOINTER_REG_26_, n46542 );
and U129702 ( n42218, n42201, P3_ADDR_REG_1_ );
and U129703 ( n42199, n42201, P3_ADDR_REG_0_ );
nand U129704 ( n37897, n39853, n39854 );
nand U129705 ( n39854, n39855, P4_IR_REG_31_ );
nand U129706 ( n39853, P4_IR_REG_12_, n76794 );
and U129707 ( n39855, n39856, n39857 );
xnor U129708 ( n46079, n47155, n47156 );
xor U129709 ( n47155, n76342, P2_P1_INSTADDRPOINTER_REG_10_ );
nor U129710 ( n47156, n7543, n47121 );
not U129711 ( n7543, n47124 );
nand U129712 ( n15581, n47140, n47141 );
nand U129713 ( n47141, n76860, P2_P1_INSTADDRPOINTER_REG_10_ );
nor U129714 ( n47140, n47142, n47143 );
nor U129715 ( n47143, n74769, n76332 );
xnor U129716 ( n67043, n68186, n68187 );
xor U129717 ( n68186, n76198, P2_P3_INSTADDRPOINTER_REG_10_ );
nor U129718 ( n68187, n5757, n68152 );
not U129719 ( n5757, n68155 );
xnor U129720 ( n25143, n26185, n26186 );
xor U129721 ( n26185, n76522, P1_P2_INSTADDRPOINTER_REG_10_ );
nor U129722 ( n26186, n3999, n26151 );
not U129723 ( n3999, n26154 );
xnor U129724 ( n58281, n59324, n59325 );
xor U129725 ( n59324, n76264, P2_P2_INSTADDRPOINTER_REG_10_ );
nor U129726 ( n59325, n6632, n59290 );
not U129727 ( n6632, n59293 );
nand U129728 ( n11091, n68171, n68172 );
nand U129729 ( n68172, n76195, P2_P3_INSTADDRPOINTER_REG_10_ );
nor U129730 ( n68171, n68173, n68174 );
nor U129731 ( n68174, n74745, n76871 );
nand U129732 ( n6601, n26170, n26171 );
nand U129733 ( n26171, n76519, P1_P2_INSTADDRPOINTER_REG_10_ );
nor U129734 ( n26170, n26172, n26173 );
nor U129735 ( n26173, n74744, n76906 );
nand U129736 ( n13336, n59309, n59310 );
nand U129737 ( n59310, n76261, P2_P2_INSTADDRPOINTER_REG_10_ );
nor U129738 ( n59309, n59311, n59312 );
nor U129739 ( n59312, n74743, n76880 );
nand U129740 ( n39627, P4_IR_REG_16_, n40571 );
nand U129741 ( n40571, n2202, n74391 );
nand U129742 ( n4356, n33424, n33425 );
nand U129743 ( n33425, n76468, P1_P3_INSTADDRPOINTER_REG_10_ );
nor U129744 ( n33424, n33426, n33427 );
nor U129745 ( n33427, n74746, n76897 );
nand U129746 ( n40049, n40095, P4_REG3_REG_6_ );
nand U129747 ( n39970, n40004, P4_REG3_REG_8_ );
nand U129748 ( n39857, P4_IR_REG_12_, n40593 );
nand U129749 ( n40593, n2204, n74335 );
xnor U129750 ( n36654, n74062, P4_REG3_REG_3_ );
nand U129751 ( n17928, n8214, P4_DATAO_REG_1_ );
nand U129752 ( n50031, DIN_26_, n76929 );
nand U129753 ( n13087, P1_P1_INSTADDRPOINTER_REG_23_, n76606 );
nor U129754 ( n13977, n14192, P1_P1_INSTADDRPOINTER_REG_4_ );
nor U129755 ( n72067, n74388, n71104 );
xor U129756 ( n49259, n65323, P3_REG3_REG_11_ );
nand U129757 ( n66278, P3_REG3_REG_4_, P3_REG3_REG_3_ );
nand U129758 ( n66096, n66185, P3_REG3_REG_6_ );
nand U129759 ( n65930, n66010, P3_REG3_REG_8_ );
nand U129760 ( n65323, P3_REG3_REG_10_, n65806 );
nand U129761 ( n13613, n13682, n13683 );
nand U129762 ( n13682, P1_P1_INSTADDRPOINTER_REG_11_, n76606 );
nand U129763 ( n13683, n13588, n13525 );
and U129764 ( n12344, n13605, n13607 );
nand U129765 ( n13605, n13617, n13618 );
nand U129766 ( n13607, n13608, n13609 );
nand U129767 ( n13618, P1_P1_INSTADDRPOINTER_REG_13_, n76606 );
nand U129768 ( n8861, n13594, n13595 );
nand U129769 ( n13595, n76887, P1_P1_INSTADDRPOINTER_REG_13_ );
nor U129770 ( n13594, n13597, n13598 );
nor U129771 ( n13598, n73240, n76599 );
xor U129772 ( n31984, n32006, P1_P3_INSTADDRPOINTER_REG_27_ );
nor U129773 ( n13678, P1_P1_INSTADDRPOINTER_REG_12_, n13679 );
xor U129774 ( n13679, n13613, n76603 );
nand U129775 ( n8856, n13653, n13654 );
nand U129776 ( n13654, n76887, P1_P1_INSTADDRPOINTER_REG_12_ );
nor U129777 ( n13653, n13655, n13657 );
nor U129778 ( n13657, n74816, n76599 );
xor U129779 ( n24752, n24774, P1_P2_INSTADDRPOINTER_REG_27_ );
xor U129780 ( n66587, n66609, P2_P3_INSTADDRPOINTER_REG_27_ );
xor U129781 ( n57886, n57908, P2_P2_INSTADDRPOINTER_REG_27_ );
nand U129782 ( n15744, P3_IR_REG_8_, n66041 );
nand U129783 ( n66041, n889, n74225 );
nand U129784 ( n45699, n45700, n45701 );
nand U129785 ( n45700, P2_P1_PHYADDRPOINTER_REG_25_, n45704 );
nand U129786 ( n45701, n45702, n76670 );
nand U129787 ( n45704, n7428, n45705 );
nand U129788 ( n39871, P4_REG3_REG_10_, n39927 );
nand U129789 ( n39770, P4_REG3_REG_12_, n39826 );
nand U129790 ( n39640, P4_REG3_REG_14_, n39700 );
nand U129791 ( n37969, n39559, n39560 );
nand U129792 ( n39559, P4_IR_REG_17_, n76794 );
or U129793 ( n39560, n39561, n76793 );
nand U129794 ( n44857, n64236, n64237 );
nand U129795 ( n64236, P3_IR_REG_15_, n76840 );
or U129796 ( n64237, n14778, n76839 );
nand U129797 ( n46113, n47197, n47198 );
nand U129798 ( n47197, P2_P1_INSTADDRPOINTER_REG_9_, n47205 );
nand U129799 ( n47198, n47199, n73078 );
nand U129800 ( n47205, n47206, n47207 );
nand U129801 ( n47199, n47200, n47201 );
nand U129802 ( n47201, n47202, n7544 );
nand U129803 ( n47200, n47203, n76006 );
nor U129804 ( n47202, P2_P1_INSTADDRPOINTER_REG_8_, n76005 );
nand U129805 ( n15576, n47180, n47181 );
nand U129806 ( n47181, n76860, P2_P1_INSTADDRPOINTER_REG_9_ );
nor U129807 ( n47180, n47182, n47183 );
nor U129808 ( n47183, n73221, n76332 );
nand U129809 ( n67077, n68228, n68229 );
nand U129810 ( n68228, P2_P3_INSTADDRPOINTER_REG_9_, n68236 );
nand U129811 ( n68229, n68230, n73084 );
nand U129812 ( n68236, n68237, n68238 );
nand U129813 ( n25179, n26227, n26228 );
nand U129814 ( n26227, P1_P2_INSTADDRPOINTER_REG_9_, n26235 );
nand U129815 ( n26228, n26229, n73085 );
nand U129816 ( n26235, n26236, n26237 );
nand U129817 ( n58315, n59366, n59367 );
nand U129818 ( n59366, P2_P2_INSTADDRPOINTER_REG_9_, n59374 );
nand U129819 ( n59367, n59368, n73086 );
nand U129820 ( n59374, n59375, n59376 );
nand U129821 ( n68230, n68231, n68232 );
nand U129822 ( n68232, n68233, n5758 );
nand U129823 ( n68231, n68234, n75990 );
nor U129824 ( n68233, P2_P3_INSTADDRPOINTER_REG_8_, n75989 );
nand U129825 ( n26229, n26230, n26231 );
nand U129826 ( n26231, n26232, n4000 );
nand U129827 ( n26230, n26233, n76027 );
nor U129828 ( n26232, P1_P2_INSTADDRPOINTER_REG_8_, n76026 );
nand U129829 ( n59368, n59369, n59370 );
nand U129830 ( n59370, n59371, n6633 );
nand U129831 ( n59369, n59372, n75998 );
nor U129832 ( n59371, P2_P2_INSTADDRPOINTER_REG_8_, n75997 );
nand U129833 ( n11086, n68211, n68212 );
nand U129834 ( n68212, n76195, P2_P3_INSTADDRPOINTER_REG_9_ );
nor U129835 ( n68211, n68213, n68214 );
nor U129836 ( n68214, n73216, n76871 );
nand U129837 ( n6596, n26210, n26211 );
nand U129838 ( n26211, n76519, P1_P2_INSTADDRPOINTER_REG_9_ );
nor U129839 ( n26210, n26212, n26213 );
nor U129840 ( n26213, n73215, n76906 );
nand U129841 ( n13331, n59349, n59350 );
nand U129842 ( n59350, n76261, P2_P2_INSTADDRPOINTER_REG_9_ );
nor U129843 ( n59349, n59351, n59352 );
nor U129844 ( n59352, n73214, n76880 );
nand U129845 ( n37091, n40447, n40448 );
nand U129846 ( n40447, P4_IR_REG_23_, n40452 );
nand U129847 ( n40448, n40449, P4_IR_REG_31_ );
nand U129848 ( n40452, n40451, P4_IR_REG_31_ );
nand U129849 ( n45007, n64035, n64036 );
nand U129850 ( n64035, P3_IR_REG_16_, n76840 );
nand U129851 ( n64036, n64037, P3_IR_REG_31_ );
and U129852 ( n64037, n14375, n14374 );
nand U129853 ( n14374, P3_IR_REG_16_, n64038 );
nand U129854 ( n64038, n855, n74395 );
nand U129855 ( n43866, n64528, n64529 );
nand U129856 ( n64528, P3_IR_REG_13_, n76841 );
or U129857 ( n64529, n15084, n76839 );
xor U129858 ( n32064, n32882, P1_P3_INSTADDRPOINTER_REG_24_ );
xor U129859 ( n66667, n67643, P2_P3_INSTADDRPOINTER_REG_24_ );
xor U129860 ( n24832, n25638, P1_P2_INSTADDRPOINTER_REG_24_ );
xor U129861 ( n57966, n58775, P2_P2_INSTADDRPOINTER_REG_24_ );
nand U129862 ( n43666, n64817, n64818 );
nand U129863 ( n64818, n64819, P3_IR_REG_31_ );
nand U129864 ( n64817, P3_IR_REG_12_, n76840 );
and U129865 ( n64819, n15214, n15213 );
nand U129866 ( n15213, P3_IR_REG_12_, n64820 );
nand U129867 ( n64820, n869, n74301 );
xor U129868 ( n12010, n13059, P1_P1_INSTADDRPOINTER_REG_24_ );
xor U129869 ( n45741, n46597, P2_P1_INSTADDRPOINTER_REG_24_ );
xnor U129870 ( n41041, n74064, P3_REG3_REG_3_ );
nand U129871 ( n4351, n33460, n33461 );
nand U129872 ( n33461, n76468, P1_P3_INSTADDRPOINTER_REG_9_ );
nor U129873 ( n33460, n33462, n33463 );
nor U129874 ( n33463, n73217, n76897 );
xor U129875 ( n11929, n12854, P1_P1_INSTADDRPOINTER_REG_26_ );
nand U129876 ( n17668, n8213, P4_DATAO_REG_1_ );
nand U129877 ( n37930, n39752, n39753 );
nand U129878 ( n39752, P4_IR_REG_14_, n76794 );
nand U129879 ( n39753, n39754, P4_IR_REG_31_ );
and U129880 ( n39754, n39755, n39756 );
nand U129881 ( n39756, P4_IR_REG_14_, n40582 );
nand U129882 ( n40582, n2203, n74390 );
nand U129883 ( n16779, n8213, P4_DATAO_REG_7_ );
nand U129884 ( n64498, P3_REG3_REG_12_, n64789 );
nand U129885 ( n64199, P3_REG3_REG_14_, n64349 );
xor U129886 ( n37938, n37939, n37940 );
xor U129887 ( n37940, n37941, P4_REG2_REG_15_ );
and U129888 ( n49468, n50007, P3_DATAO_REG_0_ );
nand U129889 ( n32130, n73167, n33038 );
nand U129890 ( n33038, n33037, P1_P3_INSTADDRPOINTER_REG_20_ );
nand U129891 ( n45825, n73148, n46746 );
nand U129892 ( n46746, n46745, P2_P1_INSTADDRPOINTER_REG_20_ );
nand U129893 ( n12093, n73158, n13264 );
nand U129894 ( n13264, n13263, P1_P1_INSTADDRPOINTER_REG_20_ );
nand U129895 ( n66776, n73149, n67793 );
nand U129896 ( n67793, n67792, P2_P3_INSTADDRPOINTER_REG_20_ );
nand U129897 ( n24898, n73150, n25790 );
nand U129898 ( n25790, n25789, P1_P2_INSTADDRPOINTER_REG_20_ );
nand U129899 ( n58035, n73151, n58928 );
nand U129900 ( n58928, n58927, P2_P2_INSTADDRPOINTER_REG_20_ );
nand U129901 ( n44395, n64390, n64391 );
nand U129902 ( n64390, P3_IR_REG_14_, n76840 );
nand U129903 ( n64391, n64392, P3_IR_REG_31_ );
and U129904 ( n64392, n14923, n14922 );
nand U129905 ( n14922, P3_IR_REG_14_, n64393 );
nand U129906 ( n64393, n860, n74392 );
nand U129907 ( n49479, P3_DATAO_REG_1_, n49484 );
nand U129908 ( n49484, n76323, n49486 );
nand U129909 ( n49486, n76651, n76835 );
nand U129910 ( n45396, n49476, n49477 );
nand U129911 ( n49476, P2_BUF1_REG_1_, n76478 );
nand U129912 ( n49477, n49478, n76476 );
nand U129913 ( n49478, n49479, n49480 );
nand U129914 ( n1706, n42180, n42181 );
nand U129915 ( n42181, n76376, n41377 );
nand U129916 ( n42180, P3_DATAO_REG_1_, n76374 );
nand U129917 ( n1716, n42172, n42173 );
nand U129918 ( n42173, n76376, n41036 );
nand U129919 ( n42172, P3_DATAO_REG_3_, n76374 );
nand U129920 ( n1711, n42174, n42175 );
nand U129921 ( n42175, n76376, n40784 );
nand U129922 ( n42174, P3_DATAO_REG_2_, n76374 );
nand U129923 ( n1736, n42164, n42165 );
nand U129924 ( n42165, n76376, n40864 );
nand U129925 ( n42164, P3_DATAO_REG_7_, n76374 );
nand U129926 ( n1731, n42166, n42167 );
nand U129927 ( n42167, n76376, n40690 );
nand U129928 ( n42166, P3_DATAO_REG_6_, n76374 );
nand U129929 ( n1726, n42168, n42169 );
nand U129930 ( n42169, n76376, n41198 );
nand U129931 ( n42168, P3_DATAO_REG_5_, n76374 );
nand U129932 ( n1721, n42170, n42171 );
nand U129933 ( n42171, n76376, n40984 );
nand U129934 ( n42170, P3_DATAO_REG_4_, n76374 );
nand U129935 ( n1766, n42148, n42149 );
nand U129936 ( n42149, n76376, n40727 );
nand U129937 ( n42148, P3_DATAO_REG_13_, n76374 );
nand U129938 ( n1756, n42156, n42157 );
nand U129939 ( n42157, n76376, n40930 );
nand U129940 ( n42156, P3_DATAO_REG_11_, n76374 );
nand U129941 ( n1741, n42162, n42163 );
nand U129942 ( n42163, n76376, n41054 );
nand U129943 ( n42162, P3_DATAO_REG_8_, n76374 );
nand U129944 ( n1746, n42160, n42161 );
nand U129945 ( n42161, n76376, n40760 );
nand U129946 ( n42160, P3_DATAO_REG_9_, n76374 );
nand U129947 ( n1751, n42158, n42159 );
nand U129948 ( n42159, n76376, n41145 );
nand U129949 ( n42158, P3_DATAO_REG_10_, n76374 );
nand U129950 ( n1701, n42182, n42183 );
nand U129951 ( n42183, n76376, n42184 );
nand U129952 ( n42182, P3_DATAO_REG_0_, n76374 );
nand U129953 ( n1761, n42150, n42151 );
nand U129954 ( n42151, n76376, n41114 );
nand U129955 ( n42150, P3_DATAO_REG_12_, n76374 );
nand U129956 ( n1776, n42144, n42145 );
nand U129957 ( n42145, n76376, n40967 );
nand U129958 ( n42144, P3_DATAO_REG_15_, n76374 );
nand U129959 ( n49284, n49285, n49286 );
nand U129960 ( n49286, P2_P1_INSTQUEUE_REG_13__1_, n49275 );
nand U129961 ( n49285, n7442, n252 );
nand U129962 ( n49093, n49094, n49095 );
nand U129963 ( n49095, P2_P1_INSTQUEUE_REG_11__1_, n49085 );
nand U129964 ( n49094, n7443, n252 );
nand U129965 ( n48999, n49000, n49001 );
nand U129966 ( n49001, P2_P1_INSTQUEUE_REG_10__1_, n48990 );
nand U129967 ( n49000, n7444, n252 );
nand U129968 ( n48900, n48901, n48902 );
nand U129969 ( n48902, P2_P1_INSTQUEUE_REG_9__1_, n48891 );
nand U129970 ( n48901, n7445, n252 );
nand U129971 ( n48633, n48634, n48635 );
nand U129972 ( n48635, P2_P1_INSTQUEUE_REG_6__1_, n48624 );
nand U129973 ( n48634, n7448, n252 );
nand U129974 ( n48539, n48540, n48541 );
nand U129975 ( n48541, P2_P1_INSTQUEUE_REG_5__1_, n48530 );
nand U129976 ( n48540, n7449, n252 );
nand U129977 ( n49362, n49363, n49364 );
nand U129978 ( n49364, P2_P1_INSTQUEUE_REG_14__1_, n49353 );
nand U129979 ( n49363, n7440, n252 );
nand U129980 ( n48726, n48727, n48728 );
nand U129981 ( n48728, P2_P1_INSTQUEUE_REG_7__1_, n48718 );
nand U129982 ( n48727, n7447, n252 );
nand U129983 ( n1781, n42142, n42143 );
nand U129984 ( n42143, n76376, n41006 );
nand U129985 ( n42142, P3_DATAO_REG_16_, n76374 );
nand U129986 ( n1791, n42138, n42139 );
nand U129987 ( n42139, n76375, n40801 );
nand U129988 ( n42138, P3_DATAO_REG_18_, n76374 );
nand U129989 ( n1771, n42146, n42147 );
nand U129990 ( n42147, n76376, n41329 );
nand U129991 ( n42146, P3_DATAO_REG_14_, n76374 );
nand U129992 ( n1786, n42140, n42141 );
nand U129993 ( n42141, n76375, n41178 );
nand U129994 ( n42140, P3_DATAO_REG_17_, n76374 );
nand U129995 ( n32035, n73232, n32886 );
nand U129996 ( n32886, n32885, P1_P3_INSTADDRPOINTER_REG_24_ );
nand U129997 ( n66638, n73223, n67647 );
nand U129998 ( n67647, n67646, P2_P3_INSTADDRPOINTER_REG_24_ );
nand U129999 ( n24803, n73224, n25642 );
nand U130000 ( n25642, n25641, P1_P2_INSTADDRPOINTER_REG_24_ );
nand U130001 ( n57937, n73225, n58779 );
nand U130002 ( n58779, n58778, P2_P2_INSTADDRPOINTER_REG_24_ );
nand U130003 ( n9251, n11524, n11525 );
nand U130004 ( n11525, P1_P1_UWORD_REG_3_, n76618 );
nor U130005 ( n11524, n11527, n11528 );
nor U130006 ( n11527, n74954, n76617 );
nand U130007 ( n9176, n11607, n11608 );
nand U130008 ( n11608, P1_P1_LWORD_REG_3_, n76618 );
nor U130009 ( n11607, n11609, n11528 );
nor U130010 ( n11609, n74630, n76616 );
nor U130011 ( n13608, n13614, n13615 );
nor U130012 ( n13615, n74468, n76034 );
and U130013 ( n13614, n13613, P1_P1_INSTADDRPOINTER_REG_12_ );
xor U130014 ( n38456, n39970, P4_REG3_REG_9_ );
nand U130015 ( n45712, n73220, n46599 );
nand U130016 ( n46599, n46600, P2_P1_INSTADDRPOINTER_REG_24_ );
nand U130017 ( n11972, n74774, n13063 );
nand U130018 ( n13063, n13064, P1_P1_INSTADDRPOINTER_REG_24_ );
nand U130019 ( n1811, n42126, n42127 );
nand U130020 ( n42127, n76375, n40913 );
nand U130021 ( n42126, P3_DATAO_REG_22_, n76374 );
nand U130022 ( n1826, n42120, n42121 );
nand U130023 ( n42121, n76375, n41024 );
nand U130024 ( n42120, P3_DATAO_REG_25_, n76374 );
nand U130025 ( n1806, n42132, n42133 );
nand U130026 ( n42133, n76375, n41090 );
nand U130027 ( n42132, P3_DATAO_REG_21_, n76374 );
nand U130028 ( n1846, n42112, n42113 );
nand U130029 ( n42113, n76375, n40852 );
nand U130030 ( n42112, P3_DATAO_REG_29_, n76374 );
nand U130031 ( n1801, n42134, n42135 );
nand U130032 ( n42135, n76375, n41297 );
nand U130033 ( n42134, P3_DATAO_REG_20_, n42109 );
nand U130034 ( n1851, n42110, n42111 );
nand U130035 ( n42111, n76375, n41948 );
nand U130036 ( n42110, P3_DATAO_REG_30_, n42109 );
nand U130037 ( n1816, n42124, n42125 );
nand U130038 ( n42125, n76375, n41134 );
nand U130039 ( n42124, P3_DATAO_REG_23_, n42109 );
nand U130040 ( n1821, n42122, n42123 );
nand U130041 ( n42123, n76375, n40747 );
nand U130042 ( n42122, P3_DATAO_REG_24_, n42109 );
nand U130043 ( n1831, n42118, n42119 );
nand U130044 ( n42119, n76375, n40950 );
nand U130045 ( n42118, P3_DATAO_REG_26_, n42109 );
nand U130046 ( n1841, n42114, n42115 );
nand U130047 ( n42115, n76375, n40713 );
nand U130048 ( n42114, P3_DATAO_REG_28_, n42109 );
nand U130049 ( n1836, n42116, n42117 );
nand U130050 ( n42117, n76375, n40834 );
nand U130051 ( n42116, P3_DATAO_REG_27_, n42109 );
nand U130052 ( n1796, n42136, n42137 );
nand U130053 ( n42137, n76375, n41284 );
nand U130054 ( n42136, P3_DATAO_REG_19_, n42109 );
nand U130055 ( n1856, n42107, n42108 );
nand U130056 ( n42108, n76376, n41510 );
nand U130057 ( n42107, P3_DATAO_REG_31_, n42109 );
nand U130058 ( n32020, n32021, n32022 );
nand U130059 ( n32021, P1_P3_PHYADDRPOINTER_REG_25_, n32026 );
nand U130060 ( n32022, n32023, n76784 );
nand U130061 ( n32026, n3052, n32027 );
xor U130062 ( n48794, n64199, P3_REG3_REG_15_ );
nand U130063 ( n66623, n66624, n66625 );
nand U130064 ( n66624, P2_P3_PHYADDRPOINTER_REG_25_, n66629 );
nand U130065 ( n66625, n66626, n76718 );
nand U130066 ( n66629, n5653, n66630 );
nand U130067 ( n24788, n24789, n24790 );
nand U130068 ( n24789, P1_P2_PHYADDRPOINTER_REG_25_, n24794 );
nand U130069 ( n24790, n24791, n76766 );
nand U130070 ( n24794, n3895, n24795 );
nand U130071 ( n57922, n57923, n57924 );
nand U130072 ( n57923, P2_P2_PHYADDRPOINTER_REG_25_, n57928 );
nand U130073 ( n57924, n57925, n76699 );
nand U130074 ( n57928, n6528, n57929 );
nand U130075 ( n961, n9765, n9767 );
nand U130076 ( n9767, n76638, n9768 );
nand U130077 ( n9765, P3_D_REG_0_, n76637 );
nand U130078 ( n966, n9648, n9649 );
nand U130079 ( n9649, n76638, n9650 );
nand U130080 ( n9648, P3_D_REG_1_, n76637 );
xor U130081 ( n38495, n40049, P4_REG3_REG_7_ );
xnor U130082 ( n38243, P4_REG3_REG_22_, n39215 );
nand U130083 ( n39516, P4_REG3_REG_16_, n39578 );
nand U130084 ( n39391, P4_REG3_REG_18_, n39449 );
nand U130085 ( n39273, P4_REG3_REG_20_, n39340 );
nand U130086 ( n8871, n13493, n13494 );
nand U130087 ( n13494, n76887, P1_P1_INSTADDRPOINTER_REG_15_ );
nor U130088 ( n13493, n13495, n13497 );
nor U130089 ( n13497, n74869, n76599 );
nand U130090 ( n15991, n45333, n45334 );
nand U130091 ( n45334, P2_P1_UWORD_REG_2_, n76352 );
nor U130092 ( n45333, n45335, n45336 );
nor U130093 ( n45335, n73265, n76351 );
nand U130094 ( n15916, n45397, n45398 );
nand U130095 ( n45398, P2_P1_LWORD_REG_2_, n45325 );
nor U130096 ( n45397, n45399, n45336 );
nor U130097 ( n45399, n73165, n76350 );
nand U130098 ( n45077, n63712, n63713 );
nand U130099 ( n63712, P3_IR_REG_17_, n76840 );
or U130100 ( n63713, n13652, n76839 );
xor U130101 ( n38395, n39770, P4_REG3_REG_13_ );
xor U130102 ( n38361, n39640, P4_REG3_REG_15_ );
and U130103 ( n1026, n76637, P3_D_REG_13_ );
and U130104 ( n1036, n76637, P3_D_REG_15_ );
and U130105 ( n1046, n76637, P3_D_REG_17_ );
and U130106 ( n1056, n76637, P3_D_REG_19_ );
and U130107 ( n1066, n76637, P3_D_REG_21_ );
and U130108 ( n1081, n76637, P3_D_REG_24_ );
and U130109 ( n1091, n76637, P3_D_REG_26_ );
and U130110 ( n1101, n76637, P3_D_REG_28_ );
and U130111 ( n1116, n76637, P3_D_REG_31_ );
and U130112 ( n971, n76637, P3_D_REG_2_ );
and U130113 ( n981, n76637, P3_D_REG_4_ );
and U130114 ( n991, n76637, P3_D_REG_6_ );
and U130115 ( n1001, n76637, P3_D_REG_8_ );
and U130116 ( n1031, n76637, P3_D_REG_14_ );
and U130117 ( n1041, n76637, P3_D_REG_16_ );
and U130118 ( n1051, n76637, P3_D_REG_18_ );
and U130119 ( n1061, n76637, P3_D_REG_20_ );
and U130120 ( n1076, n76637, P3_D_REG_23_ );
and U130121 ( n1086, n76637, P3_D_REG_25_ );
and U130122 ( n1096, n76637, P3_D_REG_27_ );
and U130123 ( n1106, n76637, P3_D_REG_29_ );
and U130124 ( n1111, n76637, P3_D_REG_30_ );
and U130125 ( n976, n76637, P3_D_REG_3_ );
and U130126 ( n986, n76637, P3_D_REG_5_ );
and U130127 ( n1006, n76637, P3_D_REG_9_ );
and U130128 ( n1016, n76637, P3_D_REG_11_ );
and U130129 ( n1011, n76637, P3_D_REG_10_ );
and U130130 ( n1021, n76637, P3_D_REG_12_ );
nand U130131 ( n16176, n44969, n44970 );
nor U130132 ( n44970, n44971, n44972 );
nor U130133 ( n44969, n44975, n44976 );
nor U130134 ( n44971, P2_P1_EAX_REG_2_, n44965 );
nand U130135 ( n11605, n16522, n16523 );
nand U130136 ( n16522, P1_BUF1_REG_2_, n76610 );
nand U130137 ( n16523, n16524, n76613 );
xnor U130138 ( n16524, n16525, n16527 );
nand U130139 ( n16362, n16363, n16364 );
nand U130140 ( n16364, P1_P1_INSTQUEUE_REG_14__2_, n16340 );
nand U130141 ( n16363, n4797, n11 );
nand U130142 ( n16257, n16258, n16259 );
nand U130143 ( n16259, P1_P1_INSTQUEUE_REG_13__2_, n16235 );
nand U130144 ( n16258, n4798, n11 );
nand U130145 ( n16054, n16055, n16057 );
nand U130146 ( n16057, P1_P1_INSTQUEUE_REG_11__2_, n16033 );
nand U130147 ( n16055, n4799, n11 );
nand U130148 ( n15947, n15948, n15949 );
nand U130149 ( n15949, P1_P1_INSTQUEUE_REG_10__2_, n15925 );
nand U130150 ( n15948, n4800, n11 );
nand U130151 ( n15842, n15843, n15844 );
nand U130152 ( n15844, P1_P1_INSTQUEUE_REG_9__2_, n15820 );
nand U130153 ( n15843, n4802, n11 );
nand U130154 ( n15533, n15534, n15535 );
nand U130155 ( n15535, P1_P1_INSTQUEUE_REG_6__2_, n15512 );
nand U130156 ( n15534, n4804, n11 );
nand U130157 ( n15427, n15428, n15429 );
nand U130158 ( n15429, P1_P1_INSTQUEUE_REG_5__2_, n15405 );
nand U130159 ( n15428, n4805, n11 );
nand U130160 ( n15634, n15635, n15637 );
nand U130161 ( n15637, P1_P1_INSTQUEUE_REG_7__2_, n15609 );
nand U130162 ( n15635, n4803, n11 );
nor U130163 ( n23160, n23214, n23215 );
nor U130164 ( n23215, n76539, P1_P2_EAX_REG_27_ );
nor U130165 ( n56281, n56335, n56336 );
nor U130166 ( n56336, n76281, P2_P2_EAX_REG_27_ );
nand U130167 ( n56208, n56209, n56210 );
nand U130168 ( n56210, n56211, n56212 );
nand U130169 ( n56209, P2_P2_EAX_REG_30_, n56214 );
nor U130170 ( n56211, n73393, n75203 );
nand U130171 ( n23087, n23088, n23089 );
nand U130172 ( n23089, n23090, n23091 );
nand U130173 ( n23088, P1_P2_EAX_REG_30_, n23093 );
nor U130174 ( n23090, n73394, n75205 );
nor U130175 ( n64648, n64693, n64694 );
nor U130176 ( n64694, n76215, P2_P3_EAX_REG_27_ );
nand U130177 ( n64577, n64578, n64579 );
nand U130178 ( n64579, n64580, n64581 );
nand U130179 ( n64578, P2_P3_EAX_REG_30_, n64583 );
nor U130180 ( n64580, n73390, n75204 );
nor U130181 ( n30489, n30534, n30535 );
nor U130182 ( n30535, n76482, P1_P3_EAX_REG_27_ );
nand U130183 ( n30418, n30419, n30420 );
nand U130184 ( n30420, n30421, n30422 );
nand U130185 ( n30419, P1_P3_EAX_REG_30_, n30424 );
nor U130186 ( n30421, n73395, n75206 );
nand U130187 ( n2931, n37677, n37678 );
nand U130188 ( n37678, n76451, n37023 );
nand U130189 ( n37677, P4_DATAO_REG_1_, n76449 );
nand U130190 ( n2936, n37675, n37676 );
nand U130191 ( n37676, n76451, n36381 );
nand U130192 ( n37675, P4_DATAO_REG_2_, n76449 );
nand U130193 ( n2961, n37663, n37664 );
nand U130194 ( n37664, n76451, n36462 );
nand U130195 ( n37663, P4_DATAO_REG_7_, n76449 );
nand U130196 ( n2941, n37673, n37674 );
nand U130197 ( n37674, n76451, n36649 );
nand U130198 ( n37673, P4_DATAO_REG_3_, n76449 );
nand U130199 ( n2946, n37671, n37672 );
nand U130200 ( n37672, n76451, n36589 );
nand U130201 ( n37671, P4_DATAO_REG_4_, n76449 );
nand U130202 ( n2951, n37669, n37670 );
nand U130203 ( n37670, n76451, n36817 );
nand U130204 ( n37669, P4_DATAO_REG_5_, n76449 );
nand U130205 ( n2956, n37667, n37668 );
nand U130206 ( n37668, n76451, n36286 );
nand U130207 ( n37667, P4_DATAO_REG_6_, n76449 );
nand U130208 ( n2991, n37651, n37652 );
nand U130209 ( n37652, n76451, n36322 );
nand U130210 ( n37651, P4_DATAO_REG_13_, n76449 );
nand U130211 ( n61966, n56587, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U130212 ( n28661, n23465, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U130213 ( n2971, n37659, n37660 );
nand U130214 ( n37660, n76451, n36355 );
nand U130215 ( n37659, P4_DATAO_REG_9_, n76449 );
nand U130216 ( n2981, n37655, n37656 );
nand U130217 ( n37656, n76451, n36532 );
nand U130218 ( n37655, P4_DATAO_REG_11_, n76449 );
nand U130219 ( n2966, n37661, n37662 );
nand U130220 ( n37662, n76451, n36667 );
nand U130221 ( n37661, P4_DATAO_REG_8_, n76449 );
nand U130222 ( n3001, n37647, n37648 );
nand U130223 ( n37648, n76451, n36572 );
nand U130224 ( n37647, P4_DATAO_REG_15_, n76449 );
nand U130225 ( n2926, n37679, n37680 );
nand U130226 ( n37680, n76451, n37288 );
nand U130227 ( n37679, P4_DATAO_REG_0_, n76449 );
nand U130228 ( n2986, n37653, n37654 );
nand U130229 ( n37654, n76451, n36730 );
nand U130230 ( n37653, P4_DATAO_REG_12_, n76449 );
nand U130231 ( n2976, n37657, n37658 );
nand U130232 ( n37658, n76451, n36762 );
nand U130233 ( n37657, P4_DATAO_REG_10_, n76449 );
nand U130234 ( n3006, n37645, n37646 );
nand U130235 ( n37646, n76451, n36613 );
nand U130236 ( n37645, P4_DATAO_REG_16_, n76449 );
nand U130237 ( n70566, n64974, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U130238 ( n3016, n37639, n37640 );
nand U130239 ( n37640, n76450, n36398 );
nand U130240 ( n37639, P4_DATAO_REG_18_, n76449 );
nand U130241 ( n35840, n30772, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U130242 ( n2996, n37649, n37650 );
nand U130243 ( n37650, n76451, n36961 );
nand U130244 ( n37649, P4_DATAO_REG_14_, n76449 );
nand U130245 ( n3011, n37641, n37642 );
nand U130246 ( n37642, n76450, n36797 );
nand U130247 ( n37641, P4_DATAO_REG_17_, n76449 );
nand U130248 ( n50030, DIN_27_, n76929 );
xor U130249 ( n54672, n66278, P3_REG3_REG_5_ );
nand U130250 ( n38038, n39498, n39499 );
nand U130251 ( n39498, P4_IR_REG_18_, n39503 );
nand U130252 ( n39499, n39500, P4_IR_REG_31_ );
nand U130253 ( n39503, n39502, P4_IR_REG_31_ );
nand U130254 ( n17702, n17054, P4_DATAO_REG_4_ );
and U130255 ( n17054, DIN_24_, n76927 );
nand U130256 ( n28670, n23469, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U130257 ( n61975, n56591, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nor U130258 ( n23469, n24210, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nor U130259 ( n56591, n57332, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U130260 ( n70575, n64978, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nor U130261 ( n64978, n65754, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130262 ( n35849, n30776, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nor U130263 ( n30776, n31504, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130264 ( n3051, n37625, n37626 );
nand U130265 ( n37626, n76450, n36925 );
nand U130266 ( n37625, P4_DATAO_REG_25_, n76449 );
nand U130267 ( n3036, n37631, n37632 );
nand U130268 ( n37632, n76450, n36339 );
nand U130269 ( n37631, P4_DATAO_REG_22_, n76449 );
nand U130270 ( n3026, n37635, n37636 );
nand U130271 ( n37636, n76450, n36512 );
nand U130272 ( n37635, P4_DATAO_REG_20_, n76449 );
nand U130273 ( n3031, n37633, n37634 );
nand U130274 ( n37634, n76450, n36747 );
nand U130275 ( n37633, P4_DATAO_REG_21_, n76449 );
nand U130276 ( n3021, n37637, n37638 );
nand U130277 ( n37638, n76450, n36702 );
nand U130278 ( n37637, P4_DATAO_REG_19_, n37612 );
nand U130279 ( n3061, n37619, n37620 );
nand U130280 ( n37620, n76450, n36442 );
nand U130281 ( n37619, P4_DATAO_REG_27_, n37612 );
nand U130282 ( n3071, n37615, n37616 );
nand U130283 ( n37616, n76450, n37295 );
nand U130284 ( n37615, P4_DATAO_REG_29_, n37612 );
nand U130285 ( n3046, n37627, n37628 );
nand U130286 ( n37628, n76450, n36551 );
nand U130287 ( n37627, P4_DATAO_REG_24_, n37612 );
nand U130288 ( n3041, n37629, n37630 );
nand U130289 ( n37630, n76450, n36633 );
nand U130290 ( n37629, P4_DATAO_REG_23_, n37612 );
nand U130291 ( n3056, n37623, n37624 );
nand U130292 ( n37624, n76450, n36305 );
nand U130293 ( n37623, P4_DATAO_REG_26_, n37612 );
nand U130294 ( n3076, n37613, n37614 );
nand U130295 ( n37614, n76450, n37299 );
nand U130296 ( n37613, P4_DATAO_REG_30_, n37612 );
nand U130297 ( n3066, n37617, n37618 );
nand U130298 ( n37618, n76450, n36429 );
nand U130299 ( n37617, P4_DATAO_REG_28_, n37612 );
nand U130300 ( n3081, n37610, n37611 );
nand U130301 ( n37611, n76451, n37353 );
nand U130302 ( n37610, P4_DATAO_REG_31_, n37612 );
nand U130303 ( n23092, n23206, P1_P2_EAX_REG_27_ );
nor U130304 ( n23206, n23207, n76539 );
nand U130305 ( n56213, n56327, P2_P2_EAX_REG_27_ );
nor U130306 ( n56327, n56328, n76281 );
nor U130307 ( n23091, P1_P2_EAX_REG_30_, n23092 );
nor U130308 ( n56212, P2_P2_EAX_REG_30_, n56213 );
nand U130309 ( n64582, n64690, P2_P3_EAX_REG_27_ );
nor U130310 ( n64690, n64691, n76215 );
nor U130311 ( n64581, P2_P3_EAX_REG_30_, n64582 );
nand U130312 ( n30423, n30531, P1_P3_EAX_REG_27_ );
nor U130313 ( n30531, n30532, n76482 );
nor U130314 ( n30422, P1_P3_EAX_REG_30_, n30423 );
nand U130315 ( n17902, n17054, P4_DATAO_REG_3_ );
nand U130316 ( n23156, n23157, n23158 );
nand U130317 ( n23157, P1_P2_EAX_REG_29_, n23095 );
nand U130318 ( n23158, n23159, P1_P2_EAX_REG_28_ );
nor U130319 ( n23159, P1_P2_EAX_REG_29_, n23092 );
xor U130320 ( n32161, n33037, P1_P3_INSTADDRPOINTER_REG_20_ );
nand U130321 ( n56277, n56278, n56279 );
nand U130322 ( n56278, P2_P2_EAX_REG_29_, n56216 );
nand U130323 ( n56279, n56280, P2_P2_EAX_REG_28_ );
nor U130324 ( n56280, P2_P2_EAX_REG_29_, n56213 );
nand U130325 ( n64644, n64645, n64646 );
nand U130326 ( n64645, P2_P3_EAX_REG_29_, n64585 );
nand U130327 ( n64646, n64647, P2_P3_EAX_REG_28_ );
nor U130328 ( n64647, P2_P3_EAX_REG_29_, n64582 );
xor U130329 ( n12137, n13263, P1_P1_INSTADDRPOINTER_REG_20_ );
nand U130330 ( n30485, n30486, n30487 );
nand U130331 ( n30486, P1_P3_EAX_REG_29_, n30426 );
nand U130332 ( n30487, n30488, P1_P3_EAX_REG_28_ );
nor U130333 ( n30488, P1_P3_EAX_REG_29_, n30423 );
xor U130334 ( n45856, n46745, P2_P1_INSTADDRPOINTER_REG_20_ );
xor U130335 ( n32063, n32885, P1_P3_INSTADDRPOINTER_REG_24_ );
xor U130336 ( n66807, n67792, P2_P3_INSTADDRPOINTER_REG_20_ );
xor U130337 ( n24929, n25789, P1_P2_INSTADDRPOINTER_REG_20_ );
xor U130338 ( n58066, n58927, P2_P2_INSTADDRPOINTER_REG_20_ );
xor U130339 ( n66666, n67646, P2_P3_INSTADDRPOINTER_REG_24_ );
xor U130340 ( n24831, n25641, P1_P2_INSTADDRPOINTER_REG_24_ );
xor U130341 ( n57965, n58778, P2_P2_INSTADDRPOINTER_REG_24_ );
nand U130342 ( n15571, n47224, n47225 );
nand U130343 ( n47225, n76860, P2_P1_INSTADDRPOINTER_REG_8_ );
nor U130344 ( n47224, n47226, n47227 );
nor U130345 ( n47227, n75965, n76332 );
nand U130346 ( n22737, P1_P2_INSTQUEUERD_ADDR_REG_1_, n73520 );
nand U130347 ( n55853, P2_P2_INSTQUEUERD_ADDR_REG_1_, n73521 );
nand U130348 ( n11081, n68255, n68256 );
nand U130349 ( n68256, n76195, P2_P3_INSTADDRPOINTER_REG_8_ );
nor U130350 ( n68255, n68257, n68258 );
nor U130351 ( n68258, n74749, n76871 );
nand U130352 ( n6591, n26254, n26255 );
nand U130353 ( n26255, n76519, P1_P2_INSTADDRPOINTER_REG_8_ );
nor U130354 ( n26254, n26256, n26257 );
nor U130355 ( n26257, n74748, n76906 );
nand U130356 ( n13326, n59393, n59394 );
nand U130357 ( n59394, n76261, P2_P2_INSTADDRPOINTER_REG_8_ );
nor U130358 ( n59393, n59395, n59396 );
nor U130359 ( n59396, n74747, n76880 );
nand U130360 ( n64077, P2_P3_INSTQUEUERD_ADDR_REG_1_, n73518 );
nand U130361 ( n30060, P1_P3_INSTQUEUERD_ADDR_REG_1_, n73532 );
xor U130362 ( n38424, n39871, P4_REG3_REG_11_ );
xor U130363 ( n54632, n66096, P3_REG3_REG_7_ );
xor U130364 ( n12009, n13064, P1_P1_INSTADDRPOINTER_REG_24_ );
nand U130365 ( n61979, n56592, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U130366 ( n28674, n23470, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U130367 ( n22736, P1_P2_INSTQUEUERD_ADDR_REG_0_, n73055 );
nand U130368 ( n55852, P2_P2_INSTQUEUERD_ADDR_REG_0_, n73054 );
nor U130369 ( n23470, n22736, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nor U130370 ( n56592, n55852, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U130371 ( n70579, n64979, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U130372 ( n64076, P2_P3_INSTQUEUERD_ADDR_REG_0_, n73053 );
xor U130373 ( n45740, n46600, P2_P1_INSTADDRPOINTER_REG_24_ );
nor U130374 ( n64979, n64076, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130375 ( n35853, n30777, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U130376 ( n30059, P1_P3_INSTQUEUERD_ADDR_REG_0_, n73059 );
nor U130377 ( n30777, n30059, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130378 ( n8866, n13542, n13543 );
nand U130379 ( n13543, n76887, P1_P1_INSTADDRPOINTER_REG_14_ );
nor U130380 ( n13542, n13544, n13545 );
nor U130381 ( n13545, n74861, n76599 );
nor U130382 ( n23466, n22737, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nor U130383 ( n56588, n55853, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nor U130384 ( n64975, n64077, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130385 ( n2186, n40438, n40439 );
nand U130386 ( n40439, n76401, n40401 );
nand U130387 ( n40438, P4_D_REG_0_, n76400 );
nand U130388 ( n2191, n40435, n40436 );
nand U130389 ( n40436, n76401, n40406 );
nand U130390 ( n40435, P4_D_REG_1_, n76400 );
nor U130391 ( n30773, n30060, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
xnor U130392 ( n48202, P3_REG3_REG_20_, n62871 );
nand U130393 ( n63675, P3_REG3_REG_16_, n63990 );
nand U130394 ( n62945, P3_REG3_REG_18_, n63267 );
nand U130395 ( n17426, n17054, P4_DATAO_REG_5_ );
nor U130396 ( n23494, n73503, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nor U130397 ( n56616, n73504, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
xor U130398 ( n49029, n64498, P3_REG3_REG_13_ );
nand U130399 ( n28914, P1_P2_INSTQUEUERD_ADDR_REG_0_, n74423 );
nand U130400 ( n62219, P2_P2_INSTQUEUERD_ADDR_REG_0_, n74424 );
nand U130401 ( n28912, n28920, n28921 );
nand U130402 ( n28920, n28923, n73503 );
nand U130403 ( n28921, P1_P2_INSTQUEUEWR_ADDR_REG_3_, n28922 );
or U130404 ( n28922, n28923, n73503 );
nand U130405 ( n62217, n62225, n62226 );
nand U130406 ( n62225, n62228, n73504 );
nand U130407 ( n62226, P2_P2_INSTQUEUEWR_ADDR_REG_3_, n62227 );
or U130408 ( n62227, n62228, n73504 );
nand U130409 ( n28915, n28928, n28929 );
nand U130410 ( n28928, n28914, n73055 );
nand U130411 ( n28929, P1_P2_INSTQUEUEWR_ADDR_REG_1_, n28930 );
nand U130412 ( n28930, P1_P2_INSTQUEUERD_ADDR_REG_1_, n4255 );
nand U130413 ( n62220, n62233, n62234 );
nand U130414 ( n62233, n62219, n73054 );
nand U130415 ( n62234, P2_P2_INSTQUEUEWR_ADDR_REG_1_, n62235 );
nand U130416 ( n62235, P2_P2_INSTQUEUERD_ADDR_REG_1_, n6888 );
nand U130417 ( n28923, n28925, n28926 );
nand U130418 ( n28925, n28915, n73516 );
nand U130419 ( n28926, P1_P2_INSTQUEUEWR_ADDR_REG_2_, n28927 );
or U130420 ( n28927, n73516, n28915 );
nand U130421 ( n62228, n62230, n62231 );
nand U130422 ( n62230, n62220, n73517 );
nand U130423 ( n62231, P2_P2_INSTQUEUEWR_ADDR_REG_2_, n62232 );
or U130424 ( n62232, n73517, n62220 );
nor U130425 ( n28919, P1_P2_INSTQUEUERD_ADDR_REG_4_, n4230 );
nor U130426 ( n62224, P2_P2_INSTQUEUERD_ADDR_REG_4_, n6863 );
nand U130427 ( n28645, n28917, n28918 );
xnor U130428 ( n28917, n28924, n28923 );
nand U130429 ( n28918, n28919, P1_P2_INSTQUEUEWR_ADDR_REG_4_ );
xor U130430 ( n28924, n73136, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U130431 ( n61950, n62222, n62223 );
xnor U130432 ( n62222, n62229, n62228 );
nand U130433 ( n62223, n62224, P2_P2_INSTQUEUEWR_ADDR_REG_4_ );
xor U130434 ( n62229, n73137, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nor U130435 ( n65003, n73502, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nor U130436 ( n30801, n73524, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130437 ( n70819, P2_P3_INSTQUEUERD_ADDR_REG_0_, n74425 );
nand U130438 ( n70817, n70825, n70826 );
nand U130439 ( n70825, n70828, n73502 );
nand U130440 ( n70826, P2_P3_INSTQUEUEWR_ADDR_REG_3_, n70827 );
or U130441 ( n70827, n70828, n73502 );
nand U130442 ( n70820, n70833, n70834 );
nand U130443 ( n70833, n70819, n73053 );
nand U130444 ( n70834, P2_P3_INSTQUEUEWR_ADDR_REG_1_, n70835 );
nand U130445 ( n70835, P2_P3_INSTQUEUERD_ADDR_REG_1_, n6033 );
nand U130446 ( n70828, n70830, n70831 );
nand U130447 ( n70830, n70820, n73515 );
nand U130448 ( n70831, P2_P3_INSTQUEUEWR_ADDR_REG_2_, n70832 );
or U130449 ( n70832, n73515, n70820 );
nor U130450 ( n70824, P2_P3_INSTQUEUERD_ADDR_REG_4_, n6008 );
nand U130451 ( n70550, n70822, n70823 );
xnor U130452 ( n70822, n70829, n70828 );
nand U130453 ( n70823, n70824, P2_P3_INSTQUEUEWR_ADDR_REG_4_ );
xor U130454 ( n70829, n73139, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U130455 ( n36093, P1_P3_INSTQUEUERD_ADDR_REG_0_, n74426 );
nand U130456 ( n36091, n36099, n36100 );
nand U130457 ( n36099, n36102, n73524 );
nand U130458 ( n36100, P1_P3_INSTQUEUEWR_ADDR_REG_3_, n36101 );
or U130459 ( n36101, n36102, n73524 );
nand U130460 ( n36094, n36107, n36108 );
nand U130461 ( n36107, n36093, n73059 );
nand U130462 ( n36108, P1_P3_INSTQUEUEWR_ADDR_REG_1_, n36109 );
nand U130463 ( n36109, P1_P3_INSTQUEUERD_ADDR_REG_1_, n3418 );
nand U130464 ( n36102, n36104, n36105 );
nand U130465 ( n36104, n36094, n73526 );
nand U130466 ( n36105, P1_P3_INSTQUEUEWR_ADDR_REG_2_, n36106 );
or U130467 ( n36106, n73526, n36094 );
nor U130468 ( n36098, P1_P3_INSTQUEUERD_ADDR_REG_4_, n3393 );
nand U130469 ( n35824, n36096, n36097 );
xnor U130470 ( n36096, n36103, n36102 );
nand U130471 ( n36097, n36098, P1_P3_INSTQUEUEWR_ADDR_REG_4_ );
xor U130472 ( n36103, n73138, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U130473 ( n33405, P1_P3_INSTADDRPOINTER_REG_9_, n76472 );
nand U130474 ( n4346, n33500, n33501 );
nand U130475 ( n33501, n76468, P1_P3_INSTADDRPOINTER_REG_8_ );
nor U130476 ( n33500, n33502, n33503 );
nor U130477 ( n33503, n74750, n76897 );
xor U130478 ( n40914, n62738, P3_REG3_REG_21_ );
nand U130479 ( n62738, P3_REG3_REG_20_, n62871 );
and U130480 ( n2196, n76400, P4_D_REG_2_ );
and U130481 ( n2206, n76400, P4_D_REG_4_ );
and U130482 ( n2216, n76400, P4_D_REG_6_ );
and U130483 ( n2231, n76400, P4_D_REG_9_ );
and U130484 ( n2241, n76400, P4_D_REG_11_ );
and U130485 ( n2251, n76400, P4_D_REG_13_ );
and U130486 ( n2261, n76400, P4_D_REG_15_ );
and U130487 ( n2271, n76400, P4_D_REG_17_ );
and U130488 ( n2281, n76400, P4_D_REG_19_ );
and U130489 ( n2291, n76400, P4_D_REG_21_ );
and U130490 ( n2306, n76400, P4_D_REG_24_ );
and U130491 ( n2316, n76400, P4_D_REG_26_ );
and U130492 ( n2201, n76400, P4_D_REG_3_ );
and U130493 ( n2211, n76400, P4_D_REG_5_ );
and U130494 ( n2226, n76400, P4_D_REG_8_ );
and U130495 ( n2236, n76400, P4_D_REG_10_ );
and U130496 ( n2246, n76400, P4_D_REG_12_ );
and U130497 ( n2256, n76400, P4_D_REG_14_ );
and U130498 ( n2266, n76400, P4_D_REG_16_ );
and U130499 ( n2276, n76400, P4_D_REG_18_ );
and U130500 ( n2286, n76400, P4_D_REG_20_ );
and U130501 ( n2301, n76400, P4_D_REG_23_ );
and U130502 ( n2311, n76400, P4_D_REG_25_ );
and U130503 ( n2321, n76400, P4_D_REG_27_ );
nand U130504 ( n23203, n23204, n23205 );
nand U130505 ( n23204, n163, P1_BUF1_REG_28_ );
or U130506 ( n23205, n23092, P1_P2_EAX_REG_28_ );
or U130507 ( n64687, n75942, n75943 );
nor U130508 ( n75942, n73390, n64648 );
nor U130509 ( n75943, n64582, P2_P3_EAX_REG_28_ );
nand U130510 ( n56324, n56325, n56326 );
nand U130511 ( n56325, n435, P2_BUF1_REG_28_ );
or U130512 ( n56326, n56213, P2_P2_EAX_REG_28_ );
xor U130513 ( n40748, n62545, P3_REG3_REG_23_ );
nand U130514 ( n62545, P3_REG3_REG_22_, n62638 );
or U130515 ( n30528, n75944, n75945 );
nor U130516 ( n75944, n73395, n30489 );
nor U130517 ( n75945, n30423, P1_P3_EAX_REG_28_ );
nand U130518 ( n32219, n74879, n33186 );
nand U130519 ( n33186, n33185, P1_P3_INSTADDRPOINTER_REG_16_ );
nand U130520 ( n12209, n74847, n13447 );
nand U130521 ( n13447, n13445, P1_P1_INSTADDRPOINTER_REG_16_ );
xnor U130522 ( n37924, n37925, n37926 );
xor U130523 ( n37926, P4_REG2_REG_14_, n1972 );
nand U130524 ( n45911, n74841, n46895 );
nand U130525 ( n46895, n46894, P2_P1_INSTADDRPOINTER_REG_16_ );
nand U130526 ( n66862, n74872, n67942 );
nand U130527 ( n67942, n67941, P2_P3_INSTADDRPOINTER_REG_16_ );
nand U130528 ( n24986, n74873, n25939 );
nand U130529 ( n25939, n25938, P1_P2_INSTADDRPOINTER_REG_16_ );
nand U130530 ( n58121, n74874, n59077 );
nand U130531 ( n59077, n59076, P2_P2_INSTADDRPOINTER_REG_16_ );
xor U130532 ( n49568, n65930, P3_REG3_REG_9_ );
and U130533 ( n2326, n76400, P4_D_REG_28_ );
and U130534 ( n2341, n76400, P4_D_REG_31_ );
and U130535 ( n2331, n76400, P4_D_REG_29_ );
and U130536 ( n2336, n76400, P4_D_REG_30_ );
nand U130537 ( n17917, n17054, P4_DATAO_REG_2_ );
nand U130538 ( n12489, P1_P1_PHYADDRPOINTER_REG_6_, n12513 );
nand U130539 ( n12032, P1_P1_PHYADDRPOINTER_REG_20_, n12104 );
nand U130540 ( n8480, n9424, P1_P1_STATE2_REG_1_ );
nor U130541 ( n9424, n4762, n9425 );
nand U130542 ( n12238, P1_P1_PHYADDRPOINTER_REG_14_, n12282 );
nand U130543 ( n12045, P1_P1_PHYADDRPOINTER_REG_21_, n5307 );
nand U130544 ( n11830, P1_P1_PHYADDRPOINTER_REG_27_, n11865 );
nand U130545 ( n12437, P1_P1_PHYADDRPOINTER_REG_8_, n12445 );
nand U130546 ( n11980, P1_P1_PHYADDRPOINTER_REG_23_, n11993 );
nand U130547 ( n11902, P1_P1_PHYADDRPOINTER_REG_25_, n11928 );
nand U130548 ( n11760, P1_P1_PHYADDRPOINTER_REG_29_, n11802 );
nand U130549 ( n12375, P1_P1_PHYADDRPOINTER_REG_10_, n12387 );
nand U130550 ( n12537, P1_P1_PHYADDRPOINTER_REG_4_, n12563 );
nand U130551 ( n8655, n8657, n8658 );
nand U130552 ( n8657, P1_P1_EBX_REG_23_, n8662 );
nand U130553 ( n8658, n8637, n8659 );
nand U130554 ( n8662, n8428, n8663 );
nand U130555 ( n9385, n9347, n9387 );
nand U130556 ( n9387, P1_P1_PHYADDRPOINTER_REG_1_, n9388 );
nand U130557 ( n9388, n8414, n9389 );
nand U130558 ( n9389, P1_P1_PHYADDRPOINTER_REG_0_, n76742 );
xor U130559 ( n48566, n63675, P3_REG3_REG_17_ );
nand U130560 ( n15921, n45393, n45394 );
nand U130561 ( n45394, P2_P1_LWORD_REG_1_, n45325 );
nor U130562 ( n45393, n45395, n45332 );
nor U130563 ( n45395, n74609, n76350 );
nand U130564 ( n15996, n45329, n45330 );
nand U130565 ( n45330, P2_P1_UWORD_REG_1_, n45325 );
nor U130566 ( n45329, n45331, n45332 );
nor U130567 ( n45331, n74908, n76351 );
nand U130568 ( n9183, n9192, n9193 );
nand U130569 ( n9192, P1_P1_EBX_REG_7_, n9197 );
nand U130570 ( n9193, n9145, n9194 );
nand U130571 ( n9197, n8428, n9198 );
nand U130572 ( n8923, n8930, n8932 );
nand U130573 ( n8930, P1_P1_EBX_REG_15_, n8935 );
nand U130574 ( n8932, n8884, n8933 );
nand U130575 ( n8935, n8428, n8937 );
nand U130576 ( n8988, n8997, n8998 );
nand U130577 ( n8997, P1_P1_EBX_REG_13_, n9002 );
nand U130578 ( n8998, n8958, n8999 );
nand U130579 ( n9002, n8428, n9003 );
nand U130580 ( n8794, n8803, n8804 );
nand U130581 ( n8803, P1_P1_EBX_REG_19_, n8808 );
nand U130582 ( n8804, n8763, n8805 );
nand U130583 ( n8808, n8428, n8809 );
xnor U130584 ( n47958, P3_REG3_REG_22_, n62638 );
xor U130585 ( n38332, n39516, P4_REG3_REG_17_ );
nand U130586 ( n46135, P2_P1_PHYADDRPOINTER_REG_6_, n46154 );
nand U130587 ( n45776, P2_P1_PHYADDRPOINTER_REG_20_, n45834 );
nand U130588 ( n45928, P2_P1_PHYADDRPOINTER_REG_14_, n45963 );
nand U130589 ( n45787, P2_P1_PHYADDRPOINTER_REG_21_, n7962 );
nand U130590 ( n45606, P2_P1_PHYADDRPOINTER_REG_27_, n45640 );
nand U130591 ( n46093, P2_P1_PHYADDRPOINTER_REG_8_, n46100 );
nand U130592 ( n45717, P2_P1_PHYADDRPOINTER_REG_23_, n45727 );
nand U130593 ( n45650, P2_P1_PHYADDRPOINTER_REG_25_, n45694 );
nand U130594 ( n45531, P2_P1_PHYADDRPOINTER_REG_29_, n45560 );
nand U130595 ( n46049, P2_P1_PHYADDRPOINTER_REG_10_, n46058 );
nand U130596 ( n46174, P2_P1_PHYADDRPOINTER_REG_4_, n46194 );
nand U130597 ( n43338, n43366, P2_P1_STATE2_REG_1_ );
nor U130598 ( n43366, n7407, n43367 );
nand U130599 ( n42718, n42719, n42720 );
nand U130600 ( n42719, P2_P1_EBX_REG_23_, n42723 );
nand U130601 ( n42720, n42703, n42721 );
nand U130602 ( n42723, n42524, n42724 );
nand U130603 ( n32127, n73167, n33041 );
nand U130604 ( n33041, n33040, P1_P3_INSTADDRPOINTER_REG_20_ );
nand U130605 ( n16484, P4_DATAO_REG_1_, n16490 );
nand U130606 ( n16490, n76589, n16493 );
nand U130607 ( n16493, n76654, n74955 );
nand U130608 ( n11600, n16480, n16482 );
nand U130609 ( n16480, P1_BUF1_REG_1_, n76610 );
nand U130610 ( n16482, n16483, n76612 );
nand U130611 ( n16483, n16484, n16485 );
nand U130612 ( n12089, n73158, n13268 );
nand U130613 ( n13268, n13267, P1_P1_INSTADDRPOINTER_REG_20_ );
nand U130614 ( n43334, n43303, n43335 );
nand U130615 ( n43335, P2_P1_PHYADDRPOINTER_REG_1_, n43336 );
nand U130616 ( n43336, n42500, n43337 );
nand U130617 ( n43337, P2_P1_PHYADDRPOINTER_REG_0_, n76675 );
nand U130618 ( n45822, n73148, n46749 );
nand U130619 ( n46749, n46748, P2_P1_INSTADDRPOINTER_REG_20_ );
nand U130620 ( n66773, n73149, n67796 );
nand U130621 ( n67796, n67795, P2_P3_INSTADDRPOINTER_REG_20_ );
nand U130622 ( n24895, n73150, n25793 );
nand U130623 ( n25793, n25792, P1_P2_INSTADDRPOINTER_REG_20_ );
nand U130624 ( n58032, n73151, n58931 );
nand U130625 ( n58931, n58930, P2_P2_INSTADDRPOINTER_REG_20_ );
nand U130626 ( n42936, n42942, n42943 );
nand U130627 ( n42942, P2_P1_EBX_REG_15_, n42946 );
nand U130628 ( n42943, n42905, n42944 );
nand U130629 ( n42946, n42524, n42947 );
nand U130630 ( n43158, n43165, n43166 );
nand U130631 ( n43165, P2_P1_EBX_REG_7_, n43169 );
nand U130632 ( n43166, n43128, n43167 );
nand U130633 ( n43169, n42524, n43170 );
nand U130634 ( n43002, n43009, n43010 );
nand U130635 ( n43009, P2_P1_EBX_REG_13_, n43013 );
nand U130636 ( n43010, n42978, n43011 );
nand U130637 ( n43013, n42524, n43014 );
nand U130638 ( n42833, n42840, n42841 );
nand U130639 ( n42840, P2_P1_EBX_REG_19_, n42844 );
nand U130640 ( n42841, n42808, n42842 );
nand U130641 ( n42844, n42524, n42845 );
nand U130642 ( n12573, P1_P1_PHYADDRPOINTER_REG_2_, P1_P1_PHYADDRPOINTER_REG_1_ );
nand U130643 ( n16352, n16353, n16354 );
nand U130644 ( n16354, P1_P1_INSTQUEUE_REG_14__1_, n16340 );
nand U130645 ( n16353, n4797, n6 );
nand U130646 ( n16247, n16248, n16249 );
nand U130647 ( n16249, P1_P1_INSTQUEUE_REG_13__1_, n16235 );
nand U130648 ( n16248, n4798, n6 );
nand U130649 ( n16044, n16045, n16047 );
nand U130650 ( n16047, P1_P1_INSTQUEUE_REG_11__1_, n16033 );
nand U130651 ( n16045, n4799, n6 );
nand U130652 ( n15937, n15938, n15939 );
nand U130653 ( n15939, P1_P1_INSTQUEUE_REG_10__1_, n15925 );
nand U130654 ( n15938, n4800, n6 );
nand U130655 ( n15832, n15833, n15834 );
nand U130656 ( n15834, P1_P1_INSTQUEUE_REG_9__1_, n15820 );
nand U130657 ( n15833, n4802, n6 );
nand U130658 ( n15523, n15524, n15525 );
nand U130659 ( n15525, P1_P1_INSTQUEUE_REG_6__1_, n15512 );
nand U130660 ( n15524, n4804, n6 );
nand U130661 ( n15417, n15418, n15419 );
nand U130662 ( n15419, P1_P1_INSTQUEUE_REG_5__1_, n15405 );
nand U130663 ( n15418, n4805, n6 );
nand U130664 ( n15624, n15625, n15627 );
nand U130665 ( n15627, P1_P1_INSTQUEUE_REG_7__1_, n15609 );
nand U130666 ( n15625, n4803, n6 );
xor U130667 ( n48331, n62945, P3_REG3_REG_19_ );
nand U130668 ( n45270, n63315, n63316 );
nand U130669 ( n63315, P3_IR_REG_18_, n76840 );
nand U130670 ( n63316, n63317, P3_IR_REG_31_ );
and U130671 ( n63317, n13174, n13173 );
nand U130672 ( n13173, P3_IR_REG_18_, n63318 );
nand U130673 ( n63318, n848, n74418 );
nand U130674 ( n38569, n76446, P4_REG3_REG_2_ );
nor U130675 ( n57225, n57226, n74632 );
nor U130676 ( n57226, n57227, n57228 );
nor U130677 ( n57227, P2_P2_EAX_REG_9_, n76281 );
nor U130678 ( n24103, n24104, n74633 );
nor U130679 ( n24104, n24105, n24106 );
nor U130680 ( n24105, P1_P2_EAX_REG_9_, n76539 );
nor U130681 ( n31397, n31398, n74629 );
nor U130682 ( n31398, n31399, n31400 );
nor U130683 ( n31399, P1_P3_EAX_REG_9_, n76482 );
nor U130684 ( n65647, n65648, n74628 );
nor U130685 ( n65648, n65649, n65650 );
nor U130686 ( n65649, P2_P3_EAX_REG_9_, n76215 );
nor U130687 ( n31231, n31232, n75278 );
nor U130688 ( n31232, n31233, n31234 );
nor U130689 ( n31233, P1_P3_EAX_REG_13_, n76482 );
nor U130690 ( n31316, n31317, n75280 );
nor U130691 ( n31317, n31318, n31319 );
nor U130692 ( n31318, P1_P3_EAX_REG_11_, n76482 );
nor U130693 ( n57063, n57064, n75266 );
nor U130694 ( n57064, n57065, n57066 );
nor U130695 ( n57065, P2_P2_EAX_REG_13_, n76281 );
nor U130696 ( n57144, n57145, n75264 );
nor U130697 ( n57145, n57146, n57147 );
nor U130698 ( n57146, P2_P2_EAX_REG_11_, n76281 );
nor U130699 ( n57306, n57307, n75265 );
nor U130700 ( n57307, n57308, n57309 );
nor U130701 ( n57308, P2_P2_EAX_REG_7_, n76281 );
nor U130702 ( n57377, n57378, n75263 );
nor U130703 ( n57378, n57379, n57380 );
nor U130704 ( n57379, P2_P2_EAX_REG_5_, n76281 );
nor U130705 ( n57398, n57399, n75267 );
nor U130706 ( n57399, n57400, n57401 );
nor U130707 ( n57400, P2_P2_EAX_REG_3_, n76281 );
nor U130708 ( n57418, n57419, n75283 );
nor U130709 ( n57419, n57420, n57421 );
nor U130710 ( n57420, P2_P2_EAX_REG_1_, n76281 );
nor U130711 ( n31478, n31479, n75281 );
nor U130712 ( n31479, n31480, n31481 );
nor U130713 ( n31480, P1_P3_EAX_REG_7_, n76482 );
nor U130714 ( n31546, n31547, n75282 );
nor U130715 ( n31547, n31548, n31549 );
nor U130716 ( n31548, P1_P3_EAX_REG_5_, n76482 );
nor U130717 ( n31567, n31568, n75279 );
nor U130718 ( n31568, n31569, n31570 );
nor U130719 ( n31569, P1_P3_EAX_REG_3_, n76482 );
nor U130720 ( n31591, n31592, n75286 );
nor U130721 ( n31592, n31593, n31594 );
nor U130722 ( n31593, P1_P3_EAX_REG_1_, n76482 );
nor U130723 ( n24022, n24023, n75274 );
nor U130724 ( n24023, n24024, n24025 );
nor U130725 ( n24024, P1_P2_EAX_REG_11_, n76539 );
nor U130726 ( n23941, n23942, n75273 );
nor U130727 ( n23942, n23943, n23944 );
nor U130728 ( n23943, P1_P2_EAX_REG_13_, n76539 );
nor U130729 ( n24184, n24185, n75275 );
nor U130730 ( n24185, n24186, n24187 );
nor U130731 ( n24186, P1_P2_EAX_REG_7_, n76539 );
nor U130732 ( n24252, n24253, n75277 );
nor U130733 ( n24253, n24254, n24255 );
nor U130734 ( n24254, P1_P2_EAX_REG_5_, n76539 );
nor U130735 ( n24275, n24276, n75276 );
nor U130736 ( n24276, n24277, n24278 );
nor U130737 ( n24277, P1_P2_EAX_REG_3_, n76539 );
nor U130738 ( n24295, n24296, n75285 );
nor U130739 ( n24296, n24297, n24298 );
nor U130740 ( n24297, P1_P2_EAX_REG_1_, n76539 );
nor U130741 ( n65728, n65729, n75271 );
nor U130742 ( n65729, n65730, n65731 );
nor U130743 ( n65730, P2_P3_EAX_REG_7_, n76215 );
nor U130744 ( n65836, n65837, n75270 );
nor U130745 ( n65837, n65838, n65839 );
nor U130746 ( n65838, P2_P3_EAX_REG_5_, n76215 );
nor U130747 ( n65857, n65858, n75272 );
nor U130748 ( n65858, n65859, n65860 );
nor U130749 ( n65859, P2_P3_EAX_REG_3_, n76215 );
nor U130750 ( n65877, n65878, n75284 );
nor U130751 ( n65878, n65879, n65880 );
nor U130752 ( n65879, P2_P3_EAX_REG_1_, n76215 );
nor U130753 ( n65485, n65486, n75268 );
nor U130754 ( n65486, n65487, n65488 );
nor U130755 ( n65487, P2_P3_EAX_REG_13_, n76215 );
nor U130756 ( n65566, n65567, n75269 );
nor U130757 ( n65567, n65568, n65569 );
nor U130758 ( n65568, P2_P3_EAX_REG_11_, n76215 );
nand U130759 ( n38586, n76446, P4_REG3_REG_1_ );
nand U130760 ( n46202, P2_P1_PHYADDRPOINTER_REG_2_, P2_P1_PHYADDRPOINTER_REG_1_ );
nand U130761 ( n28551, P1_P2_INSTQUEUERD_ADDR_REG_3_, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U130762 ( n61856, P2_P2_INSTQUEUERD_ADDR_REG_3_, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U130763 ( n70456, P2_P3_INSTQUEUERD_ADDR_REG_3_, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130764 ( n35730, P1_P3_INSTQUEUERD_ADDR_REG_3_, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U130765 ( n32165, n32166, n32167 );
nand U130766 ( n32167, n32168, n76785 );
nand U130767 ( n32166, P1_P3_PHYADDRPOINTER_REG_19_, n32170 );
and U130768 ( n32168, n3139, n32169 );
nand U130769 ( n31869, n32578, P1_P3_STATEBS16_REG );
nor U130770 ( n32578, n3063, n73182 );
nand U130771 ( n31955, n31956, n31957 );
nand U130772 ( n31956, n3059, n29359 );
nand U130773 ( n31957, P1_P3_PHYADDRPOINTER_REG_28_, n31958 );
nand U130774 ( n31958, n3053, n31959 );
nand U130775 ( n45860, n45861, n45862 );
nand U130776 ( n45862, n45863, n76671 );
nand U130777 ( n45861, P2_P1_PHYADDRPOINTER_REG_19_, n45865 );
and U130778 ( n45863, n7525, n45864 );
nand U130779 ( n66811, n66812, n66813 );
nand U130780 ( n66813, n66814, n76719 );
nand U130781 ( n66812, P2_P3_PHYADDRPOINTER_REG_19_, n66816 );
and U130782 ( n66814, n5740, n66815 );
nand U130783 ( n24935, n24936, n24937 );
nand U130784 ( n24937, n24938, n76767 );
nand U130785 ( n24936, P1_P2_PHYADDRPOINTER_REG_19_, n24940 );
and U130786 ( n24938, n3983, n24939 );
nand U130787 ( n58070, n58071, n58072 );
nand U130788 ( n58072, n58073, n76700 );
nand U130789 ( n58071, P2_P2_PHYADDRPOINTER_REG_19_, n58075 );
and U130790 ( n58073, n6615, n58074 );
nand U130791 ( n66492, n67343, P2_P3_STATEBS16_REG );
nor U130792 ( n67343, n5664, n73183 );
nand U130793 ( n45567, n46282, P2_P1_STATEBS16_REG );
nor U130794 ( n46282, n7438, n74686 );
nand U130795 ( n24655, n25336, P1_P2_STATEBS16_REG );
nor U130796 ( n25336, n3907, n73181 );
nand U130797 ( n57791, n58475, P2_P2_STATEBS16_REG );
nor U130798 ( n58475, n6539, n73180 );
nand U130799 ( n24723, n24724, n24725 );
nand U130800 ( n24724, n3903, n22040 );
nand U130801 ( n24725, P1_P2_PHYADDRPOINTER_REG_28_, n24726 );
nand U130802 ( n24726, n3897, n24727 );
nand U130803 ( n66558, n66559, n66560 );
nand U130804 ( n66559, n5660, n63122 );
nand U130805 ( n66560, P2_P3_PHYADDRPOINTER_REG_28_, n66561 );
nand U130806 ( n66561, n5654, n66562 );
nand U130807 ( n57857, n57858, n57859 );
nand U130808 ( n57858, n6535, n55150 );
nand U130809 ( n57859, P2_P2_PHYADDRPOINTER_REG_28_, n57860 );
nand U130810 ( n57860, n6529, n57861 );
nand U130811 ( n32243, n32249, n32250 );
nand U130812 ( n32250, n32251, P1_P3_PHYADDRPOINTER_REG_15_ );
nand U130813 ( n32249, P1_P3_PHYADDRPOINTER_REG_16_, n32253 );
nor U130814 ( n32251, P1_P3_PHYADDRPOINTER_REG_16_, n3045 );
nand U130815 ( n32096, n32101, n32102 );
nand U130816 ( n32102, n32103, P1_P3_PHYADDRPOINTER_REG_21_ );
nand U130817 ( n32101, P1_P3_PHYADDRPOINTER_REG_22_, n32105 );
and U130818 ( n32103, n75239, n32104 );
nand U130819 ( n41460, n70970, n70971 );
nand U130820 ( n70970, P3_IR_REG_23_, n76842 );
nand U130821 ( n70971, n70972, P3_IR_REG_31_ );
and U130822 ( n70972, n11633, n11632 );
nand U130823 ( n45931, n45937, n45938 );
nand U130824 ( n45938, n45939, P2_P1_PHYADDRPOINTER_REG_15_ );
nand U130825 ( n45937, P2_P1_PHYADDRPOINTER_REG_16_, n45941 );
nor U130826 ( n45939, P2_P1_PHYADDRPOINTER_REG_16_, n7422 );
nand U130827 ( n66882, n66888, n66889 );
nand U130828 ( n66889, n66890, P2_P3_PHYADDRPOINTER_REG_15_ );
nand U130829 ( n66888, P2_P3_PHYADDRPOINTER_REG_16_, n66892 );
nor U130830 ( n66890, P2_P3_PHYADDRPOINTER_REG_16_, n5647 );
nand U130831 ( n25006, n25012, n25013 );
nand U130832 ( n25013, n25014, P1_P2_PHYADDRPOINTER_REG_15_ );
nand U130833 ( n25012, P1_P2_PHYADDRPOINTER_REG_16_, n25016 );
nor U130834 ( n25014, P1_P2_PHYADDRPOINTER_REG_16_, n3889 );
nand U130835 ( n58141, n58147, n58148 );
nand U130836 ( n58148, n58149, P2_P2_PHYADDRPOINTER_REG_15_ );
nand U130837 ( n58147, P2_P2_PHYADDRPOINTER_REG_16_, n58151 );
nor U130838 ( n58149, P2_P2_PHYADDRPOINTER_REG_16_, n6522 );
nand U130839 ( n45634, n45635, n45636 );
nand U130840 ( n45635, n7434, n7959 );
nand U130841 ( n45636, P2_P1_PHYADDRPOINTER_REG_28_, n45637 );
nand U130842 ( n45637, n7429, n45638 );
nand U130843 ( n66699, n66704, n66705 );
nand U130844 ( n66705, n66706, P2_P3_PHYADDRPOINTER_REG_21_ );
nand U130845 ( n66704, P2_P3_PHYADDRPOINTER_REG_22_, n66708 );
and U130846 ( n66706, n75240, n66707 );
nand U130847 ( n24864, n24869, n24870 );
nand U130848 ( n24870, n24871, P1_P2_PHYADDRPOINTER_REG_21_ );
nand U130849 ( n24869, P1_P2_PHYADDRPOINTER_REG_22_, n24873 );
and U130850 ( n24871, n75241, n24872 );
nand U130851 ( n58001, n58006, n58007 );
nand U130852 ( n58007, n58008, P2_P2_PHYADDRPOINTER_REG_21_ );
nand U130853 ( n58006, P2_P2_PHYADDRPOINTER_REG_22_, n58010 );
and U130854 ( n58008, n75242, n58009 );
nand U130855 ( n32307, n32314, n32315 );
nand U130856 ( n32315, n32316, P1_P3_PHYADDRPOINTER_REG_12_ );
nand U130857 ( n32314, P1_P3_PHYADDRPOINTER_REG_13_, n32318 );
nor U130858 ( n32316, P1_P3_PHYADDRPOINTER_REG_13_, n3044 );
nand U130859 ( n45791, n45796, n45797 );
nand U130860 ( n45797, n45798, P2_P1_PHYADDRPOINTER_REG_21_ );
nand U130861 ( n45796, P2_P1_PHYADDRPOINTER_REG_22_, n45800 );
and U130862 ( n45798, n74680, n45799 );
nand U130863 ( n66946, n66953, n66954 );
nand U130864 ( n66954, n66955, P2_P3_PHYADDRPOINTER_REG_12_ );
nand U130865 ( n66953, P2_P3_PHYADDRPOINTER_REG_13_, n66957 );
nor U130866 ( n66955, P2_P3_PHYADDRPOINTER_REG_13_, n5645 );
nand U130867 ( n46006, n46013, n46014 );
nand U130868 ( n46014, n46015, P2_P1_PHYADDRPOINTER_REG_12_ );
nand U130869 ( n46013, P2_P1_PHYADDRPOINTER_REG_13_, n46017 );
nor U130870 ( n46015, P2_P1_PHYADDRPOINTER_REG_13_, n7420 );
nand U130871 ( n25070, n25077, n25078 );
nand U130872 ( n25078, n25079, P1_P2_PHYADDRPOINTER_REG_12_ );
nand U130873 ( n25077, P1_P2_PHYADDRPOINTER_REG_13_, n25081 );
nor U130874 ( n25079, P1_P2_PHYADDRPOINTER_REG_13_, n3888 );
nand U130875 ( n58205, n58212, n58213 );
nand U130876 ( n58213, n58214, P2_P2_PHYADDRPOINTER_REG_12_ );
nand U130877 ( n58212, P2_P2_PHYADDRPOINTER_REG_13_, n58216 );
nor U130878 ( n58214, P2_P2_PHYADDRPOINTER_REG_13_, n6520 );
nor U130879 ( n44136, n44889, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nor U130880 ( n32496, n32514, n32515 );
nor U130881 ( n32515, n31869, P1_P3_PHYADDRPOINTER_REG_3_ );
nand U130882 ( n32485, n32491, n32492 );
nand U130883 ( n32492, n32493, n32494 );
nand U130884 ( n32491, P1_P3_PHYADDRPOINTER_REG_5_, n32495 );
nor U130885 ( n32493, P1_P3_PHYADDRPOINTER_REG_5_, n74478 );
nor U130886 ( n67152, n67170, n67171 );
nor U130887 ( n67171, n66492, P2_P3_PHYADDRPOINTER_REG_3_ );
nor U130888 ( n25254, n25272, n25273 );
nor U130889 ( n25273, n24655, P1_P2_PHYADDRPOINTER_REG_3_ );
nor U130890 ( n58390, n58408, n58409 );
nor U130891 ( n58409, n57791, P2_P2_PHYADDRPOINTER_REG_3_ );
nor U130892 ( n46188, n46206, n46207 );
nor U130893 ( n46207, n45567, P2_P1_PHYADDRPOINTER_REG_3_ );
nand U130894 ( n67141, n67147, n67148 );
nand U130895 ( n67148, n67149, n67150 );
nand U130896 ( n67147, P2_P3_PHYADDRPOINTER_REG_5_, n67151 );
nor U130897 ( n67149, P2_P3_PHYADDRPOINTER_REG_5_, n74479 );
nand U130898 ( n25243, n25249, n25250 );
nand U130899 ( n25250, n25251, n25252 );
nand U130900 ( n25249, P1_P2_PHYADDRPOINTER_REG_5_, n25253 );
nor U130901 ( n25251, P1_P2_PHYADDRPOINTER_REG_5_, n74480 );
nand U130902 ( n58379, n58385, n58386 );
nand U130903 ( n58386, n58387, n58388 );
nand U130904 ( n58385, P2_P2_PHYADDRPOINTER_REG_5_, n58389 );
nor U130905 ( n58387, P2_P2_PHYADDRPOINTER_REG_5_, n74481 );
nand U130906 ( n46177, n46183, n46184 );
nand U130907 ( n46184, n46185, n46186 );
nand U130908 ( n46183, P2_P1_PHYADDRPOINTER_REG_5_, n46187 );
nor U130909 ( n46185, P2_P1_PHYADDRPOINTER_REG_5_, n74473 );
nor U130910 ( n72843, n74403, n71104 );
nand U130911 ( n54347, n44136, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U130912 ( n12142, n12143, n12144 );
nand U130913 ( n12143, P1_P1_PHYADDRPOINTER_REG_19_, n12148 );
nand U130914 ( n12144, n12145, n76738 );
nand U130915 ( n12148, n4782, n12149 );
nand U130916 ( n11076, n68302, n68303 );
nand U130917 ( n68303, n76195, P2_P3_INSTADDRPOINTER_REG_7_ );
nor U130918 ( n68302, n68304, n68305 );
nor U130919 ( n68305, n72966, n76871 );
nand U130920 ( n6586, n26301, n26302 );
nand U130921 ( n26302, n76519, P1_P2_INSTADDRPOINTER_REG_7_ );
nor U130922 ( n26301, n26303, n26304 );
nor U130923 ( n26304, n73199, n76906 );
nand U130924 ( n13321, n59440, n59441 );
nand U130925 ( n59441, n76261, P2_P2_INSTADDRPOINTER_REG_7_ );
nor U130926 ( n59440, n59442, n59443 );
nor U130927 ( n59443, n73198, n76880 );
nand U130928 ( n15566, n47271, n47272 );
nand U130929 ( n47272, n76861, P2_P1_INSTADDRPOINTER_REG_7_ );
nor U130930 ( n47271, n47273, n47274 );
nor U130931 ( n47274, n73206, n76332 );
nand U130932 ( n4341, n33546, n33547 );
nand U130933 ( n33547, n76468, P1_P3_INSTADDRPOINTER_REG_7_ );
nor U130934 ( n33546, n33548, n33549 );
nor U130935 ( n33549, n72967, n76897 );
nand U130936 ( n17063, n17054, P4_DATAO_REG_6_ );
nand U130937 ( n11877, n76603, P1_P1_INSTADDRPOINTER_REG_27_ );
nand U130938 ( n54338, n44132, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U130939 ( n9308, n9309, n9310 );
nand U130940 ( n9309, P1_P1_EBX_REG_3_, n9314 );
nand U130941 ( n9310, n9287, n9312 );
nand U130942 ( n9314, n8428, n9315 );
nor U130943 ( n32436, n32460, n32461 );
nor U130944 ( n32461, n31869, P1_P3_PHYADDRPOINTER_REG_6_ );
nand U130945 ( n32425, n32431, n32432 );
nand U130946 ( n32432, n32433, n32434 );
nand U130947 ( n32431, P1_P3_PHYADDRPOINTER_REG_8_, n32435 );
nor U130948 ( n32433, P1_P3_PHYADDRPOINTER_REG_8_, n73102 );
xor U130949 ( n33479, n76471, P1_P3_INSTADDRPOINTER_REG_9_ );
nor U130950 ( n67092, n67116, n67117 );
nor U130951 ( n67117, n66492, P2_P3_PHYADDRPOINTER_REG_6_ );
nor U130952 ( n32365, n32392, n32393 );
nor U130953 ( n32393, n31869, P1_P3_PHYADDRPOINTER_REG_9_ );
nor U130954 ( n46128, n46152, n46153 );
nor U130955 ( n46153, n45567, P2_P1_PHYADDRPOINTER_REG_6_ );
nor U130956 ( n25194, n25218, n25219 );
nor U130957 ( n25219, n24655, P1_P2_PHYADDRPOINTER_REG_6_ );
nor U130958 ( n58330, n58354, n58355 );
nor U130959 ( n58355, n57791, P2_P2_PHYADDRPOINTER_REG_6_ );
nand U130960 ( n67081, n67087, n67088 );
nand U130961 ( n67088, n67089, n67090 );
nand U130962 ( n67087, P2_P3_PHYADDRPOINTER_REG_8_, n67091 );
nor U130963 ( n67089, P2_P3_PHYADDRPOINTER_REG_8_, n73100 );
nand U130964 ( n25183, n25189, n25190 );
nand U130965 ( n25190, n25191, n25192 );
nand U130966 ( n25189, P1_P2_PHYADDRPOINTER_REG_8_, n25193 );
nor U130967 ( n25191, P1_P2_PHYADDRPOINTER_REG_8_, n73103 );
nand U130968 ( n58319, n58325, n58326 );
nand U130969 ( n58326, n58327, n58328 );
nand U130970 ( n58325, P2_P2_PHYADDRPOINTER_REG_8_, n58329 );
nor U130971 ( n58327, P2_P2_PHYADDRPOINTER_REG_8_, n73101 );
nand U130972 ( n32354, n32360, n32361 );
nand U130973 ( n32361, n32362, n32363 );
nand U130974 ( n32360, P1_P3_PHYADDRPOINTER_REG_11_, n32364 );
nor U130975 ( n32362, P1_P3_PHYADDRPOINTER_REG_11_, n74557 );
nand U130976 ( n46117, n46123, n46124 );
nand U130977 ( n46124, n46125, n46126 );
nand U130978 ( n46123, P2_P1_PHYADDRPOINTER_REG_8_, n46127 );
nor U130979 ( n46125, P2_P1_PHYADDRPOINTER_REG_8_, n73098 );
nor U130980 ( n67028, n67055, n67056 );
nor U130981 ( n67056, n66492, P2_P3_PHYADDRPOINTER_REG_9_ );
nor U130982 ( n46064, n46091, n46092 );
nor U130983 ( n46092, n45567, P2_P1_PHYADDRPOINTER_REG_9_ );
nor U130984 ( n25128, n25155, n25156 );
nor U130985 ( n25156, n24655, P1_P2_PHYADDRPOINTER_REG_9_ );
nor U130986 ( n58266, n58293, n58294 );
nor U130987 ( n58294, n57791, P2_P2_PHYADDRPOINTER_REG_9_ );
nand U130988 ( n46053, n46059, n46060 );
nand U130989 ( n46060, n46061, n46062 );
nand U130990 ( n46059, P2_P1_PHYADDRPOINTER_REG_11_, n46063 );
nor U130991 ( n46061, P2_P1_PHYADDRPOINTER_REG_11_, n74554 );
nand U130992 ( n67017, n67023, n67024 );
nand U130993 ( n67024, n67025, n67026 );
nand U130994 ( n67023, P2_P3_PHYADDRPOINTER_REG_11_, n67027 );
nor U130995 ( n67025, P2_P3_PHYADDRPOINTER_REG_11_, n74558 );
nand U130996 ( n25117, n25123, n25124 );
nand U130997 ( n25124, n25125, n25126 );
nand U130998 ( n25123, P1_P2_PHYADDRPOINTER_REG_11_, n25127 );
nor U130999 ( n25125, P1_P2_PHYADDRPOINTER_REG_11_, n74559 );
nand U131000 ( n58255, n58261, n58262 );
nand U131001 ( n58262, n58263, n58264 );
nand U131002 ( n58261, P2_P2_PHYADDRPOINTER_REG_11_, n58265 );
nor U131003 ( n58263, P2_P2_PHYADDRPOINTER_REG_11_, n74560 );
nand U131004 ( n43331, P2_P1_INSTQUEUERD_ADDR_REG_1_, n73512 );
nand U131005 ( n11810, n12667, P1_P1_STATEBS16_REG );
nor U131006 ( n12667, n4794, n74685 );
nand U131007 ( n11858, n11859, n11860 );
nand U131008 ( n11859, n4790, n5304 );
nand U131009 ( n11860, P1_P1_PHYADDRPOINTER_REG_28_, n11862 );
nand U131010 ( n11862, n4785, n11863 );
nand U131011 ( n9050, n9060, n9062 );
nand U131012 ( n9060, P1_P1_EBX_REG_11_, n9065 );
nand U131013 ( n9062, n9025, n9063 );
nand U131014 ( n9065, n8428, n9067 );
nand U131015 ( n9245, n9254, n9255 );
nand U131016 ( n9254, P1_P1_EBX_REG_5_, n9259 );
nand U131017 ( n9255, n9220, n9257 );
nand U131018 ( n9259, n8428, n9260 );
xor U131019 ( n38259, n39273, P4_REG3_REG_21_ );
nand U131020 ( n32174, n32175, P1_P3_PHYADDRPOINTER_REG_18_ );
nor U131021 ( n32175, P1_P3_PHYADDRPOINTER_REG_19_, n3048 );
not U131022 ( n3048, n32176 );
nand U131023 ( n11632, P3_IR_REG_23_, n67314 );
nand U131024 ( n66820, n66821, P2_P3_PHYADDRPOINTER_REG_18_ );
nor U131025 ( n66821, P2_P3_PHYADDRPOINTER_REG_19_, n5649 );
not U131026 ( n5649, n66822 );
nand U131027 ( n24944, n24945, P1_P2_PHYADDRPOINTER_REG_18_ );
nor U131028 ( n24945, P1_P2_PHYADDRPOINTER_REG_19_, n3892 );
not U131029 ( n3892, n24946 );
nand U131030 ( n58079, n58080, P2_P2_PHYADDRPOINTER_REG_18_ );
nor U131031 ( n58080, P2_P2_PHYADDRPOINTER_REG_19_, n6524 );
not U131032 ( n6524, n58081 );
nand U131033 ( n43272, n43273, n43274 );
nand U131034 ( n43273, P2_P1_EBX_REG_3_, n43277 );
nand U131035 ( n43274, n43255, n43275 );
nand U131036 ( n43277, n42524, n43278 );
nand U131037 ( n45869, n45870, P2_P1_PHYADDRPOINTER_REG_18_ );
nor U131038 ( n45870, P2_P1_PHYADDRPOINTER_REG_19_, n7424 );
not U131039 ( n7424, n45871 );
nand U131040 ( n11959, P1_P1_PHYADDRPOINTER_REG_25_, n11964 );
nand U131041 ( n11964, n4784, n11965 );
nand U131042 ( n11965, n11772, n74737 );
not U131043 ( n4784, n11967 );
nand U131044 ( n12242, n12249, n12250 );
nand U131045 ( n12250, n12252, P1_P1_PHYADDRPOINTER_REG_15_ );
nand U131046 ( n12249, P1_P1_PHYADDRPOINTER_REG_16_, n12254 );
nor U131047 ( n12252, P1_P1_PHYADDRPOINTER_REG_16_, n4778 );
nand U131048 ( n12050, n12057, n12058 );
nand U131049 ( n12058, n12059, P1_P1_PHYADDRPOINTER_REG_21_ );
nand U131050 ( n12057, P1_P1_PHYADDRPOINTER_REG_22_, n12062 );
and U131051 ( n12059, n74677, n12060 );
nand U131052 ( n12322, n12330, n12332 );
nand U131053 ( n12332, n12333, P1_P1_PHYADDRPOINTER_REG_12_ );
nand U131054 ( n12330, P1_P1_PHYADDRPOINTER_REG_13_, n12335 );
nor U131055 ( n12333, P1_P1_PHYADDRPOINTER_REG_13_, n4777 );
nor U131056 ( n10265, n11178, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131057 ( n28638, n28909, n28910 );
nand U131058 ( n28909, n28912, n74612 );
nand U131059 ( n28910, P1_P2_INSTQUEUEWR_ADDR_REG_4_, n28911 );
nand U131060 ( n28911, P1_P2_INSTQUEUERD_ADDR_REG_4_, n4230 );
nand U131061 ( n61943, n62214, n62215 );
nand U131062 ( n62214, n62217, n74614 );
nand U131063 ( n62215, P2_P2_INSTQUEUEWR_ADDR_REG_4_, n62216 );
nand U131064 ( n62216, P2_P2_INSTQUEUERD_ADDR_REG_4_, n6863 );
nand U131065 ( n43052, n43060, n43061 );
nand U131066 ( n43060, P2_P1_EBX_REG_11_, n43064 );
nand U131067 ( n43061, n43032, n43062 );
nand U131068 ( n43064, n42524, n43065 );
nand U131069 ( n43208, n43215, n43216 );
nand U131070 ( n43215, P2_P1_EBX_REG_5_, n43219 );
nand U131071 ( n43216, n43188, n43217 );
nand U131072 ( n43219, n42524, n43220 );
nand U131073 ( n70543, n70814, n70815 );
nand U131074 ( n70814, n70817, n74613 );
nand U131075 ( n70815, P2_P3_INSTQUEUEWR_ADDR_REG_4_, n70816 );
nand U131076 ( n70816, P2_P3_INSTQUEUERD_ADDR_REG_4_, n6008 );
nand U131077 ( n35817, n36088, n36089 );
nand U131078 ( n36088, n36091, n74611 );
nand U131079 ( n36089, P1_P3_INSTQUEUEWR_ADDR_REG_4_, n36090 );
nand U131080 ( n36090, P1_P3_INSTQUEUERD_ADDR_REG_4_, n3393 );
nand U131081 ( n8422, n8432, n8433 );
nand U131082 ( n8433, n8434, P1_P1_REIP_REG_29_ );
nand U131083 ( n8432, n5305, n8437 );
nor U131084 ( n8434, P1_P1_REIP_REG_30_, n237 );
nand U131085 ( n21364, n10265, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U131086 ( n9256, n11519, n11520 );
nand U131087 ( n11520, P1_P1_UWORD_REG_2_, n76618 );
nor U131088 ( n11519, n11522, n11523 );
nor U131089 ( n11522, n73266, n76617 );
nand U131090 ( n9181, n11602, n11603 );
nand U131091 ( n11603, P1_P1_LWORD_REG_2_, n76618 );
nor U131092 ( n11602, n11604, n11523 );
nor U131093 ( n11604, n73166, n76616 );
nor U131094 ( n12555, n12578, n12579 );
nor U131095 ( n12579, n11810, P1_P1_PHYADDRPOINTER_REG_3_ );
nand U131096 ( n12542, n12549, n12550 );
nand U131097 ( n12550, n12552, n12553 );
nand U131098 ( n12549, P1_P1_PHYADDRPOINTER_REG_5_, n12554 );
nor U131099 ( n12552, P1_P1_PHYADDRPOINTER_REG_5_, n74484 );
nand U131100 ( n9367, n9368, n9369 );
nand U131101 ( n9369, P1_P1_EBX_REG_1_, n9370 );
nand U131102 ( n9368, n9373, n74477 );
nand U131103 ( n9370, n8428, n9372 );
nand U131104 ( n23633, n23634, n23635 );
nand U131105 ( n23634, P1_P2_EAX_REG_20_, n23638 );
nand U131106 ( n23635, n23636, n23637 );
nand U131107 ( n23638, n154, n23639 );
nand U131108 ( n23722, n23723, n23724 );
nand U131109 ( n23723, P1_P2_EAX_REG_18_, n23727 );
nand U131110 ( n23724, n23725, n23726 );
nand U131111 ( n23727, n153, n23728 );
nand U131112 ( n23544, n23545, n23546 );
nand U131113 ( n23545, P1_P2_EAX_REG_22_, n23549 );
nand U131114 ( n23546, n23547, n23548 );
nand U131115 ( n23549, n155, n23550 );
nand U131116 ( n56755, n56756, n56757 );
nand U131117 ( n56756, P2_P2_EAX_REG_20_, n56760 );
nand U131118 ( n56757, n56758, n56759 );
nand U131119 ( n56760, n427, n56761 );
nand U131120 ( n56666, n56667, n56668 );
nand U131121 ( n56667, P2_P2_EAX_REG_22_, n56671 );
nand U131122 ( n56668, n56669, n56670 );
nand U131123 ( n56671, n428, n56672 );
nand U131124 ( n56844, n56845, n56846 );
nand U131125 ( n56845, P2_P2_EAX_REG_18_, n56849 );
nand U131126 ( n56846, n56847, n56848 );
nand U131127 ( n56849, n425, n56850 );
nand U131128 ( n23811, n23812, n23813 );
nand U131129 ( n23812, P1_P2_EAX_REG_16_, n23816 );
nand U131130 ( n23813, n23814, n23815 );
nand U131131 ( n23816, n23817, n23818 );
nand U131132 ( n56936, n56937, n56938 );
nand U131133 ( n56937, P2_P2_EAX_REG_16_, n56941 );
nand U131134 ( n56938, n56939, n56940 );
nand U131135 ( n56941, n56942, n56943 );
nand U131136 ( n23300, n23301, n23302 );
nand U131137 ( n23301, P1_P2_EAX_REG_26_, n23305 );
nand U131138 ( n23302, n23303, n23304 );
nand U131139 ( n23305, n158, n23306 );
nand U131140 ( n23397, n23398, n23399 );
nand U131141 ( n23398, P1_P2_EAX_REG_24_, n23402 );
nand U131142 ( n23399, n23400, n23401 );
nand U131143 ( n23402, n157, n23403 );
nand U131144 ( n31108, n31109, n31110 );
nand U131145 ( n31109, P1_P3_EAX_REG_16_, n31113 );
nand U131146 ( n31110, n31111, n31112 );
nand U131147 ( n31113, n31114, n31115 );
nand U131148 ( n56424, n56425, n56426 );
nand U131149 ( n56425, P2_P2_EAX_REG_26_, n56429 );
nand U131150 ( n56426, n56427, n56428 );
nand U131151 ( n56429, n430, n56430 );
nand U131152 ( n65362, n65363, n65364 );
nand U131153 ( n65363, P2_P3_EAX_REG_16_, n65367 );
nand U131154 ( n65364, n65365, n65366 );
nand U131155 ( n65367, n65368, n65369 );
nand U131156 ( n56519, n56520, n56521 );
nand U131157 ( n56520, P2_P2_EAX_REG_24_, n56524 );
nand U131158 ( n56521, n56522, n56523 );
nand U131159 ( n56524, n429, n56525 );
nand U131160 ( n65055, n65056, n65057 );
nand U131161 ( n65056, P2_P3_EAX_REG_22_, n65060 );
nand U131162 ( n65057, n65058, n65059 );
nand U131163 ( n65060, n464, n65061 );
nand U131164 ( n65140, n65141, n65142 );
nand U131165 ( n65141, P2_P3_EAX_REG_20_, n65145 );
nand U131166 ( n65142, n65143, n65144 );
nand U131167 ( n65145, n463, n65146 );
nand U131168 ( n65225, n65226, n65227 );
nand U131169 ( n65226, P2_P3_EAX_REG_18_, n65230 );
nand U131170 ( n65227, n65228, n65229 );
nand U131171 ( n65230, n462, n65231 );
nand U131172 ( n31023, n31024, n31025 );
nand U131173 ( n31024, P1_P3_EAX_REG_18_, n31028 );
nand U131174 ( n31025, n31026, n31027 );
nand U131175 ( n31028, n190, n31029 );
nand U131176 ( n30938, n30939, n30940 );
nand U131177 ( n30939, P1_P3_EAX_REG_20_, n30943 );
nand U131178 ( n30940, n30941, n30942 );
nand U131179 ( n30943, n192, n30944 );
nand U131180 ( n30853, n30854, n30855 );
nand U131181 ( n30854, P1_P3_EAX_REG_22_, n30858 );
nand U131182 ( n30855, n30856, n30857 );
nand U131183 ( n30858, n193, n30859 );
nand U131184 ( n64824, n64825, n64826 );
nand U131185 ( n64825, P2_P3_EAX_REG_26_, n64829 );
nand U131186 ( n64826, n64827, n64828 );
nand U131187 ( n64829, n467, n64830 );
nand U131188 ( n64913, n64914, n64915 );
nand U131189 ( n64914, P2_P3_EAX_REG_24_, n64918 );
nand U131190 ( n64915, n64916, n64917 );
nand U131191 ( n64918, n465, n64919 );
nand U131192 ( n30618, n30619, n30620 );
nand U131193 ( n30619, P1_P3_EAX_REG_26_, n30623 );
nand U131194 ( n30620, n30621, n30622 );
nand U131195 ( n30623, n195, n30624 );
nand U131196 ( n30707, n30708, n30709 );
nand U131197 ( n30708, P1_P3_EAX_REG_24_, n30712 );
nand U131198 ( n30709, n30710, n30711 );
nand U131199 ( n30712, n194, n30713 );
nand U131200 ( n21355, n10260, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
xnor U131201 ( n38275, P4_REG3_REG_20_, n39340 );
nor U131202 ( n44133, n43331, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131203 ( n49730, n50007, P3_DATAO_REG_7_ );
nand U131204 ( n43319, n43320, n43321 );
nand U131205 ( n43321, P2_P1_EBX_REG_1_, n43322 );
nand U131206 ( n43320, n43324, n74467 );
nand U131207 ( n43322, n42524, n43323 );
nand U131208 ( n9382, P1_P1_INSTQUEUERD_ADDR_REG_1_, n73533 );
nor U131209 ( n12480, n12510, n12512 );
nor U131210 ( n12512, n11810, P1_P1_PHYADDRPOINTER_REG_6_ );
nand U131211 ( n12467, n12474, n12475 );
nand U131212 ( n12475, n12477, n12478 );
nand U131213 ( n12474, P1_P1_PHYADDRPOINTER_REG_8_, n12479 );
nor U131214 ( n12477, P1_P1_PHYADDRPOINTER_REG_8_, n73097 );
nor U131215 ( n12394, n12434, n12435 );
nor U131216 ( n12435, n11810, P1_P1_PHYADDRPOINTER_REG_9_ );
nand U131217 ( n12380, n12388, n12389 );
nand U131218 ( n12389, n12390, n12392 );
nand U131219 ( n12388, P1_P1_PHYADDRPOINTER_REG_11_, n12393 );
nor U131220 ( n12390, P1_P1_PHYADDRPOINTER_REG_11_, n74577 );
nand U131221 ( n17129, DIN_25_, n76928 );
nand U131222 ( n17697, n8212, P4_DATAO_REG_2_ );
nand U131223 ( n9238, n9239, n9240 );
nand U131224 ( n9239, n9243, n76890 );
nand U131225 ( n9240, n9242, n76744 );
nor U131226 ( n9243, P1_P1_EBX_REG_5_, n5464 );
nand U131227 ( n8849, n8850, n8852 );
nand U131228 ( n8850, P1_P1_EBX_REG_17_, n8854 );
nand U131229 ( n8852, n8853, n76743 );
nand U131230 ( n8854, n8428, n8855 );
nand U131231 ( n12153, n12154, P1_P1_PHYADDRPOINTER_REG_18_ );
nor U131232 ( n12154, P1_P1_PHYADDRPOINTER_REG_19_, n4780 );
not U131233 ( n4780, n12155 );
nand U131234 ( n43330, P2_P1_INSTQUEUERD_ADDR_REG_0_, n73052 );
nor U131235 ( n44137, n43330, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131236 ( n9307, n9317, n9318 );
nand U131237 ( n9318, n9319, n76890 );
nand U131238 ( n9317, n9320, n76744 );
nor U131239 ( n9319, P1_P1_EBX_REG_3_, n5465 );
nand U131240 ( n9337, n9348, n9349 );
nand U131241 ( n9349, n9333, P1_P1_REIP_REG_1_ );
nand U131242 ( n9348, n9350, n76744 );
nor U131243 ( n9350, n5285, n9352 );
nand U131244 ( n8914, n8915, n8917 );
nand U131245 ( n8917, n8918, n76889 );
nand U131246 ( n8915, n8919, n76743 );
nor U131247 ( n8918, P1_P1_EBX_REG_15_, n5458 );
nand U131248 ( n9173, n9174, n9175 );
nand U131249 ( n9175, n9177, n76890 );
nand U131250 ( n9174, n9178, n76743 );
nor U131251 ( n9177, P1_P1_EBX_REG_7_, n5463 );
nand U131252 ( n9043, n9044, n9045 );
nand U131253 ( n9045, n9047, n76889 );
nand U131254 ( n9044, n9048, n76743 );
nor U131255 ( n9047, P1_P1_EBX_REG_11_, n5460 );
nand U131256 ( n8978, n8979, n8980 );
nand U131257 ( n8980, n8982, n76889 );
nand U131258 ( n8979, n8983, n76743 );
nor U131259 ( n8982, P1_P1_EBX_REG_13_, n5459 );
nand U131260 ( n8782, n8783, n8784 );
nand U131261 ( n8784, n8785, n76889 );
nand U131262 ( n8783, n8787, n76742 );
nor U131263 ( n8785, P1_P1_EBX_REG_19_, n5455 );
nand U131264 ( n8654, n8664, n8665 );
nand U131265 ( n8665, n8667, n76889 );
nand U131266 ( n8664, n8668, n76742 );
nor U131267 ( n8667, P1_P1_EBX_REG_23_, n5453 );
nand U131268 ( n54351, n44137, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U131269 ( n8489, n8504, n8505 );
nand U131270 ( n8505, n8507, n8508 );
nand U131271 ( n8504, n8510, n76742 );
nor U131272 ( n8508, P1_P1_REIP_REG_28_, n73309 );
nand U131273 ( n8682, n8697, n8698 );
nand U131274 ( n8698, n8699, n8700 );
nand U131275 ( n8697, n8703, n76742 );
nor U131276 ( n8700, P1_P1_REIP_REG_22_, n74952 );
nand U131277 ( n8851, n13702, n13703 );
nand U131278 ( n13703, n76887, P1_P1_INSTADDRPOINTER_REG_11_ );
nor U131279 ( n13702, n13704, n13705 );
nor U131280 ( n13705, n74812, n76598 );
nand U131281 ( n31835, P1_P3_PHYADDRPOINTER_REG_31_, n31839 );
nand U131282 ( n31839, n3057, n31840 );
nand U131283 ( n31840, n31841, n75185 );
not U131284 ( n3057, n31842 );
nand U131285 ( n43202, n43203, n43204 );
nand U131286 ( n43203, n43206, n76863 );
nand U131287 ( n43204, n43205, n76677 );
nor U131288 ( n43206, P2_P1_EBX_REG_5_, n8118 );
nand U131289 ( n24621, P1_P2_PHYADDRPOINTER_REG_31_, n24625 );
nand U131290 ( n24625, n3900, n24626 );
nand U131291 ( n24626, n24627, n75186 );
not U131292 ( n3900, n24628 );
nand U131293 ( n57753, P2_P2_PHYADDRPOINTER_REG_31_, n57757 );
nand U131294 ( n57757, n6533, n57758 );
nand U131295 ( n57758, n57759, n75187 );
not U131296 ( n6533, n57760 );
nand U131297 ( n66458, P2_P3_PHYADDRPOINTER_REG_31_, n66462 );
nand U131298 ( n66462, n5658, n66463 );
nand U131299 ( n66463, n66464, n75188 );
not U131300 ( n5658, n66465 );
nand U131301 ( n9441, n11284, n11285 );
nor U131302 ( n11285, n11287, n11288 );
nor U131303 ( n11284, n11292, n11293 );
nor U131304 ( n11287, P1_P1_EAX_REG_2_, n11279 );
nor U131305 ( n10262, n9382, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131306 ( n42877, n42878, n42879 );
nand U131307 ( n42878, P2_P1_EBX_REG_17_, n42881 );
nand U131308 ( n42879, n42880, n76676 );
nand U131309 ( n42881, n42524, n42882 );
nand U131310 ( n31990, P1_P3_PHYADDRPOINTER_REG_26_, n31997 );
nand U131311 ( n31997, n31998, n31999 );
nor U131312 ( n31998, n32000, n32001 );
nor U131313 ( n32001, n31977, n31861 );
nand U131314 ( n45534, P2_P1_PHYADDRPOINTER_REG_31_, n45538 );
nand U131315 ( n45538, n7432, n45539 );
nand U131316 ( n45539, n45540, n74931 );
not U131317 ( n7432, n45541 );
nand U131318 ( n43150, n43151, n43152 );
nand U131319 ( n43152, n43153, n76862 );
nand U131320 ( n43151, n43154, n76677 );
nor U131321 ( n43153, P2_P1_EBX_REG_7_, n8117 );
nand U131322 ( n66593, P2_P3_PHYADDRPOINTER_REG_26_, n66600 );
nand U131323 ( n66600, n66601, n66602 );
nor U131324 ( n66601, n66603, n66604 );
nor U131325 ( n66604, n66580, n66484 );
nand U131326 ( n24758, P1_P2_PHYADDRPOINTER_REG_26_, n24765 );
nand U131327 ( n24765, n24766, n24767 );
nor U131328 ( n24766, n24768, n24769 );
nor U131329 ( n24769, n24745, n24647 );
nand U131330 ( n57892, P2_P2_PHYADDRPOINTER_REG_26_, n57899 );
nand U131331 ( n57899, n57900, n57901 );
nor U131332 ( n57900, n57902, n57903 );
nor U131333 ( n57903, n57879, n57783 );
nand U131334 ( n45764, P2_P1_PHYADDRPOINTER_REG_23_, n45771 );
nand U131335 ( n45771, n45772, n45773 );
nor U131336 ( n45772, n45774, n45775 );
nor U131337 ( n45775, n45733, n45559 );
nand U131338 ( n46316, P2_P1_INSTADDRPOINTER_REG_31_, n76342 );
nand U131339 ( n31882, P1_P3_PHYADDRPOINTER_REG_29_, n31889 );
nand U131340 ( n31889, n31890, n31891 );
nor U131341 ( n31890, n31892, n31893 );
nor U131342 ( n31893, n31868, n31861 );
nand U131343 ( n45669, P2_P1_PHYADDRPOINTER_REG_26_, n45676 );
nand U131344 ( n45676, n45677, n45678 );
nor U131345 ( n45677, n45679, n45680 );
nor U131346 ( n45680, n45656, n45559 );
nand U131347 ( n43271, n43279, n43280 );
nand U131348 ( n43280, n43281, n76863 );
nand U131349 ( n43279, n43282, n76677 );
nor U131350 ( n43281, P2_P1_EBX_REG_3_, n8119 );
nand U131351 ( n32069, P1_P3_PHYADDRPOINTER_REG_23_, n32076 );
nand U131352 ( n32076, n32077, n32078 );
nor U131353 ( n32077, n32079, n32080 );
nor U131354 ( n32080, n32056, n31861 );
nand U131355 ( n43295, n43304, n43305 );
nand U131356 ( n43305, n43292, P2_P1_REIP_REG_1_ );
nand U131357 ( n43304, n43306, n76677 );
nor U131358 ( n43306, n7940, n43307 );
nand U131359 ( n66505, P2_P3_PHYADDRPOINTER_REG_29_, n66512 );
nand U131360 ( n66512, n66513, n66514 );
nor U131361 ( n66513, n66515, n66516 );
nor U131362 ( n66516, n66491, n66484 );
nand U131363 ( n24670, P1_P2_PHYADDRPOINTER_REG_29_, n24677 );
nand U131364 ( n24677, n24678, n24679 );
nor U131365 ( n24678, n24680, n24681 );
nor U131366 ( n24681, n24654, n24647 );
nand U131367 ( n57804, P2_P2_PHYADDRPOINTER_REG_29_, n57811 );
nand U131368 ( n57811, n57812, n57813 );
nor U131369 ( n57812, n57814, n57815 );
nor U131370 ( n57815, n57790, n57783 );
nand U131371 ( n66672, P2_P3_PHYADDRPOINTER_REG_23_, n66679 );
nand U131372 ( n66679, n66680, n66681 );
nor U131373 ( n66680, n66682, n66683 );
nor U131374 ( n66683, n66659, n66484 );
nand U131375 ( n24837, P1_P2_PHYADDRPOINTER_REG_23_, n24844 );
nand U131376 ( n24844, n24845, n24846 );
nor U131377 ( n24845, n24847, n24848 );
nor U131378 ( n24848, n24824, n24647 );
nand U131379 ( n57971, P2_P2_PHYADDRPOINTER_REG_23_, n57978 );
nand U131380 ( n57978, n57979, n57980 );
nor U131381 ( n57979, n57981, n57982 );
nor U131382 ( n57982, n57958, n57783 );
nand U131383 ( n32189, n32190, n32191 );
nand U131384 ( n32190, n3059, n29615 );
nand U131385 ( n32191, P1_P3_PHYADDRPOINTER_REG_18_, n32172 );
nand U131386 ( n32265, n32266, n32267 );
nand U131387 ( n32266, n3059, n29658 );
nand U131388 ( n32267, P1_P3_PHYADDRPOINTER_REG_15_, n32255 );
nand U131389 ( n45580, P2_P1_PHYADDRPOINTER_REG_29_, n45587 );
nand U131390 ( n45587, n45588, n45589 );
nor U131391 ( n45588, n45590, n45591 );
nor U131392 ( n45591, n45566, n45559 );
nand U131393 ( n66835, n66836, n66837 );
nand U131394 ( n66836, n5660, n63514 );
nand U131395 ( n66837, P2_P3_PHYADDRPOINTER_REG_18_, n66818 );
nand U131396 ( n24959, n24960, n24961 );
nand U131397 ( n24960, n3903, n22294 );
nand U131398 ( n24961, P1_P2_PHYADDRPOINTER_REG_18_, n24942 );
nand U131399 ( n58094, n58095, n58096 );
nand U131400 ( n58095, n6535, n55406 );
nand U131401 ( n58096, P2_P2_PHYADDRPOINTER_REG_18_, n58077 );
nand U131402 ( n32045, n32046, n32047 );
nand U131403 ( n32046, n3059, n29455 );
nand U131404 ( n32047, P1_P3_PHYADDRPOINTER_REG_24_, n32028 );
nand U131405 ( n42929, n42930, n42931 );
nand U131406 ( n42931, n42932, n76862 );
nand U131407 ( n42930, n42933, n76676 );
nor U131408 ( n42932, P2_P1_EBX_REG_15_, n8112 );
nand U131409 ( n66904, n66905, n66906 );
nand U131410 ( n66905, n5660, n63557 );
nand U131411 ( n66906, P2_P3_PHYADDRPOINTER_REG_15_, n66894 );
nand U131412 ( n25028, n25029, n25030 );
nand U131413 ( n25029, n3903, n22337 );
nand U131414 ( n25030, P1_P2_PHYADDRPOINTER_REG_15_, n25018 );
nand U131415 ( n58163, n58164, n58165 );
nand U131416 ( n58164, n6535, n55449 );
nand U131417 ( n58165, P2_P2_PHYADDRPOINTER_REG_15_, n58153 );
nand U131418 ( n43046, n43047, n43048 );
nand U131419 ( n43048, n43049, n76863 );
nand U131420 ( n43047, n43050, n76676 );
nor U131421 ( n43049, P2_P1_EBX_REG_11_, n8114 );
nand U131422 ( n42994, n42995, n42996 );
nand U131423 ( n42996, n42997, n76862 );
nand U131424 ( n42995, n42998, n76676 );
nor U131425 ( n42997, P2_P1_EBX_REG_13_, n8113 );
nand U131426 ( n42823, n42824, n42825 );
nand U131427 ( n42825, n42826, n76862 );
nand U131428 ( n42824, n42827, n76676 );
nor U131429 ( n42826, P2_P1_EBX_REG_19_, n8109 );
nand U131430 ( n45953, n45954, n45955 );
nand U131431 ( n45954, n7434, n42905 );
nand U131432 ( n45955, P2_P1_PHYADDRPOINTER_REG_15_, n45943 );
nand U131433 ( n66648, n66649, n66650 );
nand U131434 ( n66649, n5660, n63218 );
nand U131435 ( n66650, P2_P3_PHYADDRPOINTER_REG_24_, n66631 );
nand U131436 ( n24813, n24814, n24815 );
nand U131437 ( n24814, n3903, n22136 );
nand U131438 ( n24815, P1_P2_PHYADDRPOINTER_REG_24_, n24796 );
nand U131439 ( n57947, n57948, n57949 );
nand U131440 ( n57948, n6535, n55246 );
nand U131441 ( n57949, P2_P2_PHYADDRPOINTER_REG_24_, n57930 );
nand U131442 ( n45644, n45645, n45646 );
nand U131443 ( n45645, n7434, n42582 );
nand U131444 ( n45646, P2_P1_PHYADDRPOINTER_REG_27_, n45639 );
nand U131445 ( n45884, n45885, n45886 );
nand U131446 ( n45885, n7434, n42862 );
nand U131447 ( n45886, P2_P1_PHYADDRPOINTER_REG_18_, n45867 );
nand U131448 ( n42717, n42725, n42726 );
nand U131449 ( n42726, n42727, n76862 );
nand U131450 ( n42725, n42728, n76675 );
nor U131451 ( n42727, P2_P1_EBX_REG_23_, n8107 );
nand U131452 ( n45722, n45723, n45724 );
nand U131453 ( n45723, n7434, n7957 );
nand U131454 ( n45724, P2_P1_PHYADDRPOINTER_REG_24_, n45706 );
nand U131455 ( n42561, n42573, n42574 );
nand U131456 ( n42574, n42575, n42576 );
nand U131457 ( n42573, n42578, n76675 );
nor U131458 ( n42576, P2_P1_REIP_REG_28_, n73308 );
nand U131459 ( n42743, n42755, n42756 );
nand U131460 ( n42756, n42757, n42758 );
nand U131461 ( n42755, n42760, n76675 );
nor U131462 ( n42758, P2_P1_REIP_REG_22_, n74951 );
nand U131463 ( n31965, n31966, n31967 );
nand U131464 ( n31966, n3059, n29360 );
nand U131465 ( n31967, P1_P3_PHYADDRPOINTER_REG_27_, n31960 );
nand U131466 ( n24733, n24734, n24735 );
nand U131467 ( n24734, n3903, n22041 );
nand U131468 ( n24735, P1_P2_PHYADDRPOINTER_REG_27_, n24728 );
nand U131469 ( n66568, n66569, n66570 );
nand U131470 ( n66569, n5660, n63123 );
nand U131471 ( n66570, P2_P3_PHYADDRPOINTER_REG_27_, n66563 );
nand U131472 ( n57867, n57868, n57869 );
nand U131473 ( n57868, n6535, n55151 );
nand U131474 ( n57869, P2_P2_PHYADDRPOINTER_REG_27_, n57862 );
nand U131475 ( n38120, n38748, n2082 );
nor U131476 ( n38748, n2194, n38749 );
nor U131477 ( n38749, n76459, n38750 );
nor U131478 ( n38750, P4_B_REG, n37080 );
nand U131479 ( n45827, n45828, n45829 );
nand U131480 ( n45828, n7434, n42764 );
nand U131481 ( n45829, P2_P1_PHYADDRPOINTER_REG_21_, n45802 );
xor U131482 ( n32261, P1_P3_INSTADDRPOINTER_REG_16_, n33185 );
nand U131483 ( n32132, n32133, n32134 );
nand U131484 ( n32133, n3059, n29513 );
nand U131485 ( n32134, P1_P3_PHYADDRPOINTER_REG_21_, n32107 );
xor U131486 ( n12264, P1_P1_INSTADDRPOINTER_REG_16_, n13445 );
nand U131487 ( n32330, n32331, n32332 );
nand U131488 ( n32332, n32317, n74615 );
nand U131489 ( n32331, P1_P3_PHYADDRPOINTER_REG_12_, n32320 );
nand U131490 ( n66778, n66779, n66780 );
nand U131491 ( n66779, n5660, n63342 );
nand U131492 ( n66780, P2_P3_PHYADDRPOINTER_REG_21_, n66710 );
nand U131493 ( n24900, n24901, n24902 );
nand U131494 ( n24901, n3903, n22194 );
nand U131495 ( n24902, P1_P2_PHYADDRPOINTER_REG_21_, n24875 );
nand U131496 ( n58037, n58038, n58039 );
nand U131497 ( n58038, n6535, n55308 );
nand U131498 ( n58039, P2_P2_PHYADDRPOINTER_REG_21_, n58012 );
xor U131499 ( n45949, P2_P1_INSTADDRPOINTER_REG_16_, n46894 );
nand U131500 ( n66969, n66970, n66971 );
nand U131501 ( n66971, n66956, n74616 );
nand U131502 ( n66970, P2_P3_PHYADDRPOINTER_REG_12_, n66959 );
nand U131503 ( n25093, n25094, n25095 );
nand U131504 ( n25095, n25080, n74617 );
nand U131505 ( n25094, P1_P2_PHYADDRPOINTER_REG_12_, n25083 );
nand U131506 ( n58231, n58232, n58233 );
nand U131507 ( n58233, n58215, n74618 );
nand U131508 ( n58232, P2_P2_PHYADDRPOINTER_REG_12_, n58218 );
nand U131509 ( n46029, n46030, n46031 );
nand U131510 ( n46031, n46016, n74607 );
nand U131511 ( n46030, P2_P1_PHYADDRPOINTER_REG_12_, n46019 );
xor U131512 ( n66900, P2_P3_INSTADDRPOINTER_REG_16_, n67941 );
xor U131513 ( n25024, P1_P2_INSTADDRPOINTER_REG_16_, n25938 );
xor U131514 ( n58159, P2_P2_INSTADDRPOINTER_REG_16_, n59076 );
nand U131515 ( n9380, P1_P1_INSTQUEUERD_ADDR_REG_0_, n73060 );
nor U131516 ( n10267, n9380, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nor U131517 ( n44161, n73497, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131518 ( n32030, n32031, P1_P3_PHYADDRPOINTER_REG_24_ );
and U131519 ( n32031, n74804, n32032 );
nand U131520 ( n66633, n66634, P2_P3_PHYADDRPOINTER_REG_24_ );
and U131521 ( n66634, n74805, n66635 );
nand U131522 ( n24798, n24799, P1_P2_PHYADDRPOINTER_REG_24_ );
and U131523 ( n24799, n74806, n24800 );
nand U131524 ( n57932, n57933, P2_P2_PHYADDRPOINTER_REG_24_ );
and U131525 ( n57933, n74807, n57934 );
nand U131526 ( n45708, n45709, P2_P1_PHYADDRPOINTER_REG_24_ );
and U131527 ( n45709, n75236, n45710 );
nand U131528 ( n32616, P1_P3_INSTADDRPOINTER_REG_31_, n76472 );
nand U131529 ( n32234, n32235, n32236 );
nand U131530 ( n32235, n29616, n32146 );
nand U131531 ( n32236, P1_P3_PHYADDRPOINTER_REG_17_, n32237 );
nand U131532 ( n32237, n32238, n32239 );
nand U131533 ( n21368, n10267, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U131534 ( n32142, n32148, n32149 );
nand U131535 ( n32149, n32150, n32151 );
nand U131536 ( n32148, P1_P3_PHYADDRPOINTER_REG_20_, n32153 );
nor U131537 ( n32151, P1_P3_PHYADDRPOINTER_REG_20_, n32138 );
nand U131538 ( n66788, n66794, n66795 );
nand U131539 ( n66795, n66796, n66797 );
nand U131540 ( n66794, P2_P3_PHYADDRPOINTER_REG_20_, n66799 );
nor U131541 ( n66797, P2_P3_PHYADDRPOINTER_REG_20_, n66784 );
nand U131542 ( n24910, n24916, n24917 );
nand U131543 ( n24917, n24918, n24919 );
nand U131544 ( n24916, P1_P2_PHYADDRPOINTER_REG_20_, n24921 );
nor U131545 ( n24919, P1_P2_PHYADDRPOINTER_REG_20_, n24906 );
nand U131546 ( n58047, n58053, n58054 );
nand U131547 ( n58054, n58055, n58056 );
nand U131548 ( n58053, P2_P2_PHYADDRPOINTER_REG_20_, n58058 );
nor U131549 ( n58056, P2_P2_PHYADDRPOINTER_REG_20_, n58043 );
nand U131550 ( n45906, n45907, n45908 );
nand U131551 ( n45908, n45909, n76671 );
nand U131552 ( n45907, P2_P1_PHYADDRPOINTER_REG_17_, n45912 );
and U131553 ( n45909, n45910, n45911 );
nand U131554 ( n66857, n66858, n66859 );
nand U131555 ( n66859, n66860, n76719 );
nand U131556 ( n66858, P2_P3_PHYADDRPOINTER_REG_17_, n66863 );
and U131557 ( n66860, n66861, n66862 );
nand U131558 ( n45837, n45843, n45844 );
nand U131559 ( n45844, n45845, n45846 );
nand U131560 ( n45843, P2_P1_PHYADDRPOINTER_REG_20_, n45848 );
nor U131561 ( n45846, P2_P1_PHYADDRPOINTER_REG_20_, n45833 );
nand U131562 ( n17421, n8212, P4_DATAO_REG_3_ );
nand U131563 ( n24981, n24982, n24983 );
nand U131564 ( n24983, n24984, n76767 );
nand U131565 ( n24982, P1_P2_PHYADDRPOINTER_REG_17_, n24987 );
and U131566 ( n24984, n24985, n24986 );
nand U131567 ( n58116, n58117, n58118 );
nand U131568 ( n58118, n58119, n76700 );
nand U131569 ( n58117, P2_P2_PHYADDRPOINTER_REG_17_, n58122 );
and U131570 ( n58119, n58120, n58121 );
nand U131571 ( n32286, n32291, n32292 );
nand U131572 ( n32292, n32293, n32294 );
nand U131573 ( n32291, P1_P3_PHYADDRPOINTER_REG_14_, n32296 );
nor U131574 ( n32294, P1_P3_PHYADDRPOINTER_REG_14_, n32277 );
nand U131575 ( n32557, n32558, n32559 );
nand U131576 ( n32559, P1_P3_PHYADDRPOINTER_REG_1_, n32560 );
nand U131577 ( n32558, n32561, n3060 );
nand U131578 ( n32560, n31969, n31869 );
and U131579 ( n32572, n32574, P1_P3_STATE2_REG_0_ );
nor U131580 ( n32574, n3232, n3063 );
nand U131581 ( n66925, n66930, n66931 );
nand U131582 ( n66931, n66932, n66933 );
nand U131583 ( n66930, P2_P3_PHYADDRPOINTER_REG_14_, n66935 );
nor U131584 ( n66933, P2_P3_PHYADDRPOINTER_REG_14_, n66916 );
nand U131585 ( n45974, n45979, n45980 );
nand U131586 ( n45980, n45981, n45982 );
nand U131587 ( n45979, P2_P1_PHYADDRPOINTER_REG_14_, n45984 );
nor U131588 ( n45982, P2_P1_PHYADDRPOINTER_REG_14_, n45965 );
nand U131589 ( n25049, n25054, n25055 );
nand U131590 ( n25055, n25056, n25057 );
nand U131591 ( n25054, P1_P2_PHYADDRPOINTER_REG_14_, n25059 );
nor U131592 ( n25057, P1_P2_PHYADDRPOINTER_REG_14_, n25040 );
nand U131593 ( n58184, n58189, n58190 );
nand U131594 ( n58190, n58191, n58192 );
nand U131595 ( n58189, P2_P2_PHYADDRPOINTER_REG_14_, n58194 );
nor U131596 ( n58192, P2_P2_PHYADDRPOINTER_REG_14_, n58175 );
nand U131597 ( n25376, P1_P2_INSTADDRPOINTER_REG_31_, n76522 );
nand U131598 ( n67381, P2_P3_INSTADDRPOINTER_REG_31_, n76198 );
nand U131599 ( n58513, P2_P2_INSTADDRPOINTER_REG_31_, n76264 );
xor U131600 ( n12119, n13267, P1_P1_INSTADDRPOINTER_REG_20_ );
xor U131601 ( n32147, n33040, P1_P3_INSTADDRPOINTER_REG_20_ );
nand U131602 ( n11764, P1_P1_PHYADDRPOINTER_REG_31_, n11769 );
nand U131603 ( n11769, n4788, n11770 );
nand U131604 ( n11770, n11772, n74924 );
not U131605 ( n4788, n11773 );
nand U131606 ( n12017, P1_P1_PHYADDRPOINTER_REG_23_, n12025 );
nand U131607 ( n12025, n12027, n12028 );
nor U131608 ( n12027, n12029, n12030 );
nor U131609 ( n12030, n12000, n11800 );
xor U131610 ( n45842, n46748, P2_P1_INSTADDRPOINTER_REG_20_ );
xor U131611 ( n66793, n67795, P2_P3_INSTADDRPOINTER_REG_20_ );
xor U131612 ( n24915, n25792, P1_P2_INSTADDRPOINTER_REG_20_ );
xor U131613 ( n58052, n58930, P2_P2_INSTADDRPOINTER_REG_20_ );
nand U131614 ( n11930, P1_P1_PHYADDRPOINTER_REG_26_, n11939 );
nand U131615 ( n11939, n11940, n11942 );
nor U131616 ( n11940, n11943, n11944 );
nor U131617 ( n11944, n11909, n11800 );
xor U131618 ( n38294, n39391, P4_REG3_REG_19_ );
nand U131619 ( n32304, n33267, n33268 );
nand U131620 ( n33268, P1_P3_INSTADDRPOINTER_REG_14_, n3142 );
nor U131621 ( n33267, n33269, n33270 );
nor U131622 ( n33270, n3142, n33271 );
nand U131623 ( n12318, n13553, n13554 );
nand U131624 ( n13554, P1_P1_INSTADDRPOINTER_REG_14_, n4884 );
nor U131625 ( n13553, n13555, n13557 );
nor U131626 ( n13557, n4884, n13558 );
nand U131627 ( n45992, n46991, n46992 );
nand U131628 ( n46992, P2_P1_INSTADDRPOINTER_REG_14_, n7529 );
nor U131629 ( n46991, n46993, n46994 );
nor U131630 ( n46994, n7529, n46995 );
nand U131631 ( n12269, n12270, n12272 );
nand U131632 ( n12270, n4790, n8884 );
nand U131633 ( n12272, P1_P1_PHYADDRPOINTER_REG_15_, n12257 );
nand U131634 ( n11824, n11831, n11832 );
nand U131635 ( n11832, n11833, n75170 );
nand U131636 ( n11831, P1_P1_PHYADDRPOINTER_REG_29_, n11839 );
nand U131637 ( n11833, n11834, n11835 );
nand U131638 ( n66943, n68026, n68027 );
nand U131639 ( n68027, P2_P3_INSTADDRPOINTER_REG_14_, n5743 );
nor U131640 ( n68026, n68028, n68029 );
nor U131641 ( n68029, n5743, n68030 );
nand U131642 ( n25067, n26023, n26024 );
nand U131643 ( n26024, P1_P2_INSTADDRPOINTER_REG_14_, n3985 );
nor U131644 ( n26023, n26025, n26026 );
nor U131645 ( n26026, n3985, n26027 );
nand U131646 ( n58202, n59164, n59165 );
nand U131647 ( n59165, P2_P2_INSTADDRPOINTER_REG_14_, n6618 );
nor U131648 ( n59164, n59166, n59167 );
nor U131649 ( n59167, n6618, n59168 );
nand U131650 ( n11894, n11895, n11897 );
nand U131651 ( n11895, n4790, n8515 );
nand U131652 ( n11897, P1_P1_PHYADDRPOINTER_REG_27_, n11864 );
nand U131653 ( n12172, n12173, n12174 );
nand U131654 ( n12173, n4790, n8830 );
nand U131655 ( n12174, P1_P1_PHYADDRPOINTER_REG_18_, n12150 );
nand U131656 ( n11987, n11988, n11989 );
nand U131657 ( n11988, n4790, n5302 );
nand U131658 ( n11989, P1_P1_PHYADDRPOINTER_REG_24_, n11967 );
xor U131659 ( n37910, n37911, n37912 );
xor U131660 ( n37912, n37913, P4_REG2_REG_13_ );
nand U131661 ( n49480, P3_DATAO_REG_0_, n49481 );
nand U131662 ( n49481, n49482, n49483 );
nand U131663 ( n49483, n76649, n73425 );
nand U131664 ( n12095, n12097, n12098 );
nand U131665 ( n12097, n4790, n8708 );
nand U131666 ( n12098, P1_P1_PHYADDRPOINTER_REG_21_, n12064 );
nor U131667 ( n10297, n73525, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131668 ( n12350, n12352, n12353 );
nand U131669 ( n12353, n12334, n74644 );
nand U131670 ( n12352, P1_P1_PHYADDRPOINTER_REG_12_, n12338 );
xor U131671 ( n38227, n39150, P4_REG3_REG_23_ );
nand U131672 ( n39150, P4_REG3_REG_22_, n39215 );
nand U131673 ( n67322, n67323, n67324 );
nand U131674 ( n67324, P2_P3_PHYADDRPOINTER_REG_1_, n67325 );
nand U131675 ( n67323, n67326, n5662 );
nand U131676 ( n67325, n66572, n66492 );
nand U131677 ( n25315, n25316, n25317 );
nand U131678 ( n25317, P1_P2_PHYADDRPOINTER_REG_1_, n25318 );
nand U131679 ( n25316, n25319, n3904 );
nand U131680 ( n25318, n24737, n24655 );
nand U131681 ( n58454, n58455, n58456 );
nand U131682 ( n58456, P2_P2_PHYADDRPOINTER_REG_1_, n58457 );
nand U131683 ( n58455, n58458, n6537 );
nand U131684 ( n58457, n57871, n57791 );
and U131685 ( n25330, n25332, P1_P2_STATE2_REG_0_ );
nor U131686 ( n25332, n4059, n3907 );
and U131687 ( n67337, n67339, P2_P3_STATE2_REG_0_ );
nor U131688 ( n67339, n5830, n5664 );
and U131689 ( n58469, n58471, P2_P2_STATE2_REG_0_ );
nor U131690 ( n58471, n6692, n6539 );
nand U131691 ( n11960, n11962, P1_P1_PHYADDRPOINTER_REG_24_ );
and U131692 ( n11962, n75235, n11963 );
nand U131693 ( n12230, n12232, n12233 );
nand U131694 ( n12232, n8832, n12118 );
nand U131695 ( n12233, P1_P1_PHYADDRPOINTER_REG_17_, n12234 );
nand U131696 ( n12234, n12235, n12237 );
nand U131697 ( n12113, n12120, n12122 );
nand U131698 ( n12122, n12123, n12124 );
nand U131699 ( n12120, P1_P1_PHYADDRPOINTER_REG_20_, n12127 );
nor U131700 ( n12124, P1_P1_PHYADDRPOINTER_REG_20_, n12103 );
nand U131701 ( n46261, n46262, n46263 );
nand U131702 ( n46263, P2_P1_PHYADDRPOINTER_REG_1_, n46264 );
nand U131703 ( n46262, n46265, n7435 );
nand U131704 ( n46264, n45648, n45567 );
and U131705 ( n46276, n46278, P2_P1_STATE2_REG_0_ );
nor U131706 ( n46278, n7618, n7438 );
nand U131707 ( n12295, n12302, n12303 );
nand U131708 ( n12303, n12304, n12305 );
nand U131709 ( n12302, P1_P1_PHYADDRPOINTER_REG_14_, n12308 );
nor U131710 ( n12305, P1_P1_PHYADDRPOINTER_REG_14_, n12284 );
xnor U131711 ( n38147, P4_REG3_REG_28_, n38844 );
nand U131712 ( n39036, P4_REG3_REG_24_, n39091 );
nand U131713 ( n38910, P4_REG3_REG_26_, n38969 );
xnor U131714 ( n46937, P3_REG3_REG_24_, n62429 );
nand U131715 ( n32524, n32529, n32530 );
nand U131716 ( n32530, n32531, n76778 );
nand U131717 ( n32529, P1_P3_PHYADDRPOINTER_REG_3_, n32514 );
nor U131718 ( n32531, P1_P3_PHYADDRPOINTER_REG_3_, n74699 );
nand U131719 ( n46228, n46233, n46234 );
nand U131720 ( n46234, n46235, n76664 );
nand U131721 ( n46233, P2_P1_PHYADDRPOINTER_REG_3_, n46206 );
nor U131722 ( n46235, P2_P1_PHYADDRPOINTER_REG_3_, n74717 );
nand U131723 ( n67180, n67185, n67186 );
nand U131724 ( n67186, n67187, n76712 );
nand U131725 ( n67185, P2_P3_PHYADDRPOINTER_REG_3_, n67170 );
nor U131726 ( n67187, P2_P3_PHYADDRPOINTER_REG_3_, n74700 );
nand U131727 ( n25282, n25287, n25288 );
nand U131728 ( n25288, n25289, n76760 );
nand U131729 ( n25287, P1_P2_PHYADDRPOINTER_REG_3_, n25272 );
nor U131730 ( n25289, P1_P2_PHYADDRPOINTER_REG_3_, n74701 );
nand U131731 ( n58418, n58423, n58424 );
nand U131732 ( n58424, n58425, n76693 );
nand U131733 ( n58423, P2_P2_PHYADDRPOINTER_REG_3_, n58408 );
nor U131734 ( n58425, P2_P2_PHYADDRPOINTER_REG_3_, n74702 );
nand U131735 ( n12979, n76603, P1_P1_INSTADDRPOINTER_REG_25_ );
xor U131736 ( n12462, P1_P1_INSTADDRPOINTER_REG_9_, n13808 );
nor U131737 ( n13808, n13809, n13810 );
nor U131738 ( n13809, P1_P1_INSTADDRPOINTER_REG_8_, n13763 );
nand U131739 ( n13810, n13812, n13813 );
nand U131740 ( n8841, n13790, n13792 );
nand U131741 ( n13792, n76887, P1_P1_INSTADDRPOINTER_REG_9_ );
nor U131742 ( n13790, n13793, n13794 );
nor U131743 ( n13794, n73222, n76598 );
nor U131744 ( n57440, P2_P2_EAX_REG_0_, n76281 );
nor U131745 ( n24317, P1_P2_EAX_REG_0_, n76539 );
nor U131746 ( n31613, P1_P3_EAX_REG_0_, n76482 );
nor U131747 ( n65899, P2_P3_EAX_REG_0_, n76215 );
nand U131748 ( n32465, n32471, n32472 );
nand U131749 ( n32472, n32473, n76778 );
nand U131750 ( n32471, P1_P3_PHYADDRPOINTER_REG_6_, n32460 );
nor U131751 ( n32473, P1_P3_PHYADDRPOINTER_REG_6_, n32409 );
nand U131752 ( n67121, n67127, n67128 );
nand U131753 ( n67128, n67129, n76712 );
nand U131754 ( n67127, P2_P3_PHYADDRPOINTER_REG_6_, n67116 );
nor U131755 ( n67129, P2_P3_PHYADDRPOINTER_REG_6_, n67072 );
nand U131756 ( n46157, n46163, n46164 );
nand U131757 ( n46164, n46165, n76664 );
nand U131758 ( n46163, P2_P1_PHYADDRPOINTER_REG_6_, n46152 );
nor U131759 ( n46165, P2_P1_PHYADDRPOINTER_REG_6_, n46108 );
nand U131760 ( n25223, n25229, n25230 );
nand U131761 ( n25230, n25231, n76760 );
nand U131762 ( n25229, P1_P2_PHYADDRPOINTER_REG_6_, n25218 );
nor U131763 ( n25231, P1_P2_PHYADDRPOINTER_REG_6_, n25174 );
nand U131764 ( n58359, n58365, n58366 );
nand U131765 ( n58366, n58367, n76693 );
nand U131766 ( n58365, P2_P2_PHYADDRPOINTER_REG_6_, n58354 );
nor U131767 ( n58367, P2_P2_PHYADDRPOINTER_REG_6_, n58310 );
nand U131768 ( n32397, n32403, n32404 );
nand U131769 ( n32404, n32405, n76778 );
nand U131770 ( n32403, P1_P3_PHYADDRPOINTER_REG_9_, n32392 );
nor U131771 ( n32405, P1_P3_PHYADDRPOINTER_REG_9_, n32339 );
nand U131772 ( n46096, n46102, n46103 );
nand U131773 ( n46103, n46104, n76664 );
nand U131774 ( n46102, P2_P1_PHYADDRPOINTER_REG_9_, n46091 );
nor U131775 ( n46104, P2_P1_PHYADDRPOINTER_REG_9_, n46038 );
nand U131776 ( n67060, n67066, n67067 );
nand U131777 ( n67067, n67068, n76712 );
nand U131778 ( n67066, P2_P3_PHYADDRPOINTER_REG_9_, n67055 );
nor U131779 ( n67068, P2_P3_PHYADDRPOINTER_REG_9_, n66978 );
nand U131780 ( n25162, n25168, n25169 );
nand U131781 ( n25169, n25170, n76760 );
nand U131782 ( n25168, P1_P2_PHYADDRPOINTER_REG_9_, n25155 );
nor U131783 ( n25170, P1_P2_PHYADDRPOINTER_REG_9_, n25102 );
nand U131784 ( n58298, n58304, n58305 );
nand U131785 ( n58305, n58306, n76693 );
nand U131786 ( n58304, P2_P2_PHYADDRPOINTER_REG_9_, n58293 );
nor U131787 ( n58306, P2_P2_PHYADDRPOINTER_REG_9_, n58240 );
nand U131788 ( n31853, n31854, n31855 );
nand U131789 ( n31854, n3059, n29275 );
nand U131790 ( n31855, P1_P3_PHYADDRPOINTER_REG_30_, n31842 );
nand U131791 ( n24639, n24640, n24641 );
nand U131792 ( n24640, n3903, n21958 );
nand U131793 ( n24641, P1_P2_PHYADDRPOINTER_REG_30_, n24628 );
nand U131794 ( n57775, n57776, n57777 );
nand U131795 ( n57776, n6535, n55070 );
nand U131796 ( n57777, P2_P2_PHYADDRPOINTER_REG_30_, n57760 );
nand U131797 ( n66476, n66477, n66478 );
nand U131798 ( n66477, n5660, n63042 );
nand U131799 ( n66478, P2_P3_PHYADDRPOINTER_REG_30_, n66465 );
nand U131800 ( n45551, n45552, n45553 );
nand U131801 ( n45552, n7434, n42490 );
nand U131802 ( n45553, P2_P1_PHYADDRPOINTER_REG_30_, n45541 );
xnor U131803 ( n45750, P3_REG3_REG_28_, n61596 );
nand U131804 ( n62363, P3_REG3_REG_24_, n62429 );
nand U131805 ( n62246, P3_REG3_REG_26_, n62302 );
nor U131806 ( n57004, n76281, n57008 );
or U131807 ( n57008, n56898, P2_P2_EAX_REG_15_ );
nor U131808 ( n23880, n76539, n23884 );
or U131809 ( n23884, n23773, P1_P2_EAX_REG_15_ );
nor U131810 ( n31173, n76482, n31176 );
or U131811 ( n31176, n31072, P1_P3_EAX_REG_15_ );
nor U131812 ( n65427, n76215, n65430 );
or U131813 ( n65430, n65274, P2_P3_EAX_REG_15_ );
nor U131814 ( n57428, n76281, n57431 );
nand U131815 ( n57431, P2_P2_EAX_REG_0_, n73128 );
nor U131816 ( n24305, n76539, n24308 );
nand U131817 ( n24308, P1_P2_EAX_REG_0_, n73129 );
nor U131818 ( n31601, n76482, n31604 );
nand U131819 ( n31604, P1_P3_EAX_REG_0_, n72957 );
nor U131820 ( n65887, n76215, n65890 );
nand U131821 ( n65890, P2_P3_EAX_REG_0_, n73127 );
nand U131822 ( n12632, n12633, n12634 );
nand U131823 ( n12634, P1_P1_PHYADDRPOINTER_REG_1_, n12635 );
nand U131824 ( n12633, n12637, n4792 );
nand U131825 ( n12635, n11899, n11810 );
and U131826 ( n12659, n12662, P1_P1_STATE2_REG_0_ );
nor U131827 ( n12662, n4964, n4794 );
nand U131828 ( n12590, n12597, n12598 );
nand U131829 ( n12598, n12599, n76731 );
nand U131830 ( n12597, P1_P1_PHYADDRPOINTER_REG_3_, n12578 );
nor U131831 ( n12599, P1_P1_PHYADDRPOINTER_REG_3_, n74718 );
xnor U131832 ( n38182, P4_REG3_REG_26_, n38969 );
nand U131833 ( n12517, n12524, n12525 );
nand U131834 ( n12525, n12527, n76731 );
nand U131835 ( n12524, P1_P1_PHYADDRPOINTER_REG_6_, n12510 );
nor U131836 ( n12527, P1_P1_PHYADDRPOINTER_REG_6_, n12455 );
nand U131837 ( n54228, P2_P1_INSTQUEUERD_ADDR_REG_3_, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131838 ( n12440, n12448, n12449 );
nand U131839 ( n12449, n12450, n76731 );
nand U131840 ( n12448, P1_P1_PHYADDRPOINTER_REG_9_, n12434 );
nor U131841 ( n12450, P1_P1_PHYADDRPOINTER_REG_9_, n12362 );
nand U131842 ( n49725, n8240, P3_DATAO_REG_6_ );
nand U131843 ( n11790, n11792, n11793 );
nand U131844 ( n11792, n4790, n5305 );
nand U131845 ( n11793, P1_P1_PHYADDRPOINTER_REG_30_, n11773 );
nand U131846 ( n32345, n74458, n33384 );
nand U131847 ( n33384, n3138, P1_P3_INSTADDRPOINTER_REG_11_ );
nand U131848 ( n46044, n74427, n47105 );
nand U131849 ( n47105, n7524, P2_P1_INSTADDRPOINTER_REG_11_ );
nand U131850 ( n46529, n76006, P2_P1_INSTADDRPOINTER_REG_25_ );
nand U131851 ( n66984, n74438, n68136 );
nand U131852 ( n68136, n5739, P2_P3_INSTADDRPOINTER_REG_11_ );
nand U131853 ( n12369, n74476, n13697 );
nand U131854 ( n13697, n4879, P1_P1_INSTADDRPOINTER_REG_11_ );
nand U131855 ( n25108, n74439, n26133 );
nand U131856 ( n26133, n3982, P1_P2_INSTADDRPOINTER_REG_11_ );
nand U131857 ( n58246, n74440, n59274 );
nand U131858 ( n59274, n6614, P2_P2_INSTADDRPOINTER_REG_11_ );
nand U131859 ( n67590, n75990, P2_P3_INSTADDRPOINTER_REG_25_ );
nand U131860 ( n25585, n76027, P1_P2_INSTADDRPOINTER_REG_25_ );
nand U131861 ( n58722, n75998, P2_P2_INSTADDRPOINTER_REG_25_ );
nand U131862 ( n9186, n11597, n11598 );
nand U131863 ( n11598, P1_P1_LWORD_REG_1_, n76618 );
nor U131864 ( n11597, n11599, n11513 );
nor U131865 ( n11599, n74608, n76616 );
nand U131866 ( n9261, n11509, n11510 );
nand U131867 ( n11510, P1_P1_UWORD_REG_1_, n11504 );
nor U131868 ( n11509, n11512, n11513 );
nor U131869 ( n11512, n74909, n76617 );
nand U131870 ( n32825, n76022, P1_P3_INSTADDRPOINTER_REG_25_ );
nand U131871 ( n13680, n76602, P1_P1_INSTADDRPOINTER_REG_12_ );
nand U131872 ( n32216, n74879, n33189 );
nand U131873 ( n33189, n33188, P1_P3_INSTADDRPOINTER_REG_16_ );
nand U131874 ( n21230, P1_P1_INSTQUEUERD_ADDR_REG_3_, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U131875 ( n12205, n74847, n13450 );
nand U131876 ( n13450, n13449, P1_P1_INSTADDRPOINTER_REG_16_ );
nand U131877 ( n45922, n74841, n46898 );
nand U131878 ( n46898, n46897, P2_P1_INSTADDRPOINTER_REG_16_ );
nand U131879 ( n66873, n74872, n67945 );
nand U131880 ( n67945, n67944, P2_P3_INSTADDRPOINTER_REG_16_ );
nand U131881 ( n24997, n74873, n25942 );
nand U131882 ( n25942, n25941, P1_P2_INSTADDRPOINTER_REG_16_ );
nand U131883 ( n58132, n74874, n59080 );
nand U131884 ( n59080, n59079, P2_P2_INSTADDRPOINTER_REG_16_ );
xnor U131885 ( n38211, P4_REG3_REG_24_, n39091 );
nor U131886 ( n71668, n74437, n71104 );
nand U131887 ( n8846, n13740, n13742 );
nand U131888 ( n13742, n76887, P1_P1_INSTADDRPOINTER_REG_10_ );
nor U131889 ( n13740, n13743, n13744 );
nor U131890 ( n13744, n74770, n76598 );
xor U131891 ( n38195, n39036, P4_REG3_REG_25_ );
nand U131892 ( n38128, n38844, P4_REG3_REG_28_ );
and U131893 ( n17672, n17054, P4_DATAO_REG_1_ );
xor U131894 ( n46549, n62363, P3_REG3_REG_25_ );
nand U131895 ( n50034, DIN_28_, n76929 );
xor U131896 ( n38163, n38910, P4_REG3_REG_27_ );
nand U131897 ( n68123, n75990, P2_P3_INSTADDRPOINTER_REG_12_ );
nand U131898 ( n47092, n76006, P2_P1_INSTADDRPOINTER_REG_12_ );
nand U131899 ( n26120, n76027, P1_P2_INSTADDRPOINTER_REG_12_ );
nand U131900 ( n59261, n75998, P2_P2_INSTADDRPOINTER_REG_12_ );
xnor U131901 ( n46220, P3_REG3_REG_26_, n62302 );
nand U131902 ( n17077, DIN_26_, n76928 );
xor U131903 ( n12345, P1_P1_INSTADDRPOINTER_REG_13_, n13512 );
nand U131904 ( n42231, n45265, n42216 );
nand U131905 ( n45265, n45266, P3_REG1_REG_0_ );
nor U131906 ( n45266, n45267, n73024 );
nor U131907 ( n45267, P3_REG1_REG_1_, n45201 );
nand U131908 ( n44859, n45215, n45216 );
nand U131909 ( n45215, n44393, n44395 );
nand U131910 ( n45216, P3_REG1_REG_14_, n45217 );
or U131911 ( n45217, n44393, n44395 );
nand U131912 ( n45017, n45212, n45213 );
nand U131913 ( n45212, n44859, n44857 );
nand U131914 ( n45213, P3_REG1_REG_15_, n45214 );
or U131915 ( n45214, n44859, n44857 );
nor U131916 ( n45247, n45250, n42686 );
nor U131917 ( n45250, P3_REG1_REG_7_, n42678 );
nor U131918 ( n45253, n45256, n45257 );
nor U131919 ( n45256, P3_REG1_REG_5_, n42344 );
nand U131920 ( n45257, n45258, n42308 );
nand U131921 ( n45258, n45259, n42353 );
nor U131922 ( n45228, n872, n45230 );
nor U131923 ( n45230, P3_REG1_REG_11_, n43559 );
nor U131924 ( n45241, n890, n45244 );
nor U131925 ( n45244, P3_REG1_REG_8_, n42957 );
xor U131926 ( n32326, P1_P3_INSTADDRPOINTER_REG_13_, n33238 );
xor U131927 ( n46025, P2_P1_INSTADDRPOINTER_REG_13_, n46958 );
xor U131928 ( n66965, P2_P3_INSTADDRPOINTER_REG_13_, n67993 );
xor U131929 ( n25089, P1_P2_INSTADDRPOINTER_REG_13_, n25990 );
xor U131930 ( n58224, P2_P2_INSTADDRPOINTER_REG_13_, n59128 );
nor U131931 ( n72889, n74446, n71104 );
nor U131932 ( n72888, n74444, n71105 );
nand U131933 ( n12317, n13562, n13563 );
nand U131934 ( n13563, P1_P1_INSTADDRPOINTER_REG_14_, n4910 );
nor U131935 ( n13562, n13555, n13564 );
nor U131936 ( n13564, n4910, n13558 );
nor U131937 ( n13550, n13559, n13560 );
nor U131938 ( n13559, P1_P1_INSTADDRPOINTER_REG_14_, n13540 );
and U131939 ( n13560, n12317, n4848 );
nand U131940 ( n32303, n33274, n33275 );
nand U131941 ( n33275, P1_P3_INSTADDRPOINTER_REG_14_, n3173 );
nor U131942 ( n33274, n33269, n33276 );
nor U131943 ( n33276, n3173, n33271 );
nor U131944 ( n33265, n33272, n33273 );
nor U131945 ( n33272, P1_P3_INSTADDRPOINTER_REG_14_, n33257 );
and U131946 ( n33273, n32303, n3103 );
nand U131947 ( n45991, n46998, n46999 );
nand U131948 ( n46999, P2_P1_INSTADDRPOINTER_REG_14_, n7559 );
nor U131949 ( n46998, n46993, n47000 );
nor U131950 ( n47000, n7559, n46995 );
nor U131951 ( n46989, n46996, n46997 );
nor U131952 ( n46996, P2_P1_INSTADDRPOINTER_REG_14_, n46981 );
and U131953 ( n46997, n45991, n7490 );
nand U131954 ( n66942, n68033, n68034 );
nand U131955 ( n68034, P2_P3_INSTADDRPOINTER_REG_14_, n5772 );
nor U131956 ( n68033, n68028, n68035 );
nor U131957 ( n68035, n5772, n68030 );
nand U131958 ( n25066, n26030, n26031 );
nand U131959 ( n26031, P1_P2_INSTADDRPOINTER_REG_14_, n4013 );
nor U131960 ( n26030, n26025, n26032 );
nor U131961 ( n26032, n4013, n26027 );
nand U131962 ( n58201, n59171, n59172 );
nand U131963 ( n59172, P2_P2_INSTADDRPOINTER_REG_14_, n6645 );
nor U131964 ( n59171, n59166, n59173 );
nor U131965 ( n59173, n6645, n59168 );
nor U131966 ( n68024, n68031, n68032 );
nor U131967 ( n68031, P2_P3_INSTADDRPOINTER_REG_14_, n68016 );
and U131968 ( n68032, n66942, n5704 );
nor U131969 ( n26021, n26028, n26029 );
nor U131970 ( n26028, P1_P2_INSTADDRPOINTER_REG_14_, n26013 );
and U131971 ( n26029, n25066, n3947 );
nor U131972 ( n59162, n59169, n59170 );
nor U131973 ( n59169, P2_P2_INSTADDRPOINTER_REG_14_, n59151 );
and U131974 ( n59170, n58201, n6579 );
nand U131975 ( n45009, n45147, n45148 );
nand U131976 ( n45147, n44855, n44857 );
nand U131977 ( n45148, P3_REG2_REG_15_, n45149 );
or U131978 ( n45149, n44855, n44857 );
nor U131979 ( n45188, n45191, n45192 );
nor U131980 ( n45191, P3_REG2_REG_5_, n42344 );
nand U131981 ( n45192, n45193, n42303 );
nand U131982 ( n45193, n45194, n42339 );
nor U131983 ( n45143, n45146, n45076 );
nor U131984 ( n45146, P3_REG2_REG_17_, n45077 );
nor U131985 ( n45181, n45185, n42677 );
nor U131986 ( n45185, P3_REG2_REG_7_, n42678 );
nor U131987 ( n45176, n892, n45178 );
nor U131988 ( n45178, P3_REG2_REG_8_, n42957 );
nor U131989 ( n45163, n875, n45165 );
nor U131990 ( n45165, P3_REG2_REG_11_, n43559 );
nand U131991 ( n44855, n45150, n45151 );
nand U131992 ( n45150, n44390, n44395 );
nand U131993 ( n45151, P3_REG2_REG_14_, n45152 );
or U131994 ( n45152, n44390, n44395 );
nand U131995 ( n32387, n73115, n33456 );
nand U131996 ( n33456, P1_P3_INSTADDRPOINTER_REG_9_, n33455 );
nand U131997 ( n12428, n74735, n13785 );
nand U131998 ( n13785, P1_P1_INSTADDRPOINTER_REG_9_, n13784 );
nand U131999 ( n46086, n74734, n47176 );
nand U132000 ( n47176, P2_P1_INSTADDRPOINTER_REG_9_, n47175 );
nand U132001 ( n67050, n74758, n68207 );
nand U132002 ( n68207, P2_P3_INSTADDRPOINTER_REG_9_, n68206 );
nand U132003 ( n25150, n74759, n26206 );
nand U132004 ( n26206, P1_P2_INSTADDRPOINTER_REG_9_, n26205 );
nand U132005 ( n58288, n74760, n59345 );
nand U132006 ( n59345, P2_P2_INSTADDRPOINTER_REG_9_, n59344 );
xor U132007 ( n12263, P1_P1_INSTADDRPOINTER_REG_16_, n13449 );
xor U132008 ( n32260, P1_P3_INSTADDRPOINTER_REG_16_, n33188 );
xor U132009 ( n45948, P2_P1_INSTADDRPOINTER_REG_16_, n46897 );
xor U132010 ( n32372, P1_P3_INSTADDRPOINTER_REG_11_, n3138 );
xor U132011 ( n66899, P2_P3_INSTADDRPOINTER_REG_16_, n67944 );
xor U132012 ( n46071, P2_P1_INSTADDRPOINTER_REG_11_, n7524 );
xor U132013 ( n25023, P1_P2_INSTADDRPOINTER_REG_16_, n25941 );
xor U132014 ( n58158, P2_P2_INSTADDRPOINTER_REG_16_, n59079 );
xor U132015 ( n67035, P2_P3_INSTADDRPOINTER_REG_11_, n5739 );
xor U132016 ( n25135, P1_P2_INSTADDRPOINTER_REG_11_, n3982 );
xor U132017 ( n58273, P2_P2_INSTADDRPOINTER_REG_11_, n6614 );
xor U132018 ( n12403, P1_P1_INSTADDRPOINTER_REG_11_, n4879 );
nor U132019 ( n72895, n74445, n71108 );
nand U132020 ( n8836, n13837, n13838 );
nand U132021 ( n13838, n76887, P1_P1_INSTADDRPOINTER_REG_8_ );
nor U132022 ( n13837, n13839, n13840 );
nor U132023 ( n13840, n75967, n76598 );
nand U132024 ( n35607, n35637, n35638 );
nor U132025 ( n35638, n35639, n35640 );
nor U132026 ( n35637, n35642, n74662 );
nor U132027 ( n35640, P1_P3_STATE2_REG_0_, n35641 );
nand U132028 ( n28430, n28458, n28459 );
nor U132029 ( n28459, n28460, n28461 );
nor U132030 ( n28458, n28463, n74663 );
nor U132031 ( n28461, P1_P2_STATE2_REG_0_, n28462 );
nand U132032 ( n70335, n70363, n70364 );
nor U132033 ( n70364, n70365, n70366 );
nor U132034 ( n70363, n70368, n74660 );
nor U132035 ( n70366, P2_P3_STATE2_REG_0_, n70367 );
nand U132036 ( n61735, n61763, n61764 );
nor U132037 ( n61764, n61765, n61766 );
nor U132038 ( n61763, n61768, n74661 );
nor U132039 ( n61766, P2_P2_STATE2_REG_0_, n61767 );
nand U132040 ( n35693, n35687, n35741 );
nand U132041 ( n35741, P1_P3_INSTQUEUERD_ADDR_REG_0_, n35685 );
nand U132042 ( n28514, n28508, n28562 );
nand U132043 ( n28562, P1_P2_INSTQUEUERD_ADDR_REG_0_, n28506 );
nand U132044 ( n70419, n70413, n70467 );
nand U132045 ( n70467, P2_P3_INSTQUEUERD_ADDR_REG_0_, n70411 );
nand U132046 ( n61819, n61813, n61867 );
nand U132047 ( n61867, P2_P2_INSTQUEUERD_ADDR_REG_0_, n61811 );
nor U132048 ( n35642, n35643, n74591 );
nor U132049 ( n35643, P1_P3_STATE2_REG_1_, n35610 );
nor U132050 ( n28463, n28464, n74592 );
nor U132051 ( n28464, P1_P2_STATE2_REG_1_, n28433 );
nor U132052 ( n70368, n70369, n74593 );
nor U132053 ( n70369, P2_P3_STATE2_REG_1_, n70338 );
nor U132054 ( n61768, n61769, n74594 );
nor U132055 ( n61769, P2_P2_STATE2_REG_1_, n61738 );
nor U132056 ( n35690, P1_P3_INSTQUEUERD_ADDR_REG_1_, n35692 );
nor U132057 ( n35692, n3097, n35693 );
nor U132058 ( n28511, P1_P2_INSTQUEUERD_ADDR_REG_1_, n28513 );
nor U132059 ( n28513, n3940, n28514 );
nor U132060 ( n70416, P2_P3_INSTQUEUERD_ADDR_REG_1_, n70418 );
nor U132061 ( n70418, n5698, n70419 );
nor U132062 ( n61816, P2_P2_INSTQUEUERD_ADDR_REG_1_, n61818 );
nor U132063 ( n61818, n6573, n61819 );
nand U132064 ( n35647, n35648, n35649 );
nand U132065 ( n35649, n29194, n35650 );
nand U132066 ( n35648, n35665, n75032 );
or U132067 ( n35650, P1_P3_MORE_REG, P1_P3_FLUSH_REG );
nand U132068 ( n28468, n28469, n28470 );
nand U132069 ( n28470, n21877, n28471 );
nand U132070 ( n28469, n28486, n75033 );
or U132071 ( n28471, P1_P2_MORE_REG, P1_P2_FLUSH_REG );
nand U132072 ( n70373, n70374, n70375 );
nand U132073 ( n70375, n62912, n70376 );
nand U132074 ( n70374, n70391, n75034 );
or U132075 ( n70376, P2_P3_MORE_REG, P2_P3_FLUSH_REG );
nand U132076 ( n61773, n61774, n61775 );
nand U132077 ( n61775, n54968, n61776 );
nand U132078 ( n61774, n61791, n75035 );
or U132079 ( n61776, P2_P2_MORE_REG, P2_P2_FLUSH_REG );
nand U132080 ( n54107, n54135, n54136 );
nor U132081 ( n54136, n54137, n54138 );
nor U132082 ( n54135, n54140, n73190 );
nor U132083 ( n54138, P2_P1_STATE2_REG_0_, n54139 );
nor U132084 ( n54140, n54141, n74648 );
nor U132085 ( n54141, P2_P1_STATE2_REG_1_, n54110 );
nand U132086 ( n54191, n54185, n54239 );
nand U132087 ( n54239, P2_P1_INSTQUEUERD_ADDR_REG_0_, n54183 );
nor U132088 ( n54188, P2_P1_INSTQUEUERD_ADDR_REG_1_, n54190 );
nor U132089 ( n54190, n7484, n54191 );
nand U132090 ( n54145, n54146, n54147 );
nand U132091 ( n54147, n42403, n54148 );
nand U132092 ( n54146, n54163, n75030 );
or U132093 ( n54148, P2_P1_MORE_REG, P2_P1_FLUSH_REG );
nand U132094 ( n67809, n75990, P2_P3_INSTADDRPOINTER_REG_20_ );
nand U132095 ( n46762, n76006, P2_P1_INSTADDRPOINTER_REG_20_ );
nand U132096 ( n25806, n76027, P1_P2_INSTADDRPOINTER_REG_20_ );
nand U132097 ( n58944, n75998, P2_P2_INSTADDRPOINTER_REG_20_ );
not U132098 ( n76924, P4_STATE_REG );
nand U132099 ( n45491, n61596, P3_REG3_REG_28_ );
nand U132100 ( n32549, n32550, n32551 );
nand U132101 ( n32550, n32553, P1_P3_REIP_REG_2_ );
nand U132102 ( n32551, n76785, n32552 );
nand U132103 ( n46253, n46254, n46255 );
nand U132104 ( n46254, n46257, P2_P1_REIP_REG_2_ );
nand U132105 ( n46255, n76671, n46256 );
nand U132106 ( n67205, n67206, n67207 );
nand U132107 ( n67206, n67209, P2_P3_REIP_REG_2_ );
nand U132108 ( n67207, n76719, n67208 );
nand U132109 ( n25307, n25308, n25309 );
nand U132110 ( n25308, n25311, P1_P2_REIP_REG_2_ );
nand U132111 ( n25309, n76767, n25310 );
nand U132112 ( n58446, n58447, n58448 );
nand U132113 ( n58447, n58450, P2_P2_REIP_REG_2_ );
nand U132114 ( n58448, n76700, n58449 );
xor U132115 ( n40715, n62246, P3_REG3_REG_27_ );
nand U132116 ( n54169, n54201, n54202 );
nand U132117 ( n54201, n494, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U132118 ( n54202, n47996, n54176 );
nand U132119 ( n35671, n35703, n35704 );
nand U132120 ( n35703, n189, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U132121 ( n35704, n34250, n35678 );
nand U132122 ( n28492, n28524, n28525 );
nand U132123 ( n28524, n152, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U132124 ( n28525, n27005, n28499 );
nand U132125 ( n70397, n70429, n70430 );
nand U132126 ( n70429, n460, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U132127 ( n70430, n69004, n70404 );
nand U132128 ( n61797, n61829, n61830 );
nand U132129 ( n61829, n424, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U132130 ( n61830, n60148, n61804 );
nand U132131 ( n61745, P2_P2_STATE2_REG_0_, n61735 );
nand U132132 ( n28440, P1_P2_STATE2_REG_0_, n28430 );
nand U132133 ( n35619, P1_P3_STATE2_REG_0_, n35607 );
nand U132134 ( n70345, P2_P3_STATE2_REG_0_, n70335 );
nand U132135 ( n54117, P2_P1_STATE2_REG_0_, n54107 );
nand U132136 ( n796, n31921, n31922 );
nor U132137 ( n31922, n31923, n31924 );
nor U132138 ( n31921, n31926, n31927 );
or U132139 ( n31924, P2_P1_BE_N_REG_0_, P2_P1_BE_N_REG_1_ );
not U132140 ( n76479, n31928 );
nand U132141 ( n31928, P2_P1_ADDRESS_REG_29_, n54064 );
nand U132142 ( n54064, n54065, n54066 );
nor U132143 ( n54065, n54080, n54081 );
nor U132144 ( n54066, n54067, n54068 );
nand U132145 ( n54068, n54069, n54070 );
nand U132146 ( n54067, n54074, n54075 );
nor U132147 ( n54069, P2_P1_ADDRESS_REG_22_, n54073 );
or U132148 ( n31926, n76476, P2_P1_ADS_N_REG );
nand U132149 ( n616, n27746, n27747 );
nand U132150 ( n27747, P2_P1_DATAO_REG_31_, n76682 );
nor U132151 ( n27746, n27748, n27749 );
nor U132152 ( n27749, n76514, n75445 );
nor U132153 ( n28155, n75587, n76512 );
nor U132154 ( n28057, n75588, n76512 );
nor U132155 ( n28252, n75589, n76512 );
nor U132156 ( n27956, n75590, n76512 );
nor U132157 ( n28933, n75591, n76512 );
nor U132158 ( n28420, n75592, n76512 );
nand U132159 ( n611, n27847, n27848 );
nand U132160 ( n27848, P2_P1_DATAO_REG_30_, n76682 );
nor U132161 ( n27847, n27849, n27850 );
nor U132162 ( n27850, n76514, n75406 );
nand U132163 ( n596, n28153, n28154 );
nand U132164 ( n28154, P2_P1_DATAO_REG_27_, n76682 );
nor U132165 ( n28153, n28155, n28156 );
nor U132166 ( n28156, n76514, n75407 );
nand U132167 ( n601, n28055, n28056 );
nand U132168 ( n28056, P2_P1_DATAO_REG_28_, n76682 );
nor U132169 ( n28055, n28057, n28058 );
nor U132170 ( n28058, n76514, n75408 );
nand U132171 ( n591, n28250, n28251 );
nand U132172 ( n28251, P2_P1_DATAO_REG_26_, n76682 );
nor U132173 ( n28250, n28252, n28253 );
nor U132174 ( n28253, n76514, n75366 );
nand U132175 ( n606, n27954, n27955 );
nand U132176 ( n27955, P2_P1_DATAO_REG_29_, n76682 );
nor U132177 ( n27954, n27956, n27957 );
nor U132178 ( n27957, n76514, n75367 );
nand U132179 ( n581, n28931, n28932 );
nand U132180 ( n28932, P2_P1_DATAO_REG_24_, n76682 );
nor U132181 ( n28931, n28933, n28934 );
nor U132182 ( n28934, n76514, n75409 );
nand U132183 ( n586, n28418, n28419 );
nand U132184 ( n28419, P2_P1_DATAO_REG_25_, n76682 );
nor U132185 ( n28418, n28420, n28421 );
nor U132186 ( n28421, n76514, n75368 );
nor U132187 ( n31577, n75504, n76510 );
nor U132188 ( n29837, n75505, n76511 );
nor U132189 ( n30395, n75506, n76510 );
nor U132190 ( n29086, n75507, n76511 );
nor U132191 ( n29042, n75508, n76511 );
nor U132192 ( n30203, n75509, n76511 );
nor U132193 ( n30302, n75510, n76510 );
nor U132194 ( n29128, n75511, n76511 );
nor U132195 ( n31649, n75512, n76510 );
nor U132196 ( n31271, n75513, n76510 );
nor U132197 ( n30106, n75514, n76511 );
nor U132198 ( n31747, n75515, n76510 );
nor U132199 ( n29306, n75516, n76511 );
nor U132200 ( n30751, n75517, n76510 );
nor U132201 ( n29180, n75518, n76511 );
nor U132202 ( n28941, n75519, n76511 );
nor U132203 ( n31628, n75520, n76510 );
nor U132204 ( n31743, n75521, n76510 );
nor U132205 ( n28998, n75522, n76511 );
nor U132206 ( n31788, n75523, n76510 );
nor U132207 ( n31693, n75524, n76510 );
nor U132208 ( n29571, n75525, n76511 );
nor U132209 ( n28937, n75526, n76511 );
nor U132210 ( n31911, n75527, n76510 );
nand U132211 ( n12622, n12623, n12624 );
nand U132212 ( n12623, n12627, P1_P1_REIP_REG_2_ );
nand U132213 ( n12624, n76738, n12625 );
nand U132214 ( n496, n31575, n31576 );
nand U132215 ( n31576, P2_P1_DATAO_REG_7_, n76683 );
nor U132216 ( n31575, n31577, n31578 );
nor U132217 ( n31578, n76516, n75448 );
nand U132218 ( n531, n29835, n29836 );
nand U132219 ( n29836, P2_P1_DATAO_REG_14_, n76682 );
nor U132220 ( n29835, n29837, n29838 );
nor U132221 ( n29838, n76515, n75429 );
nand U132222 ( n511, n30393, n30394 );
nand U132223 ( n30394, P2_P1_DATAO_REG_10_, n76683 );
nor U132224 ( n30393, n30395, n30396 );
nor U132225 ( n30396, n76515, n75430 );
nand U132226 ( n556, n29084, n29085 );
nand U132227 ( n29085, P2_P1_DATAO_REG_19_, n76682 );
nor U132228 ( n29084, n29086, n29087 );
nor U132229 ( n29087, n76515, n75369 );
nand U132230 ( n561, n29040, n29041 );
nand U132231 ( n29041, P2_P1_DATAO_REG_20_, n76682 );
nor U132232 ( n29040, n29042, n29043 );
nor U132233 ( n29043, n76514, n75370 );
nand U132234 ( n521, n30201, n30202 );
nand U132235 ( n30202, P2_P1_DATAO_REG_12_, n76683 );
nor U132236 ( n30201, n30203, n30204 );
nor U132237 ( n30204, n76515, n75431 );
nand U132238 ( n516, n30300, n30301 );
nand U132239 ( n30301, P2_P1_DATAO_REG_11_, n76683 );
nor U132240 ( n30300, n30302, n30303 );
nor U132241 ( n30303, n76515, n75432 );
nand U132242 ( n551, n29126, n29127 );
nand U132243 ( n29127, P2_P1_DATAO_REG_18_, n76682 );
nor U132244 ( n29126, n29128, n29129 );
nor U132245 ( n29129, n76515, n75371 );
nand U132246 ( n486, n31647, n31648 );
nand U132247 ( n31648, P2_P1_DATAO_REG_5_, n76683 );
nor U132248 ( n31647, n31649, n31650 );
nor U132249 ( n31650, n76516, n75449 );
nand U132250 ( n501, n31269, n31270 );
nand U132251 ( n31270, P2_P1_DATAO_REG_8_, n76683 );
nor U132252 ( n31269, n31271, n31272 );
nor U132253 ( n31272, n76515, n75433 );
nand U132254 ( n526, n30104, n30105 );
nand U132255 ( n30105, P2_P1_DATAO_REG_13_, n76682 );
nor U132256 ( n30104, n30106, n30107 );
nor U132257 ( n30107, n76515, n75434 );
nand U132258 ( n471, n31745, n31746 );
nand U132259 ( n31746, P2_P1_DATAO_REG_2_, n76683 );
nor U132260 ( n31745, n31747, n31748 );
nor U132261 ( n31748, n76516, n75450 );
nand U132262 ( n541, n29304, n29305 );
nand U132263 ( n29305, P2_P1_DATAO_REG_16_, n76682 );
nor U132264 ( n29304, n29306, n29307 );
nor U132265 ( n29307, n76515, n75372 );
nand U132266 ( n506, n30749, n30750 );
nand U132267 ( n30750, P2_P1_DATAO_REG_9_, n76683 );
nor U132268 ( n30749, n30751, n30752 );
nor U132269 ( n30752, n76515, n75435 );
nand U132270 ( n546, n29178, n29179 );
nand U132271 ( n29179, P2_P1_DATAO_REG_17_, n76682 );
nor U132272 ( n29178, n29180, n29181 );
nor U132273 ( n29181, n76515, n75373 );
nand U132274 ( n571, n28939, n28940 );
nand U132275 ( n28940, P2_P1_DATAO_REG_22_, n76682 );
nor U132276 ( n28939, n28941, n28942 );
nor U132277 ( n28942, n76514, n75374 );
nand U132278 ( n491, n31626, n31627 );
nand U132279 ( n31627, P2_P1_DATAO_REG_6_, n76683 );
nor U132280 ( n31626, n31628, n31629 );
nor U132281 ( n31629, n76516, n75451 );
nand U132282 ( n476, n31741, n31742 );
nand U132283 ( n31742, P2_P1_DATAO_REG_3_, n76683 );
nor U132284 ( n31741, n31743, n31744 );
nor U132285 ( n31744, n76516, n75452 );
nand U132286 ( n566, n28996, n28997 );
nand U132287 ( n28997, P2_P1_DATAO_REG_21_, n76682 );
nor U132288 ( n28996, n28998, n28999 );
nor U132289 ( n28999, n76514, n75375 );
nand U132290 ( n466, n31786, n31787 );
nand U132291 ( n31787, P2_P1_DATAO_REG_1_, n76683 );
nor U132292 ( n31786, n31788, n31789 );
nor U132293 ( n31789, n76516, n75453 );
nand U132294 ( n481, n31691, n31692 );
nand U132295 ( n31692, P2_P1_DATAO_REG_4_, n76683 );
nor U132296 ( n31691, n31693, n31694 );
nor U132297 ( n31694, n76516, n75454 );
nand U132298 ( n536, n29569, n29570 );
nand U132299 ( n29570, P2_P1_DATAO_REG_15_, n76682 );
nor U132300 ( n29569, n29571, n29572 );
nor U132301 ( n29572, n76515, n75436 );
nand U132302 ( n576, n28935, n28936 );
nand U132303 ( n28936, P2_P1_DATAO_REG_23_, n76682 );
nor U132304 ( n28935, n28937, n28938 );
nor U132305 ( n28938, n76514, n75376 );
nand U132306 ( n461, n31909, n31910 );
nand U132307 ( n31910, P2_P1_DATAO_REG_0_, n76683 );
nor U132308 ( n31909, n31911, n31912 );
nor U132309 ( n31912, n76516, n75455 );
nand U132310 ( n21124, n21152, n21153 );
nor U132311 ( n21153, n21154, n21155 );
nor U132312 ( n21152, n21157, n73191 );
nor U132313 ( n21155, P1_P1_STATE2_REG_0_, n21156 );
nor U132314 ( n21157, n21158, n74649 );
nor U132315 ( n21158, P1_P1_STATE2_REG_1_, n21127 );
nand U132316 ( n21208, n21201, n21260 );
nand U132317 ( n21260, P1_P1_INSTQUEUERD_ADDR_REG_0_, n21199 );
nor U132318 ( n21205, P1_P1_INSTQUEUERD_ADDR_REG_1_, n21207 );
nor U132319 ( n21207, n4842, n21208 );
nand U132320 ( n21162, n21163, n21164 );
nand U132321 ( n21164, n8320, n21165 );
nand U132322 ( n21163, n21180, n75031 );
or U132323 ( n21165, P1_P1_MORE_REG, P1_P1_FLUSH_REG );
xor U132324 ( n13288, n76035, P1_P1_INSTADDRPOINTER_REG_20_ );
xor U132325 ( n12973, n76035, P1_P1_INSTADDRPOINTER_REG_26_ );
nand U132326 ( n35634, n185, P1_P3_STATE2_REG_1_ );
nand U132327 ( n28455, n148, P1_P2_STATE2_REG_1_ );
nand U132328 ( n70360, n457, P2_P3_STATE2_REG_1_ );
nand U132329 ( n61760, n420, P2_P2_STATE2_REG_1_ );
nand U132330 ( n3601, n35628, n35629 );
nand U132331 ( n35629, P1_P3_STATE2_REG_1_, n35630 );
nand U132332 ( n35628, P1_P3_STATE2_REG_2_, n35634 );
nand U132333 ( n35630, n35631, n35632 );
nand U132334 ( n5846, n28449, n28450 );
nand U132335 ( n28450, P1_P2_STATE2_REG_1_, n28451 );
nand U132336 ( n28449, P1_P2_STATE2_REG_2_, n28455 );
nand U132337 ( n28451, n28452, n28453 );
nand U132338 ( n10336, n70354, n70355 );
nand U132339 ( n70355, P2_P3_STATE2_REG_1_, n70356 );
nand U132340 ( n70354, P2_P3_STATE2_REG_2_, n70360 );
nand U132341 ( n70356, n70357, n70358 );
nand U132342 ( n12581, n61754, n61755 );
nand U132343 ( n61755, P2_P2_STATE2_REG_1_, n61756 );
nand U132344 ( n61754, P2_P2_STATE2_REG_2_, n61760 );
nand U132345 ( n61756, n61757, n61758 );
nand U132346 ( n54132, n490, P2_P1_STATE2_REG_1_ );
nand U132347 ( n14826, n54126, n54127 );
nand U132348 ( n54127, P2_P1_STATE2_REG_1_, n54128 );
nand U132349 ( n54126, P2_P1_STATE2_REG_2_, n54132 );
nand U132350 ( n54128, n54129, n54130 );
nand U132351 ( n54081, n54082, n54083 );
nor U132352 ( n54082, P2_P1_ADDRESS_REG_0_, n54086 );
nor U132353 ( n54083, n54084, n54085 );
nand U132354 ( n54086, n73064, n74273 );
nand U132355 ( n42216, P3_REG1_REG_1_, n45201 );
nand U132356 ( n54080, n54087, n54088 );
nor U132357 ( n54088, n54089, n54090 );
nor U132358 ( n54087, P2_P1_ADDRESS_REG_16_, n54091 );
or U132359 ( n54089, P2_P1_ADDRESS_REG_20_, P2_P1_ADDRESS_REG_21_ );
nand U132360 ( n42211, P3_REG2_REG_1_, n45201 );
and U132361 ( n16470, n17054, P4_DATAO_REG_0_ );
xnor U132362 ( n28641, n28915, n28916 );
xor U132363 ( n28916, P1_P2_INSTQUEUEWR_ADDR_REG_2_, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
xnor U132364 ( n61946, n62220, n62221 );
xor U132365 ( n62221, P2_P2_INSTQUEUEWR_ADDR_REG_2_, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
xnor U132366 ( n70546, n70820, n70821 );
xor U132367 ( n70821, P2_P3_INSTQUEUEWR_ADDR_REG_2_, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
xnor U132368 ( n35820, n36094, n36095 );
xor U132369 ( n36095, P1_P3_INSTQUEUEWR_ADDR_REG_2_, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nor U132370 ( n30195, n30196, n74979 );
nor U132371 ( n30196, n30197, n30198 );
nor U132372 ( n30197, P1_P3_EBX_REG_21_, n76489 );
nor U132373 ( n30218, n30219, n74933 );
nor U132374 ( n30219, n30220, n30221 );
nor U132375 ( n30220, P1_P3_EBX_REG_19_, n76489 );
nor U132376 ( n30237, n30238, n74893 );
nor U132377 ( n30238, n30239, n30240 );
nor U132378 ( n30239, P1_P3_EBX_REG_17_, n76489 );
nor U132379 ( n30256, n30257, n74832 );
nor U132380 ( n30257, n30258, n30259 );
nor U132381 ( n30258, P1_P3_EBX_REG_15_, n76489 );
nand U132382 ( n21188, n21249, n21250 );
nand U132383 ( n21249, n223, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U132384 ( n21250, n14785, n21202 );
nor U132385 ( n30157, n30158, n75072 );
nor U132386 ( n30158, n30159, n30160 );
nor U132387 ( n30159, P1_P3_EBX_REG_25_, n76489 );
nor U132388 ( n30176, n30177, n75022 );
nor U132389 ( n30177, n30178, n30179 );
nor U132390 ( n30178, P1_P3_EBX_REG_23_, n76489 );
nor U132391 ( n30131, n30132, n75181 );
nor U132392 ( n30132, n30133, n30134 );
nor U132393 ( n30133, P1_P3_EBX_REG_28_, n76489 );
nor U132394 ( n43497, n43498, n74978 );
nor U132395 ( n43498, n43499, n43500 );
nor U132396 ( n43499, P2_P1_EBX_REG_21_, n76363 );
nor U132397 ( n43516, n43517, n74932 );
nor U132398 ( n43517, n43518, n43519 );
nor U132399 ( n43518, P2_P1_EBX_REG_19_, n76363 );
nor U132400 ( n43535, n43536, n74892 );
nor U132401 ( n43536, n43537, n43538 );
nor U132402 ( n43537, P2_P1_EBX_REG_17_, n76363 );
nor U132403 ( n43567, n43568, n74831 );
nor U132404 ( n43568, n43569, n43570 );
nor U132405 ( n43569, P2_P1_EBX_REG_15_, n76363 );
nor U132406 ( n9547, n9548, n74981 );
nor U132407 ( n9548, n9549, n9550 );
nor U132408 ( n9549, P1_P1_EBX_REG_21_, n76633 );
nor U132409 ( n9570, n9572, n74935 );
nor U132410 ( n9572, n9573, n9574 );
nor U132411 ( n9573, P1_P1_EBX_REG_19_, n76633 );
nor U132412 ( n9593, n9594, n74895 );
nor U132413 ( n9594, n9595, n9597 );
nor U132414 ( n9595, P1_P1_EBX_REG_17_, n76633 );
nor U132415 ( n9617, n9618, n74834 );
nor U132416 ( n9618, n9619, n9620 );
nor U132417 ( n9619, P1_P1_EBX_REG_15_, n76633 );
nor U132418 ( n64261, n64262, n74980 );
nor U132419 ( n64262, n64263, n64264 );
nor U132420 ( n64263, P2_P3_EBX_REG_21_, n76222 );
nor U132421 ( n64280, n64281, n74934 );
nor U132422 ( n64281, n64282, n64283 );
nor U132423 ( n64282, P2_P3_EBX_REG_19_, n76222 );
nor U132424 ( n64299, n64300, n74894 );
nor U132425 ( n64300, n64301, n64302 );
nor U132426 ( n64301, P2_P3_EBX_REG_17_, n76222 );
nor U132427 ( n64318, n64319, n74833 );
nor U132428 ( n64319, n64320, n64321 );
nor U132429 ( n64320, P2_P3_EBX_REG_15_, n76222 );
nor U132430 ( n43459, n43460, n75071 );
nor U132431 ( n43460, n43461, n43462 );
nor U132432 ( n43461, P2_P1_EBX_REG_25_, n76363 );
nor U132433 ( n43478, n43479, n75021 );
nor U132434 ( n43479, n43480, n43481 );
nor U132435 ( n43480, P2_P1_EBX_REG_23_, n76363 );
nor U132436 ( n64170, n64171, n75073 );
nor U132437 ( n64171, n64172, n64173 );
nor U132438 ( n64172, P2_P3_EBX_REG_25_, n76222 );
nor U132439 ( n55946, n55947, n75076 );
nor U132440 ( n55947, n55948, n55949 );
nor U132441 ( n55948, P2_P2_EBX_REG_25_, n76284 );
nor U132442 ( n55968, n55969, n75026 );
nor U132443 ( n55969, n55970, n55971 );
nor U132444 ( n55970, P2_P2_EBX_REG_23_, n76284 );
nor U132445 ( n9499, n9500, n75075 );
nor U132446 ( n9500, n9502, n9503 );
nor U132447 ( n9502, P1_P1_EBX_REG_25_, n76633 );
nor U132448 ( n43400, n43401, n75190 );
nor U132449 ( n43401, n43402, n43403 );
nor U132450 ( n43402, P2_P1_EBX_REG_28_, n76363 );
nor U132451 ( n64242, n64243, n75023 );
nor U132452 ( n64243, n64244, n64245 );
nor U132453 ( n64244, P2_P3_EBX_REG_23_, n76222 );
nor U132454 ( n22832, n22833, n75074 );
nor U132455 ( n22833, n22834, n22835 );
nor U132456 ( n22834, P1_P2_EBX_REG_25_, n76542 );
nor U132457 ( n9523, n9524, n75025 );
nor U132458 ( n9524, n9525, n9527 );
nor U132459 ( n9525, P1_P1_EBX_REG_23_, n76633 );
nor U132460 ( n22851, n22852, n75024 );
nor U132461 ( n22852, n22853, n22854 );
nor U132462 ( n22853, P1_P2_EBX_REG_23_, n76542 );
nor U132463 ( n22872, n22873, n74982 );
nor U132464 ( n22873, n22874, n22875 );
nor U132465 ( n22874, P1_P2_EBX_REG_21_, n76542 );
nor U132466 ( n22891, n22892, n74936 );
nor U132467 ( n22892, n22893, n22894 );
nor U132468 ( n22893, P1_P2_EBX_REG_19_, n76542 );
nor U132469 ( n22910, n22911, n74896 );
nor U132470 ( n22911, n22912, n22913 );
nor U132471 ( n22912, P1_P2_EBX_REG_17_, n76542 );
nor U132472 ( n22929, n22930, n74835 );
nor U132473 ( n22930, n22931, n22932 );
nor U132474 ( n22931, P1_P2_EBX_REG_15_, n76542 );
nor U132475 ( n64144, n64145, n75182 );
nor U132476 ( n64145, n64146, n64147 );
nor U132477 ( n64146, P2_P3_EBX_REG_28_, n76222 );
nor U132478 ( n22806, n22807, n75183 );
nor U132479 ( n22807, n22808, n22809 );
nor U132480 ( n22808, P1_P2_EBX_REG_28_, n76542 );
nor U132481 ( n9467, n9468, n75189 );
nor U132482 ( n9468, n9469, n9470 );
nor U132483 ( n9469, P1_P1_EBX_REG_28_, n76633 );
nor U132484 ( n55987, n55988, n74983 );
nor U132485 ( n55988, n55989, n55990 );
nor U132486 ( n55989, P2_P2_EBX_REG_21_, n76284 );
nor U132487 ( n56006, n56007, n74937 );
nor U132488 ( n56007, n56008, n56009 );
nor U132489 ( n56008, P2_P2_EBX_REG_19_, n76284 );
nor U132490 ( n56025, n56026, n74897 );
nor U132491 ( n56026, n56027, n56028 );
nor U132492 ( n56027, P2_P2_EBX_REG_17_, n76284 );
nor U132493 ( n56044, n56045, n74836 );
nor U132494 ( n56045, n56046, n56047 );
nor U132495 ( n56046, P2_P2_EBX_REG_15_, n76284 );
nor U132496 ( n55920, n55921, n75184 );
nor U132497 ( n55921, n55922, n55923 );
nor U132498 ( n55922, P2_P2_EBX_REG_28_, n76284 );
nor U132499 ( n30387, n30388, n74531 );
nor U132500 ( n30388, n30389, n30390 );
nor U132501 ( n30389, P1_P3_EBX_REG_1_, n76490 );
nor U132502 ( n30317, n30318, n74719 );
nor U132503 ( n30318, n30319, n30320 );
nor U132504 ( n30319, P1_P3_EBX_REG_9_, n76490 );
nor U132505 ( n30275, n30276, n74792 );
nor U132506 ( n30276, n30277, n30278 );
nor U132507 ( n30277, P1_P3_EBX_REG_13_, n76490 );
nor U132508 ( n30294, n30295, n74762 );
nor U132509 ( n30295, n30296, n30297 );
nor U132510 ( n30296, P1_P3_EBX_REG_11_, n76490 );
nor U132511 ( n30336, n30337, n74664 );
nor U132512 ( n30337, n30338, n30339 );
nor U132513 ( n30338, P1_P3_EBX_REG_7_, n76490 );
nor U132514 ( n30353, n30354, n74601 );
nor U132515 ( n30354, n30355, n30356 );
nor U132516 ( n30355, P1_P3_EBX_REG_5_, n76490 );
nor U132517 ( n30370, n30371, n74568 );
nor U132518 ( n30371, n30372, n30373 );
nor U132519 ( n30372, P1_P3_EBX_REG_3_, n76490 );
nand U132520 ( n5131, n30350, n30351 );
nand U132521 ( n30351, n3072, P1_P3_INSTQUEUE_REG_0__6_ );
nor U132522 ( n30350, n30352, n30353 );
nor U132523 ( n30352, n30357, n30358 );
nand U132524 ( n5121, n30367, n30368 );
nand U132525 ( n30368, n3072, P1_P3_INSTQUEUE_REG_0__4_ );
nor U132526 ( n30367, n30369, n30370 );
nor U132527 ( n30369, n30374, n30375 );
nand U132528 ( n5111, n30384, n30385 );
nand U132529 ( n30385, n3072, P1_P3_INSTQUEUE_REG_0__2_ );
nor U132530 ( n30384, n30386, n30387 );
nor U132531 ( n30386, n30391, n30392 );
nor U132532 ( n9640, n9642, n74794 );
nor U132533 ( n9642, n9643, n9644 );
nor U132534 ( n9643, P1_P1_EBX_REG_13_, n76634 );
nor U132535 ( n9668, n9669, n74764 );
nor U132536 ( n9669, n9670, n9672 );
nor U132537 ( n9670, P1_P1_EBX_REG_11_, n76634 );
nor U132538 ( n9715, n9717, n74665 );
nor U132539 ( n9717, n9718, n9719 );
nor U132540 ( n9718, P1_P1_EBX_REG_7_, n76634 );
nor U132541 ( n9737, n9738, n74602 );
nor U132542 ( n9738, n9739, n9740 );
nor U132543 ( n9739, P1_P1_EBX_REG_5_, n76634 );
nor U132544 ( n9758, n9759, n74569 );
nor U132545 ( n9759, n9760, n9762 );
nor U132546 ( n9760, P1_P1_EBX_REG_3_, n76634 );
nor U132547 ( n43586, n43587, n74795 );
nor U132548 ( n43587, n43588, n43589 );
nor U132549 ( n43588, P2_P1_EBX_REG_13_, n76364 );
nor U132550 ( n43605, n43606, n74765 );
nor U132551 ( n43606, n43607, n43608 );
nor U132552 ( n43607, P2_P1_EBX_REG_11_, n76364 );
nor U132553 ( n43643, n43644, n74667 );
nor U132554 ( n43644, n43645, n43646 );
nor U132555 ( n43645, P2_P1_EBX_REG_7_, n76364 );
nor U132556 ( n43674, n43675, n74604 );
nor U132557 ( n43675, n43676, n43677 );
nor U132558 ( n43676, P2_P1_EBX_REG_5_, n76364 );
nor U132559 ( n43691, n43692, n74571 );
nor U132560 ( n43692, n43693, n43694 );
nor U132561 ( n43693, P2_P1_EBX_REG_3_, n76364 );
nor U132562 ( n64550, n64551, n74534 );
nor U132563 ( n64551, n64552, n64553 );
nor U132564 ( n64552, P2_P3_EBX_REG_1_, n76223 );
nor U132565 ( n43708, n43709, n74536 );
nor U132566 ( n43709, n43710, n43711 );
nor U132567 ( n43710, P2_P1_EBX_REG_1_, n76364 );
nor U132568 ( n64436, n64437, n74720 );
nor U132569 ( n64437, n64438, n64439 );
nor U132570 ( n64438, P2_P3_EBX_REG_9_, n76223 );
nor U132571 ( n9692, n9693, n74721 );
nor U132572 ( n9693, n9694, n9695 );
nor U132573 ( n9694, P1_P1_EBX_REG_9_, n76634 );
nor U132574 ( n43624, n43625, n74722 );
nor U132575 ( n43625, n43626, n43627 );
nor U132576 ( n43626, P2_P1_EBX_REG_9_, n76364 );
nor U132577 ( n64398, n64399, n74793 );
nor U132578 ( n64399, n64400, n64401 );
nor U132579 ( n64400, P2_P3_EBX_REG_13_, n76223 );
nor U132580 ( n64417, n64418, n74763 );
nor U132581 ( n64418, n64419, n64420 );
nor U132582 ( n64419, P2_P3_EBX_REG_11_, n76223 );
nor U132583 ( n64455, n64456, n74666 );
nor U132584 ( n64456, n64457, n64458 );
nor U132585 ( n64457, P2_P3_EBX_REG_7_, n76223 );
nor U132586 ( n64472, n64473, n74603 );
nor U132587 ( n64473, n64474, n64475 );
nor U132588 ( n64474, P2_P3_EBX_REG_5_, n76223 );
nor U132589 ( n64533, n64534, n74570 );
nor U132590 ( n64534, n64535, n64536 );
nor U132591 ( n64535, P2_P3_EBX_REG_3_, n76223 );
nor U132592 ( n9783, n9784, n74533 );
nor U132593 ( n9784, n9785, n9787 );
nor U132594 ( n9785, P1_P1_EBX_REG_1_, n76634 );
nand U132595 ( n11866, n64469, n64470 );
nand U132596 ( n64470, n5673, P2_P3_INSTQUEUE_REG_0__6_ );
nor U132597 ( n64469, n64471, n64472 );
nor U132598 ( n64471, n64476, n64477 );
nand U132599 ( n11856, n64530, n64531 );
nand U132600 ( n64531, n5673, P2_P3_INSTQUEUE_REG_0__4_ );
nor U132601 ( n64530, n64532, n64533 );
nor U132602 ( n64532, n64537, n64538 );
nand U132603 ( n16356, n43671, n43672 );
nand U132604 ( n43672, n7458, P2_P1_INSTQUEUE_REG_0__6_ );
nor U132605 ( n43671, n43673, n43674 );
nor U132606 ( n43673, n43678, n43679 );
nand U132607 ( n16346, n43688, n43689 );
nand U132608 ( n43689, n7458, P2_P1_INSTQUEUE_REG_0__4_ );
nor U132609 ( n43688, n43690, n43691 );
nor U132610 ( n43690, n43695, n43696 );
nand U132611 ( n9621, n9733, n9734 );
nand U132612 ( n9734, n4814, P1_P1_INSTQUEUE_REG_0__6_ );
nor U132613 ( n9733, n9735, n9737 );
nor U132614 ( n9735, n9742, n9743 );
nand U132615 ( n9611, n9754, n9755 );
nand U132616 ( n9755, n4814, P1_P1_INSTQUEUE_REG_0__4_ );
nor U132617 ( n9754, n9757, n9758 );
nor U132618 ( n9757, n9763, n9764 );
nand U132619 ( n9601, n9779, n9780 );
nand U132620 ( n9780, n4814, P1_P1_INSTQUEUE_REG_0__2_ );
nor U132621 ( n9779, n9782, n9783 );
nor U132622 ( n9782, n9788, n9789 );
nand U132623 ( n11846, n64547, n64548 );
nand U132624 ( n64548, n5673, P2_P3_INSTQUEUE_REG_0__2_ );
nor U132625 ( n64547, n64549, n64550 );
nor U132626 ( n64549, n64554, n64555 );
nand U132627 ( n16336, n43705, n43706 );
nand U132628 ( n43706, n7458, P2_P1_INSTQUEUE_REG_0__2_ );
nor U132629 ( n43705, n43707, n43708 );
nor U132630 ( n43707, n43712, n43713 );
nor U132631 ( n23060, n23061, n74532 );
nor U132632 ( n23061, n23062, n23063 );
nor U132633 ( n23062, P1_P2_EBX_REG_1_, n76543 );
nor U132634 ( n56181, n56182, n74535 );
nor U132635 ( n56182, n56183, n56184 );
nor U132636 ( n56183, P2_P2_EBX_REG_1_, n76285 );
nor U132637 ( n22988, n22989, n74723 );
nor U132638 ( n22989, n22990, n22991 );
nor U132639 ( n22990, P1_P2_EBX_REG_9_, n76543 );
nor U132640 ( n56104, n56105, n74724 );
nor U132641 ( n56105, n56106, n56107 );
nor U132642 ( n56106, P2_P2_EBX_REG_9_, n76285 );
nor U132643 ( n22948, n22949, n74796 );
nor U132644 ( n22949, n22950, n22951 );
nor U132645 ( n22950, P1_P2_EBX_REG_13_, n76543 );
nor U132646 ( n22969, n22970, n74766 );
nor U132647 ( n22970, n22971, n22972 );
nor U132648 ( n22971, P1_P2_EBX_REG_11_, n76543 );
nor U132649 ( n23007, n23008, n74668 );
nor U132650 ( n23008, n23009, n23010 );
nor U132651 ( n23009, P1_P2_EBX_REG_7_, n76543 );
nor U132652 ( n23024, n23025, n74605 );
nor U132653 ( n23025, n23026, n23027 );
nor U132654 ( n23026, P1_P2_EBX_REG_5_, n76543 );
nor U132655 ( n23041, n23042, n74572 );
nor U132656 ( n23042, n23043, n23044 );
nor U132657 ( n23043, P1_P2_EBX_REG_3_, n76543 );
nor U132658 ( n56066, n56067, n74797 );
nor U132659 ( n56067, n56068, n56069 );
nor U132660 ( n56068, P2_P2_EBX_REG_13_, n76285 );
nor U132661 ( n56085, n56086, n74767 );
nor U132662 ( n56086, n56087, n56088 );
nor U132663 ( n56087, P2_P2_EBX_REG_11_, n76285 );
nor U132664 ( n56123, n56124, n74669 );
nor U132665 ( n56124, n56125, n56126 );
nor U132666 ( n56125, P2_P2_EBX_REG_7_, n76285 );
nor U132667 ( n56140, n56141, n74606 );
nor U132668 ( n56141, n56142, n56143 );
nor U132669 ( n56142, P2_P2_EBX_REG_5_, n76285 );
nor U132670 ( n56160, n56161, n74573 );
nor U132671 ( n56161, n56162, n56163 );
nor U132672 ( n56162, P2_P2_EBX_REG_3_, n76285 );
nand U132673 ( n7376, n23021, n23022 );
nand U132674 ( n23022, n76757, P1_P2_INSTQUEUE_REG_0__6_ );
nor U132675 ( n23021, n23023, n23024 );
nor U132676 ( n23023, n23028, n23029 );
nand U132677 ( n7366, n23038, n23039 );
nand U132678 ( n23039, n76757, P1_P2_INSTQUEUE_REG_0__4_ );
nor U132679 ( n23038, n23040, n23041 );
nor U132680 ( n23040, n23045, n23046 );
nand U132681 ( n7356, n23057, n23058 );
nand U132682 ( n23058, n76757, P1_P2_INSTQUEUE_REG_0__2_ );
nor U132683 ( n23057, n23059, n23060 );
nor U132684 ( n23059, n23064, n23065 );
nand U132685 ( n14111, n56137, n56138 );
nand U132686 ( n56138, n76690, P2_P2_INSTQUEUE_REG_0__6_ );
nor U132687 ( n56137, n56139, n56140 );
nor U132688 ( n56139, n56144, n56145 );
nand U132689 ( n14101, n56157, n56158 );
nand U132690 ( n56158, n76690, P2_P2_INSTQUEUE_REG_0__4_ );
nor U132691 ( n56157, n56159, n56160 );
nor U132692 ( n56159, n56164, n56165 );
nand U132693 ( n14091, n56178, n56179 );
nand U132694 ( n56179, n76690, P2_P2_INSTQUEUE_REG_0__2_ );
nor U132695 ( n56178, n56180, n56181 );
nor U132696 ( n56180, n56185, n56186 );
or U132697 ( n54090, P2_P1_ADDRESS_REG_19_, P2_P1_ADDRESS_REG_1_ );
nand U132698 ( n21134, P1_P1_STATE2_REG_0_, n21124 );
and U132699 ( n54070, n75946, n75947 );
nor U132700 ( n75946, P2_P1_ADDRESS_REG_27_, P2_P1_ADDRESS_REG_28_ );
nor U132701 ( n75947, P2_P1_ADDRESS_REG_25_, P2_P1_ADDRESS_REG_26_ );
nand U132702 ( n16723, n17401, DIN_30_ );
or U132703 ( n54073, P2_P1_ADDRESS_REG_23_, P2_P1_ADDRESS_REG_24_ );
nand U132704 ( n21608, P1_P1_INSTQUEUERD_ADDR_REG_0_, n74435 );
nand U132705 ( n21606, n21614, n21615 );
nand U132706 ( n21614, n21617, n73525 );
nand U132707 ( n21615, P1_P1_INSTQUEUEWR_ADDR_REG_3_, n21616 );
or U132708 ( n21616, n21617, n73525 );
nand U132709 ( n21339, n21611, n21612 );
xnor U132710 ( n21611, n21618, n21617 );
nand U132711 ( n21612, n21613, P1_P1_INSTQUEUEWR_ADDR_REG_4_ );
xor U132712 ( n21618, n74538, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U132713 ( n21609, n21622, n21623 );
nand U132714 ( n21622, n21608, n73060 );
nand U132715 ( n21623, P1_P1_INSTQUEUEWR_ADDR_REG_1_, n21624 );
nand U132716 ( n21624, P1_P1_INSTQUEUERD_ADDR_REG_1_, n5165 );
nor U132717 ( n21613, P1_P1_INSTQUEUERD_ADDR_REG_4_, n5140 );
nand U132718 ( n21617, n21619, n21620 );
nand U132719 ( n21619, n21609, n73527 );
nand U132720 ( n21620, P1_P1_INSTQUEUEWR_ADDR_REG_2_, n21621 );
or U132721 ( n21621, n73527, n21609 );
nor U132722 ( n35709, n35710, n35711 );
nor U132723 ( n35711, P1_P3_INSTQUEUERD_ADDR_REG_1_, n35687 );
nor U132724 ( n35710, n3403, n35712 );
and U132725 ( n35712, n34061, n35713 );
nor U132726 ( n28530, n28531, n28532 );
nor U132727 ( n28532, P1_P2_INSTQUEUERD_ADDR_REG_1_, n28508 );
nor U132728 ( n28531, n4240, n28533 );
and U132729 ( n28533, n26816, n28534 );
nor U132730 ( n70435, n70436, n70437 );
nor U132731 ( n70437, P2_P3_INSTQUEUERD_ADDR_REG_1_, n70413 );
nor U132732 ( n70436, n6018, n70438 );
and U132733 ( n70438, n68815, n70439 );
nor U132734 ( n61835, n61836, n61837 );
nor U132735 ( n61837, P2_P2_INSTQUEUERD_ADDR_REG_1_, n61813 );
nor U132736 ( n61836, n6873, n61838 );
and U132737 ( n61838, n59956, n61839 );
nor U132738 ( n54207, n54208, n54209 );
nor U132739 ( n54209, P2_P1_INSTQUEUERD_ADDR_REG_1_, n54185 );
nor U132740 ( n54208, n7805, n54210 );
and U132741 ( n54210, n47795, n54211 );
nand U132742 ( n21149, n219, P1_P1_STATE2_REG_1_ );
nand U132743 ( n8091, n21143, n21144 );
nand U132744 ( n21144, P1_P1_STATE2_REG_1_, n21145 );
nand U132745 ( n21143, P1_P1_STATE2_REG_2_, n21149 );
nand U132746 ( n21145, n21146, n21147 );
nand U132747 ( n8831, n13894, n13895 );
nand U132748 ( n13895, n76888, P1_P1_INSTADDRPOINTER_REG_7_ );
nor U132749 ( n13894, n13897, n13898 );
nor U132750 ( n13898, n73207, n76598 );
nand U132751 ( n35668, n35718, n35719 );
nand U132752 ( n35718, n189, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U132753 ( n35719, n34261, n35678 );
nand U132754 ( n28489, n28539, n28540 );
nand U132755 ( n28539, n152, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U132756 ( n28540, n27018, n28499 );
nand U132757 ( n70394, n70444, n70445 );
nand U132758 ( n70444, n460, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U132759 ( n70445, n69015, n70404 );
nand U132760 ( n61794, n61844, n61845 );
nand U132761 ( n61844, n424, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U132762 ( n61845, n60159, n61804 );
nor U132763 ( n35722, n31169, n35740 );
nand U132764 ( n35740, P1_P3_INSTQUEUERD_ADDR_REG_1_, n35693 );
nor U132765 ( n28543, n23877, n28561 );
nand U132766 ( n28561, P1_P2_INSTQUEUERD_ADDR_REG_1_, n28514 );
nor U132767 ( n70448, n65423, n70466 );
nand U132768 ( n70466, P2_P3_INSTQUEUERD_ADDR_REG_1_, n70419 );
nor U132769 ( n61848, n57001, n61866 );
nand U132770 ( n61866, P2_P2_INSTQUEUERD_ADDR_REG_1_, n61819 );
xor U132771 ( n12463, n13784, P1_P1_INSTADDRPOINTER_REG_9_ );
nand U132772 ( n54166, n54216, n54217 );
nand U132773 ( n54216, n494, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U132774 ( n54217, n48007, n54176 );
nor U132775 ( n54220, n44548, n54238 );
nand U132776 ( n54238, P2_P1_INSTQUEUERD_ADDR_REG_1_, n54191 );
xor U132777 ( n32415, n33455, P1_P3_INSTADDRPOINTER_REG_9_ );
xor U132778 ( n46114, n47175, P2_P1_INSTADDRPOINTER_REG_9_ );
xor U132779 ( n67078, n68206, P2_P3_INSTADDRPOINTER_REG_9_ );
xor U132780 ( n25180, n26205, P1_P2_INSTADDRPOINTER_REG_9_ );
xor U132781 ( n58316, n59344, P2_P2_INSTADDRPOINTER_REG_9_ );
nor U132782 ( n21254, n21255, n73527 );
nor U132783 ( n21255, n21256, n21257 );
nor U132784 ( n21257, P1_P1_INSTQUEUERD_ADDR_REG_1_, n21201 );
nor U132785 ( n21256, n5150, n21258 );
nand U132786 ( n54591, P2_P1_INSTQUEUERD_ADDR_REG_0_, n74442 );
nand U132787 ( n54589, n54597, n54598 );
nand U132788 ( n54597, n54600, n73497 );
nand U132789 ( n54598, P2_P1_INSTQUEUEWR_ADDR_REG_3_, n54599 );
or U132790 ( n54599, n54600, n73497 );
nand U132791 ( n54592, n54605, n54606 );
nand U132792 ( n54605, n54591, n73052 );
nand U132793 ( n54606, P2_P1_INSTQUEUEWR_ADDR_REG_1_, n54607 );
nand U132794 ( n54607, P2_P1_INSTQUEUERD_ADDR_REG_1_, n7820 );
nor U132795 ( n54596, P2_P1_INSTQUEUERD_ADDR_REG_4_, n7795 );
nand U132796 ( n54322, n54594, n54595 );
xnor U132797 ( n54594, n54601, n54600 );
nand U132798 ( n54595, n54596, P2_P1_INSTQUEUEWR_ADDR_REG_4_ );
xor U132799 ( n54601, n74525, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U132800 ( n54600, n54602, n54603 );
nand U132801 ( n54602, n54592, n73511 );
nand U132802 ( n54603, P2_P1_INSTQUEUEWR_ADDR_REG_2_, n54604 );
or U132803 ( n54604, n73511, n54592 );
nand U132804 ( n63034, n64101, n64102 );
nor U132805 ( n64102, n477, n64094 );
and U132806 ( n64101, n64092, P2_P3_EBX_REG_31_ );
nand U132807 ( n29267, n30084, n30085 );
nor U132808 ( n30085, n205, n30077 );
and U132809 ( n30084, n30075, P1_P3_EBX_REG_31_ );
nand U132810 ( n21950, n22763, n22764 );
nor U132811 ( n22764, n172, n22756 );
and U132812 ( n22763, n22754, P1_P2_EBX_REG_31_ );
nand U132813 ( n55062, n55877, n55878 );
nor U132814 ( n55878, n444, n55870 );
and U132815 ( n55877, n55868, P2_P2_EBX_REG_31_ );
nand U132816 ( n63196, n63197, n63198 );
nand U132817 ( n63197, P2_P3_REIP_REG_25_, n63201 );
nand U132818 ( n63198, P2_P3_EBX_REG_25_, n63199 );
nand U132819 ( n63201, n63202, n63203 );
nand U132820 ( n63363, n63364, n63365 );
or U132821 ( n63364, n74944, n63331 );
nand U132822 ( n63365, P2_P3_EBX_REG_21_, n63366 );
nand U132823 ( n63366, n63064, n63367 );
nand U132824 ( n29433, n29434, n29435 );
nand U132825 ( n29434, P1_P3_REIP_REG_25_, n29438 );
nand U132826 ( n29435, P1_P3_EBX_REG_25_, n29436 );
nand U132827 ( n29438, n29439, n29440 );
nand U132828 ( n29534, n29535, n29536 );
or U132829 ( n29535, n74945, n29502 );
nand U132830 ( n29536, P1_P3_EBX_REG_21_, n29537 );
nand U132831 ( n29537, n29297, n29538 );
nand U132832 ( n22215, n22216, n22217 );
or U132833 ( n22216, n74939, n22183 );
nand U132834 ( n22217, P1_P2_EBX_REG_21_, n22218 );
nand U132835 ( n22218, n21982, n22219 );
nand U132836 ( n22114, n22115, n22116 );
nand U132837 ( n22115, P1_P2_REIP_REG_25_, n22119 );
nand U132838 ( n22116, P1_P2_EBX_REG_25_, n22117 );
nand U132839 ( n22119, n22120, n22121 );
nand U132840 ( n55329, n55330, n55331 );
or U132841 ( n55330, n74938, n55297 );
nand U132842 ( n55331, P2_P2_EBX_REG_21_, n55332 );
nand U132843 ( n55332, n55092, n55333 );
nand U132844 ( n55224, n55225, n55226 );
nand U132845 ( n55225, P2_P2_REIP_REG_25_, n55229 );
nand U132846 ( n55226, P2_P2_EBX_REG_25_, n55227 );
nand U132847 ( n55229, n55230, n55231 );
nand U132848 ( n63529, n63530, n63531 );
nand U132849 ( n63531, n63532, n76226 );
nand U132850 ( n63530, P2_P3_EBX_REG_17_, n63533 );
xor U132851 ( n63532, n63516, n63515 );
nand U132852 ( n29630, n29631, n29632 );
nand U132853 ( n29632, n29633, n76493 );
nand U132854 ( n29631, P1_P3_EBX_REG_17_, n29634 );
xor U132855 ( n29633, n29617, n29616 );
nand U132856 ( n22309, n22310, n22311 );
nand U132857 ( n22311, n22312, n76546 );
nand U132858 ( n22310, P1_P2_EBX_REG_17_, n22313 );
xor U132859 ( n22312, n22296, n22295 );
nand U132860 ( n55421, n55422, n55423 );
nand U132861 ( n55423, n55424, n76292 );
nand U132862 ( n55422, P2_P2_EBX_REG_17_, n55425 );
xor U132863 ( n55424, n55408, n55407 );
nand U132864 ( n63234, n63235, n63236 );
nand U132865 ( n63236, n63219, n63237 );
nand U132866 ( n63235, P2_P3_EBX_REG_23_, n63239 );
nand U132867 ( n63237, n63052, n63238 );
nand U132868 ( n29471, n29472, n29473 );
nand U132869 ( n29473, n29456, n29474 );
nand U132870 ( n29472, P1_P3_EBX_REG_23_, n29476 );
nand U132871 ( n29474, n29285, n29475 );
nand U132872 ( n22152, n22153, n22154 );
nand U132873 ( n22154, n22137, n22155 );
nand U132874 ( n22153, P1_P2_EBX_REG_23_, n22157 );
nand U132875 ( n22155, n21970, n22156 );
nand U132876 ( n55266, n55267, n55268 );
nand U132877 ( n55268, n55247, n55269 );
nand U132878 ( n55267, P2_P2_EBX_REG_23_, n55271 );
nand U132879 ( n55269, n55080, n55270 );
nand U132880 ( n63806, n63812, n63813 );
nand U132881 ( n63812, n63785, n73216 );
nand U132882 ( n63813, P2_P3_EBX_REG_9_, n63814 );
nand U132883 ( n63814, n63064, n63815 );
nand U132884 ( n29850, n29856, n29857 );
nand U132885 ( n29856, n29825, n73217 );
nand U132886 ( n29857, P1_P3_EBX_REG_9_, n29858 );
nand U132887 ( n29858, n29297, n29859 );
nand U132888 ( n22527, n22533, n22534 );
nand U132889 ( n22533, n22506, n73215 );
nand U132890 ( n22534, P1_P2_EBX_REG_9_, n22535 );
nand U132891 ( n22535, n21982, n22536 );
nand U132892 ( n55640, n55646, n55647 );
nand U132893 ( n55646, n55619, n73214 );
nand U132894 ( n55647, P2_P2_EBX_REG_9_, n55648 );
nand U132895 ( n55648, n55092, n55649 );
nand U132896 ( n63144, n63145, n63146 );
or U132897 ( n63145, n75003, n63112 );
nand U132898 ( n63146, P2_P3_EBX_REG_27_, n63147 );
nand U132899 ( n63147, n63064, n63148 );
nand U132900 ( n29381, n29382, n29383 );
or U132901 ( n29382, n75004, n29349 );
nand U132902 ( n29383, P1_P3_EBX_REG_27_, n29384 );
nand U132903 ( n29384, n29297, n29385 );
nand U132904 ( n22062, n22063, n22064 );
or U132905 ( n22063, n74999, n22030 );
nand U132906 ( n22064, P1_P2_EBX_REG_27_, n22065 );
nand U132907 ( n22065, n21982, n22066 );
nand U132908 ( n55172, n55173, n55174 );
or U132909 ( n55173, n75000, n55140 );
nand U132910 ( n55174, P2_P2_EBX_REG_27_, n55175 );
nand U132911 ( n55175, n55092, n55176 );
nor U132912 ( n45198, P3_REG2_REG_2_, n42229 );
nor U132913 ( n45263, P3_REG1_REG_2_, n42229 );
nand U132914 ( n63588, n63594, n63595 );
nand U132915 ( n63595, n63557, n63596 );
nand U132916 ( n63594, P2_P3_EBX_REG_15_, n63598 );
nand U132917 ( n63596, n63052, n63597 );
nand U132918 ( n29689, n29695, n29696 );
nand U132919 ( n29696, n29658, n29697 );
nand U132920 ( n29695, P1_P3_EBX_REG_15_, n29699 );
nand U132921 ( n29697, n29285, n29698 );
nand U132922 ( n22368, n22374, n22375 );
nand U132923 ( n22375, n22337, n22376 );
nand U132924 ( n22374, P1_P2_EBX_REG_15_, n22378 );
nand U132925 ( n22376, n21970, n22377 );
nand U132926 ( n55480, n55486, n55487 );
nand U132927 ( n55487, n55449, n55488 );
nand U132928 ( n55486, P2_P2_EBX_REG_15_, n55490 );
nand U132929 ( n55488, n55080, n55489 );
nand U132930 ( n63751, n63759, n63760 );
nand U132931 ( n63760, n63731, n63761 );
nand U132932 ( n63759, P2_P3_EBX_REG_11_, n63763 );
nand U132933 ( n63761, n63052, n63762 );
nand U132934 ( n63857, n63864, n63865 );
nand U132935 ( n63865, n63827, n63866 );
nand U132936 ( n63864, P2_P3_EBX_REG_7_, n63868 );
nand U132937 ( n63866, n63052, n63867 );
nand U132938 ( n63907, n63914, n63915 );
nand U132939 ( n63915, n63887, n63916 );
nand U132940 ( n63914, P2_P3_EBX_REG_5_, n63918 );
nand U132941 ( n63916, n63052, n63917 );
nand U132942 ( n29791, n29799, n29800 );
nand U132943 ( n29800, n29771, n29801 );
nand U132944 ( n29799, P1_P3_EBX_REG_11_, n29803 );
nand U132945 ( n29801, n29285, n29802 );
nand U132946 ( n29901, n29908, n29909 );
nand U132947 ( n29909, n29871, n29910 );
nand U132948 ( n29908, P1_P3_EBX_REG_7_, n29912 );
nand U132949 ( n29910, n29285, n29911 );
nand U132950 ( n29951, n29958, n29959 );
nand U132951 ( n29959, n29931, n29960 );
nand U132952 ( n29958, P1_P3_EBX_REG_5_, n29962 );
nand U132953 ( n29960, n29285, n29961 );
nand U132954 ( n22578, n22585, n22586 );
nand U132955 ( n22586, n22548, n22587 );
nand U132956 ( n22585, P1_P2_EBX_REG_7_, n22589 );
nand U132957 ( n22587, n21970, n22588 );
nand U132958 ( n22470, n22478, n22479 );
nand U132959 ( n22479, n22450, n22480 );
nand U132960 ( n22478, P1_P2_EBX_REG_11_, n22482 );
nand U132961 ( n22480, n21970, n22481 );
nand U132962 ( n22628, n22635, n22636 );
nand U132963 ( n22636, n22608, n22637 );
nand U132964 ( n22635, P1_P2_EBX_REG_5_, n22639 );
nand U132965 ( n22637, n21970, n22638 );
nand U132966 ( n55691, n55698, n55699 );
nand U132967 ( n55699, n55661, n55700 );
nand U132968 ( n55698, P2_P2_EBX_REG_7_, n55702 );
nand U132969 ( n55700, n55080, n55701 );
nand U132970 ( n55585, n55593, n55594 );
nand U132971 ( n55594, n55565, n55595 );
nand U132972 ( n55593, P2_P2_EBX_REG_11_, n55597 );
nand U132973 ( n55595, n55080, n55596 );
nand U132974 ( n55741, n55748, n55749 );
nand U132975 ( n55749, n55721, n55750 );
nand U132976 ( n55748, P2_P2_EBX_REG_5_, n55752 );
nand U132977 ( n55750, n55080, n55751 );
nand U132978 ( n63485, n63492, n63493 );
nand U132979 ( n63493, n63460, n63494 );
nand U132980 ( n63492, P2_P3_EBX_REG_19_, n63496 );
nand U132981 ( n63494, n63052, n63495 );
nand U132982 ( n63640, n63647, n63648 );
nand U132983 ( n63648, n63616, n63649 );
nand U132984 ( n63647, P2_P3_EBX_REG_13_, n63651 );
nand U132985 ( n63649, n63052, n63650 );
nand U132986 ( n29586, n29593, n29594 );
nand U132987 ( n29594, n29557, n29595 );
nand U132988 ( n29593, P1_P3_EBX_REG_19_, n29597 );
nand U132989 ( n29595, n29285, n29596 );
nand U132990 ( n29741, n29748, n29749 );
nand U132991 ( n29749, n29717, n29750 );
nand U132992 ( n29748, P1_P3_EBX_REG_13_, n29752 );
nand U132993 ( n29750, n29285, n29751 );
nand U132994 ( n22420, n22427, n22428 );
nand U132995 ( n22428, n22396, n22429 );
nand U132996 ( n22427, P1_P2_EBX_REG_13_, n22431 );
nand U132997 ( n22429, n21970, n22430 );
nand U132998 ( n22265, n22272, n22273 );
nand U132999 ( n22273, n22240, n22274 );
nand U133000 ( n22272, P1_P2_EBX_REG_19_, n22276 );
nand U133001 ( n22274, n21970, n22275 );
nand U133002 ( n55535, n55542, n55543 );
nand U133003 ( n55543, n55508, n55544 );
nand U133004 ( n55542, P2_P2_EBX_REG_13_, n55546 );
nand U133005 ( n55544, n55080, n55545 );
nand U133006 ( n55377, n55384, n55385 );
nand U133007 ( n55385, n55352, n55386 );
nand U133008 ( n55384, P2_P2_EBX_REG_19_, n55388 );
nand U133009 ( n55386, n55080, n55387 );
xor U133010 ( n37884, n37885, n37886 );
xor U133011 ( n37886, n37883, P4_REG2_REG_11_ );
nand U133012 ( n45005, n45006, n858 );
xor U133013 ( n45006, n45007, P3_REG2_REG_16_ );
nand U133014 ( n5261, n30067, n30068 );
nor U133015 ( n30067, n30086, n30087 );
nor U133016 ( n30068, n30069, n30070 );
nor U133017 ( n30087, P1_P3_INSTQUEUERD_ADDR_REG_0_, n30061 );
nor U133018 ( n25359, n76519, P1_P2_STATE2_REG_2_ );
nor U133019 ( n58496, n76261, P2_P2_STATE2_REG_2_ );
nand U133020 ( n7506, n22746, n22747 );
nor U133021 ( n22746, n22765, n22766 );
nor U133022 ( n22747, n22748, n22749 );
nor U133023 ( n22766, P1_P2_INSTQUEUERD_ADDR_REG_0_, n22738 );
nand U133024 ( n14241, n55860, n55861 );
nor U133025 ( n55860, n55879, n55880 );
nor U133026 ( n55861, n55862, n55863 );
nor U133027 ( n55880, P2_P2_INSTQUEUERD_ADDR_REG_0_, n55854 );
nand U133028 ( n11996, n64084, n64085 );
nor U133029 ( n64084, n64103, n64104 );
nor U133030 ( n64085, n64086, n64087 );
nor U133031 ( n64104, P2_P3_INSTQUEUERD_ADDR_REG_0_, n64078 );
nor U133032 ( n32599, n76468, P1_P3_STATE2_REG_2_ );
nor U133033 ( n67364, n76195, P2_P3_STATE2_REG_2_ );
nand U133034 ( n4316, n33927, n33928 );
nand U133035 ( n33928, n76468, P1_P3_INSTADDRPOINTER_REG_2_ );
nor U133036 ( n33927, n33929, n33930 );
nor U133037 ( n33929, n33931, n76894 );
nand U133038 ( n11051, n68683, n68684 );
nand U133039 ( n68684, n76195, P2_P3_INSTADDRPOINTER_REG_2_ );
nor U133040 ( n68683, n68685, n68686 );
nor U133041 ( n68685, n68687, n76868 );
nand U133042 ( n6561, n26682, n26683 );
nand U133043 ( n26683, n76519, P1_P2_INSTADDRPOINTER_REG_2_ );
nor U133044 ( n26682, n26684, n26685 );
nor U133045 ( n26684, n26686, n76903 );
nand U133046 ( n13296, n59824, n59825 );
nand U133047 ( n59825, n76261, P2_P2_INSTADDRPOINTER_REG_2_ );
nor U133048 ( n59824, n59826, n59827 );
nor U133049 ( n59826, n59828, n76877 );
nand U133050 ( n4321, n33850, n33851 );
nand U133051 ( n33851, n76468, P1_P3_INSTADDRPOINTER_REG_3_ );
nor U133052 ( n33850, n33852, n33853 );
nor U133053 ( n33852, n33854, n76894 );
nand U133054 ( n11056, n68606, n68607 );
nand U133055 ( n68607, n76195, P2_P3_INSTADDRPOINTER_REG_3_ );
nor U133056 ( n68606, n68608, n68609 );
nor U133057 ( n68608, n68610, n76868 );
nand U133058 ( n6566, n26605, n26606 );
nand U133059 ( n26606, n76519, P1_P2_INSTADDRPOINTER_REG_3_ );
nor U133060 ( n26605, n26607, n26608 );
nor U133061 ( n26607, n26609, n76903 );
nand U133062 ( n13301, n59747, n59748 );
nand U133063 ( n59748, n76261, P2_P2_INSTADDRPOINTER_REG_3_ );
nor U133064 ( n59747, n59749, n59750 );
nor U133065 ( n59749, n59751, n76877 );
nand U133066 ( n4326, n33765, n33766 );
nand U133067 ( n33766, n76468, P1_P3_INSTADDRPOINTER_REG_4_ );
nor U133068 ( n33765, n33767, n33768 );
nor U133069 ( n33767, n33769, n76894 );
nand U133070 ( n6571, n26520, n26521 );
nand U133071 ( n26521, n76519, P1_P2_INSTADDRPOINTER_REG_4_ );
nor U133072 ( n26520, n26522, n26523 );
nor U133073 ( n26522, n26524, n76903 );
nand U133074 ( n13306, n59662, n59663 );
nand U133075 ( n59663, n76261, P2_P2_INSTADDRPOINTER_REG_4_ );
nor U133076 ( n59662, n59664, n59665 );
nor U133077 ( n59664, n59666, n76877 );
nand U133078 ( n4331, n33686, n33687 );
nand U133079 ( n33687, n76468, P1_P3_INSTADDRPOINTER_REG_5_ );
nor U133080 ( n33686, n33688, n33689 );
nor U133081 ( n33688, n33690, n76894 );
nand U133082 ( n11061, n68521, n68522 );
nand U133083 ( n68522, n76195, P2_P3_INSTADDRPOINTER_REG_4_ );
nor U133084 ( n68521, n68523, n68524 );
nor U133085 ( n68523, n68525, n76868 );
nand U133086 ( n11066, n68442, n68443 );
nand U133087 ( n68443, n76195, P2_P3_INSTADDRPOINTER_REG_5_ );
nor U133088 ( n68442, n68444, n68445 );
nor U133089 ( n68444, n68446, n76868 );
nand U133090 ( n6576, n26441, n26442 );
nand U133091 ( n26442, n76519, P1_P2_INSTADDRPOINTER_REG_5_ );
nor U133092 ( n26441, n26443, n26444 );
nor U133093 ( n26443, n26445, n76903 );
nand U133094 ( n13311, n59580, n59581 );
nand U133095 ( n59581, n76261, P2_P2_INSTADDRPOINTER_REG_5_ );
nor U133096 ( n59580, n59582, n59583 );
nor U133097 ( n59582, n59584, n76877 );
nand U133098 ( n4311, n34002, n34003 );
nand U133099 ( n34003, n76468, P1_P3_INSTADDRPOINTER_REG_1_ );
nor U133100 ( n34002, n34004, n34005 );
nor U133101 ( n34004, n34006, n76894 );
nand U133102 ( n6551, n26806, n26807 );
nand U133103 ( n26807, n76519, P1_P2_INSTADDRPOINTER_REG_0_ );
nor U133104 ( n26806, n26808, n26809 );
nor U133105 ( n26808, n75260, n76906 );
nand U133106 ( n13286, n59946, n59947 );
nand U133107 ( n59947, n76261, P2_P2_INSTADDRPOINTER_REG_0_ );
nor U133108 ( n59946, n59948, n59949 );
nor U133109 ( n59948, n75261, n76880 );
nand U133110 ( n4306, n34051, n34052 );
nand U133111 ( n34052, n76468, P1_P3_INSTADDRPOINTER_REG_0_ );
nor U133112 ( n34051, n34053, n34054 );
nor U133113 ( n34053, n75258, n76897 );
nand U133114 ( n11046, n68758, n68759 );
nand U133115 ( n68759, n76195, P2_P3_INSTADDRPOINTER_REG_1_ );
nor U133116 ( n68758, n68760, n68761 );
nor U133117 ( n68760, n68762, n76868 );
nand U133118 ( n6556, n26759, n26760 );
nand U133119 ( n26760, n76519, P1_P2_INSTADDRPOINTER_REG_1_ );
nor U133120 ( n26759, n26761, n26762 );
nor U133121 ( n26761, n26763, n76903 );
nand U133122 ( n13291, n59899, n59900 );
nand U133123 ( n59900, n76261, P2_P2_INSTADDRPOINTER_REG_1_ );
nor U133124 ( n59899, n59901, n59902 );
nor U133125 ( n59901, n59903, n76877 );
nand U133126 ( n4336, n33592, n33593 );
nand U133127 ( n33593, n76468, P1_P3_INSTADDRPOINTER_REG_6_ );
nor U133128 ( n33592, n33594, n33595 );
nor U133129 ( n33594, n33596, n76894 );
nand U133130 ( n11071, n68348, n68349 );
nand U133131 ( n68349, n76195, P2_P3_INSTADDRPOINTER_REG_6_ );
nor U133132 ( n68348, n68350, n68351 );
nor U133133 ( n68350, n68352, n76868 );
nand U133134 ( n6581, n26347, n26348 );
nand U133135 ( n26348, n76519, P1_P2_INSTADDRPOINTER_REG_6_ );
nor U133136 ( n26347, n26349, n26350 );
nor U133137 ( n26349, n26351, n76903 );
nand U133138 ( n13316, n59486, n59487 );
nand U133139 ( n59487, n76261, P2_P2_INSTADDRPOINTER_REG_6_ );
nor U133140 ( n59486, n59488, n59489 );
nor U133141 ( n59488, n59490, n76877 );
nand U133142 ( n11041, n68805, n68806 );
nand U133143 ( n68806, n76195, P2_P3_INSTADDRPOINTER_REG_0_ );
nor U133144 ( n68805, n68807, n68808 );
nor U133145 ( n68807, n75257, n76871 );
nand U133146 ( n35723, n35724, n35725 );
nand U133147 ( n35725, n35726, n35727 );
nand U133148 ( n35724, n35734, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nor U133149 ( n35727, n29143, n35728 );
nand U133150 ( n28544, n28545, n28546 );
nand U133151 ( n28546, n28547, n28548 );
nand U133152 ( n28545, n28555, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nor U133153 ( n28548, n21828, n28549 );
nand U133154 ( n70449, n70450, n70451 );
nand U133155 ( n70451, n70452, n70453 );
nand U133156 ( n70450, n70460, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nor U133157 ( n70453, n62810, n70454 );
nand U133158 ( n61849, n61850, n61851 );
nand U133159 ( n61851, n61852, n61853 );
nand U133160 ( n61850, n61860, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nor U133161 ( n61853, n54904, n61854 );
nand U133162 ( n54221, n54222, n54223 );
nand U133163 ( n54223, n54224, n54225 );
nand U133164 ( n54222, n54232, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nor U133165 ( n54225, n42322, n54226 );
nand U133166 ( n45559, n46283, P2_P1_STATE2_REG_2_ );
nor U133167 ( n46283, P2_P1_STATE2_REG_0_, n7438 );
nand U133168 ( n64065, n64066, n64067 );
nand U133169 ( n64066, n64070, n74469 );
nand U133170 ( n64067, P2_P3_EBX_REG_1_, n64068 );
nand U133171 ( n64070, n63052, n64071 );
nand U133172 ( n30048, n30049, n30050 );
nand U133173 ( n30049, n30053, n74470 );
nand U133174 ( n30050, P1_P3_EBX_REG_1_, n30051 );
nand U133175 ( n30053, n29285, n30054 );
nand U133176 ( n22725, n22726, n22727 );
nand U133177 ( n22726, n22730, n74471 );
nand U133178 ( n22727, P1_P2_EBX_REG_1_, n22728 );
nand U133179 ( n22730, n21970, n22731 );
nand U133180 ( n55841, n55842, n55843 );
nand U133181 ( n55842, n55846, n74472 );
nand U133182 ( n55843, P2_P2_EBX_REG_1_, n55844 );
nand U133183 ( n55846, n55080, n55847 );
nor U133184 ( n10424, n10478, n10479 );
nor U133185 ( n10479, n9908, P1_P1_EAX_REG_19_ );
nor U133186 ( n44263, n44306, n44307 );
nor U133187 ( n44307, n43808, P2_P1_EAX_REG_19_ );
nand U133188 ( n10417, n10418, n10419 );
nand U133189 ( n10419, n10420, n10422 );
nand U133190 ( n10418, P1_P1_EAX_REG_21_, n10423 );
nor U133191 ( n10420, P1_P1_EAX_REG_21_, n74966 );
nand U133192 ( n44257, n44258, n44259 );
nand U133193 ( n44259, n44260, n44261 );
nand U133194 ( n44258, P2_P1_EAX_REG_21_, n44262 );
nor U133195 ( n44260, P2_P1_EAX_REG_21_, n74965 );
nand U133196 ( n31861, n32579, P1_P3_STATE2_REG_2_ );
nor U133197 ( n32579, P1_P3_STATE2_REG_0_, n3063 );
nand U133198 ( n63957, n63958, n63959 );
nand U133199 ( n63959, n63940, n63960 );
nand U133200 ( n63958, P2_P3_EBX_REG_3_, n63962 );
nand U133201 ( n63960, n63052, n63961 );
nand U133202 ( n30001, n30002, n30003 );
nand U133203 ( n30003, n29984, n30004 );
nand U133204 ( n30002, P1_P3_EBX_REG_3_, n30006 );
nand U133205 ( n30004, n29285, n30005 );
nand U133206 ( n22678, n22679, n22680 );
nand U133207 ( n22680, n22661, n22681 );
nand U133208 ( n22679, P1_P2_EBX_REG_3_, n22683 );
nand U133209 ( n22681, n21970, n22682 );
nand U133210 ( n55794, n55795, n55796 );
nand U133211 ( n55796, n55774, n55797 );
nand U133212 ( n55795, P2_P2_EBX_REG_3_, n55799 );
nand U133213 ( n55797, n55080, n55798 );
nand U133214 ( n31836, n31837, P1_P3_PHYADDRPOINTER_REG_30_ );
nor U133215 ( n31837, P1_P3_PHYADDRPOINTER_REG_31_, n3054 );
not U133216 ( n3054, n31838 );
nand U133217 ( n24647, n25337, P1_P2_STATE2_REG_2_ );
nor U133218 ( n25337, P1_P2_STATE2_REG_0_, n3907 );
nand U133219 ( n66484, n67344, P2_P3_STATE2_REG_2_ );
nor U133220 ( n67344, P2_P3_STATE2_REG_0_, n5664 );
nand U133221 ( n57783, n58476, P2_P2_STATE2_REG_2_ );
nor U133222 ( n58476, P2_P2_STATE2_REG_0_, n6539 );
nor U133223 ( n10585, n10638, n10639 );
nor U133224 ( n10639, n9908, P1_P1_EAX_REG_16_ );
nor U133225 ( n10190, n10247, n10248 );
nor U133226 ( n10248, n9908, P1_P1_EAX_REG_22_ );
nor U133227 ( n44406, n44448, n44449 );
nor U133228 ( n44449, n43808, P2_P1_EAX_REG_16_ );
nor U133229 ( n44076, n44121, n44122 );
nor U133230 ( n44122, n43808, P2_P1_EAX_REG_22_ );
nand U133231 ( n10578, n10579, n10580 );
nand U133232 ( n10580, n10582, n10583 );
nand U133233 ( n10579, P1_P1_EAX_REG_18_, n10584 );
nor U133234 ( n10582, P1_P1_EAX_REG_18_, n74909 );
nand U133235 ( n10183, n10184, n10185 );
nand U133236 ( n10185, n10187, n10188 );
nand U133237 ( n10184, P1_P1_EAX_REG_24_, n10189 );
nor U133238 ( n10187, P1_P1_EAX_REG_24_, n75013 );
nand U133239 ( n44400, n44401, n44402 );
nand U133240 ( n44402, n44403, n44404 );
nand U133241 ( n44401, P2_P1_EAX_REG_18_, n44405 );
nor U133242 ( n44403, P2_P1_EAX_REG_18_, n74908 );
nand U133243 ( n44070, n44071, n44072 );
nand U133244 ( n44072, n44073, n44074 );
nand U133245 ( n44071, P2_P1_EAX_REG_24_, n44075 );
nor U133246 ( n44073, P2_P1_EAX_REG_24_, n75012 );
nand U133247 ( n24622, n24623, P1_P2_PHYADDRPOINTER_REG_30_ );
nor U133248 ( n24623, P1_P2_PHYADDRPOINTER_REG_31_, n3898 );
not U133249 ( n3898, n24624 );
nand U133250 ( n57754, n57755, P2_P2_PHYADDRPOINTER_REG_30_ );
nor U133251 ( n57755, P2_P2_PHYADDRPOINTER_REG_31_, n6530 );
not U133252 ( n6530, n57756 );
nand U133253 ( n66459, n66460, P2_P3_PHYADDRPOINTER_REG_30_ );
nor U133254 ( n66460, P2_P3_PHYADDRPOINTER_REG_31_, n5655 );
not U133255 ( n5655, n66461 );
nor U133256 ( n9824, n9909, n9910 );
nor U133257 ( n9910, n9908, P1_P1_EAX_REG_28_ );
nor U133258 ( n10022, n10069, n10070 );
nor U133259 ( n10070, n9908, P1_P1_EAX_REG_25_ );
nor U133260 ( n43741, n43809, n43810 );
nor U133261 ( n43810, n43808, P2_P1_EAX_REG_28_ );
nor U133262 ( n43938, n43983, n43984 );
nor U133263 ( n43984, n43808, P2_P1_EAX_REG_25_ );
nand U133264 ( n9817, n9818, n9819 );
nand U133265 ( n9819, n9820, P1_P1_EAX_REG_29_ );
nand U133266 ( n9818, P1_P1_EAX_REG_30_, n9823 );
nor U133267 ( n9820, P1_P1_EAX_REG_30_, n9822 );
nand U133268 ( n43735, n43736, n43737 );
nand U133269 ( n43737, n43738, P2_P1_EAX_REG_29_ );
nand U133270 ( n43736, P2_P1_EAX_REG_30_, n43740 );
nor U133271 ( n43738, P2_P1_EAX_REG_30_, n43739 );
nand U133272 ( n10016, n10017, n10018 );
nand U133273 ( n10018, n10019, n10020 );
nand U133274 ( n10017, P1_P1_EAX_REG_27_, n10021 );
nor U133275 ( n10019, P1_P1_EAX_REG_27_, n75085 );
nand U133276 ( n43932, n43933, n43934 );
nand U133277 ( n43934, n43935, n43936 );
nand U133278 ( n43933, P2_P1_EAX_REG_27_, n43937 );
nor U133279 ( n43935, P2_P1_EAX_REG_27_, n75084 );
nand U133280 ( n21978, n21979, n21980 );
nand U133281 ( n21979, P1_P2_REIP_REG_30_, n21984 );
nand U133282 ( n21980, P1_P2_EBX_REG_30_, n21981 );
nand U133283 ( n21984, n175, n21985 );
nand U133284 ( n29293, n29294, n29295 );
nand U133285 ( n29294, P1_P3_REIP_REG_30_, n29299 );
nand U133286 ( n29295, P1_P3_EBX_REG_30_, n29296 );
nand U133287 ( n29299, n209, n29300 );
nand U133288 ( n63060, n63061, n63062 );
nand U133289 ( n63061, P2_P3_REIP_REG_30_, n63066 );
nand U133290 ( n63062, P2_P3_EBX_REG_30_, n63063 );
nand U133291 ( n63066, n480, n63067 );
nand U133292 ( n55088, n55089, n55090 );
nand U133293 ( n55089, P2_P2_REIP_REG_30_, n55094 );
nand U133294 ( n55090, P2_P2_EBX_REG_30_, n55091 );
nand U133295 ( n55094, n447, n55095 );
xor U133296 ( n32313, n33235, P1_P3_INSTADDRPOINTER_REG_13_ );
xor U133297 ( n12329, n13508, P1_P1_INSTADDRPOINTER_REG_13_ );
xor U133298 ( n46012, n46955, P2_P1_INSTADDRPOINTER_REG_13_ );
nor U133299 ( n10947, n10948, n74802 );
nor U133300 ( n10948, n10949, n10950 );
nor U133301 ( n10949, P1_P1_EAX_REG_11_, n9908 );
nor U133302 ( n44690, n44691, n74803 );
nor U133303 ( n44691, n44692, n44693 );
nor U133304 ( n44692, P2_P1_EAX_REG_11_, n43808 );
nor U133305 ( n10774, n10775, n74864 );
nor U133306 ( n10775, n10777, n10778 );
nor U133307 ( n10777, P1_P1_EAX_REG_14_, n9908 );
nor U133308 ( n44552, n44553, n74865 );
nor U133309 ( n44553, n44554, n44555 );
nor U133310 ( n44554, P2_P1_EAX_REG_14_, n43808 );
xor U133311 ( n66952, n67990, P2_P3_INSTADDRPOINTER_REG_13_ );
xor U133312 ( n25076, n25987, P1_P2_INSTADDRPOINTER_REG_13_ );
xor U133313 ( n58211, n59125, P2_P2_INSTADDRPOINTER_REG_13_ );
nor U133314 ( n11274, n11275, n74630 );
nor U133315 ( n11275, n11277, n11278 );
nor U133316 ( n11277, P1_P1_EAX_REG_2_, n9908 );
nor U133317 ( n44961, n44962, n74631 );
nor U133318 ( n44962, n44963, n44964 );
nor U133319 ( n44963, P2_P1_EAX_REG_2_, n43808 );
nor U133320 ( n11097, n11098, n74756 );
nor U133321 ( n11098, n11099, n11100 );
nor U133322 ( n11099, P1_P1_EAX_REG_8_, n9908 );
nor U133323 ( n44810, n44811, n74757 );
nor U133324 ( n44811, n44812, n44813 );
nor U133325 ( n44812, P2_P1_EAX_REG_8_, n43808 );
nor U133326 ( n44931, n44932, n74704 );
nor U133327 ( n44932, n44933, n44934 );
nor U133328 ( n44933, P2_P1_EAX_REG_5_, n43808 );
nor U133329 ( n11230, n11232, n74705 );
nor U133330 ( n11232, n11233, n11234 );
nor U133331 ( n11233, P1_P1_EAX_REG_5_, n9908 );
nand U133332 ( n33366, n76475, P1_P3_INSTADDRPOINTER_REG_12_ );
nand U133333 ( n49679, n51657, P3_DATAO_REG_0_ );
and U133334 ( n51657, n76930, DIN_30_ );
or U133335 ( n9902, n75948, n75949 );
nor U133336 ( n75948, n75219, n9824 );
nor U133337 ( n75949, n9822, P1_P1_EAX_REG_29_ );
or U133338 ( n43803, n75950, n75951 );
nor U133339 ( n75950, n75218, n43741 );
nor U133340 ( n75951, n43739, P2_P1_EAX_REG_29_ );
nand U133341 ( n11800, n12668, P1_P1_STATE2_REG_2_ );
nor U133342 ( n12668, P1_P1_STATE2_REG_0_, n4794 );
nand U133343 ( n17076, DIN_27_, n76928 );
nor U133344 ( n30407, P1_P3_EBX_REG_0_, n76489 );
nand U133345 ( n5101, n30403, n30404 );
nand U133346 ( n30404, P1_P3_EBX_REG_0_, n30405 );
nor U133347 ( n30403, n30406, n30407 );
nor U133348 ( n30406, n73987, n30123 );
nor U133349 ( n9803, P1_P1_EBX_REG_0_, n76633 );
nor U133350 ( n23076, P1_P2_EBX_REG_0_, n76542 );
nor U133351 ( n43724, P2_P1_EBX_REG_0_, n76363 );
nor U133352 ( n56197, P2_P2_EBX_REG_0_, n76284 );
nor U133353 ( n64566, P2_P3_EBX_REG_0_, n76222 );
nand U133354 ( n9591, n9798, n9799 );
nand U133355 ( n9799, P1_P1_EBX_REG_0_, n9800 );
nor U133356 ( n9798, n9802, n9803 );
nor U133357 ( n9802, n74005, n9457 );
nand U133358 ( n7346, n23072, n23073 );
nand U133359 ( n23073, P1_P2_EBX_REG_0_, n23074 );
nor U133360 ( n23072, n23075, n23076 );
nor U133361 ( n23075, n73641, n22798 );
nand U133362 ( n16326, n43720, n43721 );
nand U133363 ( n43721, P2_P1_EBX_REG_0_, n43722 );
nor U133364 ( n43720, n43723, n43724 );
nor U133365 ( n43723, n73553, n43392 );
nand U133366 ( n14081, n56193, n56194 );
nand U133367 ( n56194, P2_P2_EBX_REG_0_, n56195 );
nor U133368 ( n56193, n56196, n56197 );
nor U133369 ( n56196, n73642, n55912 );
nand U133370 ( n11836, n64562, n64563 );
nand U133371 ( n64563, P2_P3_EBX_REG_0_, n64564 );
nor U133372 ( n64562, n64565, n64566 );
nor U133373 ( n64565, n73643, n64136 );
nand U133374 ( n456, n63409, n63410 );
nor U133375 ( n63410, n63411, n63412 );
nor U133376 ( n63409, n63414, n63415 );
or U133377 ( n63412, P1_P1_BE_N_REG_0_, P1_P1_BE_N_REG_1_ );
nand U133378 ( n63415, n76611, P1_P1_W_R_N_REG );
buf U133379 ( n76609, n11647 );
nand U133380 ( n11647, P1_P1_ADDRESS_REG_29_, n63416 );
nand U133381 ( n63416, n63417, n63418 );
nor U133382 ( n63418, n63419, n63420 );
nand U133383 ( n276, n38301, n38302 );
nand U133384 ( n38302, P1_P1_DATAO_REG_31_, n76749 );
nor U133385 ( n38301, n38303, n38304 );
nor U133386 ( n38304, n75446, n76434 );
nand U133387 ( n271, n38466, n38467 );
nand U133388 ( n38467, P1_P1_DATAO_REG_30_, n76749 );
nor U133389 ( n38466, n38468, n38469 );
nor U133390 ( n38469, n75413, n76434 );
nor U133391 ( n38654, n75593, n76432 );
nor U133392 ( n38688, n75594, n76432 );
nor U133393 ( n38722, n75595, n76432 );
nor U133394 ( n38620, n75596, n76432 );
nor U133395 ( n39811, n75597, n76432 );
nor U133396 ( n39197, n75598, n76432 );
nand U133397 ( n261, n38652, n38653 );
nand U133398 ( n38653, P1_P1_DATAO_REG_28_, n76749 );
nor U133399 ( n38652, n38654, n38655 );
nor U133400 ( n38655, n75414, n76434 );
nand U133401 ( n256, n38686, n38687 );
nand U133402 ( n38687, P1_P1_DATAO_REG_27_, n76749 );
nor U133403 ( n38686, n38688, n38689 );
nor U133404 ( n38689, n75415, n76434 );
nand U133405 ( n251, n38720, n38721 );
nand U133406 ( n38721, P1_P1_DATAO_REG_26_, n76749 );
nor U133407 ( n38720, n38722, n38723 );
nor U133408 ( n38723, n75391, n76434 );
nand U133409 ( n266, n38618, n38619 );
nand U133410 ( n38619, P1_P1_DATAO_REG_29_, n76749 );
nor U133411 ( n38618, n38620, n38621 );
nor U133412 ( n38621, n75392, n76434 );
nand U133413 ( n241, n39809, n39810 );
nand U133414 ( n39810, P1_P1_DATAO_REG_24_, n76749 );
nor U133415 ( n39809, n39811, n39812 );
nor U133416 ( n39812, n75416, n76434 );
nand U133417 ( n246, n39195, n39196 );
nand U133418 ( n39196, P1_P1_DATAO_REG_25_, n76749 );
nor U133419 ( n39195, n39197, n39198 );
nor U133420 ( n39198, n75393, n76434 );
nor U133421 ( n40245, n75528, n76431 );
nor U133422 ( n41074, n75529, n76431 );
nor U133423 ( n42739, n75530, n76430 );
nor U133424 ( n42178, n75531, n76430 );
nor U133425 ( n40433, n75532, n76431 );
nor U133426 ( n42130, n75533, n76431 );
nor U133427 ( n42154, n75534, n76430 );
nor U133428 ( n45097, n75535, n76430 );
nor U133429 ( n40563, n75536, n76431 );
nor U133430 ( n40499, n75537, n76431 );
nor U133431 ( n40429, n75538, n76431 );
nor U133432 ( n54773, n75539, n76430 );
nor U133433 ( n42105, n75540, n76431 );
nor U133434 ( n60480, n75541, n76430 );
nor U133435 ( n40668, n75542, n76431 );
nor U133436 ( n40425, n75543, n76431 );
nor U133437 ( n57770, n75544, n76430 );
nor U133438 ( n61664, n75545, n76430 );
nor U133439 ( n40622, n75546, n76431 );
nor U133440 ( n40887, n75547, n76431 );
nor U133441 ( n48939, n75548, n76430 );
nor U133442 ( n56168, n75549, n76430 );
nor U133443 ( n63372, n75550, n76430 );
nor U133444 ( n47027, n75551, n76430 );
nand U133445 ( n236, n40243, n40244 );
nand U133446 ( n40244, P1_P1_DATAO_REG_23_, n76749 );
nor U133447 ( n40243, n40245, n40246 );
nor U133448 ( n40246, n75394, n76434 );
nand U133449 ( n191, n41072, n41073 );
nand U133450 ( n41073, P1_P1_DATAO_REG_14_, n76749 );
nor U133451 ( n41072, n41074, n41075 );
nor U133452 ( n41075, n75437, n76435 );
nand U133453 ( n166, n42737, n42738 );
nand U133454 ( n42738, P1_P1_DATAO_REG_9_, n76750 );
nor U133455 ( n42737, n42739, n42740 );
nor U133456 ( n42740, n75438, n76435 );
nand U133457 ( n171, n42176, n42177 );
nand U133458 ( n42177, P1_P1_DATAO_REG_10_, n76750 );
nor U133459 ( n42176, n42178, n42179 );
nor U133460 ( n42179, n75439, n76435 );
nand U133461 ( n221, n40431, n40432 );
nand U133462 ( n40432, P1_P1_DATAO_REG_20_, n76749 );
nor U133463 ( n40431, n40433, n40434 );
nor U133464 ( n40434, n75395, n76434 );
nand U133465 ( n181, n42128, n42129 );
nand U133466 ( n42129, P1_P1_DATAO_REG_12_, n76750 );
nor U133467 ( n42128, n42130, n42131 );
nor U133468 ( n42131, n75440, n76435 );
nand U133469 ( n176, n42152, n42153 );
nand U133470 ( n42153, P1_P1_DATAO_REG_11_, n76750 );
nor U133471 ( n42152, n42154, n42155 );
nor U133472 ( n42155, n75441, n76435 );
nand U133473 ( n161, n45095, n45096 );
nand U133474 ( n45096, P1_P1_DATAO_REG_8_, n76750 );
nor U133475 ( n45095, n45097, n45098 );
nor U133476 ( n45098, n75442, n76435 );
nand U133477 ( n211, n40561, n40562 );
nand U133478 ( n40562, P1_P1_DATAO_REG_18_, n76749 );
nor U133479 ( n40561, n40563, n40564 );
nor U133480 ( n40564, n75396, n76435 );
nand U133481 ( n216, n40497, n40498 );
nand U133482 ( n40498, P1_P1_DATAO_REG_19_, n76749 );
nor U133483 ( n40497, n40499, n40500 );
nor U133484 ( n40500, n75397, n76435 );
nand U133485 ( n226, n40427, n40428 );
nand U133486 ( n40428, P1_P1_DATAO_REG_21_, n76749 );
nor U133487 ( n40427, n40429, n40430 );
nor U133488 ( n40430, n75398, n76434 );
nand U133489 ( n146, n54771, n54772 );
nand U133490 ( n54772, P1_P1_DATAO_REG_5_, n76750 );
nor U133491 ( n54771, n54773, n54774 );
nor U133492 ( n54774, n75456, n76436 );
nand U133493 ( n186, n42103, n42104 );
nand U133494 ( n42104, P1_P1_DATAO_REG_13_, n76749 );
nor U133495 ( n42103, n42105, n42106 );
nor U133496 ( n42106, n75443, n76435 );
nand U133497 ( n131, n60478, n60479 );
nand U133498 ( n60479, P1_P1_DATAO_REG_2_, n76750 );
nor U133499 ( n60478, n60480, n60481 );
nor U133500 ( n60481, n75457, n76436 );
nand U133501 ( n201, n40666, n40667 );
nand U133502 ( n40667, P1_P1_DATAO_REG_16_, n76749 );
nor U133503 ( n40666, n40668, n40669 );
nor U133504 ( n40669, n75399, n76435 );
nand U133505 ( n231, n40423, n40424 );
nand U133506 ( n40424, P1_P1_DATAO_REG_22_, n76749 );
nor U133507 ( n40423, n40425, n40426 );
nor U133508 ( n40426, n75400, n76434 );
nand U133509 ( n136, n57768, n57769 );
nand U133510 ( n57769, P1_P1_DATAO_REG_3_, n76750 );
nor U133511 ( n57768, n57770, n57771 );
nor U133512 ( n57771, n75458, n76436 );
nand U133513 ( n126, n61662, n61663 );
nand U133514 ( n61663, P1_P1_DATAO_REG_1_, n76750 );
nor U133515 ( n61662, n61664, n61665 );
nor U133516 ( n61665, n75459, n76436 );
nand U133517 ( n206, n40620, n40621 );
nand U133518 ( n40621, P1_P1_DATAO_REG_17_, n76749 );
nor U133519 ( n40620, n40622, n40623 );
nor U133520 ( n40623, n75401, n76435 );
nand U133521 ( n196, n40885, n40886 );
nand U133522 ( n40886, P1_P1_DATAO_REG_15_, n76749 );
nor U133523 ( n40885, n40887, n40888 );
nor U133524 ( n40888, n75444, n76435 );
nand U133525 ( n151, n48937, n48938 );
nand U133526 ( n48938, P1_P1_DATAO_REG_6_, n76750 );
nor U133527 ( n48937, n48939, n48940 );
nor U133528 ( n48940, n75460, n76436 );
nand U133529 ( n141, n56166, n56167 );
nand U133530 ( n56167, P1_P1_DATAO_REG_4_, n76750 );
nor U133531 ( n56166, n56168, n56169 );
nor U133532 ( n56169, n75461, n76436 );
nand U133533 ( n121, n63370, n63371 );
nand U133534 ( n63371, P1_P1_DATAO_REG_0_, n76750 );
nor U133535 ( n63370, n63372, n63373 );
nor U133536 ( n63373, n75462, n76436 );
nand U133537 ( n156, n47025, n47026 );
nand U133538 ( n47026, P1_P1_DATAO_REG_7_, n76750 );
nor U133539 ( n47025, n47027, n47028 );
nor U133540 ( n47028, n75463, n76436 );
nor U133541 ( n35749, n35753, n73524 );
nor U133542 ( n35753, n35754, n35755 );
nor U133543 ( n35754, n30782, n35713 );
nor U133544 ( n35755, P1_P3_INSTQUEUERD_ADDR_REG_0_, n34061 );
nor U133545 ( n28570, n28574, n73503 );
nor U133546 ( n28574, n28575, n28576 );
nor U133547 ( n28575, n23475, n28534 );
nor U133548 ( n28576, P1_P2_INSTQUEUERD_ADDR_REG_0_, n26816 );
nor U133549 ( n70475, n70479, n73502 );
nor U133550 ( n70479, n70480, n70481 );
nor U133551 ( n70480, n64984, n70439 );
nor U133552 ( n70481, P2_P3_INSTQUEUERD_ADDR_REG_0_, n68815 );
nor U133553 ( n61875, n61879, n73504 );
nor U133554 ( n61879, n61880, n61881 );
nor U133555 ( n61880, n56597, n61839 );
nor U133556 ( n61881, P2_P2_INSTQUEUERD_ADDR_REG_0_, n59956 );
nand U133557 ( n32343, n74458, n33386 );
nand U133558 ( n33386, n33387, P1_P3_INSTADDRPOINTER_REG_11_ );
nor U133559 ( n54247, n54251, n73497 );
nor U133560 ( n54251, n54252, n54253 );
nor U133561 ( n54252, n44142, n54211 );
nor U133562 ( n54253, P2_P1_INSTQUEUERD_ADDR_REG_0_, n47795 );
nand U133563 ( n21332, n21603, n21604 );
nand U133564 ( n21603, n21606, n74646 );
nand U133565 ( n21604, P1_P1_INSTQUEUEWR_ADDR_REG_4_, n21605 );
nand U133566 ( n21605, P1_P1_INSTQUEUERD_ADDR_REG_4_, n5140 );
nor U133567 ( n63434, P1_P1_ADDRESS_REG_0_, n63438 );
nand U133568 ( n63438, n73451, n73030 );
nor U133569 ( n21222, n10763, n21240 );
nand U133570 ( n21240, P1_P1_INSTQUEUERD_ADDR_REG_1_, n21208 );
nand U133571 ( n12367, n74476, n13699 );
nand U133572 ( n13699, n13700, P1_P1_INSTADDRPOINTER_REG_11_ );
nand U133573 ( n21183, n21218, n21219 );
nand U133574 ( n21219, n223, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U133575 ( n21218, n14799, n21202 );
nand U133576 ( n46042, n74427, n47107 );
nand U133577 ( n47107, n47108, P2_P1_INSTADDRPOINTER_REG_11_ );
nand U133578 ( n66982, n74438, n68138 );
nand U133579 ( n68138, n68139, P2_P3_INSTADDRPOINTER_REG_11_ );
nand U133580 ( n25106, n74439, n26135 );
nand U133581 ( n26135, n26136, P1_P2_INSTADDRPOINTER_REG_11_ );
nand U133582 ( n58244, n74440, n59276 );
nand U133583 ( n59276, n59277, P2_P2_INSTADDRPOINTER_REG_11_ );
and U133584 ( n16658, n17401, DIN_29_ );
nand U133585 ( n45535, n45536, P2_P1_PHYADDRPOINTER_REG_30_ );
and U133586 ( n45536, n74967, n45537 );
nand U133587 ( n63923, n63924, n63925 );
nand U133588 ( n63924, P2_P3_REIP_REG_4_, n63931 );
nand U133589 ( n63925, n63926, n76875 );
nand U133590 ( n63931, n63932, n63933 );
nand U133591 ( n64042, n64043, n64044 );
nand U133592 ( n64043, P2_P3_REIP_REG_2_, n63976 );
nand U133593 ( n64044, n64045, n76875 );
nor U133594 ( n64045, n6338, n64046 );
nand U133595 ( n29967, n29968, n29969 );
nand U133596 ( n29968, P1_P3_REIP_REG_4_, n29975 );
nand U133597 ( n29969, n29970, n76901 );
nand U133598 ( n29975, n29976, n29977 );
nand U133599 ( n30025, n30026, n30027 );
nand U133600 ( n30026, P1_P3_REIP_REG_2_, n30020 );
nand U133601 ( n30027, n30028, n76901 );
nor U133602 ( n30028, n3704, n30029 );
nand U133603 ( n22644, n22645, n22646 );
nand U133604 ( n22645, P1_P2_REIP_REG_4_, n22652 );
nand U133605 ( n22646, n22647, n76910 );
nand U133606 ( n22652, n22653, n22654 );
nand U133607 ( n22702, n22703, n22704 );
nand U133608 ( n22703, P1_P2_REIP_REG_2_, n22697 );
nand U133609 ( n22704, n22705, n76910 );
nor U133610 ( n22705, n4598, n22706 );
nand U133611 ( n55757, n55758, n55759 );
nand U133612 ( n55758, P2_P2_REIP_REG_4_, n55765 );
nand U133613 ( n55759, n55760, n76884 );
nand U133614 ( n55765, n55766, n55767 );
nand U133615 ( n55818, n55819, n55820 );
nand U133616 ( n55819, P2_P2_REIP_REG_2_, n55813 );
nand U133617 ( n55820, n55821, n76884 );
nor U133618 ( n55821, n7230, n55822 );
nand U133619 ( n63501, n63502, n63503 );
nand U133620 ( n63502, n63509, n63484 );
nand U133621 ( n63503, n63504, n76874 );
nor U133622 ( n63509, P2_P3_REIP_REG_18_, n74884 );
nand U133623 ( n29602, n29603, n29604 );
nand U133624 ( n29603, n29610, n29585 );
nand U133625 ( n29604, n29605, n76900 );
nor U133626 ( n29610, P1_P3_REIP_REG_18_, n74885 );
nand U133627 ( n22281, n22282, n22283 );
nand U133628 ( n22282, n22289, n22264 );
nand U133629 ( n22283, n22284, n76909 );
nor U133630 ( n22289, P1_P2_REIP_REG_18_, n74883 );
nand U133631 ( n55393, n55394, n55395 );
nand U133632 ( n55394, n55401, n55376 );
nand U133633 ( n55395, n55396, n76883 );
nor U133634 ( n55401, P2_P2_REIP_REG_18_, n74882 );
nor U133635 ( n30120, n76490, n30124 );
or U133636 ( n30124, n30112, P1_P3_EBX_REG_30_ );
nand U133637 ( n63322, n63323, n63324 );
nand U133638 ( n63323, P2_P3_REIP_REG_22_, n63330 );
nand U133639 ( n63324, n63325, n76874 );
nand U133640 ( n63330, n63331, n63332 );
nand U133641 ( n29493, n29494, n29495 );
nand U133642 ( n29494, P1_P3_REIP_REG_22_, n29501 );
nand U133643 ( n29495, n29496, n76900 );
nand U133644 ( n29501, n29502, n29503 );
nand U133645 ( n22174, n22175, n22176 );
nand U133646 ( n22175, P1_P2_REIP_REG_22_, n22182 );
nand U133647 ( n22176, n22177, n76909 );
nand U133648 ( n22182, n22183, n22184 );
nand U133649 ( n22021, n22022, n22023 );
nand U133650 ( n22022, P1_P2_REIP_REG_28_, n22029 );
nand U133651 ( n22023, n22024, n76909 );
nand U133652 ( n22029, n22030, n22031 );
nand U133653 ( n55288, n55289, n55290 );
nand U133654 ( n55289, P2_P2_REIP_REG_22_, n55296 );
nand U133655 ( n55290, n55291, n76883 );
nand U133656 ( n55296, n55297, n55298 );
nand U133657 ( n29340, n29341, n29342 );
nand U133658 ( n29341, P1_P3_REIP_REG_28_, n29348 );
nand U133659 ( n29342, n29343, n76900 );
nand U133660 ( n29348, n29349, n29350 );
nand U133661 ( n63103, n63104, n63105 );
nand U133662 ( n63104, P2_P3_REIP_REG_28_, n63111 );
nand U133663 ( n63105, n63106, n76874 );
nand U133664 ( n63111, n63112, n63113 );
nand U133665 ( n55131, n55132, n55133 );
nand U133666 ( n55132, P2_P2_REIP_REG_28_, n55139 );
nand U133667 ( n55133, n55134, n76883 );
nand U133668 ( n55139, n55140, n55141 );
nand U133669 ( n5251, n30117, n30118 );
nand U133670 ( n30118, P1_P3_EBX_REG_30_, n30116 );
nor U133671 ( n30117, n30120, n30121 );
nor U133672 ( n30121, n30122, n30123 );
nand U133673 ( n5206, n30205, n30206 );
nand U133674 ( n30206, n3072, n30207 );
nor U133675 ( n30205, n30208, n30209 );
and U133676 ( n30209, n30198, P1_P3_EBX_REG_21_ );
nand U133677 ( n5186, n30243, n30244 );
nand U133678 ( n30244, n3072, n30245 );
nor U133679 ( n30243, n30246, n30247 );
and U133680 ( n30247, n30240, P1_P3_EBX_REG_17_ );
nand U133681 ( n5176, n30262, n30263 );
nand U133682 ( n30263, n3072, n30264 );
nor U133683 ( n30262, n30265, n30266 );
and U133684 ( n30266, n30259, P1_P3_EBX_REG_15_ );
nor U133685 ( n30148, n76489, n30151 );
or U133686 ( n30151, n30144, P1_P3_EBX_REG_27_ );
nand U133687 ( n5196, n30224, n30225 );
nand U133688 ( n30225, n3072, n30226 );
nor U133689 ( n30224, n30227, n30228 );
and U133690 ( n30228, n30221, P1_P3_EBX_REG_19_ );
nand U133691 ( n5166, n30281, n30282 );
nand U133692 ( n30282, n3072, n30283 );
nor U133693 ( n30281, n30284, n30285 );
and U133694 ( n30285, n30278, P1_P3_EBX_REG_13_ );
nand U133695 ( n5156, n30304, n30305 );
nand U133696 ( n30305, n3072, n30306 );
nor U133697 ( n30304, n30307, n30308 );
and U133698 ( n30308, n30297, P1_P3_EBX_REG_11_ );
nand U133699 ( n5146, n30323, n30324 );
nand U133700 ( n30324, n3072, n30325 );
nor U133701 ( n30323, n30326, n30327 );
and U133702 ( n30327, n30320, P1_P3_EBX_REG_9_ );
nand U133703 ( n5136, n30342, n30343 );
nand U133704 ( n30343, n3072, P1_P3_INSTQUEUE_REG_0__7_ );
nor U133705 ( n30342, n30344, n30345 );
and U133706 ( n30345, n30339, P1_P3_EBX_REG_7_ );
nand U133707 ( n5126, n30359, n30360 );
nand U133708 ( n30360, n3072, P1_P3_INSTQUEUE_REG_0__5_ );
nor U133709 ( n30359, n30361, n30362 );
and U133710 ( n30362, n30356, P1_P3_EBX_REG_5_ );
nand U133711 ( n5116, n30376, n30377 );
nand U133712 ( n30377, n3072, P1_P3_INSTQUEUE_REG_0__3_ );
nor U133713 ( n30376, n30378, n30379 );
and U133714 ( n30379, n30373, P1_P3_EBX_REG_3_ );
nand U133715 ( n63797, n63804, n63481 );
nand U133716 ( n63804, n63805, n76875 );
nor U133717 ( n63805, P2_P3_EBX_REG_9_, n6334 );
nand U133718 ( n29841, n29848, n29582 );
nand U133719 ( n29848, n29849, n76901 );
nor U133720 ( n29849, P1_P3_EBX_REG_9_, n3700 );
nand U133721 ( n22518, n22525, n22261 );
nand U133722 ( n22525, n22526, n76910 );
nor U133723 ( n22526, P1_P2_EBX_REG_9_, n4594 );
nand U133724 ( n55631, n55638, n55373 );
nand U133725 ( n55638, n55639, n76884 );
nor U133726 ( n55639, P2_P2_EBX_REG_9_, n7227 );
nor U133727 ( n43389, n76364, n43393 );
or U133728 ( n43393, n43381, P2_P1_EBX_REG_30_ );
nor U133729 ( n64133, n76223, n64137 );
or U133730 ( n64137, n64125, P2_P3_EBX_REG_30_ );
nor U133731 ( n22795, n76543, n22799 );
or U133732 ( n22799, n22787, P1_P2_EBX_REG_30_ );
nor U133733 ( n55909, n76285, n55913 );
or U133734 ( n55913, n55901, P2_P2_EBX_REG_30_ );
nand U133735 ( n16476, n43386, n43387 );
nand U133736 ( n43387, P2_P1_EBX_REG_30_, n43385 );
nor U133737 ( n43386, n43389, n43390 );
nor U133738 ( n43390, n43391, n43392 );
nand U133739 ( n11986, n64130, n64131 );
nand U133740 ( n64131, P2_P3_EBX_REG_30_, n64129 );
nor U133741 ( n64130, n64133, n64134 );
nor U133742 ( n64134, n64135, n64136 );
nand U133743 ( n16431, n43503, n43504 );
nand U133744 ( n43504, n7458, n43505 );
nor U133745 ( n43503, n43506, n43507 );
and U133746 ( n43507, n43500, P2_P1_EBX_REG_21_ );
nand U133747 ( n16411, n43541, n43542 );
nand U133748 ( n43542, n7458, n43543 );
nor U133749 ( n43541, n43544, n43545 );
and U133750 ( n43545, n43538, P2_P1_EBX_REG_17_ );
nand U133751 ( n16401, n43573, n43574 );
nand U133752 ( n43574, n7458, n43575 );
nor U133753 ( n43573, n43576, n43577 );
and U133754 ( n43577, n43570, P2_P1_EBX_REG_15_ );
nand U133755 ( n11941, n64267, n64268 );
nand U133756 ( n64268, n5673, n64269 );
nor U133757 ( n64267, n64270, n64271 );
and U133758 ( n64271, n64264, P2_P3_EBX_REG_21_ );
nand U133759 ( n11921, n64305, n64306 );
nand U133760 ( n64306, n5673, n64307 );
nor U133761 ( n64305, n64308, n64309 );
and U133762 ( n64309, n64302, P2_P3_EBX_REG_17_ );
nand U133763 ( n11911, n64324, n64325 );
nand U133764 ( n64325, n5673, n64326 );
nor U133765 ( n64324, n64327, n64328 );
and U133766 ( n64328, n64321, P2_P3_EBX_REG_15_ );
nand U133767 ( n9696, n9554, n9555 );
nand U133768 ( n9555, n4814, n9557 );
nor U133769 ( n9554, n9558, n9559 );
and U133770 ( n9559, n9550, P1_P1_EBX_REG_21_ );
nand U133771 ( n9676, n9600, n9602 );
nand U133772 ( n9602, n4814, n9603 );
nor U133773 ( n9600, n9604, n9605 );
and U133774 ( n9605, n9597, P1_P1_EBX_REG_17_ );
nand U133775 ( n9666, n9624, n9625 );
nand U133776 ( n9625, n4814, n9627 );
nor U133777 ( n9624, n9628, n9629 );
and U133778 ( n9629, n9620, P1_P1_EBX_REG_15_ );
nand U133779 ( n14231, n55906, n55907 );
nand U133780 ( n55907, P2_P2_EBX_REG_30_, n55905 );
nor U133781 ( n55906, n55909, n55910 );
nor U133782 ( n55910, n55911, n55912 );
nand U133783 ( n5216, n30182, n30183 );
or U133784 ( n30183, n30123, n30184 );
nor U133785 ( n30182, n30185, n30186 );
and U133786 ( n30186, n30179, P1_P3_EBX_REG_23_ );
nand U133787 ( n5226, n30163, n30164 );
or U133788 ( n30164, n30165, n30123 );
nor U133789 ( n30163, n30166, n30167 );
and U133790 ( n30167, n30160, P1_P3_EBX_REG_25_ );
nor U133791 ( n30399, n76490, n30402 );
or U133792 ( n30402, n73119, P1_P3_EBX_REG_1_ );
nor U133793 ( n9453, n76634, n9458 );
or U133794 ( n9458, n9443, P1_P1_EBX_REG_30_ );
nand U133795 ( n5106, n30397, n30398 );
nand U133796 ( n30398, n3072, P1_P3_INSTQUEUE_REG_0__1_ );
nor U133797 ( n30397, n30399, n30400 );
and U133798 ( n30400, n30390, P1_P3_EBX_REG_1_ );
nor U133799 ( n43417, n76363, n43420 );
or U133800 ( n43420, n43413, P2_P1_EBX_REG_27_ );
nor U133801 ( n64161, n76222, n64164 );
or U133802 ( n64164, n64157, P2_P3_EBX_REG_27_ );
nor U133803 ( n22823, n76542, n22826 );
or U133804 ( n22826, n22819, P1_P2_EBX_REG_27_ );
nand U133805 ( n9741, n9449, n9450 );
nand U133806 ( n9450, P1_P1_EBX_REG_30_, n9448 );
nor U133807 ( n9449, n9453, n9454 );
nor U133808 ( n9454, n9455, n9457 );
nand U133809 ( n7496, n22792, n22793 );
nand U133810 ( n22793, P1_P2_EBX_REG_30_, n22791 );
nor U133811 ( n22792, n22795, n22796 );
nor U133812 ( n22796, n22797, n22798 );
nand U133813 ( n16421, n43522, n43523 );
nand U133814 ( n43523, n7458, n43524 );
nor U133815 ( n43522, n43525, n43526 );
and U133816 ( n43526, n43519, P2_P1_EBX_REG_19_ );
nand U133817 ( n11931, n64286, n64287 );
nand U133818 ( n64287, n5673, n64288 );
nor U133819 ( n64286, n64289, n64290 );
and U133820 ( n64290, n64283, P2_P3_EBX_REG_19_ );
nand U133821 ( n11901, n64404, n64405 );
nand U133822 ( n64405, n5673, n64406 );
nor U133823 ( n64404, n64407, n64408 );
and U133824 ( n64408, n64401, P2_P3_EBX_REG_13_ );
nand U133825 ( n11891, n64423, n64424 );
nand U133826 ( n64424, n5673, n64425 );
nor U133827 ( n64423, n64426, n64427 );
and U133828 ( n64427, n64420, P2_P3_EBX_REG_11_ );
nand U133829 ( n9636, n9699, n9700 );
nand U133830 ( n9700, n4814, n9702 );
nor U133831 ( n9699, n9703, n9704 );
and U133832 ( n9704, n9695, P1_P1_EBX_REG_9_ );
nand U133833 ( n11881, n64442, n64443 );
nand U133834 ( n64443, n5673, n64444 );
nor U133835 ( n64442, n64445, n64446 );
and U133836 ( n64446, n64439, P2_P3_EBX_REG_9_ );
nand U133837 ( n11871, n64461, n64462 );
nand U133838 ( n64462, n5673, P2_P3_INSTQUEUE_REG_0__7_ );
nor U133839 ( n64461, n64463, n64464 );
and U133840 ( n64464, n64458, P2_P3_EBX_REG_7_ );
nand U133841 ( n11861, n64478, n64479 );
nand U133842 ( n64479, n5673, P2_P3_INSTQUEUE_REG_0__5_ );
nor U133843 ( n64478, n64480, n64481 );
and U133844 ( n64481, n64475, P2_P3_EBX_REG_5_ );
nand U133845 ( n11851, n64539, n64540 );
nand U133846 ( n64540, n5673, P2_P3_INSTQUEUE_REG_0__3_ );
nor U133847 ( n64539, n64541, n64542 );
and U133848 ( n64542, n64536, P2_P3_EBX_REG_3_ );
nand U133849 ( n16391, n43592, n43593 );
nand U133850 ( n43593, n7458, n43594 );
nor U133851 ( n43592, n43595, n43596 );
and U133852 ( n43596, n43589, P2_P1_EBX_REG_13_ );
nand U133853 ( n16381, n43611, n43612 );
nand U133854 ( n43612, n7458, n43613 );
nor U133855 ( n43611, n43614, n43615 );
and U133856 ( n43615, n43608, P2_P1_EBX_REG_11_ );
nand U133857 ( n16371, n43630, n43631 );
nand U133858 ( n43631, n7458, n43632 );
nor U133859 ( n43630, n43633, n43634 );
and U133860 ( n43634, n43627, P2_P1_EBX_REG_9_ );
nand U133861 ( n16361, n43649, n43650 );
nand U133862 ( n43650, n7458, P2_P1_INSTQUEUE_REG_0__7_ );
nor U133863 ( n43649, n43651, n43652 );
and U133864 ( n43652, n43646, P2_P1_EBX_REG_7_ );
nand U133865 ( n16351, n43680, n43681 );
nand U133866 ( n43681, n7458, P2_P1_INSTQUEUE_REG_0__5_ );
nor U133867 ( n43680, n43682, n43683 );
and U133868 ( n43683, n43677, P2_P1_EBX_REG_5_ );
nand U133869 ( n16341, n43697, n43698 );
nand U133870 ( n43698, n7458, P2_P1_INSTQUEUE_REG_0__3_ );
nor U133871 ( n43697, n43699, n43700 );
and U133872 ( n43700, n43694, P2_P1_EBX_REG_3_ );
nor U133873 ( n9488, n76633, n9492 );
or U133874 ( n9492, n9483, P1_P1_EBX_REG_27_ );
nor U133875 ( n55937, n76284, n55940 );
or U133876 ( n55940, n55933, P2_P2_EBX_REG_27_ );
nand U133877 ( n7451, n22878, n22879 );
nand U133878 ( n22879, n76756, n22880 );
nor U133879 ( n22878, n22881, n22882 );
and U133880 ( n22882, n22875, P1_P2_EBX_REG_21_ );
nand U133881 ( n7431, n22916, n22917 );
nand U133882 ( n22917, n76756, n22918 );
nor U133883 ( n22916, n22919, n22920 );
and U133884 ( n22920, n22913, P1_P2_EBX_REG_17_ );
nand U133885 ( n7421, n22935, n22936 );
nand U133886 ( n22936, n76756, n22937 );
nor U133887 ( n22935, n22938, n22939 );
and U133888 ( n22939, n22932, P1_P2_EBX_REG_15_ );
nand U133889 ( n14186, n55993, n55994 );
nand U133890 ( n55994, n76689, n55995 );
nor U133891 ( n55993, n55996, n55997 );
and U133892 ( n55997, n55990, P2_P2_EBX_REG_21_ );
nand U133893 ( n14166, n56031, n56032 );
nand U133894 ( n56032, n76689, n56033 );
nor U133895 ( n56031, n56034, n56035 );
and U133896 ( n56035, n56028, P2_P2_EBX_REG_17_ );
nand U133897 ( n14156, n56053, n56054 );
nand U133898 ( n56054, n76689, n56055 );
nor U133899 ( n56053, n56056, n56057 );
and U133900 ( n56057, n56047, P2_P2_EBX_REG_15_ );
nand U133901 ( n9686, n9578, n9579 );
nand U133902 ( n9579, n4814, n9580 );
nor U133903 ( n9578, n9582, n9583 );
and U133904 ( n9583, n9574, P1_P1_EBX_REG_19_ );
nand U133905 ( n9656, n9652, n9653 );
nand U133906 ( n9653, n4814, n9654 );
nor U133907 ( n9652, n9655, n9657 );
and U133908 ( n9657, n9644, P1_P1_EBX_REG_13_ );
nand U133909 ( n9646, n9675, n9677 );
nand U133910 ( n9677, n4814, n9678 );
nor U133911 ( n9675, n9679, n9680 );
and U133912 ( n9680, n9672, P1_P1_EBX_REG_11_ );
nand U133913 ( n9626, n9723, n9724 );
nand U133914 ( n9724, n4814, P1_P1_INSTQUEUE_REG_0__7_ );
nor U133915 ( n9723, n9725, n9727 );
and U133916 ( n9727, n9719, P1_P1_EBX_REG_7_ );
nand U133917 ( n9616, n9744, n9745 );
nand U133918 ( n9745, n4814, P1_P1_INSTQUEUE_REG_0__5_ );
nor U133919 ( n9744, n9747, n9748 );
and U133920 ( n9748, n9740, P1_P1_EBX_REG_5_ );
nand U133921 ( n9606, n9769, n9770 );
nand U133922 ( n9770, n4814, P1_P1_INSTQUEUE_REG_0__3_ );
nor U133923 ( n9769, n9772, n9773 );
and U133924 ( n9773, n9762, P1_P1_EBX_REG_3_ );
nand U133925 ( n7471, n22838, n22839 );
nand U133926 ( n22839, n22840, n76756 );
nor U133927 ( n22838, n22841, n22842 );
and U133928 ( n22842, n22835, P1_P2_EBX_REG_25_ );
nand U133929 ( n14206, n55955, n55956 );
nand U133930 ( n55956, n55957, n76689 );
nor U133931 ( n55955, n55958, n55959 );
and U133932 ( n55959, n55949, P2_P2_EBX_REG_25_ );
nand U133933 ( n7461, n22857, n22858 );
nand U133934 ( n22858, n76756, n22859 );
nor U133935 ( n22857, n22860, n22861 );
and U133936 ( n22861, n22854, P1_P2_EBX_REG_23_ );
nand U133937 ( n14196, n55974, n55975 );
nand U133938 ( n55975, n76689, n55976 );
nor U133939 ( n55974, n55977, n55978 );
and U133940 ( n55978, n55971, P2_P2_EBX_REG_23_ );
nand U133941 ( n7381, n23013, n23014 );
nand U133942 ( n23014, n76757, P1_P2_INSTQUEUE_REG_0__7_ );
nor U133943 ( n23013, n23015, n23016 );
and U133944 ( n23016, n23010, P1_P2_EBX_REG_7_ );
nand U133945 ( n7371, n23030, n23031 );
nand U133946 ( n23031, n76757, P1_P2_INSTQUEUE_REG_0__5_ );
nor U133947 ( n23030, n23032, n23033 );
and U133948 ( n23033, n23027, P1_P2_EBX_REG_5_ );
nand U133949 ( n7361, n23047, n23048 );
nand U133950 ( n23048, n76757, P1_P2_INSTQUEUE_REG_0__3_ );
nor U133951 ( n23047, n23049, n23050 );
and U133952 ( n23050, n23044, P1_P2_EBX_REG_3_ );
nand U133953 ( n14116, n56129, n56130 );
nand U133954 ( n56130, n76690, P2_P2_INSTQUEUE_REG_0__7_ );
nor U133955 ( n56129, n56131, n56132 );
and U133956 ( n56132, n56126, P2_P2_EBX_REG_7_ );
nand U133957 ( n14106, n56149, n56150 );
nand U133958 ( n56150, n76690, P2_P2_INSTQUEUE_REG_0__5_ );
nor U133959 ( n56149, n56151, n56152 );
and U133960 ( n56152, n56143, P2_P2_EBX_REG_5_ );
nand U133961 ( n14096, n56170, n56171 );
nand U133962 ( n56171, n76690, P2_P2_INSTQUEUE_REG_0__3_ );
nor U133963 ( n56170, n56172, n56173 );
and U133964 ( n56173, n56163, P2_P2_EBX_REG_3_ );
nand U133965 ( n16441, n43484, n43485 );
or U133966 ( n43485, n43392, n43486 );
nor U133967 ( n43484, n43487, n43488 );
and U133968 ( n43488, n43481, P2_P1_EBX_REG_23_ );
nand U133969 ( n11951, n64248, n64249 );
or U133970 ( n64249, n64136, n64250 );
nor U133971 ( n64248, n64251, n64252 );
and U133972 ( n64252, n64245, P2_P3_EBX_REG_23_ );
nand U133973 ( n9706, n9530, n9532 );
or U133974 ( n9532, n9457, n9533 );
nor U133975 ( n9530, n9534, n9535 );
and U133976 ( n9535, n9527, P1_P1_EBX_REG_23_ );
nand U133977 ( n16451, n43465, n43466 );
or U133978 ( n43466, n43467, n43392 );
nor U133979 ( n43465, n43468, n43469 );
and U133980 ( n43469, n43462, P2_P1_EBX_REG_25_ );
nand U133981 ( n11961, n64176, n64177 );
or U133982 ( n64177, n64178, n64136 );
nor U133983 ( n64176, n64179, n64180 );
and U133984 ( n64180, n64173, P2_P3_EBX_REG_25_ );
nand U133985 ( n9716, n9507, n9508 );
or U133986 ( n9508, n9509, n9457 );
nor U133987 ( n9507, n9510, n9512 );
and U133988 ( n9512, n9503, P1_P1_EBX_REG_25_ );
nand U133989 ( n7441, n22897, n22898 );
nand U133990 ( n22898, n76756, n22899 );
nor U133991 ( n22897, n22900, n22901 );
and U133992 ( n22901, n22894, P1_P2_EBX_REG_19_ );
nand U133993 ( n7411, n22954, n22955 );
nand U133994 ( n22955, n76757, n22956 );
nor U133995 ( n22954, n22957, n22958 );
and U133996 ( n22958, n22951, P1_P2_EBX_REG_13_ );
nand U133997 ( n7401, n22975, n22976 );
nand U133998 ( n22976, n76757, n22977 );
nor U133999 ( n22975, n22978, n22979 );
and U134000 ( n22979, n22972, P1_P2_EBX_REG_11_ );
nand U134001 ( n7391, n22994, n22995 );
nand U134002 ( n22995, n76757, n22996 );
nor U134003 ( n22994, n22997, n22998 );
and U134004 ( n22998, n22991, P1_P2_EBX_REG_9_ );
nand U134005 ( n14176, n56012, n56013 );
nand U134006 ( n56013, n76689, n56014 );
nor U134007 ( n56012, n56015, n56016 );
and U134008 ( n56016, n56009, P2_P2_EBX_REG_19_ );
nand U134009 ( n14146, n56072, n56073 );
nand U134010 ( n56073, n76690, n56074 );
nor U134011 ( n56072, n56075, n56076 );
and U134012 ( n56076, n56069, P2_P2_EBX_REG_13_ );
nand U134013 ( n14136, n56091, n56092 );
nand U134014 ( n56092, n76690, n56093 );
nor U134015 ( n56091, n56094, n56095 );
and U134016 ( n56095, n56088, P2_P2_EBX_REG_11_ );
nand U134017 ( n14126, n56110, n56111 );
nand U134018 ( n56111, n76690, n56112 );
nor U134019 ( n56110, n56113, n56114 );
and U134020 ( n56114, n56107, P2_P2_EBX_REG_9_ );
nor U134021 ( n9793, n76634, n9797 );
or U134022 ( n9797, n73126, P1_P1_EBX_REG_1_ );
nor U134023 ( n64558, n76223, n64561 );
or U134024 ( n64561, n73121, P2_P3_EBX_REG_1_ );
nor U134025 ( n43716, n76364, n43719 );
or U134026 ( n43719, n73123, P2_P1_EBX_REG_1_ );
nand U134027 ( n21964, n21972, n21973 );
nand U134028 ( n21973, n21974, P1_P2_REIP_REG_29_ );
nand U134029 ( n21972, n21976, n76910 );
and U134030 ( n21974, n75064, n21975 );
nand U134031 ( n29279, n29287, n29288 );
nand U134032 ( n29288, n29289, P1_P3_REIP_REG_29_ );
nand U134033 ( n29287, n29291, n76901 );
and U134034 ( n29289, n75069, n29290 );
nand U134035 ( n63046, n63054, n63055 );
nand U134036 ( n63055, n63056, P2_P3_REIP_REG_29_ );
nand U134037 ( n63054, n63058, n76875 );
and U134038 ( n63056, n75070, n63057 );
nand U134039 ( n55074, n55082, n55083 );
nand U134040 ( n55083, n55084, P2_P2_REIP_REG_29_ );
nand U134041 ( n55082, n55086, n76884 );
and U134042 ( n55084, n75063, n55085 );
nand U134043 ( n9596, n9790, n9792 );
nand U134044 ( n9792, n4814, P1_P1_INSTQUEUE_REG_0__1_ );
nor U134045 ( n9790, n9793, n9794 );
and U134046 ( n9794, n9787, P1_P1_EBX_REG_1_ );
nand U134047 ( n11841, n64556, n64557 );
nand U134048 ( n64557, n5673, P2_P3_INSTQUEUE_REG_0__1_ );
nor U134049 ( n64556, n64558, n64559 );
and U134050 ( n64559, n64553, P2_P3_EBX_REG_1_ );
nand U134051 ( n16331, n43714, n43715 );
nand U134052 ( n43715, n7458, P2_P1_INSTQUEUE_REG_0__1_ );
nor U134053 ( n43714, n43716, n43717 );
and U134054 ( n43717, n43711, P2_P1_EBX_REG_1_ );
nor U134055 ( n23068, n76543, n23071 );
or U134056 ( n23071, n73120, P1_P2_EBX_REG_1_ );
nor U134057 ( n56189, n76285, n56192 );
or U134058 ( n56192, n73122, P2_P2_EBX_REG_1_ );
nand U134059 ( n7351, n23066, n23067 );
nand U134060 ( n23067, n3915, P1_P2_INSTQUEUE_REG_0__1_ );
nor U134061 ( n23066, n23068, n23069 );
nand U134062 ( n14086, n56187, n56188 );
nand U134063 ( n56188, n6548, P2_P2_INSTQUEUE_REG_0__1_ );
nor U134064 ( n56187, n56189, n56190 );
nor U134065 ( n63439, P1_P1_ADDRESS_REG_16_, n63443 );
nand U134066 ( n63443, n73049, n73508 );
nand U134067 ( n63528, n63535, n63481 );
nand U134068 ( n63535, n63536, n76874 );
nor U134069 ( n63536, P2_P3_EBX_REG_17_, n6329 );
nand U134070 ( n29629, n29636, n29582 );
nand U134071 ( n29636, n29637, n76900 );
nor U134072 ( n29637, P1_P3_EBX_REG_17_, n3695 );
nand U134073 ( n22308, n22315, n22261 );
nand U134074 ( n22315, n22316, n76909 );
nor U134075 ( n22316, P1_P2_EBX_REG_17_, n4589 );
nand U134076 ( n55420, n55427, n55373 );
nand U134077 ( n55427, n55428, n76883 );
nor U134078 ( n55428, P2_P2_EBX_REG_17_, n7222 );
nand U134079 ( n63182, n63189, n63190 );
nand U134080 ( n63190, n63191, n63192 );
nand U134081 ( n63189, n63194, n76874 );
nor U134082 ( n63192, P2_P3_REIP_REG_25_, n74987 );
nand U134083 ( n63351, n63358, n63359 );
nand U134084 ( n63359, n63360, n63337 );
nand U134085 ( n63358, n63361, n76874 );
nor U134086 ( n63360, P2_P3_REIP_REG_21_, n74928 );
nand U134087 ( n29419, n29426, n29427 );
nand U134088 ( n29427, n29428, n29429 );
nand U134089 ( n29426, n29431, n76900 );
nor U134090 ( n29429, P1_P3_REIP_REG_25_, n74988 );
nand U134091 ( n29522, n29529, n29530 );
nand U134092 ( n29530, n29531, n29508 );
nand U134093 ( n29529, n29532, n76900 );
nor U134094 ( n29531, P1_P3_REIP_REG_21_, n74929 );
nand U134095 ( n29369, n29376, n29377 );
nand U134096 ( n29377, n29378, n208 );
nand U134097 ( n29376, n29379, n76900 );
nor U134098 ( n29378, P1_P3_REIP_REG_27_, n73297 );
nand U134099 ( n22203, n22210, n22211 );
nand U134100 ( n22211, n22212, n22189 );
nand U134101 ( n22210, n22213, n76909 );
nor U134102 ( n22212, P1_P2_REIP_REG_21_, n74926 );
nand U134103 ( n22100, n22107, n22108 );
nand U134104 ( n22108, n22109, n22110 );
nand U134105 ( n22107, n22112, n76909 );
nor U134106 ( n22110, P1_P2_REIP_REG_25_, n74970 );
nand U134107 ( n55317, n55324, n55325 );
nand U134108 ( n55325, n55326, n55303 );
nand U134109 ( n55324, n55327, n76883 );
nor U134110 ( n55326, P2_P2_REIP_REG_21_, n74925 );
nand U134111 ( n55210, n55217, n55218 );
nand U134112 ( n55218, n55219, n55220 );
nand U134113 ( n55217, n55222, n76883 );
nor U134114 ( n55220, P2_P2_REIP_REG_25_, n74969 );
nand U134115 ( n63132, n63139, n63140 );
nand U134116 ( n63140, n63141, n479 );
nand U134117 ( n63139, n63142, n76874 );
nor U134118 ( n63141, P2_P3_REIP_REG_27_, n73296 );
nand U134119 ( n22050, n22057, n22058 );
nand U134120 ( n22058, n22059, n174 );
nand U134121 ( n22057, n22060, n76909 );
nor U134122 ( n22059, P1_P2_REIP_REG_27_, n73294 );
nand U134123 ( n55160, n55167, n55168 );
nand U134124 ( n55168, n55169, n446 );
nand U134125 ( n55167, n55170, n76883 );
nor U134126 ( n55169, P2_P2_REIP_REG_27_, n73295 );
nand U134127 ( n63420, n63421, n63422 );
nor U134128 ( n63421, P1_P1_ADDRESS_REG_22_, n63425 );
nor U134129 ( n63422, n63423, n63424 );
or U134130 ( n63425, P1_P1_ADDRESS_REG_23_, P1_P1_ADDRESS_REG_24_ );
or U134131 ( n63424, P1_P1_ADDRESS_REG_25_, P1_P1_ADDRESS_REG_26_ );
nand U134132 ( n5256, n30108, n30109 );
nand U134133 ( n30108, P1_P3_EBX_REG_31_, n30114 );
nand U134134 ( n30109, n30110, n30111 );
nand U134135 ( n30114, n3073, n30115 );
nand U134136 ( n11991, n64121, n64122 );
nand U134137 ( n64121, P2_P3_EBX_REG_31_, n64127 );
nand U134138 ( n64122, n64123, n64124 );
nand U134139 ( n64127, n5674, n64128 );
nand U134140 ( n7501, n22783, n22784 );
nand U134141 ( n22783, P1_P2_EBX_REG_31_, n22789 );
nand U134142 ( n22784, n22785, n22786 );
nand U134143 ( n22789, n3917, n22790 );
nand U134144 ( n14236, n55897, n55898 );
nand U134145 ( n55897, P2_P2_EBX_REG_31_, n55903 );
nand U134146 ( n55898, n55899, n55900 );
nand U134147 ( n55903, n6549, n55904 );
nand U134148 ( n16481, n43377, n43378 );
nand U134149 ( n43377, P2_P1_EBX_REG_31_, n43383 );
nand U134150 ( n43378, n43379, n43380 );
nand U134151 ( n43383, n7459, n43384 );
nand U134152 ( n9746, n9438, n9439 );
nand U134153 ( n9438, P1_P1_EBX_REG_31_, n9445 );
nand U134154 ( n9439, n9440, n9442 );
nand U134155 ( n9445, n4815, n9447 );
or U134156 ( n63442, P1_P1_ADDRESS_REG_19_, P1_P1_ADDRESS_REG_1_ );
nor U134157 ( n22774, n3875, n22773 );
nor U134158 ( n30095, n3032, n30094 );
nor U134159 ( n64112, n5633, n64111 );
nor U134160 ( n55888, n6508, n55887 );
nand U134161 ( n66684, n66785, P2_P3_PHYADDRPOINTER_REG_20_ );
nand U134162 ( n32081, n32139, P1_P3_PHYADDRPOINTER_REG_20_ );
nand U134163 ( n24849, n24907, P1_P2_PHYADDRPOINTER_REG_20_ );
nand U134164 ( n57983, n58044, P2_P2_PHYADDRPOINTER_REG_20_ );
nand U134165 ( n67099, n67118, P2_P3_PHYADDRPOINTER_REG_6_ );
nand U134166 ( n32443, n32462, P1_P3_PHYADDRPOINTER_REG_6_ );
nand U134167 ( n25201, n25220, P1_P2_PHYADDRPOINTER_REG_6_ );
nand U134168 ( n58337, n58356, P2_P2_PHYADDRPOINTER_REG_6_ );
nand U134169 ( n24783, n24808, P1_P2_PHYADDRPOINTER_REG_24_ );
nand U134170 ( n32015, n32040, P1_P3_PHYADDRPOINTER_REG_24_ );
nand U134171 ( n66618, n66643, P2_P3_PHYADDRPOINTER_REG_24_ );
nand U134172 ( n57917, n57942, P2_P2_PHYADDRPOINTER_REG_24_ );
nand U134173 ( n66878, n66914, P2_P3_PHYADDRPOINTER_REG_14_ );
nand U134174 ( n32240, n32275, P1_P3_PHYADDRPOINTER_REG_14_ );
nand U134175 ( n25002, n25038, P1_P2_PHYADDRPOINTER_REG_14_ );
nand U134176 ( n58137, n58173, P2_P2_PHYADDRPOINTER_REG_14_ );
nand U134177 ( n67057, n67064, P2_P3_PHYADDRPOINTER_REG_8_ );
nand U134178 ( n32394, n32401, P1_P3_PHYADDRPOINTER_REG_8_ );
nand U134179 ( n25157, n25166, P1_P2_PHYADDRPOINTER_REG_8_ );
nand U134180 ( n58295, n58302, P2_P2_PHYADDRPOINTER_REG_8_ );
nand U134181 ( n24729, n24739, P1_P2_PHYADDRPOINTER_REG_26_ );
nand U134182 ( n31961, n31971, P1_P3_PHYADDRPOINTER_REG_26_ );
nand U134183 ( n66564, n66574, P2_P3_PHYADDRPOINTER_REG_26_ );
nand U134184 ( n57863, n57873, P2_P2_PHYADDRPOINTER_REG_26_ );
nand U134185 ( n24818, n24860, P1_P2_PHYADDRPOINTER_REG_22_ );
nand U134186 ( n32050, n32092, P1_P3_PHYADDRPOINTER_REG_22_ );
nand U134187 ( n66653, n66695, P2_P3_PHYADDRPOINTER_REG_22_ );
nand U134188 ( n57952, n57994, P2_P2_PHYADDRPOINTER_REG_22_ );
nand U134189 ( n24648, n24696, P1_P2_PHYADDRPOINTER_REG_28_ );
nand U134190 ( n31862, n31908, P1_P3_PHYADDRPOINTER_REG_28_ );
nand U134191 ( n66485, n66531, P2_P3_PHYADDRPOINTER_REG_28_ );
nand U134192 ( n57784, n57830, P2_P2_PHYADDRPOINTER_REG_28_ );
nand U134193 ( n67138, n67158, P2_P3_PHYADDRPOINTER_REG_4_ );
nand U134194 ( n32482, n32502, P1_P3_PHYADDRPOINTER_REG_4_ );
nand U134195 ( n25240, n25260, P1_P2_PHYADDRPOINTER_REG_4_ );
nand U134196 ( n58376, n58396, P2_P2_PHYADDRPOINTER_REG_4_ );
nand U134197 ( n66989, n67022, P2_P3_PHYADDRPOINTER_REG_10_ );
nand U134198 ( n32350, n32359, P1_P3_PHYADDRPOINTER_REG_10_ );
nand U134199 ( n25113, n25122, P1_P2_PHYADDRPOINTER_REG_10_ );
nand U134200 ( n58251, n58260, P2_P2_PHYADDRPOINTER_REG_10_ );
xor U134201 ( n22773, n24617, P1_P2_PHYADDRPOINTER_REG_31_ );
nand U134202 ( n24617, n24618, P1_P2_PHYADDRPOINTER_REG_30_ );
xor U134203 ( n30094, n31831, P1_P3_PHYADDRPOINTER_REG_31_ );
nand U134204 ( n31831, n31832, P1_P3_PHYADDRPOINTER_REG_30_ );
xor U134205 ( n64111, n66454, P2_P3_PHYADDRPOINTER_REG_31_ );
nand U134206 ( n66454, n66455, P2_P3_PHYADDRPOINTER_REG_30_ );
xor U134207 ( n55887, n57749, P2_P2_PHYADDRPOINTER_REG_31_ );
nand U134208 ( n57749, n57750, P2_P2_PHYADDRPOINTER_REG_30_ );
nand U134209 ( n64080, n64049, n64081 );
nand U134210 ( n64081, P2_P3_PHYADDRPOINTER_REG_1_, n64082 );
nand U134211 ( n64082, n63070, n64083 );
nand U134212 ( n64083, P2_P3_PHYADDRPOINTER_REG_0_, n76226 );
nand U134213 ( n30063, n30032, n30064 );
nand U134214 ( n30064, P1_P3_PHYADDRPOINTER_REG_1_, n30065 );
nand U134215 ( n30065, n29303, n30066 );
nand U134216 ( n30066, P1_P3_PHYADDRPOINTER_REG_0_, n76493 );
nand U134217 ( n22740, n22709, n22741 );
nand U134218 ( n22741, P1_P2_PHYADDRPOINTER_REG_1_, n22742 );
nand U134219 ( n22742, n21988, n22743 );
nand U134220 ( n22743, P1_P2_PHYADDRPOINTER_REG_0_, n76546 );
nand U134221 ( n55856, n55825, n55857 );
nand U134222 ( n55857, P2_P2_PHYADDRPOINTER_REG_1_, n55858 );
nand U134223 ( n55858, n55098, n55859 );
nand U134224 ( n55859, P2_P2_PHYADDRPOINTER_REG_0_, n76292 );
or U134225 ( n63423, P1_P1_ADDRESS_REG_27_, P1_P1_ADDRESS_REG_28_ );
nand U134226 ( n54315, n54586, n54587 );
nand U134227 ( n54586, n54589, n74626 );
nand U134228 ( n54587, P2_P1_INSTQUEUEWR_ADDR_REG_4_, n54588 );
nand U134229 ( n54588, P2_P1_INSTQUEUERD_ADDR_REG_4_, n7795 );
nand U134230 ( n11765, n11767, P1_P1_PHYADDRPOINTER_REG_30_ );
and U134231 ( n11767, n74964, n11768 );
nand U134232 ( n45392, n49445, n49446 );
nand U134233 ( n49445, P2_BUF1_REG_0_, n76477 );
nand U134234 ( n49446, n49447, n76651 );
nor U134235 ( n49447, n76477, n76834 );
and U134236 ( n10848, n10778, P1_P1_EAX_REG_14_ );
and U134237 ( n10998, n10950, P1_P1_EAX_REG_11_ );
and U134238 ( n44731, n44693, P2_P1_EAX_REG_11_ );
and U134239 ( n44611, n44555, P2_P1_EAX_REG_14_ );
nand U134240 ( n49350, n49351, n49352 );
nand U134241 ( n49352, P2_P1_INSTQUEUE_REG_14__0_, n49353 );
nand U134242 ( n49351, n7440, n245 );
nand U134243 ( n49272, n49273, n49274 );
nand U134244 ( n49274, P2_P1_INSTQUEUE_REG_13__0_, n49275 );
nand U134245 ( n49273, n7442, n245 );
nand U134246 ( n49082, n49083, n49084 );
nand U134247 ( n49084, P2_P1_INSTQUEUE_REG_11__0_, n49085 );
nand U134248 ( n49083, n7443, n245 );
nand U134249 ( n48987, n48988, n48989 );
nand U134250 ( n48989, P2_P1_INSTQUEUE_REG_10__0_, n48990 );
nand U134251 ( n48988, n7444, n245 );
nand U134252 ( n48888, n48889, n48890 );
nand U134253 ( n48890, P2_P1_INSTQUEUE_REG_9__0_, n48891 );
nand U134254 ( n48889, n7445, n245 );
nand U134255 ( n43347, P2_P1_STATE2_REG_2_, n42617 );
nand U134256 ( n42785, n42786, n42787 );
or U134257 ( n42786, n74958, n42753 );
nand U134258 ( n42787, P2_P1_EBX_REG_21_, n42788 );
nand U134259 ( n42788, n42524, n42789 );
nand U134260 ( n42656, n42657, n42658 );
nand U134261 ( n42657, P2_P1_REIP_REG_25_, n42661 );
nand U134262 ( n42658, P2_P1_EBX_REG_25_, n42659 );
nand U134263 ( n42661, n42662, n42663 );
nand U134264 ( n48715, n48716, n48717 );
nand U134265 ( n48717, P2_P1_INSTQUEUE_REG_7__0_, n48718 );
nand U134266 ( n48716, n7447, n245 );
nand U134267 ( n48621, n48622, n48623 );
nand U134268 ( n48623, P2_P1_INSTQUEUE_REG_6__0_, n48624 );
nand U134269 ( n48622, n7448, n245 );
nand U134270 ( n48527, n48528, n48529 );
nand U134271 ( n48529, P2_P1_INSTQUEUE_REG_5__0_, n48530 );
nand U134272 ( n48528, n7449, n245 );
and U134273 ( n11288, n11278, P1_P1_EAX_REG_2_ );
and U134274 ( n44972, n44964, P2_P1_EAX_REG_2_ );
and U134275 ( n11148, n11100, P1_P1_EAX_REG_8_ );
and U134276 ( n11250, n11234, P1_P1_EAX_REG_5_ );
and U134277 ( n44865, n44813, P2_P1_EAX_REG_8_ );
and U134278 ( n44942, n44934, P2_P1_EAX_REG_5_ );
nand U134279 ( n43107, n43113, n43114 );
nand U134280 ( n43113, n43086, n73221 );
nand U134281 ( n43114, P2_P1_EBX_REG_9_, n43115 );
nand U134282 ( n43115, n42524, n43116 );
nand U134283 ( n42302, P3_REG2_REG_4_, n42299 );
nand U134284 ( n42603, n42604, n42605 );
or U134285 ( n42604, n75014, n42571 );
nand U134286 ( n42605, P2_P1_EBX_REG_27_, n42606 );
nand U134287 ( n42606, n42524, n42607 );
and U134288 ( n21194, n14758, P1_P1_INSTQUEUEWR_ADDR_REG_0_ );
and U134289 ( n14758, n21196, n21197 );
nand U134290 ( n21196, P1_P1_INSTQUEUERD_ADDR_REG_0_, n21200 );
nand U134291 ( n21197, n21198, n73533 );
nand U134292 ( n21200, n21201, n12837 );
or U134293 ( n63441, P1_P1_ADDRESS_REG_20_, P1_P1_ADDRESS_REG_21_ );
nand U134294 ( n42309, P3_REG1_REG_4_, n42299 );
nand U134295 ( n9191, n11590, n11592 );
nand U134296 ( n11592, P1_P1_LWORD_REG_0_, n76618 );
nor U134297 ( n11590, n11593, n11507 );
nor U134298 ( n11593, n73162, n76616 );
nand U134299 ( n21223, n21224, n21225 );
nand U134300 ( n21225, n21226, n21227 );
nand U134301 ( n21224, n21234, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nor U134302 ( n21227, n8262, n21228 );
nor U134303 ( n71332, n74486, n71104 );
nand U134304 ( n9266, n11502, n11503 );
nand U134305 ( n11503, P1_P1_UWORD_REG_0_, n76618 );
nor U134306 ( n11502, n11505, n11507 );
nor U134307 ( n11505, n74903, n76617 );
nand U134308 ( n6891, n24577, n24578 );
nand U134309 ( n24578, P1_P2_LWORD_REG_11_, n76532 );
nor U134310 ( n24577, n24511, n24579 );
nor U134311 ( n24579, n74679, n76529 );
nand U134312 ( n6881, n24587, n24588 );
nand U134313 ( n24588, P1_P2_LWORD_REG_13_, n76532 );
nor U134314 ( n24587, n24521, n24589 );
nor U134315 ( n24589, n74733, n76529 );
nand U134316 ( n13616, n57716, n57717 );
nand U134317 ( n57717, P2_P2_LWORD_REG_13_, n76274 );
nor U134318 ( n57716, n57649, n57718 );
nor U134319 ( n57718, n74732, n76271 );
nand U134320 ( n13626, n57706, n57707 );
nand U134321 ( n57707, P2_P2_LWORD_REG_11_, n76274 );
nor U134322 ( n57706, n57641, n57708 );
nor U134323 ( n57708, n74678, n76271 );
nand U134324 ( n6961, n24513, n24514 );
nand U134325 ( n24514, P1_P2_UWORD_REG_12_, n76532 );
nor U134326 ( n24513, n24515, n24516 );
nor U134327 ( n24516, n73394, n76530 );
nand U134328 ( n13696, n57643, n57644 );
nand U134329 ( n57644, P2_P2_UWORD_REG_12_, n76274 );
nor U134330 ( n57643, n57645, n57646 );
nor U134331 ( n57646, n73393, n76272 );
nand U134332 ( n13631, n57701, n57702 );
nand U134333 ( n57702, P2_P2_LWORD_REG_10_, n76274 );
nor U134334 ( n57701, n57637, n57703 );
nor U134335 ( n57703, n74632, n76271 );
nand U134336 ( n6896, n24572, n24573 );
nand U134337 ( n24573, P1_P2_LWORD_REG_10_, n76532 );
nor U134338 ( n24572, n24507, n24574 );
nor U134339 ( n24574, n74633, n76529 );
nand U134340 ( n6876, n24592, n24593 );
nand U134341 ( n24593, P1_P2_LWORD_REG_14_, n76532 );
nor U134342 ( n24592, n24525, n24594 );
nor U134343 ( n24594, n75273, n76529 );
nand U134344 ( n6901, n24567, n24568 );
nand U134345 ( n24568, P1_P2_LWORD_REG_9_, n76532 );
nor U134346 ( n24567, n24503, n24569 );
nor U134347 ( n24569, n75251, n76529 );
nand U134348 ( n6886, n24582, n24583 );
nand U134349 ( n24583, P1_P2_LWORD_REG_12_, n76532 );
nor U134350 ( n24582, n24515, n24584 );
nor U134351 ( n24584, n75274, n76529 );
nand U134352 ( n6966, n24509, n24510 );
nand U134353 ( n24510, P1_P2_UWORD_REG_11_, n76532 );
nor U134354 ( n24509, n24511, n24512 );
nor U134355 ( n24512, n75323, n76530 );
nand U134356 ( n6906, n24562, n24563 );
nand U134357 ( n24563, P1_P2_LWORD_REG_8_, n76532 );
nor U134358 ( n24562, n24499, n24564 );
nor U134359 ( n24564, n75275, n76529 );
nand U134360 ( n6981, n24497, n24498 );
nand U134361 ( n24498, P1_P2_UWORD_REG_8_, n76532 );
nor U134362 ( n24497, n24499, n24500 );
nor U134363 ( n24500, n75344, n76530 );
nand U134364 ( n6951, n24523, n24524 );
nand U134365 ( n24524, P1_P2_UWORD_REG_14_, n76532 );
nor U134366 ( n24523, n24525, n24526 );
nor U134367 ( n24526, n75403, n76530 );
nand U134368 ( n6956, n24519, n24520 );
nand U134369 ( n24520, P1_P2_UWORD_REG_13_, n76532 );
nor U134370 ( n24519, n24521, n24522 );
nor U134371 ( n24522, n75205, n76530 );
nand U134372 ( n13636, n57696, n57697 );
nand U134373 ( n57697, P2_P2_LWORD_REG_9_, n76274 );
nor U134374 ( n57696, n57630, n57698 );
nor U134375 ( n57698, n75249, n76271 );
nand U134376 ( n13701, n57639, n57640 );
nand U134377 ( n57640, P2_P2_UWORD_REG_11_, n76274 );
nor U134378 ( n57639, n57641, n57642 );
nor U134379 ( n57642, n75322, n76272 );
nand U134380 ( n6976, n24501, n24502 );
nand U134381 ( n24502, P1_P2_UWORD_REG_9_, n76532 );
nor U134382 ( n24501, n24503, n24504 );
nor U134383 ( n24504, n75037, n76530 );
nand U134384 ( n13621, n57711, n57712 );
nand U134385 ( n57712, P2_P2_LWORD_REG_12_, n76274 );
nor U134386 ( n57711, n57645, n57713 );
nor U134387 ( n57713, n75264, n76271 );
nand U134388 ( n13641, n57691, n57692 );
nand U134389 ( n57692, P2_P2_LWORD_REG_8_, n76274 );
nor U134390 ( n57691, n57626, n57693 );
nor U134391 ( n57693, n75265, n76271 );
nand U134392 ( n13716, n57624, n57625 );
nand U134393 ( n57625, P2_P2_UWORD_REG_8_, n76274 );
nor U134394 ( n57624, n57626, n57627 );
nor U134395 ( n57627, n75342, n76272 );
nand U134396 ( n13691, n57647, n57648 );
nand U134397 ( n57648, P2_P2_UWORD_REG_13_, n76274 );
nor U134398 ( n57647, n57649, n57650 );
nor U134399 ( n57650, n75203, n76272 );
nand U134400 ( n13711, n57628, n57629 );
nand U134401 ( n57629, P2_P2_UWORD_REG_9_, n76274 );
nor U134402 ( n57628, n57630, n57631 );
nor U134403 ( n57631, n75036, n76272 );
nand U134404 ( n13686, n57651, n57652 );
nand U134405 ( n57652, P2_P2_UWORD_REG_14_, n76274 );
nor U134406 ( n57651, n57653, n57654 );
nor U134407 ( n57654, n75402, n76272 );
nand U134408 ( n13611, n57721, n57722 );
nand U134409 ( n57722, P2_P2_LWORD_REG_14_, n76274 );
nor U134410 ( n57721, n57653, n57723 );
nor U134411 ( n57723, n75266, n76271 );
nand U134412 ( n13706, n57635, n57636 );
nand U134413 ( n57636, P2_P2_UWORD_REG_10_, n76274 );
nor U134414 ( n57635, n57637, n57638 );
nor U134415 ( n57638, n75343, n76272 );
nand U134416 ( n6971, n24505, n24506 );
nand U134417 ( n24506, P1_P2_UWORD_REG_10_, n76532 );
nor U134418 ( n24505, n24507, n24508 );
nor U134419 ( n24508, n75345, n76530 );
nand U134420 ( n6871, n24597, n24598 );
nand U134421 ( n24598, P1_P2_LWORD_REG_15_, n24463 );
nor U134422 ( n24597, n24599, n24600 );
nor U134423 ( n24599, n23882, n24530 );
nand U134424 ( n13606, n57729, n57730 );
nand U134425 ( n57730, P2_P2_LWORD_REG_15_, n57592 );
nor U134426 ( n57729, n57731, n57732 );
nor U134427 ( n57731, n57006, n57658 );
nand U134428 ( n13681, n57655, n57656 );
nand U134429 ( n57656, P2_P2_LWORD_REG_0_, n76274 );
nor U134430 ( n57655, n57657, n57594 );
nor U134431 ( n57657, n74490, n76272 );
nand U134432 ( n6946, n24527, n24528 );
nand U134433 ( n24528, P1_P2_LWORD_REG_0_, n76532 );
nor U134434 ( n24527, n24529, n24465 );
nor U134435 ( n24529, n74491, n76530 );
nand U134436 ( n11436, n66320, n66321 );
nand U134437 ( n66321, P2_P3_LWORD_REG_0_, n76208 );
nor U134438 ( n66320, n66322, n66167 );
nor U134439 ( n66322, n74487, n76206 );
nand U134440 ( n11391, n66387, n66388 );
nand U134441 ( n66388, P2_P3_LWORD_REG_9_, n76208 );
nor U134442 ( n66387, n66389, n66261 );
nor U134443 ( n66389, n75250, n76205 );
nand U134444 ( n11456, n66304, n66305 );
nand U134445 ( n66305, P2_P3_UWORD_REG_11_, n76208 );
nor U134446 ( n66304, n66306, n66307 );
nor U134447 ( n66306, n75346, n76206 );
nand U134448 ( n11446, n66312, n66313 );
nand U134449 ( n66313, P2_P3_UWORD_REG_13_, n76208 );
nor U134450 ( n66312, n66314, n66315 );
nor U134451 ( n66314, n75204, n76206 );
nand U134452 ( n11451, n66308, n66309 );
nand U134453 ( n66309, P2_P3_UWORD_REG_12_, n76208 );
nor U134454 ( n66308, n66310, n66311 );
nor U134455 ( n66310, n73390, n76206 );
nand U134456 ( n11366, n66402, n66403 );
nand U134457 ( n66403, P2_P3_LWORD_REG_14_, n76208 );
nor U134458 ( n66402, n66404, n66319 );
nor U134459 ( n66404, n75268, n76205 );
nand U134460 ( n11376, n66396, n66397 );
nand U134461 ( n66397, P2_P3_LWORD_REG_12_, n76208 );
nor U134462 ( n66396, n66398, n66311 );
nor U134463 ( n66398, n75269, n76205 );
nand U134464 ( n11396, n66384, n66385 );
nand U134465 ( n66385, P2_P3_LWORD_REG_8_, n76208 );
nor U134466 ( n66384, n66386, n66257 );
nor U134467 ( n66386, n75271, n76205 );
nand U134468 ( n13661, n57672, n57673 );
nand U134469 ( n57673, P2_P2_LWORD_REG_4_, n57592 );
nor U134470 ( n57672, n57674, n57611 );
nor U134471 ( n57674, n75267, n76271 );
nand U134472 ( n11441, n66316, n66317 );
nand U134473 ( n66317, P2_P3_UWORD_REG_14_, n76208 );
nor U134474 ( n66316, n66318, n66319 );
nor U134475 ( n66318, n75426, n76206 );
nand U134476 ( n6986, n24493, n24494 );
nand U134477 ( n24494, P1_P2_UWORD_REG_7_, n76532 );
nor U134478 ( n24493, n24495, n24496 );
nor U134479 ( n24495, n74972, n76530 );
nand U134480 ( n6921, n24548, n24549 );
nand U134481 ( n24549, P1_P2_LWORD_REG_5_, n24463 );
nor U134482 ( n24548, n24550, n24488 );
nor U134483 ( n24550, n74543, n76529 );
nand U134484 ( n6931, n24540, n24541 );
nand U134485 ( n24541, P1_P2_LWORD_REG_3_, n76532 );
nor U134486 ( n24540, n24542, n24480 );
nor U134487 ( n24542, n74510, n76530 );
nand U134488 ( n11466, n66258, n66259 );
nand U134489 ( n66259, P2_P3_UWORD_REG_9_, n76208 );
nor U134490 ( n66258, n66260, n66261 );
nor U134491 ( n66260, n75028, n76206 );
nand U134492 ( n11431, n66324, n66325 );
nand U134493 ( n66325, P2_P3_LWORD_REG_1_, n76208 );
nor U134494 ( n66324, n66326, n66229 );
nor U134495 ( n66326, n73127, n76206 );
nand U134496 ( n11371, n66399, n66400 );
nand U134497 ( n66400, P2_P3_LWORD_REG_13_, n76208 );
nor U134498 ( n66399, n66401, n66315 );
nor U134499 ( n66401, n74730, n76205 );
nand U134500 ( n11381, n66393, n66394 );
nand U134501 ( n66394, P2_P3_LWORD_REG_11_, n76208 );
nor U134502 ( n66393, n66395, n66307 );
nor U134503 ( n66395, n74675, n76205 );
nand U134504 ( n13721, n57620, n57621 );
nand U134505 ( n57621, P2_P2_UWORD_REG_7_, n76274 );
nor U134506 ( n57620, n57622, n57623 );
nor U134507 ( n57622, n74971, n76272 );
nand U134508 ( n11411, n66336, n66337 );
nand U134509 ( n66337, P2_P3_LWORD_REG_5_, n66165 );
nor U134510 ( n66336, n66338, n66245 );
nor U134511 ( n66338, n74539, n76205 );
nand U134512 ( n13656, n57679, n57680 );
nand U134513 ( n57680, P2_P2_LWORD_REG_5_, n57592 );
nor U134514 ( n57679, n57681, n57615 );
nor U134515 ( n57681, n74542, n76271 );
nand U134516 ( n11401, n66381, n66382 );
nand U134517 ( n66382, P2_P3_LWORD_REG_7_, n66165 );
nor U134518 ( n66381, n66383, n66253 );
nor U134519 ( n66383, n74581, n76205 );
nand U134520 ( n13646, n57687, n57688 );
nand U134521 ( n57688, P2_P2_LWORD_REG_7_, n57592 );
nor U134522 ( n57687, n57689, n57623 );
nor U134523 ( n57689, n74583, n76271 );
nand U134524 ( n13676, n57660, n57661 );
nand U134525 ( n57661, P2_P2_LWORD_REG_1_, n76274 );
nor U134526 ( n57660, n57662, n57599 );
nor U134527 ( n57662, n73128, n76272 );
nand U134528 ( n6941, n24532, n24533 );
nand U134529 ( n24533, P1_P2_LWORD_REG_1_, n76532 );
nor U134530 ( n24532, n24534, n24470 );
nor U134531 ( n24534, n73129, n76530 );
nand U134532 ( n11476, n66250, n66251 );
nand U134533 ( n66251, P2_P3_UWORD_REG_7_, n76208 );
nor U134534 ( n66250, n66252, n66253 );
nor U134535 ( n66252, n74968, n76206 );
nand U134536 ( n6936, n24536, n24537 );
nand U134537 ( n24537, P1_P2_LWORD_REG_2_, n76532 );
nor U134538 ( n24536, n24538, n24474 );
nor U134539 ( n24538, n75285, n76530 );
nand U134540 ( n11406, n66378, n66379 );
nand U134541 ( n66379, P2_P3_LWORD_REG_6_, n66165 );
nor U134542 ( n66378, n66380, n66249 );
nor U134543 ( n66380, n75270, n76205 );
nand U134544 ( n13651, n57683, n57684 );
nand U134545 ( n57684, P2_P2_LWORD_REG_6_, n57592 );
nor U134546 ( n57683, n57685, n57619 );
nor U134547 ( n57685, n75263, n76271 );
nand U134548 ( n13671, n57664, n57665 );
nand U134549 ( n57665, P2_P2_LWORD_REG_2_, n76274 );
nor U134550 ( n57664, n57666, n57603 );
nor U134551 ( n57666, n75283, n76272 );
nand U134552 ( n11426, n66327, n66328 );
nand U134553 ( n66328, P2_P3_LWORD_REG_2_, n76208 );
nor U134554 ( n66327, n66329, n66233 );
nor U134555 ( n66329, n75284, n76206 );
nand U134556 ( n11416, n66333, n66334 );
nand U134557 ( n66334, P2_P3_LWORD_REG_4_, n66165 );
nor U134558 ( n66333, n66335, n66241 );
nor U134559 ( n66335, n75272, n76205 );
nand U134560 ( n6916, n24552, n24553 );
nand U134561 ( n24553, P1_P2_LWORD_REG_6_, n24463 );
nor U134562 ( n24552, n24554, n24492 );
nor U134563 ( n24554, n75277, n76529 );
nand U134564 ( n6926, n24544, n24545 );
nand U134565 ( n24545, P1_P2_LWORD_REG_4_, n24463 );
nor U134566 ( n24544, n24546, n24484 );
nor U134567 ( n24546, n75276, n76529 );
nand U134568 ( n11421, n66330, n66331 );
nand U134569 ( n66331, P2_P3_LWORD_REG_3_, n76208 );
nor U134570 ( n66330, n66332, n66237 );
nor U134571 ( n66332, n74507, n76206 );
nand U134572 ( n13666, n57668, n57669 );
nand U134573 ( n57669, P2_P2_LWORD_REG_3_, n76274 );
nor U134574 ( n57668, n57670, n57607 );
nor U134575 ( n57670, n74509, n76272 );
nand U134576 ( n6911, n24556, n24557 );
nand U134577 ( n24557, P1_P2_LWORD_REG_7_, n24463 );
nor U134578 ( n24556, n24558, n24496 );
nor U134579 ( n24558, n74584, n76529 );
nand U134580 ( n11461, n66262, n66263 );
nand U134581 ( n66263, P2_P3_UWORD_REG_10_, n76208 );
nor U134582 ( n66262, n66264, n66265 );
nor U134583 ( n66264, n75389, n76206 );
nand U134584 ( n11471, n66254, n66255 );
nand U134585 ( n66255, P2_P3_UWORD_REG_8_, n76208 );
nor U134586 ( n66254, n66256, n66257 );
nor U134587 ( n66256, n75390, n76206 );
nand U134588 ( n11386, n66390, n66391 );
nand U134589 ( n66391, P2_P3_LWORD_REG_10_, n66165 );
nor U134590 ( n66390, n66392, n66265 );
nor U134591 ( n66392, n74628, n76205 );
nand U134592 ( n11361, n66405, n66406 );
nand U134593 ( n66406, P2_P3_LWORD_REG_15_, n66165 );
nor U134594 ( n66405, n66407, n66408 );
nor U134595 ( n66408, n75364, n66323 );
nand U134596 ( n9400, P1_P1_STATE2_REG_2_, n8559 );
nand U134597 ( n8734, n8735, n8737 );
or U134598 ( n8735, n74959, n8694 );
nand U134599 ( n8737, P1_P1_EBX_REG_21_, n8738 );
nand U134600 ( n8738, n8428, n8739 );
nand U134601 ( n8608, n8609, n8610 );
nand U134602 ( n8609, P1_P1_REIP_REG_25_, n8614 );
nand U134603 ( n8610, P1_P1_EBX_REG_25_, n8612 );
nand U134604 ( n8614, n8615, n8617 );
nand U134605 ( n7001, n24481, n24482 );
nand U134606 ( n24482, P1_P2_UWORD_REG_4_, n76532 );
nor U134607 ( n24481, n24483, n24484 );
nor U134608 ( n24483, n75385, n76531 );
nand U134609 ( n7011, n24471, n24472 );
nand U134610 ( n24472, P1_P2_UWORD_REG_2_, n76532 );
nor U134611 ( n24471, n24473, n24474 );
nor U134612 ( n24473, n75386, n76531 );
nand U134613 ( n6991, n24489, n24490 );
nand U134614 ( n24490, P1_P2_UWORD_REG_6_, n76532 );
nor U134615 ( n24489, n24491, n24492 );
nor U134616 ( n24491, n75387, n76531 );
nand U134617 ( n11481, n66246, n66247 );
nand U134618 ( n66247, P2_P3_UWORD_REG_6_, n76208 );
nor U134619 ( n66246, n66248, n66249 );
nor U134620 ( n66248, n75381, n76207 );
nand U134621 ( n13726, n57616, n57617 );
nand U134622 ( n57617, P2_P2_UWORD_REG_6_, n76274 );
nor U134623 ( n57616, n57618, n57619 );
nor U134624 ( n57618, n75377, n76273 );
nand U134625 ( n13736, n57608, n57609 );
nand U134626 ( n57609, P2_P2_UWORD_REG_4_, n76274 );
nor U134627 ( n57608, n57610, n57611 );
nor U134628 ( n57610, n75378, n76273 );
nand U134629 ( n13746, n57600, n57601 );
nand U134630 ( n57601, P2_P2_UWORD_REG_2_, n76274 );
nor U134631 ( n57600, n57602, n57603 );
nor U134632 ( n57602, n75379, n76273 );
nand U134633 ( n11501, n66230, n66231 );
nand U134634 ( n66231, P2_P3_UWORD_REG_2_, n76208 );
nor U134635 ( n66230, n66232, n66233 );
nor U134636 ( n66232, n75382, n76207 );
nand U134637 ( n11491, n66238, n66239 );
nand U134638 ( n66239, P2_P3_UWORD_REG_4_, n76208 );
nor U134639 ( n66238, n66240, n66241 );
nor U134640 ( n66240, n75383, n76207 );
nand U134641 ( n13756, n57590, n57591 );
nand U134642 ( n57591, P2_P2_UWORD_REG_0_, n76274 );
nor U134643 ( n57590, n57593, n57594 );
nor U134644 ( n57593, n75380, n76273 );
nand U134645 ( n7021, n24461, n24462 );
nand U134646 ( n24462, P1_P2_UWORD_REG_0_, n76532 );
nor U134647 ( n24461, n24464, n24465 );
nor U134648 ( n24464, n75388, n76531 );
nand U134649 ( n11511, n66163, n66164 );
nand U134650 ( n66164, P2_P3_UWORD_REG_0_, n76208 );
nor U134651 ( n66163, n66166, n66167 );
nor U134652 ( n66166, n75384, n76207 );
nand U134653 ( n11496, n66234, n66235 );
nand U134654 ( n66235, P2_P3_UWORD_REG_3_, n76208 );
nor U134655 ( n66234, n66236, n66237 );
nor U134656 ( n66236, n74875, n76207 );
nand U134657 ( n11486, n66242, n66243 );
nand U134658 ( n66243, P2_P3_UWORD_REG_5_, n76208 );
nor U134659 ( n66242, n66244, n66245 );
nor U134660 ( n66244, n74921, n76207 );
nand U134661 ( n7006, n24477, n24478 );
nand U134662 ( n24478, P1_P2_UWORD_REG_3_, n76532 );
nor U134663 ( n24477, n24479, n24480 );
nor U134664 ( n24479, n74878, n76531 );
nand U134665 ( n6996, n24485, n24486 );
nand U134666 ( n24486, P1_P2_UWORD_REG_5_, n24463 );
nor U134667 ( n24485, n24487, n24488 );
nor U134668 ( n24487, n74923, n76531 );
nand U134669 ( n13731, n57612, n57613 );
nand U134670 ( n57613, P2_P2_UWORD_REG_5_, n76274 );
nor U134671 ( n57612, n57614, n57615 );
nor U134672 ( n57614, n74922, n76273 );
nand U134673 ( n13741, n57604, n57605 );
nand U134674 ( n57605, P2_P2_UWORD_REG_3_, n57592 );
nor U134675 ( n57604, n57606, n57607 );
nor U134676 ( n57606, n74877, n76273 );
nand U134677 ( n11506, n66226, n66227 );
nand U134678 ( n66227, P2_P3_UWORD_REG_1_, n76208 );
nor U134679 ( n66226, n66228, n66229 );
nor U134680 ( n66228, n74814, n76207 );
nand U134681 ( n7016, n24467, n24468 );
nand U134682 ( n24468, P1_P2_UWORD_REG_1_, n76532 );
nor U134683 ( n24467, n24469, n24470 );
nor U134684 ( n24469, n74820, n76531 );
nand U134685 ( n13751, n57596, n57597 );
nand U134686 ( n57597, P2_P2_UWORD_REG_1_, n76274 );
nor U134687 ( n57596, n57598, n57599 );
nor U134688 ( n57598, n74819, n76273 );
nand U134689 ( n42339, P3_REG2_REG_3_, n42251 );
nand U134690 ( n9119, n9127, n9128 );
nand U134691 ( n9127, n9093, n73222 );
nand U134692 ( n9128, P1_P1_EBX_REG_9_, n9129 );
nand U134693 ( n9129, n8428, n9130 );
nand U134694 ( n8542, n8543, n8544 );
or U134695 ( n8543, n75015, n8502 );
nand U134696 ( n8544, P1_P1_EBX_REG_27_, n8545 );
nand U134697 ( n8545, n8428, n8547 );
nand U134698 ( n8423, n8424, n8425 );
nand U134699 ( n8424, n8430, n75217 );
nand U134700 ( n8425, P1_P1_EBX_REG_30_, n8427 );
nand U134701 ( n8427, n8428, n8429 );
and U134702 ( n30141, n30134, P1_P3_EBX_REG_28_ );
nand U134703 ( n5241, n30137, n30138 );
or U134704 ( n30138, n30139, n30123 );
nor U134705 ( n30137, n30140, n30141 );
nor U134706 ( n30140, P1_P3_EBX_REG_28_, n30135 );
nand U134707 ( n16486, n43339, n43340 );
nor U134708 ( n43339, n43359, n43360 );
nor U134709 ( n43340, n43341, n43342 );
nor U134710 ( n43360, P2_P1_INSTQUEUERD_ADDR_REG_0_, n43332 );
nand U134711 ( n42353, P3_REG1_REG_3_, n42251 );
nand U134712 ( n16466, n43406, n43407 );
or U134713 ( n43407, n43408, n43392 );
nor U134714 ( n43406, n43409, n43410 );
nor U134715 ( n43409, P2_P1_EBX_REG_28_, n43404 );
and U134716 ( n43410, n43403, P2_P1_EBX_REG_28_ );
and U134717 ( n64154, n64147, P2_P3_EBX_REG_28_ );
and U134718 ( n22816, n22809, P1_P2_EBX_REG_28_ );
and U134719 ( n55930, n55923, P2_P2_EBX_REG_28_ );
nand U134720 ( n7486, n22812, n22813 );
nand U134721 ( n22813, n22814, n76756 );
nor U134722 ( n22812, n22815, n22816 );
nor U134723 ( n22815, P1_P2_EBX_REG_28_, n22810 );
nand U134724 ( n14221, n55926, n55927 );
nand U134725 ( n55927, n55928, n76689 );
nor U134726 ( n55926, n55929, n55930 );
nor U134727 ( n55929, P2_P2_EBX_REG_28_, n55924 );
nand U134728 ( n9731, n9474, n9475 );
or U134729 ( n9475, n9477, n9457 );
nor U134730 ( n9474, n9478, n9479 );
nor U134731 ( n9478, P1_P1_EBX_REG_28_, n9472 );
and U134732 ( n9479, n9470, P1_P1_EBX_REG_28_ );
nand U134733 ( n11976, n64150, n64151 );
or U134734 ( n64151, n64152, n64136 );
nor U134735 ( n64150, n64153, n64154 );
nor U134736 ( n64153, P2_P3_EBX_REG_28_, n64148 );
nand U134737 ( n13813, P1_P1_INSTADDRPOINTER_REG_8_, n76606 );
nand U134738 ( n10524, n10525, n10527 );
nand U134739 ( n10527, n10528, n76891 );
nand U134740 ( n10525, P1_P1_EAX_REG_19_, n10478 );
nor U134741 ( n10528, P1_P1_EAX_REG_19_, n10475 );
nand U134742 ( n10363, n10364, n10365 );
nand U134743 ( n10365, n10367, n76891 );
nand U134744 ( n10364, P1_P1_EAX_REG_22_, n10247 );
nor U134745 ( n10367, P1_P1_EAX_REG_22_, n10245 );
nand U134746 ( n44343, n44344, n44345 );
nand U134747 ( n44345, n44346, n76865 );
nand U134748 ( n44344, P2_P1_EAX_REG_19_, n44306 );
nor U134749 ( n44346, P2_P1_EAX_REG_19_, n44304 );
nand U134750 ( n44214, n44215, n44216 );
nand U134751 ( n44216, n44217, n76865 );
nand U134752 ( n44215, P2_P1_EAX_REG_22_, n44121 );
nor U134753 ( n44217, P2_P1_EAX_REG_22_, n44120 );
nand U134754 ( n44486, n44487, n44488 );
nand U134755 ( n44488, n44489, n76865 );
nand U134756 ( n44487, P2_P1_EAX_REG_16_, n44448 );
nor U134757 ( n44489, P2_P1_EAX_REG_16_, n44447 );
nand U134758 ( n10685, n10687, n10688 );
nand U134759 ( n10688, n10689, n76891 );
nand U134760 ( n10687, P1_P1_EAX_REG_16_, n10638 );
nor U134761 ( n10689, P1_P1_EAX_REG_16_, n10637 );
nor U134762 ( n71103, n74495, n71104 );
nand U134763 ( n9960, n9962, n9963 );
nand U134764 ( n9963, n9964, n76891 );
nand U134765 ( n9962, P1_P1_EAX_REG_28_, n9909 );
nor U134766 ( n9964, P1_P1_EAX_REG_28_, n9907 );
nand U134767 ( n43885, n43886, n43887 );
nand U134768 ( n43887, n43888, n76865 );
nand U134769 ( n43886, P2_P1_EAX_REG_28_, n43809 );
nor U134770 ( n43888, P2_P1_EAX_REG_28_, n43807 );
nand U134771 ( n10125, n10127, n10128 );
nand U134772 ( n10128, n10129, n76891 );
nand U134773 ( n10127, P1_P1_EAX_REG_25_, n10069 );
nor U134774 ( n10129, P1_P1_EAX_REG_25_, n10068 );
nand U134775 ( n44024, n44025, n44026 );
nand U134776 ( n44026, n44027, n76865 );
nand U134777 ( n44025, P2_P1_EAX_REG_25_, n43983 );
nor U134778 ( n44027, P2_P1_EAX_REG_25_, n43982 );
nand U134779 ( n67166, P2_P3_PHYADDRPOINTER_REG_1_, P2_P3_PHYADDRPOINTER_REG_2_ );
nand U134780 ( n32510, P1_P3_PHYADDRPOINTER_REG_1_, P1_P3_PHYADDRPOINTER_REG_2_ );
nand U134781 ( n25268, P1_P2_PHYADDRPOINTER_REG_1_, P1_P2_PHYADDRPOINTER_REG_2_ );
nand U134782 ( n58404, P2_P2_PHYADDRPOINTER_REG_1_, P2_P2_PHYADDRPOINTER_REG_2_ );
nand U134783 ( n15926, n45388, n45389 );
nand U134784 ( n45389, P2_P1_LWORD_REG_0_, n45325 );
nor U134785 ( n45388, n45390, n45327 );
nor U134786 ( n45390, n73161, n76350 );
nor U134787 ( n63741, P2_P3_REIP_REG_11_, n478 );
nor U134788 ( n63897, P2_P3_REIP_REG_5_, n478 );
nor U134789 ( n29781, P1_P3_REIP_REG_11_, n207 );
nor U134790 ( n29941, P1_P3_REIP_REG_5_, n207 );
nor U134791 ( n22460, P1_P2_REIP_REG_11_, n173 );
nor U134792 ( n22618, P1_P2_REIP_REG_5_, n173 );
nor U134793 ( n55575, P2_P2_REIP_REG_11_, n445 );
nor U134794 ( n55731, P2_P2_REIP_REG_5_, n445 );
nand U134795 ( n63641, n63642, n63643 );
nand U134796 ( n63642, P2_P3_PHYADDRPOINTER_REG_13_, n5629 );
nand U134797 ( n63643, P2_P3_REIP_REG_13_, n63644 );
nand U134798 ( n63644, n63645, n63646 );
nand U134799 ( n63858, n63859, n63860 );
nand U134800 ( n63859, P2_P3_PHYADDRPOINTER_REG_7_, n5629 );
nand U134801 ( n63860, P2_P3_REIP_REG_7_, n63861 );
nand U134802 ( n63861, n63862, n63863 );
nand U134803 ( n29742, n29743, n29744 );
nand U134804 ( n29743, P1_P3_PHYADDRPOINTER_REG_13_, n3028 );
nand U134805 ( n29744, P1_P3_REIP_REG_13_, n29745 );
nand U134806 ( n29745, n29746, n29747 );
nand U134807 ( n29902, n29903, n29904 );
nand U134808 ( n29903, P1_P3_PHYADDRPOINTER_REG_7_, n3028 );
nand U134809 ( n29904, P1_P3_REIP_REG_7_, n29905 );
nand U134810 ( n29905, n29906, n29907 );
nand U134811 ( n22421, n22422, n22423 );
nand U134812 ( n22422, P1_P2_PHYADDRPOINTER_REG_13_, n3872 );
nand U134813 ( n22423, P1_P2_REIP_REG_13_, n22424 );
nand U134814 ( n22424, n22425, n22426 );
nand U134815 ( n22579, n22580, n22581 );
nand U134816 ( n22580, P1_P2_PHYADDRPOINTER_REG_7_, n3872 );
nand U134817 ( n22581, P1_P2_REIP_REG_7_, n22582 );
nand U134818 ( n22582, n22583, n22584 );
nand U134819 ( n55536, n55537, n55538 );
nand U134820 ( n55537, P2_P2_PHYADDRPOINTER_REG_13_, n6504 );
nand U134821 ( n55538, P2_P2_REIP_REG_13_, n55539 );
nand U134822 ( n55539, n55540, n55541 );
nand U134823 ( n55692, n55693, n55694 );
nand U134824 ( n55693, P2_P2_PHYADDRPOINTER_REG_7_, n6504 );
nand U134825 ( n55694, P2_P2_REIP_REG_7_, n55695 );
nand U134826 ( n55695, n55696, n55697 );
nor U134827 ( n63977, P2_P3_REIP_REG_2_, n478 );
nor U134828 ( n30021, P1_P3_REIP_REG_2_, n207 );
nor U134829 ( n55814, P2_P2_REIP_REG_2_, n445 );
nor U134830 ( n22698, P1_P2_REIP_REG_2_, n173 );
nand U134831 ( n34233, n35682, n35683 );
nand U134832 ( n35682, P1_P3_INSTQUEUERD_ADDR_REG_0_, n35686 );
nand U134833 ( n35683, n35684, n73532 );
nand U134834 ( n35686, n35687, n32707 );
nand U134835 ( n26988, n28503, n28504 );
nand U134836 ( n28503, P1_P2_INSTQUEUERD_ADDR_REG_0_, n28507 );
nand U134837 ( n28504, n28505, n73520 );
nand U134838 ( n28507, n28508, n25467 );
nand U134839 ( n68987, n70408, n70409 );
nand U134840 ( n70408, P2_P3_INSTQUEUERD_ADDR_REG_0_, n70412 );
nand U134841 ( n70409, n70410, n73518 );
nand U134842 ( n70412, n70413, n67472 );
nand U134843 ( n60131, n61808, n61809 );
nand U134844 ( n61808, P2_P2_INSTQUEUERD_ADDR_REG_0_, n61812 );
nand U134845 ( n61809, n61810, n73521 );
nand U134846 ( n61812, n61813, n58604 );
nand U134847 ( n47979, n54180, n54181 );
nand U134848 ( n54180, P2_P1_INSTQUEUERD_ADDR_REG_0_, n54184 );
nand U134849 ( n54181, n54182, n73512 );
nand U134850 ( n54184, n54185, n46408 );
nand U134851 ( n16001, n45323, n45324 );
nand U134852 ( n45324, P2_P1_UWORD_REG_0_, n76352 );
nor U134853 ( n45323, n45326, n45327 );
nor U134854 ( n45326, n74902, n76351 );
nand U134855 ( n42520, n42521, n42522 );
nand U134856 ( n42521, P2_P1_REIP_REG_30_, n42503 );
nand U134857 ( n42522, P2_P1_EBX_REG_30_, n42523 );
nand U134858 ( n42523, n42524, n42525 );
nand U134859 ( n63944, n63975, P2_P3_REIP_REG_2_ );
nor U134860 ( n63975, n478, n73163 );
nand U134861 ( n29988, n30019, P1_P3_REIP_REG_2_ );
nor U134862 ( n30019, n207, n73164 );
nand U134863 ( n22665, n22696, P1_P2_REIP_REG_2_ );
nor U134864 ( n22696, n173, n72958 );
nand U134865 ( n55778, n55812, P2_P2_REIP_REG_2_ );
nor U134866 ( n55812, n445, n72959 );
nor U134867 ( n63943, n63944, n63945 );
nand U134868 ( n63945, P2_P3_REIP_REG_3_, n74642 );
nor U134869 ( n29987, n29988, n29989 );
nand U134870 ( n29989, P1_P3_REIP_REG_3_, n74643 );
nor U134871 ( n22664, n22665, n22666 );
nand U134872 ( n22666, P1_P2_REIP_REG_3_, n74641 );
nor U134873 ( n55777, n55778, n55779 );
nand U134874 ( n55779, P2_P2_REIP_REG_3_, n74640 );
nor U134875 ( n63811, P2_P3_REIP_REG_8_, n478 );
nor U134876 ( n29855, P1_P3_REIP_REG_8_, n207 );
nor U134877 ( n22532, P1_P2_REIP_REG_8_, n173 );
nor U134878 ( n55645, P2_P2_REIP_REG_8_, n445 );
nand U134879 ( n63786, n63790, n63791 );
nand U134880 ( n63790, P2_P3_EBX_REG_10_, n474 );
nand U134881 ( n63791, P2_P3_REIP_REG_10_, n63792 );
nand U134882 ( n63792, n63793, n63794 );
nand U134883 ( n29826, n29830, n29831 );
nand U134884 ( n29830, P1_P3_EBX_REG_10_, n203 );
nand U134885 ( n29831, P1_P3_REIP_REG_10_, n29832 );
nand U134886 ( n29832, n29833, n29834 );
nand U134887 ( n22507, n22511, n22512 );
nand U134888 ( n22511, P1_P2_EBX_REG_10_, n169 );
nand U134889 ( n22512, P1_P2_REIP_REG_10_, n22513 );
nand U134890 ( n22513, n22514, n22515 );
nand U134891 ( n55620, n55624, n55625 );
nand U134892 ( n55624, P2_P2_EBX_REG_10_, n442 );
nand U134893 ( n55625, P2_P2_REIP_REG_10_, n55626 );
nand U134894 ( n55626, n55627, n55628 );
nand U134895 ( n43668, n43877, n43878 );
nand U134896 ( n43877, n43880, n43559 );
nand U134897 ( n43878, P3_REG1_REG_11_, n43879 );
nand U134898 ( n43879, n872, n882 );
nor U134899 ( n63112, n63149, n63150 );
nor U134900 ( n63150, n478, P2_P3_REIP_REG_26_ );
nor U134901 ( n29349, n29386, n29387 );
nor U134902 ( n29387, n207, P1_P3_REIP_REG_26_ );
nor U134903 ( n22030, n22067, n22068 );
nor U134904 ( n22068, n173, P1_P2_REIP_REG_26_ );
nor U134905 ( n55140, n55177, n55178 );
nor U134906 ( n55178, n445, P2_P2_REIP_REG_26_ );
nor U134907 ( n63331, n63368, n63369 );
nor U134908 ( n63369, n478, P2_P3_REIP_REG_20_ );
nor U134909 ( n63490, n63524, n63525 );
nor U134910 ( n63525, n478, P2_P3_REIP_REG_17_ );
nor U134911 ( n29591, n29625, n29626 );
nor U134912 ( n29626, n207, P1_P3_REIP_REG_17_ );
nor U134913 ( n29502, n29539, n29540 );
nor U134914 ( n29540, n207, P1_P3_REIP_REG_20_ );
nor U134915 ( n22270, n22304, n22305 );
nor U134916 ( n22305, n173, P1_P2_REIP_REG_17_ );
nor U134917 ( n55382, n55416, n55417 );
nor U134918 ( n55417, n445, P2_P2_REIP_REG_17_ );
nand U134919 ( n63486, n63487, n63488 );
nand U134920 ( n63487, P2_P3_PHYADDRPOINTER_REG_19_, n5629 );
nand U134921 ( n63488, P2_P3_REIP_REG_19_, n63489 );
nand U134922 ( n63489, n63490, n63491 );
nand U134923 ( n29587, n29588, n29589 );
nand U134924 ( n29588, P1_P3_PHYADDRPOINTER_REG_19_, n3028 );
nand U134925 ( n29589, P1_P3_REIP_REG_19_, n29590 );
nand U134926 ( n29590, n29591, n29592 );
nand U134927 ( n22266, n22267, n22268 );
nand U134928 ( n22267, P1_P2_PHYADDRPOINTER_REG_19_, n3872 );
nand U134929 ( n22268, P1_P2_REIP_REG_19_, n22269 );
nand U134930 ( n22269, n22270, n22271 );
nand U134931 ( n55378, n55379, n55380 );
nand U134932 ( n55379, P2_P2_PHYADDRPOINTER_REG_19_, n6504 );
nand U134933 ( n55380, P2_P2_REIP_REG_19_, n55381 );
nand U134934 ( n55381, n55382, n55383 );
nor U134935 ( n22183, n22220, n22221 );
nor U134936 ( n22221, n173, P1_P2_REIP_REG_20_ );
nor U134937 ( n55297, n55334, n55335 );
nor U134938 ( n55335, n445, P2_P2_REIP_REG_20_ );
nor U134939 ( n63202, n63211, n63212 );
nor U134940 ( n63212, n478, P2_P3_REIP_REG_23_ );
nor U134941 ( n29439, n29448, n29449 );
nor U134942 ( n29449, n207, P1_P3_REIP_REG_23_ );
nor U134943 ( n22120, n22129, n22130 );
nor U134944 ( n22130, n173, P1_P2_REIP_REG_23_ );
nor U134945 ( n55230, n55239, n55240 );
nor U134946 ( n55240, n445, P2_P2_REIP_REG_23_ );
nor U134947 ( n21241, n21245, n73525 );
nor U134948 ( n21245, n21246, n21247 );
nor U134949 ( n21246, n10273, n21248 );
nor U134950 ( n21247, P1_P1_INSTQUEUERD_ADDR_REG_0_, n14543 );
nand U134951 ( n43875, n43876, n43874 );
nand U134952 ( n43876, P3_REG1_REG_12_, n43872 );
nor U134953 ( n63576, n63592, n63593 );
nor U134954 ( n63593, n478, P2_P3_REIP_REG_14_ );
nor U134955 ( n29677, n29693, n29694 );
nor U134956 ( n29694, n207, P1_P3_REIP_REG_14_ );
nor U134957 ( n22356, n22372, n22373 );
nor U134958 ( n22373, n173, P1_P2_REIP_REG_14_ );
nor U134959 ( n55468, n55484, n55485 );
nor U134960 ( n55485, n445, P2_P2_REIP_REG_14_ );
nand U134961 ( n63569, n63573, n63574 );
nand U134962 ( n63573, P2_P3_EBX_REG_16_, n474 );
nand U134963 ( n63574, P2_P3_REIP_REG_16_, n63575 );
nand U134964 ( n63575, n63576, n63577 );
nand U134965 ( n29670, n29674, n29675 );
nand U134966 ( n29674, P1_P3_EBX_REG_16_, n203 );
nand U134967 ( n29675, P1_P3_REIP_REG_16_, n29676 );
nand U134968 ( n29676, n29677, n29678 );
nand U134969 ( n22349, n22353, n22354 );
nand U134970 ( n22353, P1_P2_EBX_REG_16_, n169 );
nand U134971 ( n22354, P1_P2_REIP_REG_16_, n22355 );
nand U134972 ( n22355, n22356, n22357 );
nand U134973 ( n55461, n55465, n55466 );
nand U134974 ( n55465, P2_P2_EBX_REG_16_, n442 );
nand U134975 ( n55466, P2_P2_REIP_REG_16_, n55467 );
nand U134976 ( n55467, n55468, n55469 );
nand U134977 ( n63807, n63808, n63809 );
nand U134978 ( n63808, P2_P3_PHYADDRPOINTER_REG_9_, n5629 );
or U134979 ( n63809, n73216, n63793 );
nand U134980 ( n29851, n29852, n29853 );
nand U134981 ( n29852, P1_P3_PHYADDRPOINTER_REG_9_, n3028 );
or U134982 ( n29853, n73217, n29833 );
nand U134983 ( n22528, n22529, n22530 );
nand U134984 ( n22529, P1_P2_PHYADDRPOINTER_REG_9_, n3872 );
or U134985 ( n22530, n73215, n22514 );
nand U134986 ( n55641, n55642, n55643 );
nand U134987 ( n55642, P2_P2_PHYADDRPOINTER_REG_9_, n6504 );
or U134988 ( n55643, n73214, n55627 );
nand U134989 ( n43664, n43863, n43864 );
nand U134990 ( n43863, n43557, n43559 );
nand U134991 ( n43864, P3_REG2_REG_11_, n43865 );
nand U134992 ( n43865, n875, n882 );
nand U134993 ( n16739, n17386, DIN_29_ );
nor U134994 ( n17386, n76929, n73422 );
xnor U134995 ( n37866, n37867, n37868 );
xor U134996 ( n37868, P4_REG2_REG_10_, n1950 );
nand U134997 ( n63734, n63738, n63739 );
nand U134998 ( n63738, P2_P3_EBX_REG_12_, n474 );
or U134999 ( n63739, n74800, n63645 );
nand U135000 ( n63890, n63894, n63895 );
nand U135001 ( n63894, P2_P3_EBX_REG_6_, n474 );
or U135002 ( n63895, n74711, n63862 );
nand U135003 ( n29774, n29778, n29779 );
nand U135004 ( n29778, P1_P3_EBX_REG_12_, n203 );
or U135005 ( n29779, n74801, n29746 );
nand U135006 ( n29934, n29938, n29939 );
nand U135007 ( n29938, P1_P3_EBX_REG_6_, n203 );
or U135008 ( n29939, n74712, n29906 );
nand U135009 ( n22453, n22457, n22458 );
nand U135010 ( n22457, P1_P2_EBX_REG_12_, n169 );
or U135011 ( n22458, n74799, n22425 );
nand U135012 ( n22611, n22615, n22616 );
nand U135013 ( n22615, P1_P2_EBX_REG_6_, n169 );
or U135014 ( n22616, n74710, n22583 );
nand U135015 ( n55568, n55572, n55573 );
nand U135016 ( n55572, P2_P2_EBX_REG_12_, n442 );
or U135017 ( n55573, n74798, n55540 );
nand U135018 ( n55724, n55728, n55729 );
nand U135019 ( n55728, P2_P2_EBX_REG_6_, n442 );
or U135020 ( n55729, n74709, n55696 );
xor U135021 ( n12402, P1_P1_INSTADDRPOINTER_REG_11_, n13700 );
xor U135022 ( n32371, P1_P3_INSTADDRPOINTER_REG_11_, n33387 );
nor U135023 ( n43854, n868, n43861 );
not U135024 ( n868, n43856 );
nand U135025 ( n43861, n43862, n43860 );
nand U135026 ( n43862, P3_REG2_REG_12_, n43858 );
xor U135027 ( n46070, P2_P1_INSTADDRPOINTER_REG_11_, n47108 );
nand U135028 ( n22020, n22032, n22033 );
nand U135029 ( n22033, n22034, n22035 );
nand U135030 ( n22032, n22037, n76547 );
nor U135031 ( n22035, P1_P2_REIP_REG_28_, n73294 );
nand U135032 ( n55130, n55142, n55143 );
nand U135033 ( n55143, n55144, n55145 );
nand U135034 ( n55142, n55147, n76293 );
nor U135035 ( n55145, P2_P2_REIP_REG_28_, n73295 );
nand U135036 ( n29339, n29351, n29352 );
nand U135037 ( n29352, n29353, n29354 );
nand U135038 ( n29351, n29356, n76494 );
nor U135039 ( n29354, P1_P3_REIP_REG_28_, n73297 );
nand U135040 ( n63102, n63114, n63115 );
nand U135041 ( n63115, n63116, n63117 );
nand U135042 ( n63114, n63119, n76227 );
nor U135043 ( n63117, P2_P3_REIP_REG_28_, n73296 );
nand U135044 ( n63321, n63333, n63334 );
nand U135045 ( n63334, n63335, n63336 );
nand U135046 ( n63333, n63338, n76227 );
nor U135047 ( n63336, P2_P3_REIP_REG_22_, n74928 );
nand U135048 ( n29492, n29504, n29505 );
nand U135049 ( n29505, n29506, n29507 );
nand U135050 ( n29504, n29509, n76494 );
nor U135051 ( n29507, P1_P3_REIP_REG_22_, n74929 );
nand U135052 ( n22173, n22185, n22186 );
nand U135053 ( n22186, n22187, n22188 );
nand U135054 ( n22185, n22190, n76547 );
nor U135055 ( n22188, P1_P2_REIP_REG_22_, n74926 );
nand U135056 ( n55287, n55299, n55300 );
nand U135057 ( n55300, n55301, n55302 );
nand U135058 ( n55299, n55304, n76293 );
nor U135059 ( n55302, P2_P2_REIP_REG_22_, n74925 );
xor U135060 ( n67034, P2_P3_INSTADDRPOINTER_REG_11_, n68139 );
xor U135061 ( n25134, P1_P2_INSTADDRPOINTER_REG_11_, n26136 );
xor U135062 ( n58272, P2_P2_INSTADDRPOINTER_REG_11_, n59277 );
and U135063 ( n23069, n23063, P1_P2_EBX_REG_1_ );
and U135064 ( n56190, n56184, P2_P2_EBX_REG_1_ );
or U135065 ( n63968, n75952, n75953 );
nor U135066 ( n75952, n73168, n63932 );
nor U135067 ( n75953, n63944, P2_P3_REIP_REG_3_ );
or U135068 ( n30012, n75954, n75955 );
nor U135069 ( n75954, n73169, n29976 );
nor U135070 ( n75955, n29988, P1_P3_REIP_REG_3_ );
or U135071 ( n22689, n75956, n75957 );
nor U135072 ( n75956, n72961, n22653 );
nor U135073 ( n75957, n22665, P1_P2_REIP_REG_3_ );
or U135074 ( n55805, n75958, n75959 );
nor U135075 ( n75958, n72960, n55766 );
nor U135076 ( n75959, n55778, P2_P2_REIP_REG_3_ );
nand U135077 ( n64041, n64050, n64051 );
nand U135078 ( n64051, n63977, P2_P3_REIP_REG_1_ );
nand U135079 ( n64050, n64052, n76226 );
nor U135080 ( n64052, n6153, n64053 );
nand U135081 ( n30024, n30033, n30034 );
nand U135082 ( n30034, n30021, P1_P3_REIP_REG_1_ );
nand U135083 ( n30033, n30035, n76493 );
nor U135084 ( n30035, n3538, n30036 );
nand U135085 ( n22701, n22710, n22711 );
nand U135086 ( n22711, n22698, P1_P2_REIP_REG_1_ );
nand U135087 ( n22710, n22712, n76546 );
nor U135088 ( n22712, n4375, n22713 );
nand U135089 ( n55817, n55826, n55827 );
nand U135090 ( n55827, n55814, P2_P2_REIP_REG_1_ );
nand U135091 ( n55826, n55828, n76292 );
nor U135092 ( n55828, n7008, n55829 );
nand U135093 ( n22125, n22126, n22127 );
nand U135094 ( n22127, n22128, n22111 );
or U135095 ( n22126, n74991, n22120 );
nor U135096 ( n22128, P1_P2_REIP_REG_24_, n74970 );
nand U135097 ( n55235, n55236, n55237 );
nand U135098 ( n55237, n55238, n55221 );
or U135099 ( n55236, n74990, n55230 );
nor U135100 ( n55238, P2_P2_REIP_REG_24_, n74969 );
nand U135101 ( n63589, n63590, n63591 );
nand U135102 ( n63590, P2_P3_PHYADDRPOINTER_REG_15_, n5629 );
or U135103 ( n63591, n74840, n63576 );
nand U135104 ( n29690, n29691, n29692 );
nand U135105 ( n29691, P1_P3_PHYADDRPOINTER_REG_15_, n3028 );
or U135106 ( n29692, n74839, n29677 );
nand U135107 ( n22369, n22370, n22371 );
nand U135108 ( n22370, P1_P2_PHYADDRPOINTER_REG_15_, n3872 );
or U135109 ( n22371, n74838, n22356 );
nand U135110 ( n55481, n55482, n55483 );
nand U135111 ( n55482, P2_P2_PHYADDRPOINTER_REG_15_, n6504 );
or U135112 ( n55483, n74837, n55468 );
nand U135113 ( n63207, n63208, n63209 );
nand U135114 ( n63209, n63210, n63193 );
or U135115 ( n63208, n74993, n63202 );
nor U135116 ( n63210, P2_P3_REIP_REG_24_, n74987 );
nand U135117 ( n29444, n29445, n29446 );
nand U135118 ( n29446, n29447, n29430 );
or U135119 ( n29445, n74994, n29439 );
nor U135120 ( n29447, P1_P3_REIP_REG_24_, n74988 );
nand U135121 ( n43238, n43239, n43240 );
nand U135122 ( n43239, P2_P1_REIP_REG_4_, n43246 );
nand U135123 ( n43240, n43241, n76863 );
nand U135124 ( n43246, n43247, n43248 );
nand U135125 ( n43296, n43297, n43298 );
nand U135126 ( n43297, P2_P1_REIP_REG_2_, n43291 );
nand U135127 ( n43298, n43299, n76863 );
nor U135128 ( n43299, n8119, n43300 );
nand U135129 ( n42849, n42850, n42851 );
nand U135130 ( n42850, n42857, n42832 );
nand U135131 ( n42851, n42852, n76862 );
nor U135132 ( n42857, P2_P1_REIP_REG_18_, n74904 );
nor U135133 ( n28630, n4255, n28644 );
nor U135134 ( n28644, n74423, P1_P2_INSTQUEUERD_ADDR_REG_0_ );
nor U135135 ( n61935, n6888, n61949 );
nor U135136 ( n61949, n74424, P2_P2_INSTQUEUERD_ADDR_REG_0_ );
nand U135137 ( n42744, n42745, n42746 );
nand U135138 ( n42745, P2_P1_REIP_REG_22_, n42752 );
nand U135139 ( n42746, n42747, n76862 );
nand U135140 ( n42752, n42753, n42754 );
nand U135141 ( n42562, n42563, n42564 );
nand U135142 ( n42563, P2_P1_REIP_REG_28_, n42570 );
nand U135143 ( n42564, n42565, n76862 );
nand U135144 ( n42570, n42571, n42572 );
nor U135145 ( n70535, n6033, n70549 );
nor U135146 ( n70549, n74425, P2_P3_INSTQUEUERD_ADDR_REG_0_ );
nor U135147 ( n35809, n3418, n35823 );
nor U135148 ( n35823, n74426, P1_P3_INSTQUEUERD_ADDR_REG_0_ );
nand U135149 ( n43098, n43105, n42829 );
nand U135150 ( n43105, n43106, n76863 );
nor U135151 ( n43106, P2_P1_EBX_REG_9_, n8115 );
nand U135152 ( n8963, n8964, n8965 );
nand U135153 ( n8964, n4751, P1_P1_PHYADDRPOINTER_REG_14_ );
nand U135154 ( n8965, n4759, n8957 );
nand U135155 ( n9030, n9032, n9033 );
nand U135156 ( n9032, n4751, P1_P1_PHYADDRPOINTER_REG_12_ );
nand U135157 ( n9033, n4759, n9024 );
nand U135158 ( n9095, n9097, n9098 );
nand U135159 ( n9097, n4751, P1_P1_PHYADDRPOINTER_REG_10_ );
nand U135160 ( n9098, n4759, n5292 );
nand U135161 ( n9158, n9159, n9160 );
nand U135162 ( n9159, n4751, P1_P1_PHYADDRPOINTER_REG_8_ );
nand U135163 ( n9160, n4759, n5290 );
nand U135164 ( n9295, n9297, n9298 );
nand U135165 ( n9297, n4751, P1_P1_PHYADDRPOINTER_REG_4_ );
nand U135166 ( n9298, n4759, n5288 );
nand U135167 ( n9357, n9358, n9359 );
nand U135168 ( n9358, n4751, P1_P1_PHYADDRPOINTER_REG_2_ );
nand U135169 ( n9359, n4759, n9354 );
nand U135170 ( n8837, n8838, n8839 );
nand U135171 ( n8838, n4751, P1_P1_PHYADDRPOINTER_REG_18_ );
nand U135172 ( n8839, n4759, n8830 );
nand U135173 ( n8900, n8902, n8903 );
nand U135174 ( n8902, n4751, P1_P1_PHYADDRPOINTER_REG_16_ );
nand U135175 ( n8903, n4759, n5295 );
nand U135176 ( n9225, n9227, n9228 );
nand U135177 ( n9227, n4751, P1_P1_PHYADDRPOINTER_REG_6_ );
nand U135178 ( n9228, n4759, n5289 );
nand U135179 ( n42506, n42514, n42515 );
nand U135180 ( n42515, n42516, P2_P1_REIP_REG_29_ );
nand U135181 ( n42514, n42518, n76863 );
nor U135182 ( n42516, P2_P1_REIP_REG_30_, n508 );
nand U135183 ( n42982, n42983, n42984 );
nand U135184 ( n42983, n7393, P2_P1_PHYADDRPOINTER_REG_14_ );
nand U135185 ( n42984, n7404, n42977 );
nand U135186 ( n43036, n43037, n43038 );
nand U135187 ( n43037, n7393, P2_P1_PHYADDRPOINTER_REG_12_ );
nand U135188 ( n43038, n7404, n43031 );
nand U135189 ( n43088, n43089, n43090 );
nand U135190 ( n43089, n7393, P2_P1_PHYADDRPOINTER_REG_10_ );
nand U135191 ( n43090, n7404, n7947 );
nand U135192 ( n43138, n43139, n43140 );
nand U135193 ( n43139, n7393, P2_P1_PHYADDRPOINTER_REG_8_ );
nand U135194 ( n43140, n7404, n7945 );
nand U135195 ( n43262, n43263, n43264 );
nand U135196 ( n43263, n7393, P2_P1_PHYADDRPOINTER_REG_4_ );
nand U135197 ( n43264, n7404, n7943 );
nand U135198 ( n43311, n43312, n43313 );
nand U135199 ( n43312, n7393, P2_P1_PHYADDRPOINTER_REG_2_ );
nand U135200 ( n43313, n7404, n43309 );
nand U135201 ( n42867, n42868, n42869 );
nand U135202 ( n42868, n7393, P2_P1_PHYADDRPOINTER_REG_18_ );
nand U135203 ( n42869, n7404, n42862 );
nand U135204 ( n42918, n42919, n42920 );
nand U135205 ( n42919, n7393, P2_P1_PHYADDRPOINTER_REG_16_ );
nand U135206 ( n42920, n7404, n7950 );
nand U135207 ( n43192, n43193, n43194 );
nand U135208 ( n43193, n7393, P2_P1_PHYADDRPOINTER_REG_6_ );
nand U135209 ( n43194, n7404, n7944 );
nand U135210 ( n42876, n42883, n42829 );
nand U135211 ( n42883, n42884, n76862 );
nor U135212 ( n42884, P2_P1_EBX_REG_17_, n8110 );
nand U135213 ( n42773, n42780, n42781 );
nand U135214 ( n42781, n42782, n42759 );
nand U135215 ( n42780, n42783, n76862 );
nor U135216 ( n42782, P2_P1_REIP_REG_21_, n74951 );
nand U135217 ( n42642, n42649, n42650 );
nand U135218 ( n42650, n42651, n42652 );
nand U135219 ( n42649, n42654, n76862 );
nor U135220 ( n42652, P2_P1_REIP_REG_25_, n74995 );
nand U135221 ( n42591, n42598, n42599 );
nand U135222 ( n42599, n42600, n505 );
nand U135223 ( n42598, n42601, n76862 );
nor U135224 ( n42600, P2_P1_REIP_REG_27_, n73308 );
nand U135225 ( n63518, n63522, n63523 );
nand U135226 ( n63522, P2_P3_EBX_REG_18_, n474 );
or U135227 ( n63523, n74900, n63490 );
nand U135228 ( n29619, n29623, n29624 );
nand U135229 ( n29623, P1_P3_EBX_REG_18_, n203 );
or U135230 ( n29624, n74901, n29591 );
nand U135231 ( n22298, n22302, n22303 );
nand U135232 ( n22302, P1_P2_EBX_REG_18_, n169 );
or U135233 ( n22303, n74899, n22270 );
nand U135234 ( n55410, n55414, n55415 );
nand U135235 ( n55414, P2_P2_EBX_REG_18_, n442 );
or U135236 ( n55415, n74898, n55382 );
nand U135237 ( n8483, n8484, n8485 );
nand U135238 ( n8485, n229, P1_P1_EBX_REG_29_ );
nand U135239 ( n8484, n4759, n8478 );
nand U135240 ( n8520, n8522, n8523 );
nand U135241 ( n8523, P1_P1_EBX_REG_28_, n229 );
nand U135242 ( n8522, n4759, n5304 );
nand U135243 ( n8713, n8714, n8715 );
nand U135244 ( n8715, P1_P1_EBX_REG_22_, n229 );
nand U135245 ( n8714, n4759, n5300 );
nand U135246 ( n8774, n8775, n8777 );
nand U135247 ( n8777, P1_P1_EBX_REG_20_, n229 );
nand U135248 ( n8775, n4759, n8762 );
nand U135249 ( n8584, n8585, n8587 );
nand U135250 ( n8587, P1_P1_EBX_REG_26_, n229 );
nand U135251 ( n8585, n4759, n5303 );
nand U135252 ( n8648, n8649, n8650 );
nand U135253 ( n8650, P1_P1_EBX_REG_24_, n229 );
nand U135254 ( n8649, n4759, n5302 );
nand U135255 ( n42556, n42557, n42558 );
nand U135256 ( n42558, n500, P2_P1_EBX_REG_29_ );
nand U135257 ( n42557, n7404, n7960 );
nand U135258 ( n42586, n42587, n42588 );
nand U135259 ( n42588, P2_P1_EBX_REG_28_, n500 );
nand U135260 ( n42587, n7404, n7959 );
nand U135261 ( n42817, n42818, n42819 );
nand U135262 ( n42819, P2_P1_EBX_REG_20_, n500 );
nand U135263 ( n42818, n7404, n42807 );
nand U135264 ( n42637, n42638, n42639 );
nand U135265 ( n42639, P2_P1_EBX_REG_26_, n500 );
nand U135266 ( n42638, n7404, n7958 );
nand U135267 ( n42712, n42713, n42714 );
nand U135268 ( n42714, P2_P1_EBX_REG_24_, n500 );
nand U135269 ( n42713, n7404, n7957 );
nand U135270 ( n42768, n42769, n42770 );
nand U135271 ( n42770, P2_P1_EBX_REG_22_, n500 );
nand U135272 ( n42769, n7404, n7955 );
nand U135273 ( n9265, n9267, n9268 );
nand U135274 ( n9267, P1_P1_REIP_REG_4_, n9275 );
nand U135275 ( n9268, n9269, n76890 );
nand U135276 ( n9275, n9277, n9278 );
nand U135277 ( n9338, n9339, n9340 );
nand U135278 ( n9339, P1_P1_REIP_REG_2_, n9332 );
nand U135279 ( n9340, n9342, n76890 );
nor U135280 ( n9342, n5465, n9343 );
nand U135281 ( n9108, n9117, n8789 );
nand U135282 ( n9117, n9118, n76890 );
nor U135283 ( n9118, P1_P1_EBX_REG_9_, n5462 );
nand U135284 ( n23252, n23253, n23254 );
nand U135285 ( n23254, n23255, n76540 );
nand U135286 ( n23253, P1_P2_EAX_REG_27_, n23214 );
nor U135287 ( n23255, P1_P2_EAX_REG_27_, n23207 );
nand U135288 ( n56376, n56377, n56378 );
nand U135289 ( n56378, n56379, n76282 );
nand U135290 ( n56377, P2_P2_EAX_REG_27_, n56335 );
nor U135291 ( n56379, P2_P2_EAX_REG_27_, n56328 );
nand U135292 ( n8814, n8815, n8817 );
nand U135293 ( n8815, n8824, n8793 );
nand U135294 ( n8817, n8818, n76889 );
nor U135295 ( n8824, P1_P1_REIP_REG_18_, n74905 );
nand U135296 ( n8490, n8492, n8493 );
nand U135297 ( n8492, P1_P1_REIP_REG_28_, n8500 );
nand U135298 ( n8493, n8494, n76889 );
nand U135299 ( n8500, n8502, n8503 );
nand U135300 ( n8683, n8684, n8685 );
nand U135301 ( n8684, P1_P1_REIP_REG_22_, n8693 );
nand U135302 ( n8685, n8687, n76889 );
nand U135303 ( n8693, n8694, n8695 );
nand U135304 ( n64732, n64733, n64734 );
nand U135305 ( n64734, n64735, n76216 );
nand U135306 ( n64733, P2_P3_EAX_REG_27_, n64693 );
nor U135307 ( n64735, P2_P3_EAX_REG_27_, n64691 );
nand U135308 ( n30573, n30574, n30575 );
nand U135309 ( n30575, n30576, n76483 );
nand U135310 ( n30574, P1_P3_EAX_REG_27_, n30534 );
nor U135311 ( n30576, P1_P3_EAX_REG_27_, n30532 );
nand U135312 ( n49698, n49704, n76929 );
xor U135313 ( n49704, n49705, n49706 );
nand U135314 ( n49706, P3_DATAO_REG_1_, DIN_30_ );
nand U135315 ( n49705, P3_DATAO_REG_2_, DIN_29_ );
nand U135316 ( n30392, n76024, P1_P3_EBX_REG_1_ );
nand U135317 ( n8848, n8857, n8789 );
nand U135318 ( n8857, n8858, n76889 );
nor U135319 ( n8858, P1_P1_EBX_REG_17_, n5457 );
nand U135320 ( n9789, n76037, P1_P1_EBX_REG_1_ );
nand U135321 ( n64555, n75992, P2_P3_EBX_REG_1_ );
nand U135322 ( n43713, n76008, P2_P1_EBX_REG_1_ );
nand U135323 ( n23065, n76029, P1_P2_EBX_REG_1_ );
nand U135324 ( n56186, n76000, P2_P2_EBX_REG_1_ );
nand U135325 ( n8719, n8728, n8729 );
nand U135326 ( n8729, n8730, n8702 );
nand U135327 ( n8728, n8732, n76889 );
nor U135328 ( n8730, P1_P1_REIP_REG_21_, n74952 );
nand U135329 ( n63549, n63565, n63481 );
nand U135330 ( n63565, n63566, n63567 );
nor U135331 ( n63567, P2_P3_REIP_REG_16_, n74830 );
and U135332 ( n63566, P2_P3_REIP_REG_15_, n63568 );
nand U135333 ( n29650, n29666, n29582 );
nand U135334 ( n29666, n29667, n29668 );
nor U135335 ( n29668, P1_P3_REIP_REG_16_, n74829 );
and U135336 ( n29667, P1_P3_REIP_REG_15_, n29669 );
nand U135337 ( n22329, n22345, n22261 );
nand U135338 ( n22345, n22346, n22347 );
nor U135339 ( n22347, P1_P2_REIP_REG_16_, n74828 );
and U135340 ( n22346, P1_P2_REIP_REG_15_, n22348 );
nand U135341 ( n55441, n55457, n55373 );
nand U135342 ( n55457, n55458, n55459 );
nor U135343 ( n55459, P2_P2_REIP_REG_16_, n74827 );
and U135344 ( n55458, P2_P2_REIP_REG_15_, n55460 );
nand U135345 ( n8590, n8599, n8600 );
nand U135346 ( n8600, n8602, n8603 );
nand U135347 ( n8599, n8605, n76889 );
nor U135348 ( n8603, P1_P1_REIP_REG_25_, n74996 );
nand U135349 ( n8527, n8535, n8537 );
nand U135350 ( n8537, n8538, n234 );
nand U135351 ( n8535, n8539, n76889 );
nor U135352 ( n8538, P1_P1_REIP_REG_27_, n73309 );
nand U135353 ( n29581, n29583, n29584 );
nor U135354 ( n29584, P1_P3_REIP_REG_19_, n74885 );
and U135355 ( n29583, P1_P3_REIP_REG_18_, n29585 );
nand U135356 ( n22260, n22262, n22263 );
nor U135357 ( n22263, P1_P2_REIP_REG_19_, n74883 );
and U135358 ( n22262, P1_P2_REIP_REG_18_, n22264 );
nand U135359 ( n55372, n55374, n55375 );
nor U135360 ( n55375, P2_P2_REIP_REG_19_, n74882 );
and U135361 ( n55374, P2_P2_REIP_REG_18_, n55376 );
and U135362 ( n63191, P2_P3_REIP_REG_24_, n63193 );
and U135363 ( n63335, P2_P3_REIP_REG_21_, n63337 );
and U135364 ( n29428, P1_P3_REIP_REG_24_, n29430 );
and U135365 ( n29506, P1_P3_REIP_REG_21_, n29508 );
and U135366 ( n22109, P1_P2_REIP_REG_24_, n22111 );
and U135367 ( n22187, P1_P2_REIP_REG_21_, n22189 );
and U135368 ( n55219, P2_P2_REIP_REG_24_, n55221 );
and U135369 ( n55301, P2_P2_REIP_REG_21_, n55303 );
nand U135370 ( n63480, n63482, n63483 );
nor U135371 ( n63483, P2_P3_REIP_REG_19_, n74884 );
and U135372 ( n63482, P2_P3_REIP_REG_18_, n63484 );
nand U135373 ( n56711, n56712, n56713 );
nand U135374 ( n56713, n56714, n76282 );
nand U135375 ( n56712, P2_P2_EAX_REG_21_, n56673 );
nor U135376 ( n56714, P2_P2_EAX_REG_21_, n56573 );
nand U135377 ( n56800, n56801, n56802 );
nand U135378 ( n56802, n56803, n76282 );
nand U135379 ( n56801, P2_P2_EAX_REG_19_, n56762 );
nor U135380 ( n56803, P2_P2_EAX_REG_19_, n56717 );
nand U135381 ( n56892, n56893, n56894 );
nand U135382 ( n56894, n56895, n76282 );
nand U135383 ( n56893, P2_P2_EAX_REG_17_, n56851 );
nor U135384 ( n56895, P2_P2_EAX_REG_17_, n56806 );
nand U135385 ( n23678, n23679, n23680 );
nand U135386 ( n23680, n23681, n76540 );
nand U135387 ( n23679, P1_P2_EAX_REG_19_, n23640 );
nor U135388 ( n23681, P1_P2_EAX_REG_19_, n23595 );
nand U135389 ( n23589, n23590, n23591 );
nand U135390 ( n23591, n23592, n76540 );
nand U135391 ( n23590, P1_P2_EAX_REG_21_, n23551 );
nor U135392 ( n23592, P1_P2_EAX_REG_21_, n23451 );
nand U135393 ( n23767, n23768, n23769 );
nand U135394 ( n23769, n23770, n76540 );
nand U135395 ( n23768, P1_P2_EAX_REG_17_, n23729 );
nor U135396 ( n23770, P1_P2_EAX_REG_17_, n23684 );
nand U135397 ( n31066, n31067, n31068 );
nand U135398 ( n31068, n31069, n76483 );
nand U135399 ( n31067, P1_P3_EAX_REG_17_, n31030 );
nor U135400 ( n31069, P1_P3_EAX_REG_17_, n30987 );
nand U135401 ( n30896, n30897, n30898 );
nand U135402 ( n30898, n30899, n76483 );
nand U135403 ( n30897, P1_P3_EAX_REG_21_, n30860 );
nor U135404 ( n30899, P1_P3_EAX_REG_21_, n30762 );
nand U135405 ( n65098, n65099, n65100 );
nand U135406 ( n65100, n65101, n76216 );
nand U135407 ( n65099, P2_P3_EAX_REG_21_, n65062 );
nor U135408 ( n65101, P2_P3_EAX_REG_21_, n64964 );
nand U135409 ( n65183, n65184, n65185 );
nand U135410 ( n65185, n65186, n76216 );
nand U135411 ( n65184, P2_P3_EAX_REG_19_, n65147 );
nor U135412 ( n65186, P2_P3_EAX_REG_19_, n65104 );
nand U135413 ( n30981, n30982, n30983 );
nand U135414 ( n30983, n30984, n76483 );
nand U135415 ( n30982, P1_P3_EAX_REG_19_, n30945 );
nor U135416 ( n30984, P1_P3_EAX_REG_19_, n30902 );
nand U135417 ( n65268, n65269, n65270 );
nand U135418 ( n65270, n65271, n76216 );
nand U135419 ( n65269, P2_P3_EAX_REG_17_, n65232 );
nor U135420 ( n65271, P2_P3_EAX_REG_17_, n65189 );
nand U135421 ( n16774, n17054, P4_DATAO_REG_7_ );
nand U135422 ( n56472, n56473, n56474 );
nand U135423 ( n56474, n56475, n76282 );
nand U135424 ( n56473, P2_P2_EAX_REG_25_, n56431 );
nor U135425 ( n56475, P2_P2_EAX_REG_25_, n56383 );
nand U135426 ( n56567, n56568, n56569 );
nand U135427 ( n56569, n56570, n76282 );
nand U135428 ( n56568, P2_P2_EAX_REG_23_, n56526 );
nor U135429 ( n56570, P2_P2_EAX_REG_23_, n56478 );
nand U135430 ( n23445, n23446, n23447 );
nand U135431 ( n23447, n23448, n76540 );
nand U135432 ( n23446, P1_P2_EAX_REG_23_, n23404 );
nor U135433 ( n23448, P1_P2_EAX_REG_23_, n23354 );
nand U135434 ( n23348, n23349, n23350 );
nand U135435 ( n23350, n23351, n76540 );
nand U135436 ( n23349, P1_P2_EAX_REG_25_, n23307 );
nor U135437 ( n23351, P1_P2_EAX_REG_25_, n23259 );
nand U135438 ( n30663, n30664, n30665 );
nand U135439 ( n30665, n30666, n76483 );
nand U135440 ( n30664, P1_P3_EAX_REG_25_, n30625 );
nor U135441 ( n30666, P1_P3_EAX_REG_25_, n30580 );
nand U135442 ( n30756, n30757, n30758 );
nand U135443 ( n30758, n30759, n76483 );
nand U135444 ( n30757, P1_P3_EAX_REG_23_, n30714 );
nor U135445 ( n30759, P1_P3_EAX_REG_23_, n30669 );
nand U135446 ( n64869, n64870, n64871 );
nand U135447 ( n64871, n64872, n76216 );
nand U135448 ( n64870, P2_P3_EAX_REG_25_, n64831 );
nor U135449 ( n64872, P2_P3_EAX_REG_25_, n64739 );
nand U135450 ( n64958, n64959, n64960 );
nand U135451 ( n64960, n64961, n76216 );
nand U135452 ( n64959, P2_P3_EAX_REG_23_, n64920 );
nor U135453 ( n64961, P2_P3_EAX_REG_23_, n64875 );
nor U135454 ( n43042, P2_P1_REIP_REG_11_, n504 );
nor U135455 ( n43198, P2_P1_REIP_REG_5_, n504 );
nand U135456 ( n43003, n43004, n43005 );
nand U135457 ( n43004, n7393, P2_P1_PHYADDRPOINTER_REG_13_ );
nand U135458 ( n43005, P2_P1_REIP_REG_13_, n43006 );
nand U135459 ( n43006, n43007, n43008 );
nand U135460 ( n43159, n43160, n43161 );
nand U135461 ( n43160, n7393, P2_P1_PHYADDRPOINTER_REG_7_ );
nand U135462 ( n43161, P2_P1_REIP_REG_7_, n43162 );
nand U135463 ( n43162, n43163, n43164 );
nor U135464 ( n43292, P2_P1_REIP_REG_2_, n504 );
nand U135465 ( n12284, P1_P1_PHYADDRPOINTER_REG_13_, P1_P1_PHYADDRPOINTER_REG_12_ );
nand U135466 ( n43259, n43290, P2_P1_REIP_REG_2_ );
nor U135467 ( n43290, n504, n72962 );
nor U135468 ( n43258, n43259, n43260 );
nand U135469 ( n43260, P2_P1_REIP_REG_3_, n74672 );
and U135470 ( n63639, n63725, P2_P3_REIP_REG_11_ );
nor U135471 ( n63725, n478, n63628 );
and U135472 ( n63856, n63881, P2_P3_REIP_REG_5_ );
nor U135473 ( n63881, n478, n63845 );
and U135474 ( n29740, n29765, P1_P3_REIP_REG_11_ );
nor U135475 ( n29765, n207, n29729 );
and U135476 ( n29900, n29925, P1_P3_REIP_REG_5_ );
nor U135477 ( n29925, n207, n29889 );
and U135478 ( n22419, n22444, P1_P2_REIP_REG_11_ );
nor U135479 ( n22444, n173, n22408 );
and U135480 ( n22577, n22602, P1_P2_REIP_REG_5_ );
nor U135481 ( n22602, n173, n22566 );
and U135482 ( n55534, n55559, P2_P2_REIP_REG_11_ );
nor U135483 ( n55559, n445, n55520 );
and U135484 ( n55690, n55715, P2_P2_REIP_REG_5_ );
nor U135485 ( n55715, n445, n55679 );
nor U135486 ( n43112, P2_P1_REIP_REG_8_, n504 );
nand U135487 ( n43092, P2_P1_REIP_REG_10_, n43093 );
nand U135488 ( n43093, n43094, n43095 );
nand U135489 ( n43095, n76102, n73221 );
nor U135490 ( n9038, P1_P1_REIP_REG_11_, n233 );
nor U135491 ( n9233, P1_P1_REIP_REG_5_, n233 );
nand U135492 ( n8989, n8990, n8992 );
nand U135493 ( n8990, n4751, P1_P1_PHYADDRPOINTER_REG_13_ );
nand U135494 ( n8992, P1_P1_REIP_REG_13_, n8993 );
nand U135495 ( n8993, n8994, n8995 );
nand U135496 ( n9184, n9185, n9187 );
nand U135497 ( n9185, n4751, P1_P1_PHYADDRPOINTER_REG_7_ );
nand U135498 ( n9187, P1_P1_REIP_REG_7_, n9188 );
nand U135499 ( n9188, n9189, n9190 );
nor U135500 ( n9333, P1_P1_REIP_REG_2_, n233 );
and U135501 ( n63785, n63816, P2_P3_REIP_REG_8_ );
nor U135502 ( n63816, n478, n63758 );
and U135503 ( n29825, n29860, P1_P3_REIP_REG_8_ );
nor U135504 ( n29860, n207, n29798 );
and U135505 ( n22506, n22537, P1_P2_REIP_REG_8_ );
nor U135506 ( n22537, n173, n22477 );
and U135507 ( n55619, n55650, P2_P2_REIP_REG_8_ );
nor U135508 ( n55650, n445, n55592 );
nand U135509 ( n63767, n63783, n63481 );
nand U135510 ( n63783, n63784, n63785 );
nor U135511 ( n63784, P2_P3_REIP_REG_10_, n73216 );
nand U135512 ( n29807, n29823, n29582 );
nand U135513 ( n29823, n29824, n29825 );
nor U135514 ( n29824, P1_P3_REIP_REG_10_, n73217 );
nand U135515 ( n22488, n22504, n22261 );
nand U135516 ( n22504, n22505, n22506 );
nor U135517 ( n22505, P1_P2_REIP_REG_10_, n73215 );
nand U135518 ( n55601, n55617, n55373 );
nand U135519 ( n55617, n55618, n55619 );
nor U135520 ( n55618, P2_P2_REIP_REG_10_, n73214 );
nand U135521 ( n63637, n63638, n63639 );
nor U135522 ( n63638, P2_P3_REIP_REG_13_, n74800 );
nand U135523 ( n63854, n63855, n63856 );
nor U135524 ( n63855, P2_P3_REIP_REG_7_, n74711 );
nand U135525 ( n29738, n29739, n29740 );
nor U135526 ( n29739, P1_P3_REIP_REG_13_, n74801 );
nand U135527 ( n29898, n29899, n29900 );
nor U135528 ( n29899, P1_P3_REIP_REG_7_, n74712 );
nand U135529 ( n22417, n22418, n22419 );
nor U135530 ( n22418, P1_P2_REIP_REG_13_, n74799 );
nand U135531 ( n22575, n22576, n22577 );
nor U135532 ( n22576, P1_P2_REIP_REG_7_, n74710 );
nand U135533 ( n55532, n55533, n55534 );
nor U135534 ( n55533, P2_P2_REIP_REG_13_, n74798 );
nand U135535 ( n55688, n55689, n55690 );
nor U135536 ( n55689, P2_P2_REIP_REG_7_, n74709 );
nand U135537 ( n45965, P2_P1_PHYADDRPOINTER_REG_13_, P2_P1_PHYADDRPOINTER_REG_12_ );
nor U135538 ( n42571, n42608, n42609 );
nor U135539 ( n42609, n504, P2_P1_REIP_REG_26_ );
nor U135540 ( n42838, n42872, n42873 );
nor U135541 ( n42873, n504, P2_P1_REIP_REG_17_ );
nor U135542 ( n42753, n42790, n42791 );
nor U135543 ( n42791, n504, P2_P1_REIP_REG_20_ );
nand U135544 ( n42834, n42835, n42836 );
nand U135545 ( n42835, n7393, P2_P1_PHYADDRPOINTER_REG_19_ );
nand U135546 ( n42836, P2_P1_REIP_REG_19_, n42837 );
nand U135547 ( n42837, n42838, n42839 );
nor U135548 ( n42662, n42695, n42696 );
nor U135549 ( n42696, n504, P2_P1_REIP_REG_23_ );
and U135550 ( n57266, n57228, P2_P2_EAX_REG_9_ );
and U135551 ( n24144, n24106, P1_P2_EAX_REG_9_ );
and U135552 ( n31438, n31400, P1_P3_EAX_REG_9_ );
and U135553 ( n65688, n65650, P2_P3_EAX_REG_9_ );
and U135554 ( n31276, n31234, P1_P3_EAX_REG_13_ );
and U135555 ( n31357, n31319, P1_P3_EAX_REG_11_ );
and U135556 ( n23982, n23944, P1_P2_EAX_REG_13_ );
and U135557 ( n24063, n24025, P1_P2_EAX_REG_11_ );
and U135558 ( n65526, n65488, P2_P3_EAX_REG_13_ );
and U135559 ( n65607, n65569, P2_P3_EAX_REG_11_ );
and U135560 ( n57104, n57066, P2_P2_EAX_REG_13_ );
and U135561 ( n57185, n57147, P2_P2_EAX_REG_11_ );
and U135562 ( n57367, n57309, P2_P2_EAX_REG_7_ );
and U135563 ( n57388, n57380, P2_P2_EAX_REG_5_ );
and U135564 ( n57409, n57401, P2_P2_EAX_REG_3_ );
and U135565 ( n24242, n24187, P1_P2_EAX_REG_7_ );
and U135566 ( n24263, n24255, P1_P2_EAX_REG_5_ );
and U135567 ( n24286, n24278, P1_P2_EAX_REG_3_ );
and U135568 ( n31536, n31481, P1_P3_EAX_REG_7_ );
and U135569 ( n31557, n31549, P1_P3_EAX_REG_5_ );
and U135570 ( n31582, n31570, P1_P3_EAX_REG_3_ );
and U135571 ( n65786, n65731, P2_P3_EAX_REG_7_ );
and U135572 ( n65847, n65839, P2_P3_EAX_REG_5_ );
and U135573 ( n65868, n65860, P2_P3_EAX_REG_3_ );
nand U135574 ( n9292, n9330, P1_P1_REIP_REG_2_ );
nor U135575 ( n9330, n233, n72963 );
nor U135576 ( n9290, n9292, n9293 );
nand U135577 ( n9293, P1_P1_REIP_REG_3_, n74673 );
and U135578 ( n57429, n57421, P2_P2_EAX_REG_1_ );
and U135579 ( n24306, n24298, P1_P2_EAX_REG_1_ );
and U135580 ( n31602, n31594, P1_P3_EAX_REG_1_ );
and U135581 ( n65888, n65880, P2_P3_EAX_REG_1_ );
nor U135582 ( n9125, P1_P1_REIP_REG_8_, n233 );
nand U135583 ( n9100, P1_P1_REIP_REG_10_, n9102 );
nand U135584 ( n9102, n9103, n9104 );
nand U135585 ( n9104, n76172, n73222 );
nand U135586 ( n31830, n32577, P1_P3_STATE2_REG_1_ );
nor U135587 ( n32577, P1_P3_STATEBS16_REG, n3063 );
nor U135588 ( n42924, n42940, n42941 );
nor U135589 ( n42941, n504, P2_P1_REIP_REG_14_ );
nand U135590 ( n42922, P2_P1_REIP_REG_16_, n42923 );
nand U135591 ( n42923, n42924, n42925 );
nand U135592 ( n42925, n76102, n74868 );
nand U135593 ( n24616, n25335, P1_P2_STATE2_REG_1_ );
nor U135594 ( n25335, P1_P2_STATEBS16_REG, n3907 );
nand U135595 ( n45529, n46281, P2_P1_STATE2_REG_1_ );
nor U135596 ( n46281, P2_P1_STATEBS16_REG, n7438 );
nand U135597 ( n66453, n67342, P2_P3_STATE2_REG_1_ );
nor U135598 ( n67342, P2_P3_STATEBS16_REG, n5664 );
nand U135599 ( n57748, n58474, P2_P2_STATE2_REG_1_ );
nor U135600 ( n58474, P2_P2_STATEBS16_REG, n6539 );
nor U135601 ( n8502, n8548, n8549 );
nor U135602 ( n8549, n233, P1_P1_REIP_REG_26_ );
nor U135603 ( n8694, n8740, n8742 );
nor U135604 ( n8742, n233, P1_P1_REIP_REG_20_ );
nor U135605 ( n8800, n8843, n8844 );
nor U135606 ( n8844, n233, P1_P1_REIP_REG_17_ );
nand U135607 ( n8795, n8797, n8798 );
nand U135608 ( n8797, n4751, P1_P1_PHYADDRPOINTER_REG_19_ );
nand U135609 ( n8798, P1_P1_REIP_REG_19_, n8799 );
nand U135610 ( n8799, n8800, n8802 );
nor U135611 ( n8615, n8627, n8628 );
nor U135612 ( n8628, n233, P1_P1_REIP_REG_23_ );
nand U135613 ( n22227, n22228, n22229 );
nand U135614 ( n22228, P1_P2_REIP_REG_20_, n22220 );
nand U135615 ( n22229, n22189, n74926 );
nand U135616 ( n55339, n55340, n55341 );
nand U135617 ( n55340, P2_P2_REIP_REG_20_, n55334 );
nand U135618 ( n55341, n55303, n74925 );
nand U135619 ( n63447, n63448, n63449 );
nand U135620 ( n63448, P2_P3_REIP_REG_20_, n63368 );
nand U135621 ( n63449, n63337, n74928 );
nand U135622 ( n29544, n29545, n29546 );
nand U135623 ( n29545, P1_P3_REIP_REG_20_, n29539 );
nand U135624 ( n29546, n29508, n74929 );
nand U135625 ( n22164, n22165, n22166 );
nand U135626 ( n22165, P1_P2_REIP_REG_23_, n22129 );
nand U135627 ( n22166, n22111, n74970 );
nand U135628 ( n55278, n55279, n55280 );
nand U135629 ( n55279, P2_P2_REIP_REG_23_, n55239 );
nand U135630 ( n55280, n55221, n74969 );
nand U135631 ( n63246, n63247, n63248 );
nand U135632 ( n63247, P2_P3_REIP_REG_23_, n63211 );
nand U135633 ( n63248, n63193, n74987 );
nand U135634 ( n29483, n29484, n29485 );
nand U135635 ( n29484, P1_P3_REIP_REG_23_, n29448 );
nand U135636 ( n29485, n29430, n74988 );
nor U135637 ( n8908, n8928, n8929 );
nor U135638 ( n8929, n233, P1_P1_REIP_REG_14_ );
nand U135639 ( n63586, n63587, n63568 );
nor U135640 ( n63587, P2_P3_REIP_REG_15_, n74830 );
nand U135641 ( n29687, n29688, n29669 );
nor U135642 ( n29688, P1_P3_REIP_REG_15_, n74829 );
nand U135643 ( n22366, n22367, n22348 );
nor U135644 ( n22367, P1_P2_REIP_REG_15_, n74828 );
nand U135645 ( n55478, n55479, n55460 );
nor U135646 ( n55479, P2_P2_REIP_REG_15_, n74827 );
nand U135647 ( n8905, P1_P1_REIP_REG_16_, n8907 );
nand U135648 ( n8907, n8908, n8909 );
nand U135649 ( n8909, n76172, n74869 );
xnor U135650 ( n28643, n73055, P1_P2_INSTQUEUEWR_ADDR_REG_1_ );
xnor U135651 ( n61948, n73054, P2_P2_INSTQUEUEWR_ADDR_REG_1_ );
xnor U135652 ( n70548, n73053, P2_P3_INSTQUEUEWR_ADDR_REG_1_ );
xnor U135653 ( n35822, n73059, P1_P3_INSTQUEUEWR_ADDR_REG_1_ );
nand U135654 ( n12713, P1_P1_INSTADDRPOINTER_REG_31_, n76606 );
or U135655 ( n43283, n75960, n75961 );
nor U135656 ( n75960, n72964, n43247 );
nor U135657 ( n75961, n43259, P2_P1_REIP_REG_3_ );
nand U135658 ( n42691, n42692, n42693 );
nand U135659 ( n42693, n42694, n42653 );
or U135660 ( n42692, n75005, n42662 );
nor U135661 ( n42694, P2_P1_REIP_REG_24_, n74995 );
nand U135662 ( n42937, n42938, n42939 );
nand U135663 ( n42938, n7393, P2_P1_PHYADDRPOINTER_REG_15_ );
or U135664 ( n42939, n74868, n42924 );
nor U135665 ( n24102, n24107, n24108 );
nand U135666 ( n24107, n4525, n74633 );
nand U135667 ( n24108, n76541, P1_P2_EAX_REG_9_ );
nor U135668 ( n57224, n57229, n57230 );
nand U135669 ( n57229, n7158, n74632 );
nand U135670 ( n57230, n76283, P2_P2_EAX_REG_9_ );
nor U135671 ( n31396, n31401, n31402 );
nand U135672 ( n31401, n3638, n74629 );
nand U135673 ( n31402, n76484, P1_P3_EAX_REG_9_ );
nor U135674 ( n65646, n65651, n65652 );
nand U135675 ( n65651, n6265, n74628 );
nand U135676 ( n65652, n76217, P2_P3_EAX_REG_9_ );
nor U135677 ( n24021, n24026, n24027 );
nand U135678 ( n24026, n4527, n75274 );
nand U135679 ( n24027, n76541, P1_P2_EAX_REG_11_ );
nor U135680 ( n23940, n23945, n23946 );
nand U135681 ( n23945, n4528, n75273 );
nand U135682 ( n23946, n76541, P1_P2_EAX_REG_13_ );
nor U135683 ( n24183, n24188, n24189 );
nand U135684 ( n24188, n4524, n75275 );
nand U135685 ( n24189, n76541, P1_P2_EAX_REG_7_ );
nor U135686 ( n24251, n24256, n24257 );
nand U135687 ( n24256, n4523, n75277 );
nand U135688 ( n24257, n76541, P1_P2_EAX_REG_5_ );
nor U135689 ( n24274, n24279, n24280 );
nand U135690 ( n24279, n4522, n75276 );
nand U135691 ( n24280, n76541, P1_P2_EAX_REG_3_ );
nor U135692 ( n31230, n31235, n31236 );
nand U135693 ( n31235, n3640, n75278 );
nand U135694 ( n31236, n76484, P1_P3_EAX_REG_13_ );
nor U135695 ( n31315, n31320, n31321 );
nand U135696 ( n31320, n3639, n75280 );
nand U135697 ( n31321, n76484, P1_P3_EAX_REG_11_ );
nor U135698 ( n65484, n65489, n65490 );
nand U135699 ( n65489, n6268, n75268 );
nand U135700 ( n65490, n76217, P2_P3_EAX_REG_13_ );
nor U135701 ( n65565, n65570, n65571 );
nand U135702 ( n65570, n6267, n75269 );
nand U135703 ( n65571, n76217, P2_P3_EAX_REG_11_ );
nor U135704 ( n57062, n57067, n57068 );
nand U135705 ( n57067, n7160, n75266 );
nand U135706 ( n57068, n76283, P2_P2_EAX_REG_13_ );
nor U135707 ( n57143, n57148, n57149 );
nand U135708 ( n57148, n7159, n75264 );
nand U135709 ( n57149, n76283, P2_P2_EAX_REG_11_ );
nor U135710 ( n57305, n57310, n57311 );
nand U135711 ( n57310, n7157, n75265 );
nand U135712 ( n57311, n76283, P2_P2_EAX_REG_7_ );
nor U135713 ( n57376, n57381, n57382 );
nand U135714 ( n57381, n7155, n75263 );
nand U135715 ( n57382, n76283, P2_P2_EAX_REG_5_ );
nor U135716 ( n57397, n57402, n57403 );
nand U135717 ( n57402, n7154, n75267 );
nand U135718 ( n57403, n76283, P2_P2_EAX_REG_3_ );
nor U135719 ( n31477, n31482, n31483 );
nand U135720 ( n31482, n3637, n75281 );
nand U135721 ( n31483, n76484, P1_P3_EAX_REG_7_ );
nor U135722 ( n31545, n31550, n31551 );
nand U135723 ( n31550, n3635, n75282 );
nand U135724 ( n31551, n76484, P1_P3_EAX_REG_5_ );
nor U135725 ( n31566, n31571, n31572 );
nand U135726 ( n31571, n3634, n75279 );
nand U135727 ( n31572, n76484, P1_P3_EAX_REG_3_ );
nor U135728 ( n65727, n65732, n65733 );
nand U135729 ( n65732, n6264, n75271 );
nand U135730 ( n65733, n76217, P2_P3_EAX_REG_7_ );
nor U135731 ( n65835, n65840, n65841 );
nand U135732 ( n65840, n6263, n75270 );
nand U135733 ( n65841, n76217, P2_P3_EAX_REG_5_ );
nor U135734 ( n65856, n65861, n65862 );
nand U135735 ( n65861, n6262, n75272 );
nand U135736 ( n65862, n76217, P2_P3_EAX_REG_3_ );
nand U135737 ( n11758, n12665, P1_P1_STATE2_REG_1_ );
nor U135738 ( n12665, P1_P1_STATEBS16_REG, n4794 );
nor U135739 ( n24294, n24299, n24300 );
nand U135740 ( n24299, P1_P2_EAX_REG_0_, n75285 );
nand U135741 ( n24300, n76540, P1_P2_EAX_REG_1_ );
nor U135742 ( n57417, n57422, n57423 );
nand U135743 ( n57422, P2_P2_EAX_REG_0_, n75283 );
nand U135744 ( n57423, n76282, P2_P2_EAX_REG_1_ );
nor U135745 ( n31590, n31595, n31596 );
nand U135746 ( n31595, P1_P3_EAX_REG_0_, n75286 );
nand U135747 ( n31596, n76483, P1_P3_EAX_REG_1_ );
nor U135748 ( n65876, n65881, n65882 );
nand U135749 ( n65881, P2_P3_EAX_REG_0_, n75284 );
nand U135750 ( n65882, n76216, P2_P3_EAX_REG_1_ );
nand U135751 ( n45916, n45917, n45918 );
nor U135752 ( n45918, P2_P1_PHYADDRPOINTER_REG_17_, n45896 );
nor U135753 ( n45917, n45919, n45567 );
nand U135754 ( n66867, n66868, n66869 );
nor U135755 ( n66869, P2_P3_PHYADDRPOINTER_REG_17_, n66847 );
nor U135756 ( n66868, n66870, n66492 );
nand U135757 ( n24991, n24992, n24993 );
nor U135758 ( n24993, P1_P2_PHYADDRPOINTER_REG_17_, n24971 );
nor U135759 ( n24992, n24994, n24655 );
nand U135760 ( n58126, n58127, n58128 );
nor U135761 ( n58128, P2_P2_PHYADDRPOINTER_REG_17_, n58106 );
nor U135762 ( n58127, n58129, n57791 );
or U135763 ( n9322, n75962, n75963 );
nor U135764 ( n75962, n72965, n9277 );
nor U135765 ( n75963, n9292, P1_P1_REIP_REG_3_ );
nand U135766 ( n8622, n8623, n8624 );
nand U135767 ( n8624, n8625, n8604 );
or U135768 ( n8623, n75006, n8615 );
nor U135769 ( n8625, P1_P1_REIP_REG_24_, n74996 );
nand U135770 ( n8924, n8925, n8927 );
nand U135771 ( n8925, n4751, P1_P1_PHYADDRPOINTER_REG_15_ );
or U135772 ( n8927, n74869, n8908 );
nand U135773 ( n8442, n8443, n8444 );
nand U135774 ( n8443, P1_P1_REIP_REG_30_, n8418 );
nand U135775 ( n8444, n8445, n8402 );
nand U135776 ( n42897, n42913, n42829 );
nand U135777 ( n42913, n42914, n42915 );
nor U135778 ( n42915, P2_P1_REIP_REG_16_, n74860 );
and U135779 ( n42914, P2_P1_REIP_REG_15_, n42916 );
nand U135780 ( n42828, n42830, n42831 );
nor U135781 ( n42831, P2_P1_REIP_REG_19_, n74904 );
and U135782 ( n42830, P2_P1_REIP_REG_18_, n42832 );
and U135783 ( n42651, P2_P1_REIP_REG_24_, n42653 );
and U135784 ( n42757, P2_P1_REIP_REG_21_, n42759 );
nand U135785 ( n8453, n8472, n8473 );
nand U135786 ( n8473, n8430, n8474 );
nand U135787 ( n8472, n8445, n8477 );
nand U135788 ( n8474, P1_P1_EBX_REG_29_, n8475 );
nand U135789 ( n8874, n8894, n8789 );
nand U135790 ( n8894, n8895, n8897 );
nor U135791 ( n8897, P1_P1_REIP_REG_16_, n74861 );
and U135792 ( n8895, P1_P1_REIP_REG_15_, n8898 );
nand U135793 ( n8788, n8790, n8792 );
nor U135794 ( n8792, P1_P1_REIP_REG_19_, n74905 );
and U135795 ( n8790, P1_P1_REIP_REG_18_, n8793 );
and U135796 ( n8699, P1_P1_REIP_REG_21_, n8702 );
and U135797 ( n8602, P1_P1_REIP_REG_24_, n8604 );
nand U135798 ( n12870, n12872, n12817 );
nor U135799 ( n12872, n12873, n12874 );
nor U135800 ( n12873, P1_P1_INSTADDRPOINTER_REG_26_, n4832 );
nor U135801 ( n12874, P1_P1_INSTADDRPOINTER_REG_27_, n4827 );
and U135802 ( n43001, n43026, P2_P1_REIP_REG_11_ );
nor U135803 ( n43026, n504, n42990 );
and U135804 ( n43157, n43182, P2_P1_REIP_REG_5_ );
nor U135805 ( n43182, n504, n43146 );
nand U135806 ( n43068, n43084, n42829 );
nand U135807 ( n43084, n43085, n43086 );
nor U135808 ( n43085, P2_P1_REIP_REG_10_, n73221 );
nand U135809 ( n42999, n43000, n43001 );
nor U135810 ( n43000, P2_P1_REIP_REG_13_, n74815 );
nand U135811 ( n43155, n43156, n43157 );
nor U135812 ( n43156, P2_P1_REIP_REG_7_, n74728 );
nor U135813 ( n43086, n75964, n75965 );
or U135814 ( n75964, n504, n43059 );
nand U135815 ( n63038, n63039, n63040 );
nand U135816 ( n63039, P2_P3_PHYADDRPOINTER_REG_31_, n5629 );
nand U135817 ( n63040, n474, P2_P3_EBX_REG_31_ );
nand U135818 ( n29271, n29272, n29273 );
nand U135819 ( n29272, P1_P3_PHYADDRPOINTER_REG_31_, n3028 );
nand U135820 ( n29273, n203, P1_P3_EBX_REG_31_ );
nand U135821 ( n21954, n21955, n21956 );
nand U135822 ( n21955, P1_P2_PHYADDRPOINTER_REG_31_, n3872 );
nand U135823 ( n21956, n169, P1_P2_EBX_REG_31_ );
nand U135824 ( n55066, n55067, n55068 );
nand U135825 ( n55067, P2_P2_PHYADDRPOINTER_REG_31_, n6504 );
nand U135826 ( n55068, n442, P2_P2_EBX_REG_31_ );
nor U135827 ( n42498, n42501, n75328 );
nor U135828 ( n42501, n42502, n42503 );
nor U135829 ( n42502, P2_P1_REIP_REG_30_, n504 );
nand U135830 ( n8826, n13950, n13952 );
nand U135831 ( n13952, n76888, P1_P1_INSTADDRPOINTER_REG_6_ );
nor U135832 ( n13950, n13953, n13954 );
nor U135833 ( n13954, n74729, n76598 );
xor U135834 ( n37856, n37857, n37858 );
xor U135835 ( n37858, n37855, P4_REG2_REG_9_ );
and U135836 ( n8987, n9018, P1_P1_REIP_REG_11_ );
nor U135837 ( n9018, n233, n8973 );
and U135838 ( n9182, n9213, P1_P1_REIP_REG_5_ );
nor U135839 ( n9213, n233, n9168 );
nand U135840 ( n15561, n47316, n47317 );
nand U135841 ( n47317, n76861, P2_P1_INSTADDRPOINTER_REG_6_ );
nor U135842 ( n47316, n47318, n47319 );
nor U135843 ( n47319, n74728, n76332 );
xor U135844 ( n42581, n45606, P2_P1_PHYADDRPOINTER_REG_28_ );
nand U135845 ( n16769, n8212, P4_DATAO_REG_6_ );
nand U135846 ( n9070, n9090, n8789 );
nand U135847 ( n9090, n9092, n9093 );
nor U135848 ( n9092, P1_P1_REIP_REG_10_, n73222 );
nand U135849 ( n8984, n8985, n8987 );
nor U135850 ( n8985, P1_P1_REIP_REG_13_, n74816 );
nand U135851 ( n9179, n9180, n9182 );
nor U135852 ( n9180, P1_P1_REIP_REG_7_, n74729 );
nor U135853 ( n9093, n75966, n75967 );
or U135854 ( n75966, n233, n9059 );
nor U135855 ( n8412, n8415, n75329 );
nor U135856 ( n8415, n8417, n8418 );
nor U135857 ( n8417, P1_P1_REIP_REG_30_, n233 );
nand U135858 ( n42795, n42796, n42797 );
nand U135859 ( n42796, P2_P1_REIP_REG_20_, n42790 );
nand U135860 ( n42797, n42759, n74951 );
nor U135861 ( n12727, n12728, n12729 );
nor U135862 ( n12728, P1_P1_INSTADDRPOINTER_REG_30_, n12730 );
nor U135863 ( n12730, n12732, n12733 );
nand U135864 ( n42730, n42731, n42732 );
nand U135865 ( n42731, P2_P1_REIP_REG_23_, n42695 );
nand U135866 ( n42732, n42653, n74995 );
nand U135867 ( n42934, n42935, n42916 );
nor U135868 ( n42935, P2_P1_REIP_REG_15_, n74860 );
nand U135869 ( n17080, DIN_28_, n76928 );
nor U135870 ( n46327, n46328, n46329 );
nor U135871 ( n46328, P2_P1_INSTADDRPOINTER_REG_30_, n46330 );
nor U135872 ( n46330, n46331, n46332 );
nand U135873 ( n8747, n8748, n8749 );
nand U135874 ( n8748, P1_P1_REIP_REG_20_, n8740 );
nand U135875 ( n8749, n8702, n74952 );
nand U135876 ( n43232, n43451, n43452 );
nand U135877 ( n43451, n42959, n42957 );
nand U135878 ( n43452, P3_REG1_REG_8_, n43453 );
nand U135879 ( n43453, n890, n887 );
not U135880 ( n76913, P2_P2_STATE2_REG_3_ );
not U135881 ( n76917, P1_P2_STATE2_REG_3_ );
not U135882 ( n76919, P1_P3_STATE2_REG_3_ );
not U135883 ( n76915, P2_P3_STATE2_REG_3_ );
xor U135884 ( n43667, n43668, n43669 );
xor U135885 ( n43669, n43666, P3_REG1_REG_12_ );
nand U135886 ( n12187, P1_P1_PHYADDRPOINTER_REG_16_, P1_P1_PHYADDRPOINTER_REG_15_ );
nand U135887 ( n8670, n8672, n8673 );
nand U135888 ( n8672, P1_P1_REIP_REG_23_, n8627 );
nand U135889 ( n8673, n8604, n74996 );
nand U135890 ( n8920, n8922, n8898 );
nor U135891 ( n8922, P1_P1_REIP_REG_15_, n74861 );
nand U135892 ( n43449, n43450, n43448 );
nand U135893 ( n43450, P3_REG1_REG_9_, n43446 );
and U135894 ( n49682, DIN_31_, n76929 );
xor U135895 ( n42627, n45650, P2_P1_PHYADDRPOINTER_REG_26_ );
nand U135896 ( n42424, P3_REG2_REG_6_, n45184 );
nand U135897 ( n45896, P2_P1_PHYADDRPOINTER_REG_16_, P2_P1_PHYADDRPOINTER_REG_15_ );
xor U135898 ( n8514, n11830, P1_P1_PHYADDRPOINTER_REG_28_ );
nand U135899 ( n42432, P3_REG1_REG_6_, n45184 );
nand U135900 ( n43228, n43438, n43439 );
nand U135901 ( n43438, n42955, n42957 );
nand U135902 ( n43439, P3_REG2_REG_8_, n43440 );
nand U135903 ( n43440, n892, n887 );
xnor U135904 ( n21335, n21609, n21610 );
xor U135905 ( n21610, P1_P1_INSTQUEUEWR_ADDR_REG_2_, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
xor U135906 ( n42702, n45717, P2_P1_PHYADDRPOINTER_REG_24_ );
nor U135907 ( n43429, n879, n43436 );
not U135908 ( n879, n43431 );
nand U135909 ( n43436, n43437, n43435 );
nand U135910 ( n43437, P3_REG2_REG_9_, n43433 );
nand U135911 ( n63620, n63621, n63622 );
nand U135912 ( n63621, P2_P3_PHYADDRPOINTER_REG_14_, n5629 );
nand U135913 ( n63622, n5630, n63615 );
nand U135914 ( n63837, n63838, n63839 );
nand U135915 ( n63838, P2_P3_PHYADDRPOINTER_REG_8_, n5629 );
nand U135916 ( n63839, n5630, n6158 );
nand U135917 ( n63947, n63948, n63949 );
nand U135918 ( n63948, P2_P3_PHYADDRPOINTER_REG_4_, n5629 );
nand U135919 ( n63949, n5630, n6155 );
nand U135920 ( n64057, n64058, n64059 );
nand U135921 ( n64058, P2_P3_PHYADDRPOINTER_REG_2_, n5629 );
nand U135922 ( n64059, n5630, n64055 );
nand U135923 ( n29721, n29722, n29723 );
nand U135924 ( n29722, P1_P3_PHYADDRPOINTER_REG_14_, n3028 );
nand U135925 ( n29723, n3029, n29716 );
nand U135926 ( n29881, n29882, n29883 );
nand U135927 ( n29882, P1_P3_PHYADDRPOINTER_REG_8_, n3028 );
nand U135928 ( n29883, n3029, n3543 );
nand U135929 ( n29991, n29992, n29993 );
nand U135930 ( n29992, P1_P3_PHYADDRPOINTER_REG_4_, n3028 );
nand U135931 ( n29993, n3029, n3540 );
nand U135932 ( n30040, n30041, n30042 );
nand U135933 ( n30041, P1_P3_PHYADDRPOINTER_REG_2_, n3028 );
nand U135934 ( n30042, n3029, n30038 );
nand U135935 ( n22400, n22401, n22402 );
nand U135936 ( n22401, P1_P2_PHYADDRPOINTER_REG_14_, n3872 );
nand U135937 ( n22402, n3873, n22395 );
nand U135938 ( n22558, n22559, n22560 );
nand U135939 ( n22559, P1_P2_PHYADDRPOINTER_REG_8_, n3872 );
nand U135940 ( n22560, n3873, n4380 );
nand U135941 ( n22668, n22669, n22670 );
nand U135942 ( n22669, P1_P2_PHYADDRPOINTER_REG_4_, n3872 );
nand U135943 ( n22670, n3873, n4378 );
nand U135944 ( n22717, n22718, n22719 );
nand U135945 ( n22718, P1_P2_PHYADDRPOINTER_REG_2_, n3872 );
nand U135946 ( n22719, n3873, n22715 );
nand U135947 ( n55512, n55513, n55514 );
nand U135948 ( n55513, P2_P2_PHYADDRPOINTER_REG_14_, n6504 );
nand U135949 ( n55514, n6505, n55507 );
nand U135950 ( n55671, n55672, n55673 );
nand U135951 ( n55672, P2_P2_PHYADDRPOINTER_REG_8_, n6504 );
nand U135952 ( n55673, n6505, n7013 );
nand U135953 ( n55781, n55782, n55783 );
nand U135954 ( n55782, P2_P2_PHYADDRPOINTER_REG_4_, n6504 );
nand U135955 ( n55783, n6505, n7010 );
nand U135956 ( n55833, n55834, n55835 );
nand U135957 ( n55834, P2_P2_PHYADDRPOINTER_REG_2_, n6504 );
nand U135958 ( n55835, n6505, n55831 );
nand U135959 ( n926, n11514, n11515 );
nand U135960 ( n11515, n933, P3_IR_REG_25_ );
nor U135961 ( n11514, n1834, n11517 );
nor U135962 ( n11517, n11518, n76626 );
nand U135963 ( n931, n11452, n11453 );
nand U135964 ( n11453, n933, P3_IR_REG_26_ );
nor U135965 ( n11452, n1834, n11454 );
nor U135966 ( n11454, n11455, n76626 );
nand U135967 ( n22045, n22046, n22047 );
nand U135968 ( n22047, P1_P2_EBX_REG_28_, n169 );
nand U135969 ( n22046, n3873, n22040 );
nand U135970 ( n29364, n29365, n29366 );
nand U135971 ( n29366, P1_P3_EBX_REG_28_, n203 );
nand U135972 ( n29365, n3029, n29359 );
nand U135973 ( n63127, n63128, n63129 );
nand U135974 ( n63129, P2_P3_EBX_REG_28_, n474 );
nand U135975 ( n63128, n5630, n63122 );
nand U135976 ( n55155, n55156, n55157 );
nand U135977 ( n55157, P2_P2_EBX_REG_28_, n442 );
nand U135978 ( n55156, n6505, n55150 );
nand U135979 ( n63177, n63178, n63179 );
nand U135980 ( n63179, P2_P3_EBX_REG_26_, n474 );
nand U135981 ( n63178, n5630, n63167 );
nand U135982 ( n63228, n63229, n63230 );
nand U135983 ( n63230, P2_P3_EBX_REG_24_, n474 );
nand U135984 ( n63229, n5630, n63218 );
nand U135985 ( n63346, n63347, n63348 );
nand U135986 ( n63348, P2_P3_EBX_REG_22_, n474 );
nand U135987 ( n63347, n5630, n63341 );
nand U135988 ( n63469, n63470, n63471 );
nand U135989 ( n63471, P2_P3_EBX_REG_20_, n474 );
nand U135990 ( n63470, n5630, n63459 );
nand U135991 ( n29414, n29415, n29416 );
nand U135992 ( n29416, P1_P3_EBX_REG_26_, n203 );
nand U135993 ( n29415, n3029, n29404 );
nand U135994 ( n29465, n29466, n29467 );
nand U135995 ( n29467, P1_P3_EBX_REG_24_, n203 );
nand U135996 ( n29466, n3029, n29455 );
nand U135997 ( n29517, n29518, n29519 );
nand U135998 ( n29519, P1_P3_EBX_REG_22_, n203 );
nand U135999 ( n29518, n3029, n29512 );
nand U136000 ( n29566, n29567, n29568 );
nand U136001 ( n29568, P1_P3_EBX_REG_20_, n203 );
nand U136002 ( n29567, n3029, n29556 );
nand U136003 ( n22095, n22096, n22097 );
nand U136004 ( n22097, P1_P2_EBX_REG_26_, n169 );
nand U136005 ( n22096, n3873, n22085 );
nand U136006 ( n22249, n22250, n22251 );
nand U136007 ( n22251, P1_P2_EBX_REG_20_, n169 );
nand U136008 ( n22250, n3873, n22239 );
nand U136009 ( n22146, n22147, n22148 );
nand U136010 ( n22148, P1_P2_EBX_REG_24_, n169 );
nand U136011 ( n22147, n3873, n22136 );
nand U136012 ( n22198, n22199, n22200 );
nand U136013 ( n22200, P1_P2_EBX_REG_22_, n169 );
nand U136014 ( n22199, n3873, n22193 );
nand U136015 ( n55205, n55206, n55207 );
nand U136016 ( n55207, P2_P2_EBX_REG_26_, n442 );
nand U136017 ( n55206, n6505, n55195 );
nand U136018 ( n55361, n55362, n55363 );
nand U136019 ( n55363, P2_P2_EBX_REG_20_, n442 );
nand U136020 ( n55362, n6505, n55351 );
nand U136021 ( n22015, n22016, n22017 );
nand U136022 ( n22017, P1_P2_EBX_REG_29_, n169 );
nand U136023 ( n22016, n3873, n4395 );
nand U136024 ( n55256, n55257, n55258 );
nand U136025 ( n55258, P2_P2_EBX_REG_24_, n442 );
nand U136026 ( n55257, n6505, n55246 );
nand U136027 ( n55312, n55313, n55314 );
nand U136028 ( n55314, P2_P2_EBX_REG_22_, n442 );
nand U136029 ( n55313, n6505, n55307 );
nand U136030 ( n29334, n29335, n29336 );
nand U136031 ( n29336, P1_P3_EBX_REG_29_, n203 );
nand U136032 ( n29335, n3029, n3558 );
nand U136033 ( n63097, n63098, n63099 );
nand U136034 ( n63099, P2_P3_EBX_REG_29_, n474 );
nand U136035 ( n63098, n5630, n6173 );
nand U136036 ( n55125, n55126, n55127 );
nand U136037 ( n55127, P2_P2_EBX_REG_29_, n442 );
nand U136038 ( n55126, n6505, n7028 );
nand U136039 ( n2156, n40501, n40502 );
nand U136040 ( n40502, P2_P3_DATAO_REG_26_, n76039 );
nor U136041 ( n40501, n40503, n40504 );
nor U136042 ( n40504, n73505, n76393 );
nand U136043 ( n2176, n40473, n40474 );
nand U136044 ( n40474, P2_P3_DATAO_REG_30_, n76039 );
nor U136045 ( n40473, n40475, n40476 );
nor U136046 ( n40476, n75299, n76393 );
nand U136047 ( n2041, n40642, n40643 );
nand U136048 ( n40643, P2_P3_DATAO_REG_3_, n76040 );
nor U136049 ( n40642, n40644, n40645 );
nor U136050 ( n40645, n73803, n76395 );
nand U136051 ( n2031, n40653, n40654 );
nand U136052 ( n40654, P2_P3_DATAO_REG_1_, n76922 );
nor U136053 ( n40653, n40655, n40656 );
nor U136054 ( n40656, n73535, n76395 );
nand U136055 ( n2146, n40519, n40520 );
nand U136056 ( n40520, P2_P3_DATAO_REG_24_, n76039 );
nor U136057 ( n40519, n40521, n40522 );
nor U136058 ( n40522, n73050, n76393 );
nand U136059 ( n2171, n40480, n40481 );
nand U136060 ( n40481, P2_P3_DATAO_REG_29_, n76039 );
nor U136061 ( n40480, n40482, n40483 );
nor U136062 ( n40483, n73058, n76393 );
nand U136063 ( n2166, n40484, n40485 );
nand U136064 ( n40485, P2_P3_DATAO_REG_28_, n76039 );
nor U136065 ( n40484, n40486, n40487 );
nor U136066 ( n40487, n73519, n76393 );
nand U136067 ( n916, n11627, n11628 );
nand U136068 ( n11628, n933, P3_IR_REG_23_ );
nor U136069 ( n11627, n1834, n11629 );
nor U136070 ( n11629, n76625, n11630 );
nand U136071 ( n921, n11569, n11570 );
nand U136072 ( n11570, n933, P3_IR_REG_24_ );
nor U136073 ( n11569, n1834, n11572 );
nor U136074 ( n11572, n76625, n11573 );
nand U136075 ( n951, n10764, n10765 );
nand U136076 ( n10765, n933, P3_IR_REG_30_ );
nor U136077 ( n10764, n1834, n10767 );
nor U136078 ( n10767, n76625, n10769 );
nand U136079 ( n906, n12105, n12107 );
nand U136080 ( n12107, P3_IR_REG_21_, n933 );
nor U136081 ( n12105, n1834, n12108 );
nor U136082 ( n12108, n76625, n12109 );
nand U136083 ( n901, n12404, n12405 );
nand U136084 ( n12405, P3_IR_REG_20_, n933 );
nor U136085 ( n12404, n1834, n12407 );
nor U136086 ( n12407, n76626, n12408 );
nand U136087 ( n911, n11782, n11783 );
nand U136088 ( n11783, P3_IR_REG_22_, n933 );
nor U136089 ( n11782, n1834, n11784 );
nor U136090 ( n11784, n76625, n11785 );
nand U136091 ( n941, n11337, n11338 );
nand U136092 ( n11338, P3_IR_REG_28_, n933 );
nor U136093 ( n11337, n1834, n11339 );
nor U136094 ( n11339, n76626, n11340 );
nand U136095 ( n946, n11240, n11242 );
nand U136096 ( n11242, P3_IR_REG_29_, n933 );
nor U136097 ( n11240, n1834, n11243 );
nor U136098 ( n11243, n76625, n11244 );
nand U136099 ( n2091, n40583, n40584 );
nand U136100 ( n40584, P2_P3_DATAO_REG_13_, n76040 );
nor U136101 ( n40583, n40585, n40586 );
nor U136102 ( n40586, n74390, n76394 );
nand U136103 ( n2081, n40594, n40595 );
nand U136104 ( n40595, P2_P3_DATAO_REG_11_, n76040 );
nor U136105 ( n40594, n40596, n40597 );
nor U136106 ( n40597, n74335, n76394 );
nand U136107 ( n2071, n40605, n40606 );
nand U136108 ( n40606, P2_P3_DATAO_REG_9_, n76040 );
nor U136109 ( n40605, n40607, n40608 );
nor U136110 ( n40608, n74298, n76394 );
nand U136111 ( n2061, n40616, n40617 );
nand U136112 ( n40617, P2_P3_DATAO_REG_7_, n76040 );
nor U136113 ( n40616, n40618, n40619 );
nor U136114 ( n40619, n74257, n76394 );
nand U136115 ( n2051, n40631, n40632 );
nand U136116 ( n40632, P2_P3_DATAO_REG_5_, n76040 );
nor U136117 ( n40631, n40633, n40634 );
nor U136118 ( n40634, n73948, n76395 );
nand U136119 ( n2136, n40531, n40532 );
nand U136120 ( n40532, P2_P3_DATAO_REG_22_, n76039 );
nor U136121 ( n40531, n40533, n40534 );
nor U136122 ( n40534, n73047, n76393 );
nand U136123 ( n2131, n40535, n40536 );
nand U136124 ( n40536, P2_P3_DATAO_REG_21_, n76039 );
nor U136125 ( n40535, n40537, n40538 );
nor U136126 ( n40538, n73494, n76393 );
nand U136127 ( n2126, n40543, n40544 );
nand U136128 ( n40544, P2_P3_DATAO_REG_20_, n76039 );
nor U136129 ( n40543, n40545, n40546 );
nor U136130 ( n40546, n73042, n76393 );
nand U136131 ( n2121, n40548, n40549 );
nand U136132 ( n40549, P2_P3_DATAO_REG_19_, n76039 );
nor U136133 ( n40548, n40550, n40551 );
nor U136134 ( n40551, n73479, n76393 );
nand U136135 ( n2111, n40557, n40558 );
nand U136136 ( n40558, P2_P3_DATAO_REG_17_, n76040 );
nor U136137 ( n40557, n40559, n40560 );
nor U136138 ( n40560, n73495, n76394 );
nand U136139 ( n2101, n40572, n40573 );
nand U136140 ( n40573, P2_P3_DATAO_REG_15_, n76040 );
nor U136141 ( n40572, n40574, n40575 );
nor U136142 ( n40575, n74391, n76394 );
xor U136143 ( n42763, n45787, P2_P1_PHYADDRPOINTER_REG_22_ );
nand U136144 ( n886, n13645, n13647 );
nand U136145 ( n13647, P1_P3_DATAO_REG_17_, n76041 );
nor U136146 ( n13645, n13648, n13649 );
nor U136147 ( n13649, n13650, n74418 );
nand U136148 ( n876, n14773, n14774 );
nand U136149 ( n14774, P1_P3_DATAO_REG_15_, n76041 );
nor U136150 ( n14773, n14775, n14777 );
nor U136151 ( n14777, n13650, n74395 );
nand U136152 ( n866, n15079, n15080 );
nand U136153 ( n15080, P1_P3_DATAO_REG_13_, n76041 );
nor U136154 ( n15079, n15082, n15083 );
nor U136155 ( n15083, n13650, n74392 );
nand U136156 ( n856, n15343, n15344 );
nand U136157 ( n15344, P1_P3_DATAO_REG_11_, n76041 );
nor U136158 ( n15343, n15345, n15347 );
nor U136159 ( n15347, n13650, n74301 );
nand U136160 ( n846, n15614, n15615 );
nand U136161 ( n15615, P1_P3_DATAO_REG_9_, n76041 );
nor U136162 ( n15614, n15617, n15618 );
nor U136163 ( n15618, n13650, n74300 );
nand U136164 ( n836, n15868, n15869 );
nand U136165 ( n15869, P1_P3_DATAO_REG_7_, n76041 );
nor U136166 ( n15868, n15870, n15872 );
nor U136167 ( n15872, n13650, n74225 );
nand U136168 ( n826, n16137, n16138 );
nand U136169 ( n16138, P1_P3_DATAO_REG_5_, n76041 );
nor U136170 ( n16137, n16139, n16140 );
nor U136171 ( n16140, n13650, n74105 );
nand U136172 ( n2106, n40565, n40566 );
nand U136173 ( n40566, P2_P3_DATAO_REG_16_, n76040 );
nor U136174 ( n40565, n40567, n40568 );
nor U136175 ( n40568, n75417, n76394 );
nand U136176 ( n891, n13167, n13168 );
nand U136177 ( n13168, P1_P3_DATAO_REG_18_, n76041 );
nor U136178 ( n13167, n13169, n13170 );
and U136179 ( n13170, n933, P3_IR_REG_18_ );
nand U136180 ( n881, n14368, n14369 );
nand U136181 ( n14369, P1_P3_DATAO_REG_16_, n76041 );
nor U136182 ( n14368, n14370, n14372 );
and U136183 ( n14372, n933, P3_IR_REG_16_ );
nand U136184 ( n871, n14915, n14917 );
nand U136185 ( n14917, P1_P3_DATAO_REG_14_, n76041 );
nor U136186 ( n14915, n14918, n14919 );
and U136187 ( n14919, n933, P3_IR_REG_14_ );
nand U136188 ( n861, n15207, n15208 );
nand U136189 ( n15208, P1_P3_DATAO_REG_12_, n76041 );
nor U136190 ( n15207, n15209, n15210 );
and U136191 ( n15210, n933, P3_IR_REG_12_ );
nand U136192 ( n851, n15474, n15475 );
nand U136193 ( n15475, P1_P3_DATAO_REG_10_, n76041 );
nor U136194 ( n15474, n15477, n15478 );
and U136195 ( n15478, n933, P3_IR_REG_10_ );
nand U136196 ( n841, n15738, n15739 );
nand U136197 ( n15739, P1_P3_DATAO_REG_8_, n76041 );
nor U136198 ( n15738, n15740, n15742 );
and U136199 ( n15742, n933, P3_IR_REG_8_ );
nand U136200 ( n831, n15994, n15995 );
nand U136201 ( n15995, P1_P3_DATAO_REG_6_, n76041 );
nor U136202 ( n15994, n15997, n15998 );
and U136203 ( n15998, n933, P3_IR_REG_6_ );
nand U136204 ( n821, n16263, n16264 );
nand U136205 ( n16264, P1_P3_DATAO_REG_4_, n76041 );
nor U136206 ( n16263, n16265, n16267 );
and U136207 ( n16267, n933, P3_IR_REG_4_ );
nand U136208 ( n2036, n40646, n40647 );
nand U136209 ( n40647, P2_P3_DATAO_REG_2_, n76040 );
nor U136210 ( n40646, n40648, n40649 );
nor U136211 ( n40649, n75423, n76395 );
nand U136212 ( n2046, n40635, n40636 );
nand U136213 ( n40636, P2_P3_DATAO_REG_4_, n76040 );
nor U136214 ( n40635, n40637, n40638 );
nor U136215 ( n40638, n75424, n76395 );
nand U136216 ( n2056, n40624, n40625 );
nand U136217 ( n40625, P2_P3_DATAO_REG_6_, n76039 );
nor U136218 ( n40624, n40626, n40627 );
nor U136219 ( n40627, n75425, n76395 );
nand U136220 ( n2066, n40609, n40610 );
nand U136221 ( n40610, P2_P3_DATAO_REG_8_, n76040 );
nor U136222 ( n40609, n40611, n40612 );
nor U136223 ( n40612, n75418, n76394 );
nand U136224 ( n2086, n40587, n40588 );
nand U136225 ( n40588, P2_P3_DATAO_REG_12_, n76040 );
nor U136226 ( n40587, n40589, n40590 );
nor U136227 ( n40590, n75419, n76394 );
nand U136228 ( n2096, n40576, n40577 );
nand U136229 ( n40577, P2_P3_DATAO_REG_14_, n76040 );
nor U136230 ( n40576, n40578, n40579 );
nor U136231 ( n40579, n75420, n76394 );
nand U136232 ( n2151, n40505, n40506 );
nand U136233 ( n40506, P2_P3_DATAO_REG_25_, n76039 );
nor U136234 ( n40505, n40507, n40508 );
nor U136235 ( n40508, n75365, n76393 );
nand U136236 ( n896, n12644, n12645 );
nand U136237 ( n12645, P1_P3_DATAO_REG_19_, n76041 );
nor U136238 ( n12644, n12647, n12648 );
and U136239 ( n12648, n933, P3_IR_REG_19_ );
nand U136240 ( n2116, n40552, n40553 );
nand U136241 ( n40553, P2_P3_DATAO_REG_18_, n76039 );
nor U136242 ( n40552, n40554, n40555 );
nor U136243 ( n40555, n73035, n76394 );
nand U136244 ( n2076, n40598, n40599 );
nand U136245 ( n40599, P2_P3_DATAO_REG_10_, n76040 );
nor U136246 ( n40598, n40600, n40601 );
nor U136247 ( n40601, n75410, n76394 );
nand U136248 ( n2161, n40490, n40491 );
nand U136249 ( n40491, P2_P3_DATAO_REG_27_, n76039 );
nor U136250 ( n40490, n40492, n40493 );
nor U136251 ( n40493, n73051, n76393 );
nand U136252 ( n2141, n40525, n40526 );
nand U136253 ( n40526, P2_P3_DATAO_REG_23_, n76039 );
nor U136254 ( n40525, n40527, n40528 );
nor U136255 ( n40528, n73496, n76393 );
xor U136256 ( n8572, n11902, P1_P1_PHYADDRPOINTER_REG_26_ );
xor U136257 ( n42904, n45936, P2_P1_PHYADDRPOINTER_REG_16_ );
nand U136258 ( n45936, n7952, P2_P1_PHYADDRPOINTER_REG_15_ );
xnor U136259 ( n54318, n54592, n54593 );
xor U136260 ( n54593, P2_P1_INSTQUEUEWR_ADDR_REG_2_, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U136261 ( n816, n16388, n16389 );
nand U136262 ( n16389, P1_P3_DATAO_REG_3_, n76042 );
nor U136263 ( n16388, n16390, n16392 );
nor U136264 ( n16392, n13650, n73797 );
nand U136265 ( n811, n16695, n16697 );
nand U136266 ( n16697, P1_P3_DATAO_REG_2_, n76042 );
nor U136267 ( n16695, n16698, n16699 );
and U136268 ( n16699, n933, P3_IR_REG_2_ );
nand U136269 ( n46300, P2_P1_STATE2_REG_2_, n47786 );
nand U136270 ( n12689, P1_P1_STATE2_REG_2_, n14532 );
nand U136271 ( n15531, n47784, n47785 );
nand U136272 ( n47785, n76861, P2_P1_INSTADDRPOINTER_REG_0_ );
nor U136273 ( n47784, n47787, n47788 );
nor U136274 ( n47787, n75259, n76332 );
nand U136275 ( n8796, n14529, n14530 );
nand U136276 ( n14530, n76888, P1_P1_INSTADDRPOINTER_REG_0_ );
nor U136277 ( n14529, n14533, n14534 );
nor U136278 ( n14533, n75262, n76598 );
nor U136279 ( n40467, n76397, n40472 );
or U136280 ( n40472, n40457, P4_IR_REG_26_ );
nand U136281 ( n2181, n40465, n40466 );
nand U136282 ( n40465, P2_P3_DATAO_REG_31_, n76039 );
nand U136283 ( n40466, n40467, n40468 );
nor U136284 ( n40468, n40469, n40470 );
nor U136285 ( n67451, P2_P3_INSTADDRPOINTER_REG_28_, n5708 );
nor U136286 ( n32686, P1_P3_INSTADDRPOINTER_REG_28_, n3107 );
nor U136287 ( n25446, P1_P2_INSTADDRPOINTER_REG_28_, n3950 );
nor U136288 ( n58583, P2_P2_INSTADDRPOINTER_REG_28_, n6583 );
nand U136289 ( n67446, P2_P3_INSTADDRPOINTER_REG_29_, n67447 );
nand U136290 ( n67447, n67448, n67449 );
nor U136291 ( n67448, n67432, n67452 );
nor U136292 ( n67449, n67450, n67451 );
nand U136293 ( n32681, P1_P3_INSTADDRPOINTER_REG_29_, n32682 );
nand U136294 ( n32682, n32683, n32684 );
nor U136295 ( n32683, n32667, n32687 );
nor U136296 ( n32684, n32685, n32686 );
nand U136297 ( n25441, P1_P2_INSTADDRPOINTER_REG_29_, n25442 );
nand U136298 ( n25442, n25443, n25444 );
nor U136299 ( n25443, n25427, n25447 );
nor U136300 ( n25444, n25445, n25446 );
nand U136301 ( n58578, P2_P2_INSTADDRPOINTER_REG_29_, n58579 );
nand U136302 ( n58579, n58580, n58581 );
nor U136303 ( n58580, n58564, n58584 );
nor U136304 ( n58581, n58582, n58583 );
nand U136305 ( n8806, n14377, n14378 );
nand U136306 ( n14378, n76888, P1_P1_INSTADDRPOINTER_REG_2_ );
nor U136307 ( n14377, n14379, n14380 );
nor U136308 ( n14379, n14382, n76594 );
nand U136309 ( n15541, n47662, n47663 );
nand U136310 ( n47663, n76861, P2_P1_INSTADDRPOINTER_REG_2_ );
nor U136311 ( n47662, n47664, n47665 );
nor U136312 ( n47664, n47666, n76328 );
nand U136313 ( n15546, n47585, n47586 );
nand U136314 ( n47586, n76861, P2_P1_INSTADDRPOINTER_REG_3_ );
nor U136315 ( n47585, n47587, n47588 );
nor U136316 ( n47587, n47589, n76328 );
nand U136317 ( n8811, n14272, n14273 );
nand U136318 ( n14273, n76888, P1_P1_INSTADDRPOINTER_REG_3_ );
nor U136319 ( n14272, n14274, n14275 );
nor U136320 ( n14274, n14277, n76594 );
nor U136321 ( n37754, P4_IR_REG_0_, n37755 );
nor U136322 ( n37755, n37756, n2153 );
nor U136323 ( n37756, P4_REG2_REG_0_, n2197 );
nand U136324 ( n8816, n14165, n14167 );
nand U136325 ( n14167, n76888, P1_P1_INSTADDRPOINTER_REG_4_ );
nor U136326 ( n14165, n14168, n14169 );
nor U136327 ( n14168, n14170, n76594 );
nand U136328 ( n15551, n47500, n47501 );
nand U136329 ( n47501, n76861, P2_P1_INSTADDRPOINTER_REG_4_ );
nor U136330 ( n47500, n47502, n47503 );
nor U136331 ( n47502, n47504, n76328 );
nand U136332 ( n8821, n14068, n14069 );
nand U136333 ( n14069, n76888, P1_P1_INSTADDRPOINTER_REG_5_ );
nor U136334 ( n14068, n14070, n14072 );
nor U136335 ( n14070, n14073, n76594 );
nand U136336 ( n15556, n47421, n47422 );
nand U136337 ( n47422, n76861, P2_P1_INSTADDRPOINTER_REG_5_ );
nor U136338 ( n47421, n47423, n47424 );
nor U136339 ( n47423, n47425, n76328 );
nand U136340 ( n15536, n47737, n47738 );
nand U136341 ( n47738, n76861, P2_P1_INSTADDRPOINTER_REG_1_ );
nor U136342 ( n47737, n47739, n47740 );
nor U136343 ( n47739, n47741, n76328 );
nand U136344 ( n8801, n14470, n14472 );
nand U136345 ( n14472, n76888, P1_P1_INSTADDRPOINTER_REG_1_ );
nor U136346 ( n14470, n14473, n14474 );
nor U136347 ( n14473, n14475, n76594 );
nand U136348 ( n35701, n189, P1_P3_INSTQUEUERD_ADDR_REG_4_ );
nand U136349 ( n28522, n152, P1_P2_INSTQUEUERD_ADDR_REG_4_ );
nand U136350 ( n70427, n460, P2_P3_INSTQUEUERD_ADDR_REG_4_ );
nand U136351 ( n61827, n424, P2_P2_INSTQUEUERD_ADDR_REG_4_ );
nor U136352 ( n32626, n32627, n32628 );
nor U136353 ( n32627, P1_P3_INSTADDRPOINTER_REG_30_, n32629 );
nor U136354 ( n32629, n32630, n32631 );
nor U136355 ( n25386, n25387, n25388 );
nor U136356 ( n25387, P1_P2_INSTADDRPOINTER_REG_30_, n25389 );
nor U136357 ( n25389, n25390, n25391 );
nor U136358 ( n67391, n67392, n67393 );
nor U136359 ( n67392, P2_P3_INSTADDRPOINTER_REG_30_, n67394 );
nor U136360 ( n67394, n67395, n67396 );
nor U136361 ( n58523, n58524, n58525 );
nor U136362 ( n58524, P2_P2_INSTADDRPOINTER_REG_30_, n58526 );
nor U136363 ( n58526, n58527, n58528 );
xor U136364 ( n8635, n11980, P1_P1_PHYADDRPOINTER_REG_24_ );
nand U136365 ( n54199, n494, P2_P1_INSTQUEUERD_ADDR_REG_4_ );
nand U136366 ( n21216, n223, P1_P1_INSTQUEUERD_ADDR_REG_4_ );
nor U136367 ( n32896, n32905, n32906 );
nor U136368 ( n32905, P1_P3_INSTADDRPOINTER_REG_24_, n32914 );
nor U136369 ( n32906, n32907, n74671 );
nor U136370 ( n32914, n32915, n3128 );
nor U136371 ( n67657, n67666, n67667 );
nor U136372 ( n67666, P2_P3_INSTADDRPOINTER_REG_24_, n67675 );
nor U136373 ( n67667, n67668, n74916 );
nor U136374 ( n67675, n67676, n5729 );
nor U136375 ( n25652, n25661, n25662 );
nor U136376 ( n25661, P1_P2_INSTADDRPOINTER_REG_24_, n25670 );
nor U136377 ( n25662, n25663, n74917 );
nor U136378 ( n25670, n25671, n3972 );
nor U136379 ( n58792, n58801, n58802 );
nor U136380 ( n58801, P2_P2_INSTADDRPOINTER_REG_24_, n58810 );
nor U136381 ( n58802, n58803, n74918 );
nor U136382 ( n58810, n58811, n6604 );
nor U136383 ( n33239, n33246, n33247 );
nor U136384 ( n33247, n33248, n74855 );
nor U136385 ( n33246, P1_P3_INSTADDRPOINTER_REG_15_, n33254 );
nor U136386 ( n33248, n33249, n33250 );
and U136387 ( n33257, n33222, n33277 );
nand U136388 ( n33277, n33278, P1_P3_INSTADDRPOINTER_REG_13_ );
nand U136389 ( n16485, P4_DATAO_REG_0_, n16487 );
nand U136390 ( n16487, n16488, n16489 );
nand U136391 ( n16489, n8222, n73422 );
nor U136392 ( n67994, n68005, n68006 );
nor U136393 ( n68006, n68007, n74852 );
nor U136394 ( n68005, P2_P3_INSTADDRPOINTER_REG_15_, n68013 );
nor U136395 ( n68007, n68008, n68009 );
nor U136396 ( n25991, n26002, n26003 );
nor U136397 ( n26003, n26004, n74853 );
nor U136398 ( n26002, P1_P2_INSTADDRPOINTER_REG_15_, n26010 );
nor U136399 ( n26004, n26005, n26006 );
nor U136400 ( n59129, n59140, n59141 );
nor U136401 ( n59141, n59142, n74854 );
nor U136402 ( n59140, P2_P2_INSTADDRPOINTER_REG_15_, n59148 );
nor U136403 ( n59142, n59143, n59144 );
and U136404 ( n68016, n67977, n68036 );
nand U136405 ( n68036, n68037, P2_P3_INSTADDRPOINTER_REG_13_ );
and U136406 ( n26013, n25974, n26033 );
nand U136407 ( n26033, n26034, P1_P2_INSTADDRPOINTER_REG_13_ );
and U136408 ( n59151, n59112, n59174 );
nand U136409 ( n59174, n59175, P2_P2_INSTADDRPOINTER_REG_13_ );
nor U136410 ( n13293, n13295, n13297 );
nor U136411 ( n13295, P1_P1_INSTADDRPOINTER_REG_20_, n13305 );
nor U136412 ( n13297, n13298, n75053 );
nor U136413 ( n13305, n13307, n13255 );
nor U136414 ( n67692, P2_P3_INSTADDRPOINTER_REG_22_, n5708 );
nor U136415 ( n25687, P1_P2_INSTADDRPOINTER_REG_22_, n3950 );
nor U136416 ( n58827, P2_P2_INSTADDRPOINTER_REG_22_, n6583 );
nand U136417 ( n67687, P2_P3_INSTADDRPOINTER_REG_23_, n67688 );
nand U136418 ( n67688, n67689, n67690 );
nor U136419 ( n67690, n5728, n67691 );
nor U136420 ( n67689, n67692, n67672 );
nand U136421 ( n25682, P1_P2_INSTADDRPOINTER_REG_23_, n25683 );
nand U136422 ( n25683, n25684, n25685 );
nor U136423 ( n25685, n3970, n25686 );
nor U136424 ( n25684, n25687, n25667 );
nand U136425 ( n58822, P2_P2_INSTADDRPOINTER_REG_23_, n58823 );
nand U136426 ( n58823, n58824, n58825 );
nor U136427 ( n58825, n6603, n58826 );
nor U136428 ( n58824, n58827, n58807 );
nor U136429 ( n33163, P1_P3_INSTADDRPOINTER_REG_16_, n3107 );
nand U136430 ( n32926, P1_P3_INSTADDRPOINTER_REG_23_, n32927 );
nand U136431 ( n32927, n32928, n32929 );
nor U136432 ( n32929, n3127, n32930 );
nor U136433 ( n32928, n32931, n32911 );
nor U136434 ( n32931, P1_P3_INSTADDRPOINTER_REG_22_, n3107 );
nand U136435 ( n67908, P2_P3_INSTADDRPOINTER_REG_17_, n67909 );
nand U136436 ( n67909, n67910, n67911 );
nor U136437 ( n67911, n5724, n67912 );
nor U136438 ( n67910, n67914, n67893 );
nand U136439 ( n25905, P1_P2_INSTADDRPOINTER_REG_17_, n25906 );
nand U136440 ( n25906, n25907, n25908 );
nor U136441 ( n25908, n3967, n25909 );
nor U136442 ( n25907, n25911, n25890 );
nand U136443 ( n59043, P2_P2_INSTADDRPOINTER_REG_17_, n59044 );
nand U136444 ( n59044, n59045, n59046 );
nor U136445 ( n59046, n6599, n59047 );
nor U136446 ( n59045, n59049, n59028 );
nor U136447 ( n67914, P2_P3_INSTADDRPOINTER_REG_16_, n5708 );
nor U136448 ( n25911, P1_P2_INSTADDRPOINTER_REG_16_, n3950 );
nor U136449 ( n59049, P2_P2_INSTADDRPOINTER_REG_16_, n6583 );
nor U136450 ( n25532, n25541, n25542 );
nor U136451 ( n25542, n25543, n74960 );
nor U136452 ( n25541, P1_P2_INSTADDRPOINTER_REG_27_, n25552 );
nor U136453 ( n25543, n25544, n25545 );
nor U136454 ( n32772, n32781, n32782 );
nor U136455 ( n32782, n32783, n74961 );
nor U136456 ( n32781, P1_P3_INSTADDRPOINTER_REG_27_, n32792 );
nor U136457 ( n32783, n32784, n32785 );
nor U136458 ( n67537, n67546, n67547 );
nor U136459 ( n67547, n67548, n74962 );
nor U136460 ( n67546, P2_P3_INSTADDRPOINTER_REG_27_, n67557 );
nor U136461 ( n67548, n67549, n67550 );
nor U136462 ( n58669, n58678, n58679 );
nor U136463 ( n58679, n58680, n74963 );
nor U136464 ( n58678, P2_P2_INSTADDRPOINTER_REG_27_, n58689 );
nor U136465 ( n58680, n58681, n58682 );
nor U136466 ( n67577, P2_P3_INSTADDRPOINTER_REG_25_, n5708 );
nor U136467 ( n32812, P1_P3_INSTADDRPOINTER_REG_25_, n3107 );
nor U136468 ( n25572, P1_P2_INSTADDRPOINTER_REG_25_, n3950 );
nor U136469 ( n58709, P2_P2_INSTADDRPOINTER_REG_25_, n6583 );
and U136470 ( n25558, n25515, n25590 );
nand U136471 ( n25590, n25591, P1_P2_INSTADDRPOINTER_REG_25_ );
and U136472 ( n32798, n32755, n32830 );
nand U136473 ( n32830, n32831, P1_P3_INSTADDRPOINTER_REG_25_ );
and U136474 ( n67563, n67520, n67595 );
nand U136475 ( n67595, n67596, P2_P3_INSTADDRPOINTER_REG_25_ );
and U136476 ( n58695, n58652, n58727 );
nand U136477 ( n58727, n58728, P2_P2_INSTADDRPOINTER_REG_25_ );
nand U136478 ( n67572, P2_P3_INSTADDRPOINTER_REG_26_, n67573 );
nand U136479 ( n67573, n67574, n67575 );
nor U136480 ( n67575, n5730, n67576 );
nor U136481 ( n67574, n67577, n67551 );
nand U136482 ( n32807, P1_P3_INSTADDRPOINTER_REG_26_, n32808 );
nand U136483 ( n32808, n32809, n32810 );
nor U136484 ( n32810, n3129, n32811 );
nor U136485 ( n32809, n32812, n32786 );
nand U136486 ( n25567, P1_P2_INSTADDRPOINTER_REG_26_, n25568 );
nand U136487 ( n25568, n25569, n25570 );
nor U136488 ( n25570, n3973, n25571 );
nor U136489 ( n25569, n25572, n25546 );
nand U136490 ( n58704, P2_P2_INSTADDRPOINTER_REG_26_, n58705 );
nand U136491 ( n58705, n58706, n58707 );
nor U136492 ( n58707, n6605, n58708 );
nor U136493 ( n58706, n58709, n58683 );
nor U136494 ( n13463, n13473, n13474 );
nor U136495 ( n13474, n13475, n74818 );
nor U136496 ( n13473, P1_P1_INSTADDRPOINTER_REG_16_, n13484 );
nor U136497 ( n13475, n13477, n13478 );
and U136498 ( n32422, P1_P3_M_IO_N_REG, n75968 );
nand U136499 ( n29171, P1_READY22_REG, n36164 );
nand U136500 ( n36164, n36165, n36166 );
and U136501 ( n36165, P3_RD_REG, P1_P3_W_R_N_REG );
and U136502 ( n36166, P1_P3_D_C_N_REG, n32422 );
nor U136503 ( n46474, n46483, n46484 );
nor U136504 ( n46484, n46485, n74930 );
nor U136505 ( n46483, P2_P1_INSTADDRPOINTER_REG_27_, n46494 );
nor U136506 ( n46485, n46486, n46487 );
nor U136507 ( n46387, P2_P1_INSTADDRPOINTER_REG_28_, n7494 );
nand U136508 ( n46382, P2_P1_INSTADDRPOINTER_REG_29_, n46383 );
nand U136509 ( n46383, n46384, n46385 );
nor U136510 ( n46384, n46368, n46388 );
nor U136511 ( n46385, n46386, n46387 );
nand U136512 ( n801, n21630, n21631 );
nand U136513 ( n21630, P1_P3_DATAO_REG_0_, n76042 );
nand U136514 ( n21631, P3_IR_REG_0_, n21632 );
nand U136515 ( n21632, n13650, n76626 );
xor U136516 ( n8707, n12045, P1_P1_PHYADDRPOINTER_REG_22_ );
nand U136517 ( n2026, n40657, n40658 );
nand U136518 ( n40657, P2_P3_DATAO_REG_0_, n76922 );
nand U136519 ( n40658, P4_IR_REG_0_, n40659 );
nand U136520 ( n40659, n76395, n76399 );
nor U136521 ( n12980, n12983, n12984 );
nor U136522 ( n12984, n12985, n74886 );
nor U136523 ( n12983, P1_P1_INSTADDRPOINTER_REG_26_, n12994 );
nor U136524 ( n12985, n12987, n12988 );
nand U136525 ( n32593, n32597, n32598 );
nand U136526 ( n32597, n76469, P1_P3_INSTADDRPOINTER_REG_31_ );
nand U136527 ( n32598, n32599, P1_P3_REIP_REG_31_ );
nand U136528 ( n25353, n25357, n25358 );
nand U136529 ( n25357, n76520, P1_P2_INSTADDRPOINTER_REG_31_ );
nand U136530 ( n25358, n25359, P1_P2_REIP_REG_31_ );
nand U136531 ( n67358, n67362, n67363 );
nand U136532 ( n67362, n76196, P2_P3_INSTADDRPOINTER_REG_31_ );
nand U136533 ( n67363, n67364, P2_P3_REIP_REG_31_ );
nand U136534 ( n58490, n58494, n58495 );
nand U136535 ( n58494, n76262, P2_P2_INSTADDRPOINTER_REG_31_ );
nand U136536 ( n58495, n58496, P2_P2_REIP_REG_31_ );
nor U136537 ( n13077, n13088, n13089 );
nor U136538 ( n13088, P1_P1_INSTADDRPOINTER_REG_24_, n13099 );
nor U136539 ( n13089, n13090, n74653 );
nor U136540 ( n13099, n13100, n4869 );
nor U136541 ( n46610, n46619, n46620 );
nor U136542 ( n46619, P2_P1_INSTADDRPOINTER_REG_24_, n46628 );
nor U136543 ( n46620, n46621, n74881 );
nor U136544 ( n46628, n46629, n46589 );
nor U136545 ( n68226, n68240, n68241 );
nor U136546 ( n68240, P2_P3_INSTADDRPOINTER_REG_9_, n68250 );
nor U136547 ( n68241, n68242, n73084 );
nor U136548 ( n68250, n68251, n68199 );
nor U136549 ( n26225, n26239, n26240 );
nor U136550 ( n26239, P1_P2_INSTADDRPOINTER_REG_9_, n26249 );
nor U136551 ( n26240, n26241, n73085 );
nor U136552 ( n26249, n26250, n26198 );
nor U136553 ( n59364, n59378, n59379 );
nor U136554 ( n59378, P2_P2_INSTADDRPOINTER_REG_9_, n59388 );
nor U136555 ( n59379, n59380, n73086 );
nor U136556 ( n59388, n59389, n59337 );
nor U136557 ( n13513, n13527, n13528 );
nor U136558 ( n13528, n13529, n74823 );
nor U136559 ( n13527, P1_P1_INSTADDRPOINTER_REG_15_, n13537 );
nor U136560 ( n13529, n13530, n13532 );
and U136561 ( n13540, n13492, n13565 );
nand U136562 ( n13565, n13567, P1_P1_INSTADDRPOINTER_REG_13_ );
nor U136563 ( n33125, n33131, n33132 );
nor U136564 ( n33131, P1_P3_INSTADDRPOINTER_REG_18_, n33139 );
nor U136565 ( n33132, n33133, n74635 );
nor U136566 ( n33139, n33140, n3124 );
nor U136567 ( n33475, n33485, n33486 );
nor U136568 ( n33485, P1_P3_INSTADDRPOINTER_REG_9_, n33495 );
nor U136569 ( n33486, n33487, n73114 );
nor U136570 ( n33495, n33496, n33448 );
xor U136571 ( n8883, n12248, P1_P1_PHYADDRPOINTER_REG_16_ );
nand U136572 ( n12248, n5297, P1_P1_PHYADDRPOINTER_REG_15_ );
nor U136573 ( n67881, n67887, n67888 );
nor U136574 ( n67887, P2_P3_INSTADDRPOINTER_REG_18_, n67895 );
nor U136575 ( n67888, n67889, n74546 );
nor U136576 ( n67895, n67896, n5725 );
nor U136577 ( n25878, n25884, n25885 );
nor U136578 ( n25884, P1_P2_INSTADDRPOINTER_REG_18_, n25892 );
nor U136579 ( n25885, n25886, n74547 );
nor U136580 ( n25892, n25893, n3968 );
nor U136581 ( n59016, n59022, n59023 );
nor U136582 ( n59022, P2_P2_INSTADDRPOINTER_REG_18_, n59030 );
nor U136583 ( n59023, n59024, n74548 );
nor U136584 ( n59030, n59031, n6600 );
nand U136585 ( n22072, n22073, n22074 );
nand U136586 ( n22073, P1_P2_REIP_REG_26_, n22067 );
nand U136587 ( n22074, n174, n73294 );
nand U136588 ( n55182, n55183, n55184 );
nand U136589 ( n55183, P2_P2_REIP_REG_26_, n55177 );
nand U136590 ( n55184, n446, n73295 );
nor U136591 ( n46959, n46970, n46971 );
nor U136592 ( n46971, n46972, n74822 );
nor U136593 ( n46970, P2_P1_INSTADDRPOINTER_REG_15_, n46978 );
nor U136594 ( n46972, n46973, n46974 );
nand U136595 ( n63154, n63155, n63156 );
nand U136596 ( n63155, P2_P3_REIP_REG_26_, n63149 );
nand U136597 ( n63156, n479, n73296 );
nand U136598 ( n29391, n29392, n29393 );
nand U136599 ( n29392, P1_P3_REIP_REG_26_, n29386 );
nand U136600 ( n29393, n208, n73297 );
and U136601 ( n46981, n46930, n47001 );
nand U136602 ( n47001, n47002, P2_P1_INSTADDRPOINTER_REG_13_ );
nor U136603 ( n45170, n45172, n45173 );
nor U136604 ( n45173, n880, n74381 );
nor U136605 ( n45172, n45174, n45175 );
nand U136606 ( n45175, P3_REG2_REG_8_, n42957 );
nand U136607 ( n63752, n63753, n63754 );
nand U136608 ( n63753, P2_P3_PHYADDRPOINTER_REG_11_, n5629 );
nand U136609 ( n63754, P2_P3_REIP_REG_11_, n63740 );
nand U136610 ( n63908, n63909, n63910 );
nand U136611 ( n63909, P2_P3_PHYADDRPOINTER_REG_5_, n5629 );
nand U136612 ( n63910, P2_P3_REIP_REG_5_, n63896 );
nand U136613 ( n29792, n29793, n29794 );
nand U136614 ( n29793, P1_P3_PHYADDRPOINTER_REG_11_, n3028 );
nand U136615 ( n29794, P1_P3_REIP_REG_11_, n29780 );
nand U136616 ( n29952, n29953, n29954 );
nand U136617 ( n29953, P1_P3_PHYADDRPOINTER_REG_5_, n3028 );
nand U136618 ( n29954, P1_P3_REIP_REG_5_, n29940 );
nand U136619 ( n22471, n22472, n22473 );
nand U136620 ( n22472, P1_P2_PHYADDRPOINTER_REG_11_, n3872 );
nand U136621 ( n22473, P1_P2_REIP_REG_11_, n22459 );
nand U136622 ( n22629, n22630, n22631 );
nand U136623 ( n22630, P1_P2_PHYADDRPOINTER_REG_5_, n3872 );
nand U136624 ( n22631, P1_P2_REIP_REG_5_, n22617 );
nand U136625 ( n55586, n55587, n55588 );
nand U136626 ( n55587, P2_P2_PHYADDRPOINTER_REG_11_, n6504 );
nand U136627 ( n55588, P2_P2_REIP_REG_11_, n55574 );
nand U136628 ( n55742, n55743, n55744 );
nand U136629 ( n55743, P2_P2_PHYADDRPOINTER_REG_5_, n6504 );
nand U136630 ( n55744, P2_P2_REIP_REG_5_, n55730 );
nor U136631 ( n68633, n68672, n68673 );
nor U136632 ( n68672, P2_P3_INSTADDRPOINTER_REG_3_, n68678 );
nor U136633 ( n68673, n68674, n74408 );
nor U136634 ( n68678, n68679, n68605 );
nor U136635 ( n33877, n33916, n33917 );
nor U136636 ( n33916, P1_P3_INSTADDRPOINTER_REG_3_, n33922 );
nor U136637 ( n33917, n33918, n74412 );
nor U136638 ( n33922, n33923, n33849 );
nor U136639 ( n26632, n26671, n26672 );
nor U136640 ( n26671, P1_P2_INSTADDRPOINTER_REG_3_, n26677 );
nor U136641 ( n26672, n26673, n74409 );
nor U136642 ( n26677, n26678, n26604 );
nor U136643 ( n59774, n59813, n59814 );
nor U136644 ( n59813, P2_P2_INSTADDRPOINTER_REG_3_, n59819 );
nor U136645 ( n59814, n59815, n74410 );
nor U136646 ( n59819, n59820, n59746 );
nand U136647 ( n62893, P2_READY22_REG, n70883 );
nand U136648 ( n70883, n70884, n70885 );
and U136649 ( n70884, P4_RD_REG, P2_P3_W_R_N_REG );
and U136650 ( n70885, n21687, P2_P3_D_C_N_REG );
and U136651 ( n21687, P2_P3_M_IO_N_REG, n75969 );
nand U136652 ( n63841, P2_P3_REIP_REG_8_, n63810 );
nand U136653 ( n29885, P1_P3_REIP_REG_8_, n29854 );
nand U136654 ( n22562, P1_P2_REIP_REG_8_, n22531 );
nand U136655 ( n55675, P2_P2_REIP_REG_8_, n55644 );
nand U136656 ( n63540, P2_P3_REIP_REG_17_, n63524 );
nand U136657 ( n29641, P1_P3_REIP_REG_17_, n29625 );
nand U136658 ( n22320, P1_P2_REIP_REG_17_, n22304 );
nand U136659 ( n55432, P2_P2_REIP_REG_17_, n55416 );
nor U136660 ( n45235, n45237, n45238 );
nor U136661 ( n45238, n880, n74380 );
nor U136662 ( n45237, n45239, n45240 );
nand U136663 ( n45240, P3_REG1_REG_8_, n42957 );
nand U136664 ( n63624, P2_P3_REIP_REG_14_, n63592 );
nand U136665 ( n29725, P1_P3_REIP_REG_14_, n29693 );
nand U136666 ( n22404, P1_P2_REIP_REG_14_, n22372 );
nand U136667 ( n55516, P2_P2_REIP_REG_14_, n55484 );
nor U136668 ( n68376, n68429, n68430 );
nor U136669 ( n68429, P2_P3_INSTADDRPOINTER_REG_6_, n68437 );
nor U136670 ( n68430, n68431, n73066 );
nor U136671 ( n68437, n68346, n68438 );
nor U136672 ( n33620, n33673, n33674 );
nor U136673 ( n33673, P1_P3_INSTADDRPOINTER_REG_6_, n33681 );
nor U136674 ( n33674, n33675, n73088 );
nor U136675 ( n33681, n33590, n33682 );
nor U136676 ( n26375, n26428, n26429 );
nor U136677 ( n26428, P1_P2_INSTADDRPOINTER_REG_6_, n26436 );
nor U136678 ( n26429, n26430, n73067 );
nor U136679 ( n26436, n26345, n26437 );
nor U136680 ( n59514, n59567, n59568 );
nor U136681 ( n59567, P2_P2_INSTADDRPOINTER_REG_6_, n59575 );
nor U136682 ( n59568, n59569, n73068 );
nor U136683 ( n59575, n59484, n59576 );
nor U136684 ( n46645, P2_P1_INSTADDRPOINTER_REG_22_, n7494 );
nand U136685 ( n46640, P2_P1_INSTADDRPOINTER_REG_23_, n46641 );
nand U136686 ( n46641, n46642, n46643 );
nor U136687 ( n46643, n7514, n46644 );
nor U136688 ( n46642, n46645, n46625 );
nor U136689 ( n46516, P2_P1_INSTADDRPOINTER_REG_25_, n7494 );
nand U136690 ( n46511, P2_P1_INSTADDRPOINTER_REG_26_, n46512 );
nand U136691 ( n46512, n46513, n46514 );
nor U136692 ( n46514, n7515, n46515 );
nor U136693 ( n46513, n46516, n46488 );
nand U136694 ( n46861, P2_P1_INSTADDRPOINTER_REG_17_, n46862 );
nand U136695 ( n46862, n46863, n46864 );
nor U136696 ( n46864, n7510, n46865 );
nor U136697 ( n46863, n46867, n46846 );
nor U136698 ( n46867, P2_P1_INSTADDRPOINTER_REG_16_, n7494 );
nor U136699 ( n42271, P3_IR_REG_0_, n42272 );
nor U136700 ( n42272, n42273, n812 );
nor U136701 ( n42273, P3_REG2_REG_0_, n814 );
xor U136702 ( n63556, n66887, P2_P3_PHYADDRPOINTER_REG_16_ );
nand U136703 ( n66887, n6164, P2_P3_PHYADDRPOINTER_REG_15_ );
xor U136704 ( n29657, n32248, P1_P3_PHYADDRPOINTER_REG_16_ );
nand U136705 ( n32248, n3549, P1_P3_PHYADDRPOINTER_REG_15_ );
xor U136706 ( n22336, n25011, P1_P2_PHYADDRPOINTER_REG_16_ );
nand U136707 ( n25011, n4387, P1_P2_PHYADDRPOINTER_REG_15_ );
xor U136708 ( n55448, n58146, P2_P2_PHYADDRPOINTER_REG_16_ );
nand U136709 ( n58146, n7019, P2_P2_PHYADDRPOINTER_REG_15_ );
nor U136710 ( n33358, P1_P3_INSTADDRPOINTER_REG_11_, n3083 );
nor U136711 ( n68115, P2_P3_INSTADDRPOINTER_REG_11_, n5684 );
nor U136712 ( n26112, P1_P2_INSTADDRPOINTER_REG_11_, n3927 );
nor U136713 ( n59253, P2_P2_INSTADDRPOINTER_REG_11_, n6559 );
nand U136714 ( n33352, P1_P3_INSTADDRPOINTER_REG_12_, n33353 );
nand U136715 ( n33353, n33354, n33355 );
nor U136716 ( n33355, n33356, n33357 );
nor U136717 ( n33354, n33358, n33333 );
nand U136718 ( n68109, P2_P3_INSTADDRPOINTER_REG_12_, n68110 );
nand U136719 ( n68110, n68111, n68112 );
nor U136720 ( n68112, n68113, n68114 );
nor U136721 ( n68111, n68115, n68090 );
nand U136722 ( n26106, P1_P2_INSTADDRPOINTER_REG_12_, n26107 );
nand U136723 ( n26107, n26108, n26109 );
nor U136724 ( n26109, n26110, n26111 );
nor U136725 ( n26108, n26112, n26087 );
nand U136726 ( n59247, P2_P2_INSTADDRPOINTER_REG_12_, n59248 );
nand U136727 ( n59248, n59249, n59250 );
nor U136728 ( n59250, n59251, n59252 );
nor U136729 ( n59249, n59253, n59228 );
nor U136730 ( n33017, P1_P3_INSTADDRPOINTER_REG_20_, n3083 );
nor U136731 ( n67773, P2_P3_INSTADDRPOINTER_REG_20_, n5684 );
nor U136732 ( n25770, P1_P2_INSTADDRPOINTER_REG_20_, n3927 );
nor U136733 ( n58908, P2_P2_INSTADDRPOINTER_REG_20_, n6559 );
nand U136734 ( n67767, P2_P3_INSTADDRPOINTER_REG_21_, n67768 );
nand U136735 ( n67768, n67769, n67770 );
nor U136736 ( n67770, n5728, n67771 );
nor U136737 ( n67769, n67773, n67774 );
nand U136738 ( n33011, P1_P3_INSTADDRPOINTER_REG_21_, n33012 );
nand U136739 ( n33012, n33013, n33014 );
nor U136740 ( n33014, n3127, n33015 );
nor U136741 ( n33013, n33017, n33018 );
nand U136742 ( n25764, P1_P2_INSTADDRPOINTER_REG_21_, n25765 );
nand U136743 ( n25765, n25766, n25767 );
nor U136744 ( n25767, n3970, n25768 );
nor U136745 ( n25766, n25770, n25771 );
nand U136746 ( n58902, P2_P2_INSTADDRPOINTER_REG_21_, n58903 );
nand U136747 ( n58903, n58904, n58905 );
nor U136748 ( n58905, n6603, n58906 );
nor U136749 ( n58904, n58908, n58909 );
nor U136750 ( n13814, n13818, n13819 );
nor U136751 ( n13818, P1_P1_INSTADDRPOINTER_REG_9_, n13830 );
nor U136752 ( n13819, n13820, n73109 );
nor U136753 ( n13830, n13832, n13775 );
nor U136754 ( n13370, n13378, n13379 );
nor U136755 ( n13378, P1_P1_INSTADDRPOINTER_REG_18_, n13388 );
nor U136756 ( n13379, n13380, n74599 );
nor U136757 ( n13388, n13389, n4865 );
nor U136758 ( n68467, n68505, n68506 );
nor U136759 ( n68505, P2_P3_INSTADDRPOINTER_REG_5_, n68513 );
nor U136760 ( n68506, n68507, n74452 );
nor U136761 ( n68513, n68514, n68439 );
nor U136762 ( n33711, n33749, n33750 );
nor U136763 ( n33749, P1_P3_INSTADDRPOINTER_REG_5_, n33757 );
nor U136764 ( n33750, n33751, n74455 );
nor U136765 ( n33757, n33758, n33683 );
nor U136766 ( n26466, n26504, n26505 );
nor U136767 ( n26504, P1_P2_INSTADDRPOINTER_REG_5_, n26512 );
nor U136768 ( n26505, n26506, n74453 );
nor U136769 ( n26512, n26513, n26438 );
nor U136770 ( n59605, n59643, n59644 );
nor U136771 ( n59643, P2_P2_INSTADDRPOINTER_REG_5_, n59651 );
nor U136772 ( n59644, n59645, n74454 );
nor U136773 ( n59651, n59652, n59577 );
nor U136774 ( n14305, n14354, n14355 );
nor U136775 ( n14354, P1_P1_INSTADDRPOINTER_REG_3_, n14362 );
nor U136776 ( n14355, n14357, n74429 );
nor U136777 ( n14362, n14363, n14270 );
nor U136778 ( n67818, n67820, n67821 );
nor U136779 ( n67820, P2_P3_INSTADDRPOINTER_REG_20_, n67829 );
nor U136780 ( n67821, n67822, n75017 );
nor U136781 ( n67829, n67830, n67786 );
nor U136782 ( n25815, n25817, n25818 );
nor U136783 ( n25817, P1_P2_INSTADDRPOINTER_REG_20_, n25826 );
nor U136784 ( n25818, n25819, n75018 );
nor U136785 ( n25826, n25827, n25783 );
nor U136786 ( n58953, n58955, n58956 );
nor U136787 ( n58955, P2_P2_INSTADDRPOINTER_REG_20_, n58964 );
nor U136788 ( n58956, n58957, n75019 );
nor U136789 ( n58964, n58965, n58921 );
xor U136790 ( n22040, n24696, P1_P2_PHYADDRPOINTER_REG_28_ );
xor U136791 ( n29359, n31908, P1_P3_PHYADDRPOINTER_REG_28_ );
xor U136792 ( n63122, n66531, P2_P3_PHYADDRPOINTER_REG_28_ );
xor U136793 ( n55150, n57830, P2_P2_PHYADDRPOINTER_REG_28_ );
nor U136794 ( n68277, n68284, n68285 );
nor U136795 ( n68284, P2_P3_INSTADDRPOINTER_REG_8_, n68292 );
nor U136796 ( n68285, n68286, n73187 );
nor U136797 ( n68292, n68293, n68254 );
nor U136798 ( n26276, n26283, n26284 );
nor U136799 ( n26283, P1_P2_INSTADDRPOINTER_REG_8_, n26291 );
nor U136800 ( n26284, n26285, n73188 );
nor U136801 ( n26291, n26292, n26253 );
nor U136802 ( n59415, n59422, n59423 );
nor U136803 ( n59422, P2_P2_INSTADDRPOINTER_REG_8_, n59430 );
nor U136804 ( n59423, n59424, n73189 );
nor U136805 ( n59430, n59431, n59392 );
nor U136806 ( n33062, n33064, n33065 );
nor U136807 ( n33064, P1_P3_INSTADDRPOINTER_REG_20_, n33073 );
nor U136808 ( n33065, n33066, n75060 );
nor U136809 ( n33073, n33074, n33031 );
nor U136810 ( n13985, n14052, n14053 );
nor U136811 ( n14052, P1_P1_INSTADDRPOINTER_REG_6_, n14062 );
nor U136812 ( n14053, n14054, n73090 );
nor U136813 ( n14062, n13948, n14063 );
nor U136814 ( n13335, P1_P1_INSTADDRPOINTER_REG_18_, n4827 );
nor U136815 ( n68149, n68156, n68157 );
nor U136816 ( n68156, P2_P3_INSTADDRPOINTER_REG_11_, n68164 );
nor U136817 ( n68157, n68158, n72950 );
nor U136818 ( n68164, n68165, n68130 );
nor U136819 ( n26148, n26155, n26156 );
nor U136820 ( n26155, P1_P2_INSTADDRPOINTER_REG_11_, n26163 );
nor U136821 ( n26156, n26157, n72951 );
nor U136822 ( n26163, n26164, n26127 );
nor U136823 ( n59287, n59294, n59295 );
nor U136824 ( n59294, P2_P2_INSTADDRPOINTER_REG_11_, n59302 );
nor U136825 ( n59295, n59296, n72952 );
nor U136826 ( n59302, n59303, n59268 );
nand U136827 ( n13325, P1_P1_INSTADDRPOINTER_REG_19_, n13327 );
nand U136828 ( n13327, n13328, n13329 );
nor U136829 ( n13329, n13330, n13332 );
nor U136830 ( n13328, n13334, n13335 );
nor U136831 ( n33522, n33528, n33529 );
nor U136832 ( n33528, P1_P3_INSTADDRPOINTER_REG_8_, n33536 );
nor U136833 ( n33529, n33530, n73197 );
nor U136834 ( n33536, n33537, n33499 );
nor U136835 ( n13023, P1_P1_INSTADDRPOINTER_REG_24_, n4827 );
nor U136836 ( n33397, n33406, n33407 );
nor U136837 ( n33406, P1_P3_INSTADDRPOINTER_REG_11_, n33414 );
nor U136838 ( n33407, n33408, n74755 );
nor U136839 ( n33414, n33415, n33378 );
nand U136840 ( n13014, P1_P1_INSTADDRPOINTER_REG_25_, n13015 );
nand U136841 ( n13015, n13017, n13018 );
nor U136842 ( n13018, n4870, n13019 );
nor U136843 ( n13017, n13022, n13023 );
nor U136844 ( n47195, n47209, n47210 );
nor U136845 ( n47209, P2_P1_INSTADDRPOINTER_REG_9_, n47219 );
nor U136846 ( n47210, n47211, n73078 );
nor U136847 ( n47219, n47220, n47168 );
nor U136848 ( n46834, n46840, n46841 );
nor U136849 ( n46840, P2_P1_INSTADDRPOINTER_REG_18_, n46848 );
nor U136850 ( n46841, n46842, n74524 );
nor U136851 ( n46848, n46849, n7512 );
xor U136852 ( n49673, P3_DATAO_REG_31_, n49682 );
nor U136853 ( n13393, n13347, n13427 );
and U136854 ( n13427, n13428, P1_P1_INSTADDRPOINTER_REG_16_ );
nor U136855 ( n47612, n47651, n47652 );
nor U136856 ( n47651, P2_P1_INSTADDRPOINTER_REG_3_, n47657 );
nor U136857 ( n47652, n47653, n74400 );
nor U136858 ( n47657, n47658, n47584 );
nor U136859 ( n13418, P1_P1_INSTADDRPOINTER_REG_16_, n4850 );
nor U136860 ( n13120, P1_P1_INSTADDRPOINTER_REG_22_, n4850 );
nand U136861 ( n13835, n13884, n13885 );
nand U136862 ( n13885, n5224, n12999 );
nand U136863 ( n13884, n13890, P1_P1_INSTADDRPOINTER_REG_7_ );
and U136864 ( n13832, n13835, P1_P1_INSTADDRPOINTER_REG_8_ );
nand U136865 ( n47223, n47263, n47264 );
nand U136866 ( n47264, n7878, n76101 );
nand U136867 ( n47263, n47268, P2_P1_INSTADDRPOINTER_REG_7_ );
nand U136868 ( n13114, P1_P1_INSTADDRPOINTER_REG_23_, n13115 );
nand U136869 ( n13115, n13117, n13118 );
nor U136870 ( n13118, n4868, n13119 );
nor U136871 ( n13117, n13120, n13095 );
and U136872 ( n47220, n47223, P2_P1_INSTADDRPOINTER_REG_8_ );
xnor U136873 ( n63514, n6175, P2_P3_PHYADDRPOINTER_REG_18_ );
xnor U136874 ( n29615, n3560, P1_P3_PHYADDRPOINTER_REG_18_ );
xnor U136875 ( n22294, n4398, P1_P2_PHYADDRPOINTER_REG_18_ );
xnor U136876 ( n55406, n7030, P2_P2_PHYADDRPOINTER_REG_18_ );
nor U136877 ( n13238, P1_P1_INSTADDRPOINTER_REG_20_, n4825 );
nand U136878 ( n13230, P1_P1_INSTADDRPOINTER_REG_21_, n13232 );
nand U136879 ( n13232, n13233, n13234 );
nor U136880 ( n13234, n4868, n13235 );
nor U136881 ( n13233, n13238, n13239 );
nor U136882 ( n47344, n47397, n47398 );
nor U136883 ( n47397, P2_P1_INSTADDRPOINTER_REG_6_, n47405 );
nor U136884 ( n47398, n47399, n73065 );
nor U136885 ( n47405, n47314, n47406 );
nand U136886 ( n13663, P1_P1_INSTADDRPOINTER_REG_12_, n13664 );
nand U136887 ( n13664, n13665, n13667 );
nor U136888 ( n13667, n13668, n13669 );
nor U136889 ( n13665, n13670, n13632 );
nor U136890 ( n13670, P1_P1_INSTADDRPOINTER_REG_11_, n4825 );
nor U136891 ( n14098, n14145, n14147 );
nor U136892 ( n14145, P1_P1_INSTADDRPOINTER_REG_5_, n14155 );
nor U136893 ( n14147, n14148, n74461 );
nor U136894 ( n14155, n14157, n14064 );
and U136895 ( n33496, n33499, P1_P3_INSTADDRPOINTER_REG_8_ );
and U136896 ( n68251, n68254, P2_P3_INSTADDRPOINTER_REG_8_ );
and U136897 ( n26250, n26253, P1_P2_INSTADDRPOINTER_REG_8_ );
and U136898 ( n59389, n59392, P2_P2_INSTADDRPOINTER_REG_8_ );
nor U136899 ( n13864, n13872, n13873 );
nor U136900 ( n13872, P1_P1_INSTADDRPOINTER_REG_8_, n13882 );
nor U136901 ( n13873, n13874, n73176 );
nor U136902 ( n13882, n13883, n13835 );
nand U136903 ( n11595, n16443, n16444 );
nand U136904 ( n16443, P1_BUF1_REG_0_, n76610 );
nand U136905 ( n16444, n16445, n76654 );
nor U136906 ( n16445, n76610, n76789 );
nand U136907 ( n63623, P2_P3_EBX_REG_14_, n474 );
nand U136908 ( n63840, P2_P3_EBX_REG_8_, n474 );
nand U136909 ( n55515, P2_P2_EBX_REG_14_, n442 );
xor U136910 ( n63167, n66574, P2_P3_PHYADDRPOINTER_REG_26_ );
xor U136911 ( n29404, n31971, P1_P3_PHYADDRPOINTER_REG_26_ );
xor U136912 ( n22085, n24739, P1_P2_PHYADDRPOINTER_REG_26_ );
xor U136913 ( n55195, n57873, P2_P2_PHYADDRPOINTER_REG_26_ );
nand U136914 ( n63950, P2_P3_EBX_REG_4_, n474 );
nand U136915 ( n64060, P2_P3_EBX_REG_2_, n474 );
nand U136916 ( n29724, P1_P3_EBX_REG_14_, n203 );
nand U136917 ( n29884, P1_P3_EBX_REG_8_, n203 );
nand U136918 ( n29994, P1_P3_EBX_REG_4_, n203 );
nand U136919 ( n30043, P1_P3_EBX_REG_2_, n203 );
nand U136920 ( n22403, P1_P2_EBX_REG_14_, n169 );
nand U136921 ( n22561, P1_P2_EBX_REG_8_, n169 );
nand U136922 ( n22671, P1_P2_EBX_REG_4_, n169 );
nand U136923 ( n22720, P1_P2_EBX_REG_2_, n169 );
nand U136924 ( n55674, P2_P2_EBX_REG_8_, n442 );
nand U136925 ( n55784, P2_P2_EBX_REG_4_, n442 );
nand U136926 ( n55836, P2_P2_EBX_REG_2_, n442 );
nor U136927 ( n13713, n13722, n13723 );
nor U136928 ( n13722, P1_P1_INSTADDRPOINTER_REG_11_, n13732 );
nor U136929 ( n13723, n13724, n73116 );
nor U136930 ( n13732, n13733, n13689 );
nor U136931 ( n13757, P1_P1_INSTADDRPOINTER_REG_9_, n4827 );
nand U136932 ( n13750, P1_P1_INSTADDRPOINTER_REG_10_, n13752 );
nand U136933 ( n13752, n13753, n13754 );
nor U136934 ( n13754, n13668, n13755 );
nor U136935 ( n13753, n13757, n13758 );
nand U136936 ( n47078, P2_P1_INSTADDRPOINTER_REG_12_, n47079 );
nand U136937 ( n47079, n47080, n47081 );
nor U136938 ( n47081, n47082, n47083 );
nor U136939 ( n47080, n47084, n47059 );
nor U136940 ( n47084, P2_P1_INSTADDRPOINTER_REG_11_, n7469 );
nor U136941 ( n46726, P2_P1_INSTADDRPOINTER_REG_20_, n7469 );
nand U136942 ( n46720, P2_P1_INSTADDRPOINTER_REG_21_, n46721 );
nand U136943 ( n46721, n46722, n46723 );
nor U136944 ( n46723, n7514, n46724 );
nor U136945 ( n46722, n46726, n46727 );
nand U136946 ( n16337, n16338, n16339 );
nand U136947 ( n16339, P1_P1_INSTQUEUE_REG_14__0_, n16340 );
nand U136948 ( n16338, n4797, n1 );
nand U136949 ( n16232, n16233, n16234 );
nand U136950 ( n16234, P1_P1_INSTQUEUE_REG_13__0_, n16235 );
nand U136951 ( n16233, n4798, n1 );
nand U136952 ( n16029, n16030, n16032 );
nand U136953 ( n16032, P1_P1_INSTQUEUE_REG_11__0_, n16033 );
nand U136954 ( n16030, n4799, n1 );
nand U136955 ( n15922, n15923, n15924 );
nand U136956 ( n15924, P1_P1_INSTQUEUE_REG_10__0_, n15925 );
nand U136957 ( n15923, n4800, n1 );
nand U136958 ( n15817, n15818, n15819 );
nand U136959 ( n15819, P1_P1_INSTQUEUE_REG_9__0_, n15820 );
nand U136960 ( n15818, n4802, n1 );
nand U136961 ( n15508, n15509, n15510 );
nand U136962 ( n15510, P1_P1_INSTQUEUE_REG_6__0_, n15512 );
nand U136963 ( n15509, n4804, n1 );
nand U136964 ( n15402, n15403, n15404 );
nand U136965 ( n15404, P1_P1_INSTQUEUE_REG_5__0_, n15405 );
nand U136966 ( n15403, n4805, n1 );
nand U136967 ( n15605, n15607, n15608 );
nand U136968 ( n15608, P1_P1_INSTQUEUE_REG_7__0_, n15609 );
nand U136969 ( n15607, n4803, n1 );
nor U136970 ( n47446, n47484, n47485 );
nor U136971 ( n47484, P2_P1_INSTADDRPOINTER_REG_5_, n47492 );
nor U136972 ( n47485, n47486, n74443 );
nor U136973 ( n47492, n47493, n47407 );
nor U136974 ( n46771, n46773, n46774 );
nor U136975 ( n46773, P2_P1_INSTADDRPOINTER_REG_20_, n46782 );
nor U136976 ( n46774, n46775, n75020 );
nor U136977 ( n46782, n46783, n46739 );
nor U136978 ( n47246, n47253, n47254 );
nor U136979 ( n47253, P2_P1_INSTADDRPOINTER_REG_8_, n47261 );
nor U136980 ( n47254, n47255, n73178 );
nor U136981 ( n47261, n47262, n47223 );
nor U136982 ( n47118, n47125, n47126 );
nor U136983 ( n47125, P2_P1_INSTADDRPOINTER_REG_11_, n47133 );
nor U136984 ( n47126, n47127, n72948 );
nor U136985 ( n47133, n47134, n47099 );
nor U136986 ( n61288, P3_B_REG, n41449 );
nor U136987 ( n12802, n12810, n12812 );
nor U136988 ( n12810, P1_P1_INSTADDRPOINTER_REG_29_, n12829 );
nor U136989 ( n12812, n12813, n73279 );
nor U136990 ( n12829, n12830, n12763 );
nor U136991 ( n13622, n13624, n13625 );
nor U136992 ( n13624, P1_P1_INSTADDRPOINTER_REG_13_, n13634 );
nor U136993 ( n13625, n13627, n74468 );
nor U136994 ( n13634, n13635, n13567 );
xor U136995 ( n42977, n45963, P2_P1_PHYADDRPOINTER_REG_14_ );
xor U136996 ( n63218, n66643, P2_P3_PHYADDRPOINTER_REG_24_ );
xor U136997 ( n29455, n32040, P1_P3_PHYADDRPOINTER_REG_24_ );
xor U136998 ( n22136, n24808, P1_P2_PHYADDRPOINTER_REG_24_ );
xor U136999 ( n55246, n57942, P2_P2_PHYADDRPOINTER_REG_24_ );
nor U137000 ( n13923, n13932, n13933 );
nor U137001 ( n13932, P1_P1_INSTADDRPOINTER_REG_7_, n13942 );
nor U137002 ( n13933, n13934, n74658 );
nor U137003 ( n13942, n13943, n13890 );
nand U137004 ( n67786, n67749, n67831 );
nand U137005 ( n67831, n67832, P2_P3_INSTADDRPOINTER_REG_19_ );
nand U137006 ( n33031, n32993, n33075 );
nand U137007 ( n33075, n33076, P1_P3_INSTADDRPOINTER_REG_19_ );
nand U137008 ( n25783, n25744, n25828 );
nand U137009 ( n25828, n25829, P1_P2_INSTADDRPOINTER_REG_19_ );
nand U137010 ( n58921, n58884, n58966 );
nand U137011 ( n58966, n58967, P2_P2_INSTADDRPOINTER_REG_19_ );
nor U137012 ( n14208, n14254, n14255 );
nor U137013 ( n14254, P1_P1_INSTADDRPOINTER_REG_4_, n14265 );
nor U137014 ( n14255, n14257, n75941 );
nor U137015 ( n14265, n14267, n14268 );
nor U137016 ( n33199, n33207, n33208 );
nor U137017 ( n33208, n33209, n74845 );
nor U137018 ( n33207, P1_P3_INSTADDRPOINTER_REG_16_, n33216 );
nor U137019 ( n33209, n33210, n33211 );
nand U137020 ( n71005, n71006, n71007 );
nor U137021 ( n71006, n71010, n71011 );
nor U137022 ( n71007, n2359, n71008 );
nor U137023 ( n71011, P1_P1_ADDRESS_REG_2_, n71012 );
nor U137024 ( n67955, n67962, n67963 );
nor U137025 ( n67963, n67964, n73130 );
nor U137026 ( n67962, P2_P3_INSTADDRPOINTER_REG_16_, n67971 );
nor U137027 ( n67964, n67965, n67966 );
nor U137028 ( n46908, n46915, n46916 );
nor U137029 ( n46916, n46917, n73118 );
nor U137030 ( n46915, P2_P1_INSTADDRPOINTER_REG_16_, n46924 );
nor U137031 ( n46917, n46918, n46919 );
nor U137032 ( n25952, n25959, n25960 );
nor U137033 ( n25960, n25961, n73131 );
nor U137034 ( n25959, P1_P2_INSTADDRPOINTER_REG_16_, n25968 );
nor U137035 ( n25961, n25962, n25963 );
nor U137036 ( n59090, n59097, n59098 );
nor U137037 ( n59098, n59099, n73132 );
nor U137038 ( n59097, P2_P2_INSTADDRPOINTER_REG_16_, n59106 );
nor U137039 ( n59099, n59100, n59101 );
nor U137040 ( n13187, n13199, n13200 );
nor U137041 ( n13200, P1_P1_INSTADDRPOINTER_REG_22_, n13202 );
nor U137042 ( n13199, n13208, n74625 );
nor U137043 ( n13202, n13203, n13204 );
nand U137044 ( n29193, n35625, P1_P3_STATE2_REG_2_ );
nor U137045 ( n35625, P1_P3_STATE2_REG_1_, n74591 );
nor U137046 ( n32977, n32987, n32988 );
nor U137047 ( n32988, P1_P3_INSTADDRPOINTER_REG_22_, n32989 );
nor U137048 ( n32987, n32994, n74652 );
nor U137049 ( n32989, n32990, n32991 );
nor U137050 ( n67731, n67743, n67744 );
nor U137051 ( n67744, P2_P3_INSTADDRPOINTER_REG_22_, n67745 );
nor U137052 ( n67743, n67750, n74595 );
nor U137053 ( n67745, n67746, n67747 );
nor U137054 ( n25726, n25738, n25739 );
nor U137055 ( n25739, P1_P2_INSTADDRPOINTER_REG_22_, n25740 );
nor U137056 ( n25738, n25745, n74596 );
nor U137057 ( n25740, n25741, n25742 );
nor U137058 ( n58866, n58878, n58879 );
nor U137059 ( n58879, P2_P2_INSTADDRPOINTER_REG_22_, n58880 );
nor U137060 ( n58878, n58885, n74597 );
nor U137061 ( n58880, n58881, n58882 );
nand U137062 ( n71004, n71014, n71015 );
nor U137063 ( n71014, n71019, n71020 );
nor U137064 ( n71015, n1220, n71016 );
nor U137065 ( n71020, P2_P1_ADDRESS_REG_2_, n71021 );
nand U137066 ( n21992, n21993, n21994 );
nand U137067 ( n21994, n21975, n73317 );
nand U137068 ( n21993, P1_P2_REIP_REG_29_, n21987 );
nand U137069 ( n55102, n55103, n55104 );
nand U137070 ( n55104, n55085, n73316 );
nand U137071 ( n55103, P2_P2_REIP_REG_29_, n55097 );
nand U137072 ( n29311, n29312, n29313 );
nand U137073 ( n29313, n29290, n73318 );
nand U137074 ( n29312, P1_P3_REIP_REG_29_, n29302 );
nand U137075 ( n63074, n63075, n63076 );
nand U137076 ( n63076, n63057, n73319 );
nand U137077 ( n63075, P2_P3_REIP_REG_29_, n63069 );
xor U137078 ( n63341, n66695, P2_P3_PHYADDRPOINTER_REG_22_ );
xor U137079 ( n29512, n32092, P1_P3_PHYADDRPOINTER_REG_22_ );
xor U137080 ( n22193, n24860, P1_P2_PHYADDRPOINTER_REG_22_ );
xor U137081 ( n55307, n57994, P2_P2_PHYADDRPOINTER_REG_22_ );
nand U137082 ( n21876, n28446, P1_P2_STATE2_REG_2_ );
nor U137083 ( n28446, P1_P2_STATE2_REG_1_, n74592 );
nand U137084 ( n54967, n61751, P2_P2_STATE2_REG_2_ );
nor U137085 ( n61751, P2_P2_STATE2_REG_1_, n74594 );
nand U137086 ( n62911, n70351, P2_P3_STATE2_REG_2_ );
nor U137087 ( n70351, P2_P3_STATE2_REG_1_, n74593 );
xor U137088 ( n8402, n11760, P1_P1_PHYADDRPOINTER_REG_30_ );
xor U137089 ( n42807, n45834, P2_P1_PHYADDRPOINTER_REG_20_ );
nor U137090 ( n46572, P2_P1_INSTADDRPOINTER_REG_24_, n7470 );
nor U137091 ( n67619, P2_P3_INSTADDRPOINTER_REG_24_, n5685 );
nor U137092 ( n25614, P1_P2_INSTADDRPOINTER_REG_24_, n3928 );
nor U137093 ( n58751, P2_P2_INSTADDRPOINTER_REG_24_, n6560 );
nor U137094 ( n33312, n33327, n33328 );
nor U137095 ( n33328, n33329, n74460 );
nor U137096 ( n33327, P1_P3_INSTADDRPOINTER_REG_13_, n33335 );
nor U137097 ( n33329, n33330, n33331 );
nand U137098 ( n67611, P2_P3_INSTADDRPOINTER_REG_25_, n67612 );
nand U137099 ( n67612, n67613, n67614 );
nor U137100 ( n67614, n5730, n67615 );
nor U137101 ( n67613, n67618, n67619 );
nand U137102 ( n25606, P1_P2_INSTADDRPOINTER_REG_25_, n25607 );
nand U137103 ( n25607, n25608, n25609 );
nor U137104 ( n25609, n3973, n25610 );
nor U137105 ( n25608, n25613, n25614 );
nand U137106 ( n58743, P2_P2_INSTADDRPOINTER_REG_25_, n58744 );
nand U137107 ( n58744, n58745, n58746 );
nor U137108 ( n58746, n6605, n58747 );
nor U137109 ( n58745, n58750, n58751 );
nand U137110 ( n46564, P2_P1_INSTADDRPOINTER_REG_25_, n46565 );
nand U137111 ( n46565, n46566, n46567 );
nor U137112 ( n46567, n7515, n46568 );
nor U137113 ( n46566, n46571, n46572 );
nor U137114 ( n67853, P2_P3_INSTADDRPOINTER_REG_18_, n5685 );
nor U137115 ( n46806, P2_P1_INSTADDRPOINTER_REG_18_, n7470 );
nor U137116 ( n25850, P1_P2_INSTADDRPOINTER_REG_18_, n3928 );
nor U137117 ( n58988, P2_P2_INSTADDRPOINTER_REG_18_, n6560 );
nor U137118 ( n32854, P1_P3_INSTADDRPOINTER_REG_24_, n3084 );
nand U137119 ( n32846, P1_P3_INSTADDRPOINTER_REG_25_, n32847 );
nand U137120 ( n32847, n32848, n32849 );
nor U137121 ( n32849, n3129, n32850 );
nor U137122 ( n32848, n32853, n32854 );
nor U137123 ( n68069, n68084, n68085 );
nor U137124 ( n68085, n68086, n73104 );
nor U137125 ( n68084, P2_P3_INSTADDRPOINTER_REG_13_, n68092 );
nor U137126 ( n68086, n68087, n68088 );
nor U137127 ( n47038, n47053, n47054 );
nor U137128 ( n47054, n47055, n73099 );
nor U137129 ( n47053, P2_P1_INSTADDRPOINTER_REG_13_, n47061 );
nor U137130 ( n47055, n47056, n47057 );
nor U137131 ( n26066, n26081, n26082 );
nor U137132 ( n26082, n26083, n73105 );
nor U137133 ( n26081, P1_P2_INSTADDRPOINTER_REG_13_, n26089 );
nor U137134 ( n26083, n26084, n26085 );
nor U137135 ( n59207, n59222, n59223 );
nor U137136 ( n59223, n59224, n73106 );
nor U137137 ( n59222, P2_P2_INSTADDRPOINTER_REG_13_, n59230 );
nor U137138 ( n59224, n59225, n59226 );
nand U137139 ( n46798, P2_P1_INSTADDRPOINTER_REG_19_, n46799 );
nand U137140 ( n46799, n46800, n46801 );
nor U137141 ( n46801, n46802, n46803 );
nor U137142 ( n46800, n46805, n46806 );
nand U137143 ( n67845, P2_P3_INSTADDRPOINTER_REG_19_, n67846 );
nand U137144 ( n67846, n67847, n67848 );
nor U137145 ( n67848, n67849, n67850 );
nor U137146 ( n67847, n67852, n67853 );
nand U137147 ( n25842, P1_P2_INSTADDRPOINTER_REG_19_, n25843 );
nand U137148 ( n25843, n25844, n25845 );
nor U137149 ( n25845, n25846, n25847 );
nor U137150 ( n25844, n25849, n25850 );
nand U137151 ( n58980, P2_P2_INSTADDRPOINTER_REG_19_, n58981 );
nand U137152 ( n58981, n58982, n58983 );
nor U137153 ( n58983, n58984, n58985 );
nor U137154 ( n58982, n58987, n58988 );
nor U137155 ( n33097, P1_P3_INSTADDRPOINTER_REG_18_, n3084 );
nand U137156 ( n13255, n13207, n13308 );
nand U137157 ( n13308, n13309, P1_P1_INSTADDRPOINTER_REG_19_ );
nand U137158 ( n33089, P1_P3_INSTADDRPOINTER_REG_19_, n33090 );
nand U137159 ( n33090, n33091, n33092 );
nor U137160 ( n33092, n33093, n33094 );
nor U137161 ( n33091, n33096, n33097 );
nand U137162 ( n46739, n46702, n46784 );
nand U137163 ( n46784, n46785, P2_P1_INSTADDRPOINTER_REG_19_ );
nor U137164 ( n47294, n47301, n47302 );
nor U137165 ( n47302, n47303, n74659 );
nor U137166 ( n47301, P2_P1_INSTADDRPOINTER_REG_7_, n47309 );
nor U137167 ( n47303, n47304, n47305 );
nor U137168 ( n68325, n68332, n68333 );
nor U137169 ( n68333, n68334, n74695 );
nor U137170 ( n68332, P2_P3_INSTADDRPOINTER_REG_7_, n68340 );
nor U137171 ( n68334, n68335, n68336 );
nor U137172 ( n33569, n33576, n33577 );
nor U137173 ( n33577, n33578, n74696 );
nor U137174 ( n33576, P1_P3_INSTADDRPOINTER_REG_7_, n33584 );
nor U137175 ( n33578, n33579, n33580 );
nor U137176 ( n26324, n26331, n26332 );
nor U137177 ( n26332, n26333, n74697 );
nor U137178 ( n26331, P1_P2_INSTADDRPOINTER_REG_7_, n26339 );
nor U137179 ( n26333, n26334, n26335 );
nor U137180 ( n59463, n59470, n59471 );
nor U137181 ( n59471, n59472, n74698 );
nor U137182 ( n59470, P2_P2_INSTADDRPOINTER_REG_7_, n59478 );
nor U137183 ( n59472, n59473, n59474 );
nor U137184 ( n46684, n46696, n46697 );
nor U137185 ( n46697, P2_P1_INSTADDRPOINTER_REG_22_, n46698 );
nor U137186 ( n46696, n46703, n74585 );
nor U137187 ( n46698, n46699, n46700 );
nor U137188 ( n42492, P2_P1_REIP_REG_31_, n508 );
nand U137189 ( n46010, n46011, P2_P1_PHYADDRPOINTER_REG_12_ );
nand U137190 ( n33432, P1_P3_INSTADDRPOINTER_REG_10_, n33433 );
nand U137191 ( n33433, n33434, n33435 );
nor U137192 ( n33435, n33356, n33436 );
nor U137193 ( n33434, n33437, n33438 );
nor U137194 ( n33437, P1_P3_INSTADDRPOINTER_REG_9_, n3084 );
and U137195 ( n14063, n14064, P1_P1_INSTADDRPOINTER_REG_5_ );
nor U137196 ( n47153, P2_P1_INSTADDRPOINTER_REG_9_, n7470 );
nor U137197 ( n68184, P2_P3_INSTADDRPOINTER_REG_9_, n5685 );
nor U137198 ( n26183, P1_P2_INSTADDRPOINTER_REG_9_, n3928 );
nor U137199 ( n59322, P2_P2_INSTADDRPOINTER_REG_9_, n6560 );
nand U137200 ( n68179, P2_P3_INSTADDRPOINTER_REG_10_, n68180 );
nand U137201 ( n68180, n68181, n68182 );
nor U137202 ( n68182, n68113, n68183 );
nor U137203 ( n68181, n68184, n68185 );
nand U137204 ( n26178, P1_P2_INSTADDRPOINTER_REG_10_, n26179 );
nand U137205 ( n26179, n26180, n26181 );
nor U137206 ( n26181, n26110, n26182 );
nor U137207 ( n26180, n26183, n26184 );
nand U137208 ( n59317, P2_P2_INSTADDRPOINTER_REG_10_, n59318 );
nand U137209 ( n59318, n59319, n59320 );
nor U137210 ( n59320, n59251, n59321 );
nor U137211 ( n59319, n59322, n59323 );
nand U137212 ( n47148, P2_P1_INSTADDRPOINTER_REG_10_, n47149 );
nand U137213 ( n47149, n47150, n47151 );
nor U137214 ( n47151, n47082, n47152 );
nor U137215 ( n47150, n47153, n47154 );
and U137216 ( n68690, n75970, n75971 );
nand U137217 ( n75970, n68675, P2_P3_INSTADDRPOINTER_REG_2_ );
nand U137218 ( n75971, n67200, n76705 );
and U137219 ( n33934, n75972, n75973 );
nand U137220 ( n75972, n33919, P1_P3_INSTADDRPOINTER_REG_2_ );
nand U137221 ( n75973, n32544, n76772 );
and U137222 ( n26689, n75974, n75975 );
nand U137223 ( n75974, n26674, P1_P2_INSTADDRPOINTER_REG_2_ );
nand U137224 ( n75975, n25302, n76751 );
and U137225 ( n59831, n75976, n75977 );
nand U137226 ( n75976, n59816, P2_P2_INSTADDRPOINTER_REG_2_ );
nand U137227 ( n75977, n58441, n76684 );
nor U137228 ( n8404, P1_P1_REIP_REG_31_, n237 );
nor U137229 ( n68555, n68592, n68593 );
nor U137230 ( n68592, P2_P3_INSTADDRPOINTER_REG_4_, n68601 );
nor U137231 ( n68593, n68594, n75937 );
nor U137232 ( n68601, n68602, n68603 );
nor U137233 ( n33799, n33836, n33837 );
nor U137234 ( n33836, P1_P3_INSTADDRPOINTER_REG_4_, n33845 );
nor U137235 ( n33837, n33838, n75940 );
nor U137236 ( n33845, n33846, n33847 );
nor U137237 ( n47534, n47571, n47572 );
nor U137238 ( n47571, P2_P1_INSTADDRPOINTER_REG_4_, n47580 );
nor U137239 ( n47572, n47573, n75934 );
nor U137240 ( n47580, n47581, n47582 );
nor U137241 ( n26554, n26591, n26592 );
nor U137242 ( n26591, P1_P2_INSTADDRPOINTER_REG_4_, n26600 );
nor U137243 ( n26592, n26593, n75938 );
nor U137244 ( n26600, n26601, n26602 );
nor U137245 ( n59696, n59733, n59734 );
nor U137246 ( n59733, P2_P2_INSTADDRPOINTER_REG_4_, n59742 );
nor U137247 ( n59734, n59735, n75939 );
nor U137248 ( n59742, n59743, n59744 );
nor U137249 ( n13635, n13639, n74476 );
nor U137250 ( n13639, n13640, n13642 );
nor U137251 ( n13640, n13643, n13644 );
nand U137252 ( n13644, P1_P1_INSTADDRPOINTER_REG_11_, n12999 );
nor U137253 ( n13943, n13945, n73090 );
nor U137254 ( n13945, n13947, n13948 );
nor U137255 ( n13947, n13889, n13949 );
nand U137256 ( n13949, P1_P1_INSTADDRPOINTER_REG_5_, n12999 );
xor U137257 ( n8957, n12282, P1_P1_PHYADDRPOINTER_REG_14_ );
xor U137258 ( n63615, n66914, P2_P3_PHYADDRPOINTER_REG_14_ );
xor U137259 ( n29716, n32275, P1_P3_PHYADDRPOINTER_REG_14_ );
xor U137260 ( n22395, n25038, P1_P2_PHYADDRPOINTER_REG_14_ );
xor U137261 ( n55507, n58173, P2_P2_PHYADDRPOINTER_REG_14_ );
and U137262 ( n14385, n75978, n75979 );
nand U137263 ( n75978, n14358, P1_P1_INSTADDRPOINTER_REG_2_ );
nand U137264 ( n75979, n12625, n76727 );
nand U137265 ( n45879, n45880, P2_P1_PHYADDRPOINTER_REG_18_ );
xor U137266 ( n43231, n43232, n43233 );
xor U137267 ( n43233, n43230, P3_REG1_REG_9_ );
nor U137268 ( n33143, n33106, n33170 );
and U137269 ( n33170, n33171, P1_P3_INSTADDRPOINTER_REG_16_ );
nor U137270 ( n67899, n67862, n67933 );
and U137271 ( n67933, n67934, P2_P3_INSTADDRPOINTER_REG_16_ );
nor U137272 ( n46852, n46815, n46886 );
and U137273 ( n46886, n46887, P2_P1_INSTADDRPOINTER_REG_16_ );
nor U137274 ( n25896, n25859, n25930 );
and U137275 ( n25930, n25931, P1_P2_INSTADDRPOINTER_REG_16_ );
nor U137276 ( n59034, n58997, n59068 );
and U137277 ( n59068, n59069, P2_P2_INSTADDRPOINTER_REG_16_ );
nand U137278 ( n42985, P2_P1_EBX_REG_14_, n500 );
nand U137279 ( n43039, P2_P1_EBX_REG_12_, n500 );
nand U137280 ( n43091, P2_P1_EBX_REG_10_, n500 );
nand U137281 ( n43141, P2_P1_EBX_REG_8_, n500 );
nand U137282 ( n43265, P2_P1_EBX_REG_4_, n500 );
nand U137283 ( n43314, P2_P1_EBX_REG_2_, n500 );
nand U137284 ( n42870, P2_P1_EBX_REG_18_, n500 );
nand U137285 ( n42921, P2_P1_EBX_REG_16_, n500 );
nand U137286 ( n43195, P2_P1_EBX_REG_6_, n500 );
xor U137287 ( n63459, n66785, P2_P3_PHYADDRPOINTER_REG_20_ );
xor U137288 ( n29556, n32139, P1_P3_PHYADDRPOINTER_REG_20_ );
xor U137289 ( n22239, n24907, P1_P2_PHYADDRPOINTER_REG_20_ );
xor U137290 ( n55351, n58044, P2_P2_PHYADDRPOINTER_REG_20_ );
xnor U137291 ( n43309, n74467, P2_P1_PHYADDRPOINTER_REG_2_ );
nor U137292 ( n21324, n5165, n21338 );
nor U137293 ( n21338, n74435, P1_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U137294 ( n68801, n68802, P2_P3_INSTADDRPOINTER_REG_1_ );
nor U137295 ( n68802, P2_P3_INSTADDRPOINTER_REG_0_, n5708 );
nand U137296 ( n34045, n34046, P1_P3_INSTADDRPOINTER_REG_1_ );
nor U137297 ( n34046, P1_P3_INSTADDRPOINTER_REG_0_, n3107 );
nand U137298 ( n26802, n26803, P1_P2_INSTADDRPOINTER_REG_1_ );
nor U137299 ( n26803, P1_P2_INSTADDRPOINTER_REG_0_, n3950 );
nand U137300 ( n59942, n59943, P2_P2_INSTADDRPOINTER_REG_1_ );
nor U137301 ( n59943, P2_P2_INSTADDRPOINTER_REG_0_, n6583 );
and U137302 ( n47669, n75980, n75981 );
nand U137303 ( n75980, n47654, P2_P1_INSTADDRPOINTER_REG_2_ );
nand U137304 ( n75981, n46248, n76657 );
xnor U137305 ( n64055, n74469, P2_P3_PHYADDRPOINTER_REG_2_ );
xnor U137306 ( n30038, n74470, P1_P3_PHYADDRPOINTER_REG_2_ );
xnor U137307 ( n22715, n74471, P1_P2_PHYADDRPOINTER_REG_2_ );
xnor U137308 ( n55831, n74472, P2_P2_PHYADDRPOINTER_REG_2_ );
nand U137309 ( n8967, P1_P1_EBX_REG_14_, n229 );
nand U137310 ( n9034, P1_P1_EBX_REG_12_, n229 );
nand U137311 ( n9099, P1_P1_EBX_REG_10_, n229 );
nand U137312 ( n9162, P1_P1_EBX_REG_8_, n229 );
nand U137313 ( n9299, P1_P1_EBX_REG_4_, n229 );
nand U137314 ( n9360, P1_P1_EBX_REG_2_, n229 );
nand U137315 ( n8840, P1_P1_EBX_REG_18_, n229 );
nand U137316 ( n8904, P1_P1_EBX_REG_16_, n229 );
nand U137317 ( n9229, P1_P1_EBX_REG_6_, n229 );
nand U137318 ( n42613, n42614, n42615 );
nand U137319 ( n42614, P2_P1_REIP_REG_26_, n42608 );
nand U137320 ( n42615, n505, n73308 );
nand U137321 ( n43053, n43054, n43055 );
nand U137322 ( n43054, n7393, P2_P1_PHYADDRPOINTER_REG_11_ );
nand U137323 ( n43055, P2_P1_REIP_REG_11_, n43041 );
nand U137324 ( n43209, n43210, n43211 );
nand U137325 ( n43210, n7393, P2_P1_PHYADDRPOINTER_REG_5_ );
nand U137326 ( n43211, P2_P1_REIP_REG_5_, n43197 );
xor U137327 ( n8762, n12104, P1_P1_PHYADDRPOINTER_REG_20_ );
nand U137328 ( n43142, P2_P1_REIP_REG_8_, n43111 );
nand U137329 ( n42888, P2_P1_REIP_REG_17_, n42872 );
nand U137330 ( n42986, P2_P1_REIP_REG_14_, n42940 );
nand U137331 ( n8554, n8555, n8557 );
nand U137332 ( n8555, P1_P1_REIP_REG_26_, n8548 );
nand U137333 ( n8557, n234, n73309 );
nand U137334 ( n9052, n9053, n9054 );
nand U137335 ( n9053, n4751, P1_P1_PHYADDRPOINTER_REG_11_ );
nand U137336 ( n9054, P1_P1_REIP_REG_11_, n9037 );
nand U137337 ( n9247, n9248, n9249 );
nand U137338 ( n9248, n4751, P1_P1_PHYADDRPOINTER_REG_5_ );
nand U137339 ( n9249, P1_P1_REIP_REG_5_, n9232 );
xor U137340 ( n22013, n24648, P1_P2_PHYADDRPOINTER_REG_29_ );
xor U137341 ( n29332, n31862, P1_P3_PHYADDRPOINTER_REG_29_ );
xor U137342 ( n63095, n66485, P2_P3_PHYADDRPOINTER_REG_29_ );
xor U137343 ( n55123, n57784, P2_P2_PHYADDRPOINTER_REG_29_ );
nand U137344 ( n9163, P1_P1_REIP_REG_8_, n9124 );
nor U137345 ( n54307, n7820, n54321 );
nor U137346 ( n54321, n74442, P2_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U137347 ( n8863, P1_P1_REIP_REG_17_, n8843 );
nand U137348 ( n8968, P1_P1_REIP_REG_14_, n8928 );
nand U137349 ( n12327, n12328, P1_P1_PHYADDRPOINTER_REG_12_ );
nand U137350 ( n47780, n47781, P2_P1_INSTADDRPOINTER_REG_1_ );
nor U137351 ( n47781, P2_P1_INSTADDRPOINTER_REG_0_, n7494 );
nand U137352 ( n23354, n23450, P1_P2_EAX_REG_22_ );
nor U137353 ( n23450, n23451, n74923 );
nand U137354 ( n23595, n23683, P1_P2_EAX_REG_18_ );
nor U137355 ( n23683, n23684, n74820 );
nand U137356 ( n23451, n23594, P1_P2_EAX_REG_20_ );
nor U137357 ( n23594, n23595, n74878 );
nand U137358 ( n56573, n56716, P2_P2_EAX_REG_20_ );
nor U137359 ( n56716, n56717, n74877 );
nand U137360 ( n56383, n56477, P2_P2_EAX_REG_24_ );
nor U137361 ( n56477, n56478, n74971 );
nand U137362 ( n56478, n56572, P2_P2_EAX_REG_22_ );
nor U137363 ( n56572, n56573, n74922 );
nand U137364 ( n56717, n56805, P2_P2_EAX_REG_18_ );
nor U137365 ( n56805, n56806, n74819 );
nand U137366 ( n23259, n23353, P1_P2_EAX_REG_24_ );
nor U137367 ( n23353, n23354, n74972 );
nand U137368 ( n23684, n23772, P1_P2_EAX_REG_16_ );
nor U137369 ( n23772, n23773, n74780 );
nand U137370 ( n56806, n56897, P2_P2_EAX_REG_16_ );
nor U137371 ( n56897, n56898, n74779 );
nand U137372 ( n23773, n23934, P1_P2_EAX_REG_14_ );
nor U137373 ( n23934, n23935, n74733 );
nand U137374 ( n56898, n57058, P2_P2_EAX_REG_14_ );
nor U137375 ( n57058, n57059, n74732 );
nand U137376 ( n23207, n23258, P1_P2_EAX_REG_26_ );
nor U137377 ( n23258, n23259, n75037 );
nand U137378 ( n56328, n56382, P2_P2_EAX_REG_26_ );
nor U137379 ( n56382, n56383, n75036 );
nand U137380 ( n57108, n57188, P2_P2_EAX_REG_9_ );
nor U137381 ( n57188, n57189, n74632 );
nand U137382 ( n23986, n24066, P1_P2_EAX_REG_9_ );
nor U137383 ( n24066, n24067, n74633 );
nand U137384 ( n57392, n57412, P2_P2_EAX_REG_2_ );
nor U137385 ( n57412, n74490, n73128 );
nand U137386 ( n57371, n57391, P2_P2_EAX_REG_4_ );
nor U137387 ( n57391, n57392, n74509 );
nand U137388 ( n57270, n57370, P2_P2_EAX_REG_6_ );
nor U137389 ( n57370, n57371, n74542 );
nand U137390 ( n24267, n24289, P1_P2_EAX_REG_2_ );
nor U137391 ( n24289, n74491, n73129 );
nand U137392 ( n57189, n57269, P2_P2_EAX_REG_8_ );
nor U137393 ( n57269, n57270, n74583 );
nand U137394 ( n24246, n24266, P1_P2_EAX_REG_4_ );
nor U137395 ( n24266, n24267, n74510 );
nand U137396 ( n24148, n24245, P1_P2_EAX_REG_6_ );
nor U137397 ( n24245, n24246, n74543 );
nand U137398 ( n57059, n57107, P2_P2_EAX_REG_12_ );
nor U137399 ( n57107, n57108, n74678 );
nand U137400 ( n24067, n24147, P1_P2_EAX_REG_8_ );
nor U137401 ( n24147, n24148, n74584 );
nand U137402 ( n23935, n23985, P1_P2_EAX_REG_12_ );
nor U137403 ( n23985, n23986, n74679 );
nand U137404 ( n64739, n64874, P2_P3_EAX_REG_24_ );
nor U137405 ( n64874, n64875, n74968 );
nand U137406 ( n64875, n64963, P2_P3_EAX_REG_22_ );
nor U137407 ( n64963, n64964, n74921 );
nand U137408 ( n64964, n65103, P2_P3_EAX_REG_20_ );
nor U137409 ( n65103, n65104, n74875 );
nand U137410 ( n65104, n65188, P2_P3_EAX_REG_18_ );
nor U137411 ( n65188, n65189, n74814 );
nand U137412 ( n65189, n65273, P2_P3_EAX_REG_16_ );
nor U137413 ( n65273, n65274, n74776 );
nand U137414 ( n65274, n65431, P2_P3_EAX_REG_14_ );
nor U137415 ( n65431, n65432, n74730 );
nand U137416 ( n64691, n64738, P2_P3_EAX_REG_26_ );
nor U137417 ( n64738, n64739, n75028 );
nand U137418 ( n65530, n65610, P2_P3_EAX_REG_9_ );
nor U137419 ( n65610, n65611, n74628 );
nand U137420 ( n65851, n65871, P2_P3_EAX_REG_2_ );
nor U137421 ( n65871, n74487, n73127 );
nand U137422 ( n65790, n65850, P2_P3_EAX_REG_4_ );
nor U137423 ( n65850, n65851, n74507 );
nand U137424 ( n65692, n65789, P2_P3_EAX_REG_6_ );
nor U137425 ( n65789, n65790, n74539 );
nand U137426 ( n65611, n65691, P2_P3_EAX_REG_8_ );
nor U137427 ( n65691, n65692, n74581 );
nand U137428 ( n65432, n65529, P2_P3_EAX_REG_12_ );
nor U137429 ( n65529, n65530, n74675 );
nor U137430 ( n64074, P2_P3_EBX_REG_1_, n63034 );
nor U137431 ( n30057, P1_P3_EBX_REG_1_, n29267 );
nor U137432 ( n22734, P1_P2_EBX_REG_1_, n21950 );
nor U137433 ( n55850, P2_P2_EBX_REG_1_, n55062 );
nand U137434 ( n64064, n64072, n64073 );
nand U137435 ( n64072, n5632, n64075 );
nand U137436 ( n64073, n64074, P2_P3_EBX_REG_0_ );
nand U137437 ( n64075, n64076, n64077 );
nand U137438 ( n30047, n30055, n30056 );
nand U137439 ( n30055, n3030, n30058 );
nand U137440 ( n30056, n30057, P1_P3_EBX_REG_0_ );
nand U137441 ( n30058, n30059, n30060 );
nand U137442 ( n22724, n22732, n22733 );
nand U137443 ( n22732, n3874, n22735 );
nand U137444 ( n22733, n22734, P1_P2_EBX_REG_0_ );
nand U137445 ( n22735, n22736, n22737 );
nand U137446 ( n55840, n55848, n55849 );
nand U137447 ( n55848, n6507, n55851 );
nand U137448 ( n55849, n55850, P2_P2_EBX_REG_0_ );
nand U137449 ( n55851, n55852, n55853 );
nand U137450 ( n30987, n31071, P1_P3_EAX_REG_16_ );
nor U137451 ( n31071, n31072, n74778 );
nand U137452 ( n30902, n30986, P1_P3_EAX_REG_18_ );
nor U137453 ( n30986, n30987, n74817 );
nand U137454 ( n30580, n30668, P1_P3_EAX_REG_24_ );
nor U137455 ( n30668, n30669, n74984 );
nand U137456 ( n30669, n30761, P1_P3_EAX_REG_22_ );
nor U137457 ( n30761, n30762, n74927 );
nand U137458 ( n30762, n30901, P1_P3_EAX_REG_20_ );
nor U137459 ( n30901, n30902, n74876 );
nand U137460 ( n31072, n31177, P1_P3_EAX_REG_14_ );
nor U137461 ( n31177, n31178, n74731 );
nand U137462 ( n31280, n31360, P1_P3_EAX_REG_9_ );
nor U137463 ( n31360, n31361, n74629 );
nand U137464 ( n31561, n31585, P1_P3_EAX_REG_2_ );
nor U137465 ( n31585, n74488, n72957 );
nand U137466 ( n31540, n31560, P1_P3_EAX_REG_4_ );
nor U137467 ( n31560, n31561, n73135 );
nand U137468 ( n31442, n31539, P1_P3_EAX_REG_6_ );
nor U137469 ( n31539, n31540, n74540 );
nand U137470 ( n31361, n31441, P1_P3_EAX_REG_8_ );
nor U137471 ( n31441, n31442, n74582 );
nand U137472 ( n31178, n31279, P1_P3_EAX_REG_12_ );
nor U137473 ( n31279, n31280, n74676 );
nand U137474 ( n30532, n30579, P1_P3_EAX_REG_26_ );
nor U137475 ( n30579, n30580, n75041 );
nand U137476 ( n67783, n67784, n73149 );
nand U137477 ( n67784, n67710, n67785 );
nand U137478 ( n67785, P2_P3_INSTADDRPOINTER_REG_20_, n67786 );
nand U137479 ( n25780, n25781, n73150 );
nand U137480 ( n25781, n25705, n25782 );
nand U137481 ( n25782, P1_P2_INSTADDRPOINTER_REG_20_, n25783 );
nand U137482 ( n58918, n58919, n73151 );
nand U137483 ( n58919, n58845, n58920 );
nand U137484 ( n58920, P2_P2_INSTADDRPOINTER_REG_20_, n58921 );
nand U137485 ( n33028, n33029, n73167 );
nand U137486 ( n33029, n32956, n33030 );
nand U137487 ( n33030, P1_P3_INSTADDRPOINTER_REG_20_, n33031 );
nand U137488 ( n42532, n42533, n42534 );
nand U137489 ( n42534, n42517, n73391 );
nand U137490 ( n42533, P2_P1_REIP_REG_29_, n42528 );
nand U137491 ( n45681, n45733, P2_P1_PHYADDRPOINTER_REG_23_ );
nand U137492 ( n11945, n12000, P1_P1_PHYADDRPOINTER_REG_23_ );
nand U137493 ( n11845, n11909, P1_P1_PHYADDRPOINTER_REG_26_ );
nand U137494 ( n45592, n45656, P2_P1_PHYADDRPOINTER_REG_26_ );
nand U137495 ( n9822, n9905, P1_P1_EAX_REG_28_ );
nor U137496 ( n9905, n9907, n9908 );
nand U137497 ( n43739, n43806, P2_P1_EAX_REG_28_ );
nor U137498 ( n43806, n43807, n43808 );
nand U137499 ( n63929, n64048, n73121 );
nor U137500 ( n64048, P2_P3_EBX_REG_2_, P2_P3_EBX_REG_1_ );
nand U137501 ( n29973, n30031, n73119 );
nor U137502 ( n30031, P1_P3_EBX_REG_2_, P1_P3_EBX_REG_1_ );
nand U137503 ( n22650, n22708, n73120 );
nor U137504 ( n22708, P1_P2_EBX_REG_2_, P1_P2_EBX_REG_1_ );
nand U137505 ( n55763, n55824, n73122 );
nor U137506 ( n55824, P2_P2_EBX_REG_2_, P2_P2_EBX_REG_1_ );
nand U137507 ( n63879, n63930, n6338 );
nor U137508 ( n63930, P2_P3_EBX_REG_4_, P2_P3_EBX_REG_3_ );
nand U137509 ( n29923, n29974, n3704 );
nor U137510 ( n29974, P1_P3_EBX_REG_4_, P1_P3_EBX_REG_3_ );
nand U137511 ( n22600, n22651, n4598 );
nor U137512 ( n22651, P1_P2_EBX_REG_4_, P1_P2_EBX_REG_3_ );
nand U137513 ( n55713, n55764, n7230 );
nor U137514 ( n55764, P2_P2_EBX_REG_4_, P2_P2_EBX_REG_3_ );
nand U137515 ( n63174, n63226, n6325 );
nor U137516 ( n63226, P2_P3_EBX_REG_24_, P2_P3_EBX_REG_23_ );
nand U137517 ( n63225, n63329, n6327 );
nor U137518 ( n63329, P2_P3_EBX_REG_22_, P2_P3_EBX_REG_21_ );
nand U137519 ( n63328, n63467, n6328 );
nor U137520 ( n63467, P2_P3_EBX_REG_20_, P2_P3_EBX_REG_19_ );
nand U137521 ( n63466, n63508, n6329 );
nor U137522 ( n63508, P2_P3_EBX_REG_18_, P2_P3_EBX_REG_17_ );
nand U137523 ( n63507, n63564, n6330 );
nor U137524 ( n63564, P2_P3_EBX_REG_16_, P2_P3_EBX_REG_15_ );
nand U137525 ( n63563, n63610, n6332 );
nor U137526 ( n63610, P2_P3_EBX_REG_14_, P2_P3_EBX_REG_13_ );
nand U137527 ( n63609, n63724, n6333 );
nor U137528 ( n63724, P2_P3_EBX_REG_12_, P2_P3_EBX_REG_11_ );
nand U137529 ( n63723, n63782, n6334 );
nor U137530 ( n63782, P2_P3_EBX_REG_9_, P2_P3_EBX_REG_10_ );
nand U137531 ( n63781, n63834, n6335 );
nor U137532 ( n63834, P2_P3_EBX_REG_8_, P2_P3_EBX_REG_7_ );
nand U137533 ( n63833, n63880, n6337 );
nor U137534 ( n63880, P2_P3_EBX_REG_6_, P2_P3_EBX_REG_5_ );
nand U137535 ( n29411, n29463, n3692 );
nor U137536 ( n29463, P1_P3_EBX_REG_24_, P1_P3_EBX_REG_23_ );
nand U137537 ( n29462, n29500, n3693 );
nor U137538 ( n29500, P1_P3_EBX_REG_22_, P1_P3_EBX_REG_21_ );
nand U137539 ( n29499, n29564, n3694 );
nor U137540 ( n29564, P1_P3_EBX_REG_20_, P1_P3_EBX_REG_19_ );
nand U137541 ( n29563, n29609, n3695 );
nor U137542 ( n29609, P1_P3_EBX_REG_18_, P1_P3_EBX_REG_17_ );
nand U137543 ( n29608, n29665, n3697 );
nor U137544 ( n29665, P1_P3_EBX_REG_16_, P1_P3_EBX_REG_15_ );
nand U137545 ( n29664, n29711, n3698 );
nor U137546 ( n29711, P1_P3_EBX_REG_14_, P1_P3_EBX_REG_13_ );
nand U137547 ( n29710, n29764, n3699 );
nor U137548 ( n29764, P1_P3_EBX_REG_12_, P1_P3_EBX_REG_11_ );
nand U137549 ( n29763, n29822, n3700 );
nor U137550 ( n29822, P1_P3_EBX_REG_9_, P1_P3_EBX_REG_10_ );
nand U137551 ( n29821, n29878, n3702 );
nor U137552 ( n29878, P1_P3_EBX_REG_8_, P1_P3_EBX_REG_7_ );
nand U137553 ( n29877, n29924, n3703 );
nor U137554 ( n29924, P1_P3_EBX_REG_6_, P1_P3_EBX_REG_5_ );
nand U137555 ( n22092, n22144, n4585 );
nor U137556 ( n22144, P1_P2_EBX_REG_24_, P1_P2_EBX_REG_23_ );
nand U137557 ( n22246, n22288, n4589 );
nor U137558 ( n22288, P1_P2_EBX_REG_18_, P1_P2_EBX_REG_17_ );
nand U137559 ( n22389, n22443, n4593 );
nor U137560 ( n22443, P1_P2_EBX_REG_12_, P1_P2_EBX_REG_11_ );
nand U137561 ( n22502, n22555, n4595 );
nor U137562 ( n22555, P1_P2_EBX_REG_8_, P1_P2_EBX_REG_7_ );
nand U137563 ( n22554, n22601, n4597 );
nor U137564 ( n22601, P1_P2_EBX_REG_6_, P1_P2_EBX_REG_5_ );
nand U137565 ( n22143, n22181, n4587 );
nor U137566 ( n22181, P1_P2_EBX_REG_22_, P1_P2_EBX_REG_21_ );
nand U137567 ( n22287, n22344, n4590 );
nor U137568 ( n22344, P1_P2_EBX_REG_16_, P1_P2_EBX_REG_15_ );
nand U137569 ( n22343, n22390, n4592 );
nor U137570 ( n22390, P1_P2_EBX_REG_14_, P1_P2_EBX_REG_13_ );
nand U137571 ( n22442, n22503, n4594 );
nor U137572 ( n22503, P1_P2_EBX_REG_9_, P1_P2_EBX_REG_10_ );
nand U137573 ( n55202, n55254, n7218 );
nor U137574 ( n55254, P2_P2_EBX_REG_24_, P2_P2_EBX_REG_23_ );
nand U137575 ( n55358, n55400, n7222 );
nor U137576 ( n55400, P2_P2_EBX_REG_18_, P2_P2_EBX_REG_17_ );
nand U137577 ( n55501, n55558, n7225 );
nor U137578 ( n55558, P2_P2_EBX_REG_12_, P2_P2_EBX_REG_11_ );
nand U137579 ( n55615, n55668, n7228 );
nor U137580 ( n55668, P2_P2_EBX_REG_8_, P2_P2_EBX_REG_7_ );
nand U137581 ( n55667, n55714, n7229 );
nor U137582 ( n55714, P2_P2_EBX_REG_6_, P2_P2_EBX_REG_5_ );
nand U137583 ( n55253, n55295, n7219 );
nor U137584 ( n55295, P2_P2_EBX_REG_22_, P2_P2_EBX_REG_21_ );
nand U137585 ( n55399, n55456, n7223 );
nor U137586 ( n55456, P2_P2_EBX_REG_16_, P2_P2_EBX_REG_15_ );
nand U137587 ( n55455, n55502, n7224 );
nor U137588 ( n55502, P2_P2_EBX_REG_14_, P2_P2_EBX_REG_13_ );
nand U137589 ( n55557, n55616, n7227 );
nor U137590 ( n55616, P2_P2_EBX_REG_9_, P2_P2_EBX_REG_10_ );
nand U137591 ( n63109, n63175, n6324 );
nor U137592 ( n63175, P2_P3_EBX_REG_26_, P2_P3_EBX_REG_25_ );
nand U137593 ( n29346, n29412, n3690 );
nor U137594 ( n29412, P1_P3_EBX_REG_26_, P1_P3_EBX_REG_25_ );
nand U137595 ( n22027, n22093, n4584 );
nor U137596 ( n22093, P1_P2_EBX_REG_26_, P1_P2_EBX_REG_25_ );
nand U137597 ( n22180, n22247, n4588 );
nor U137598 ( n22247, P1_P2_EBX_REG_20_, P1_P2_EBX_REG_19_ );
nand U137599 ( n55137, n55203, n7217 );
nor U137600 ( n55203, P2_P2_EBX_REG_26_, P2_P2_EBX_REG_25_ );
nand U137601 ( n55294, n55359, n7220 );
nor U137602 ( n55359, P2_P2_EBX_REG_20_, P2_P2_EBX_REG_19_ );
and U137603 ( n22009, n22028, n4583 );
nor U137604 ( n22028, P1_P2_EBX_REG_28_, P1_P2_EBX_REG_27_ );
and U137605 ( n29328, n29347, n3689 );
nor U137606 ( n29347, P1_P3_EBX_REG_28_, P1_P3_EBX_REG_27_ );
and U137607 ( n63091, n63110, n6323 );
nor U137608 ( n63110, P2_P3_EBX_REG_28_, P2_P3_EBX_REG_27_ );
and U137609 ( n55119, n55138, n7215 );
nor U137610 ( n55138, P2_P2_EBX_REG_28_, P2_P2_EBX_REG_27_ );
nand U137611 ( n12103, P1_P1_PHYADDRPOINTER_REG_19_, P1_P1_PHYADDRPOINTER_REG_18_ );
nand U137612 ( n8455, P1_P1_REIP_REG_29_, n8449 );
nand U137613 ( n66950, n66951, P2_P3_PHYADDRPOINTER_REG_12_ );
nand U137614 ( n32311, n32312, P1_P3_PHYADDRPOINTER_REG_12_ );
nand U137615 ( n25074, n25075, P1_P2_PHYADDRPOINTER_REG_12_ );
nand U137616 ( n58209, n58210, P2_P2_PHYADDRPOINTER_REG_12_ );
nand U137617 ( n46736, n46737, n73148 );
nand U137618 ( n46737, n46663, n46738 );
nand U137619 ( n46738, P2_P1_INSTADDRPOINTER_REG_20_, n46739 );
nand U137620 ( n13252, n13253, n73158 );
nand U137621 ( n13253, n13152, n13254 );
nand U137622 ( n13254, P1_P1_INSTADDRPOINTER_REG_20_, n13255 );
nand U137623 ( n12165, n12167, P1_P1_PHYADDRPOINTER_REG_18_ );
nand U137624 ( n14524, n14525, P1_P1_INSTADDRPOINTER_REG_1_ );
nor U137625 ( n14525, P1_P1_INSTADDRPOINTER_REG_0_, n4850 );
nand U137626 ( n24682, n24745, P1_P2_PHYADDRPOINTER_REG_26_ );
nand U137627 ( n31894, n31977, P1_P3_PHYADDRPOINTER_REG_26_ );
nand U137628 ( n66517, n66580, P2_P3_PHYADDRPOINTER_REG_26_ );
nand U137629 ( n57816, n57879, P2_P2_PHYADDRPOINTER_REG_26_ );
nand U137630 ( n66605, n66659, P2_P3_PHYADDRPOINTER_REG_23_ );
nand U137631 ( n32002, n32056, P1_P3_PHYADDRPOINTER_REG_23_ );
nand U137632 ( n24770, n24824, P1_P2_PHYADDRPOINTER_REG_23_ );
nand U137633 ( n57904, n57958, P2_P2_PHYADDRPOINTER_REG_23_ );
nor U137634 ( n65993, n76213, n75464 );
nor U137635 ( n65985, n76213, n75465 );
nor U137636 ( n57483, n76279, n75466 );
nor U137637 ( n65981, n76213, n75467 );
nor U137638 ( n57487, n76279, n75468 );
nor U137639 ( n57491, n76279, n75469 );
nor U137640 ( n57495, n76279, n75470 );
nor U137641 ( n57502, n76279, n75471 );
nor U137642 ( n57506, n76279, n75472 );
nor U137643 ( n66045, n76213, n75473 );
nor U137644 ( n65989, n76213, n75474 );
nor U137645 ( n57514, n76279, n75475 );
nor U137646 ( n65977, n76213, n75476 );
nor U137647 ( n66049, n76213, n75477 );
nor U137648 ( n66053, n76213, n75478 );
nor U137649 ( n57510, n76279, n75479 );
nand U137650 ( n13876, n57480, n57481 );
nand U137651 ( n57481, n76702, P2_P2_DATAO_REG_23_ );
nor U137652 ( n57480, n57482, n57483 );
nor U137653 ( n57482, n74971, n57452 );
nand U137654 ( n13871, n57484, n57485 );
nand U137655 ( n57485, n76702, P2_P2_DATAO_REG_22_ );
nor U137656 ( n57484, n57486, n57487 );
nor U137657 ( n57486, n75377, n57452 );
nand U137658 ( n13866, n57488, n57489 );
nand U137659 ( n57489, n76702, P2_P2_DATAO_REG_21_ );
nor U137660 ( n57488, n57490, n57491 );
nor U137661 ( n57490, n74922, n57452 );
nand U137662 ( n13861, n57492, n57493 );
nand U137663 ( n57493, n76702, P2_P2_DATAO_REG_20_ );
nor U137664 ( n57492, n57494, n57495 );
nor U137665 ( n57494, n75378, n57452 );
nand U137666 ( n13856, n57499, n57500 );
nand U137667 ( n57500, n76702, P2_P2_DATAO_REG_19_ );
nor U137668 ( n57499, n57501, n57502 );
nor U137669 ( n57501, n74877, n57452 );
nand U137670 ( n13851, n57503, n57504 );
nand U137671 ( n57504, n76703, P2_P2_DATAO_REG_18_ );
nor U137672 ( n57503, n57505, n57506 );
nor U137673 ( n57505, n75379, n57452 );
nand U137674 ( n13841, n57511, n57512 );
nand U137675 ( n57512, n76703, P2_P2_DATAO_REG_16_ );
nor U137676 ( n57511, n57513, n57514 );
nor U137677 ( n57513, n75380, n57452 );
nand U137678 ( n13846, n57507, n57508 );
nand U137679 ( n57508, n76703, P2_P2_DATAO_REG_17_ );
nor U137680 ( n57507, n57509, n57510 );
nor U137681 ( n57509, n74819, n57452 );
nand U137682 ( n11611, n65990, n65991 );
nand U137683 ( n65991, n76721, P2_P3_DATAO_REG_19_ );
nor U137684 ( n65990, n65992, n65993 );
nor U137685 ( n65992, n74875, n65911 );
nand U137686 ( n11621, n65982, n65983 );
nand U137687 ( n65983, n76721, P2_P3_DATAO_REG_21_ );
nor U137688 ( n65982, n65984, n65985 );
nor U137689 ( n65984, n74921, n65911 );
nand U137690 ( n11626, n65978, n65979 );
nand U137691 ( n65979, n76721, P2_P3_DATAO_REG_22_ );
nor U137692 ( n65978, n65980, n65981 );
nor U137693 ( n65980, n75381, n65911 );
nand U137694 ( n11606, n66042, n66043 );
nand U137695 ( n66043, n76722, P2_P3_DATAO_REG_18_ );
nor U137696 ( n66042, n66044, n66045 );
nor U137697 ( n66044, n75382, n65911 );
nand U137698 ( n11616, n65986, n65987 );
nand U137699 ( n65987, n76721, P2_P3_DATAO_REG_20_ );
nor U137700 ( n65986, n65988, n65989 );
nor U137701 ( n65988, n75383, n65911 );
nand U137702 ( n11631, n65974, n65975 );
nand U137703 ( n65975, n76721, P2_P3_DATAO_REG_23_ );
nor U137704 ( n65974, n65976, n65977 );
nor U137705 ( n65976, n74968, n65911 );
nand U137706 ( n11601, n66046, n66047 );
nand U137707 ( n66047, n76722, P2_P3_DATAO_REG_17_ );
nor U137708 ( n66046, n66048, n66049 );
nor U137709 ( n66048, n74814, n65911 );
nand U137710 ( n11596, n66050, n66051 );
nand U137711 ( n66051, n76722, P2_P3_DATAO_REG_16_ );
nor U137712 ( n66050, n66052, n66053 );
nor U137713 ( n66052, n75384, n65911 );
xnor U137714 ( n9354, n74477, P1_P1_PHYADDRPOINTER_REG_2_ );
nor U137715 ( n24359, n76537, n75480 );
nor U137716 ( n24371, n76537, n75481 );
nor U137717 ( n24375, n76537, n75482 );
nor U137718 ( n24379, n76537, n75483 );
nor U137719 ( n24367, n76537, n75484 );
nor U137720 ( n24363, n76537, n75485 );
nor U137721 ( n24389, n76537, n75486 );
nor U137722 ( n24383, n76537, n75487 );
nand U137723 ( n7141, n24356, n24357 );
nand U137724 ( n24357, P1_P2_DATAO_REG_23_, n76770 );
nor U137725 ( n24356, n24358, n24359 );
nor U137726 ( n24358, n74972, n24329 );
nand U137727 ( n7126, n24368, n24369 );
nand U137728 ( n24369, P1_P2_DATAO_REG_20_, n76770 );
nor U137729 ( n24368, n24370, n24371 );
nor U137730 ( n24370, n75385, n24329 );
nand U137731 ( n7121, n24372, n24373 );
nand U137732 ( n24373, P1_P2_DATAO_REG_19_, n76770 );
nor U137733 ( n24372, n24374, n24375 );
nor U137734 ( n24374, n74878, n24329 );
nand U137735 ( n7116, n24376, n24377 );
nand U137736 ( n24377, P1_P2_DATAO_REG_18_, n76770 );
nor U137737 ( n24376, n24378, n24379 );
nor U137738 ( n24378, n75386, n24329 );
nand U137739 ( n7131, n24364, n24365 );
nand U137740 ( n24365, P1_P2_DATAO_REG_21_, n76770 );
nor U137741 ( n24364, n24366, n24367 );
nor U137742 ( n24366, n74923, n24329 );
nand U137743 ( n7136, n24360, n24361 );
nand U137744 ( n24361, P1_P2_DATAO_REG_22_, n76770 );
nor U137745 ( n24360, n24362, n24363 );
nor U137746 ( n24362, n75387, n24329 );
nand U137747 ( n7106, n24386, n24387 );
nand U137748 ( n24387, P1_P2_DATAO_REG_16_, n76770 );
nor U137749 ( n24386, n24388, n24389 );
nor U137750 ( n24388, n75388, n24329 );
nand U137751 ( n7111, n24380, n24381 );
nand U137752 ( n24381, P1_P2_DATAO_REG_17_, n76770 );
nor U137753 ( n24380, n24382, n24383 );
nor U137754 ( n24382, n74820, n24329 );
nand U137755 ( n13047, n13048, P1_P1_INSTADDRPOINTER_REG_23_ );
nand U137756 ( n13042, n13043, n74774 );
nand U137757 ( n13043, n12998, n13044 );
nand U137758 ( n13044, P1_P1_INSTADDRPOINTER_REG_24_, n13045 );
nand U137759 ( n13045, n13003, n13047 );
nand U137760 ( n45833, P2_P1_PHYADDRPOINTER_REG_19_, P2_P1_PHYADDRPOINTER_REG_18_ );
nand U137761 ( n13340, n13342, n74586 );
nand U137762 ( n13342, n4853, n13343 );
not U137763 ( n4853, n13309 );
nand U137764 ( n13343, P1_P1_INSTADDRPOINTER_REG_18_, n13344 );
nand U137765 ( n13344, n13314, n13345 );
nand U137766 ( n13345, n13347, P1_P1_INSTADDRPOINTER_REG_17_ );
nor U137767 ( n65969, n76214, n75552 );
nor U137768 ( n65915, n76214, n75553 );
nor U137769 ( n65909, n76214, n75554 );
nor U137770 ( n65957, n76214, n75555 );
nor U137771 ( n65961, n76214, n75556 );
nor U137772 ( n65965, n76214, n75557 );
nor U137773 ( n65973, n76214, n75558 );
nor U137774 ( n57463, n76280, n75559 );
nor U137775 ( n57467, n76280, n75560 );
nor U137776 ( n57479, n76280, n75561 );
nor U137777 ( n57459, n76280, n75562 );
nor U137778 ( n57475, n76280, n75563 );
nor U137779 ( n57450, n76280, n75564 );
nor U137780 ( n57471, n76280, n75565 );
nand U137781 ( n11666, n65906, n65907 );
nand U137782 ( n65907, n76721, P2_P3_DATAO_REG_30_ );
nor U137783 ( n65906, n65908, n65909 );
nor U137784 ( n65908, n75426, n65911 );
nand U137785 ( n13901, n57460, n57461 );
nand U137786 ( n57461, n76702, P2_P2_DATAO_REG_28_ );
nor U137787 ( n57460, n57462, n57463 );
nor U137788 ( n57462, n73393, n57452 );
nand U137789 ( n13896, n57464, n57465 );
nand U137790 ( n57465, n76702, P2_P2_DATAO_REG_27_ );
nor U137791 ( n57464, n57466, n57467 );
nor U137792 ( n57466, n75322, n57452 );
nand U137793 ( n13881, n57476, n57477 );
nand U137794 ( n57477, n76702, P2_P2_DATAO_REG_24_ );
nor U137795 ( n57476, n57478, n57479 );
nor U137796 ( n57478, n75342, n57452 );
nand U137797 ( n13906, n57456, n57457 );
nand U137798 ( n57457, n76702, P2_P2_DATAO_REG_29_ );
nor U137799 ( n57456, n57458, n57459 );
nor U137800 ( n57458, n75203, n57452 );
nand U137801 ( n13886, n57472, n57473 );
nand U137802 ( n57473, n76702, P2_P2_DATAO_REG_25_ );
nor U137803 ( n57472, n57474, n57475 );
nor U137804 ( n57474, n75036, n57452 );
nand U137805 ( n13911, n57447, n57448 );
nand U137806 ( n57448, n76702, P2_P2_DATAO_REG_30_ );
nor U137807 ( n57447, n57449, n57450 );
nor U137808 ( n57449, n75402, n57452 );
nand U137809 ( n13891, n57468, n57469 );
nand U137810 ( n57469, n76702, P2_P2_DATAO_REG_26_ );
nor U137811 ( n57468, n57470, n57471 );
nor U137812 ( n57470, n75343, n57452 );
nand U137813 ( n11641, n65966, n65967 );
nand U137814 ( n65967, n76721, P2_P3_DATAO_REG_25_ );
nor U137815 ( n65966, n65968, n65969 );
nor U137816 ( n65968, n75028, n65911 );
nand U137817 ( n11661, n65912, n65913 );
nand U137818 ( n65913, n76721, P2_P3_DATAO_REG_29_ );
nor U137819 ( n65912, n65914, n65915 );
nor U137820 ( n65914, n75204, n65911 );
nand U137821 ( n11656, n65954, n65955 );
nand U137822 ( n65955, n76721, P2_P3_DATAO_REG_28_ );
nor U137823 ( n65954, n65956, n65957 );
nor U137824 ( n65956, n73390, n65911 );
nand U137825 ( n11651, n65958, n65959 );
nand U137826 ( n65959, n76721, P2_P3_DATAO_REG_27_ );
nor U137827 ( n65958, n65960, n65961 );
nor U137828 ( n65960, n75346, n65911 );
nand U137829 ( n11646, n65962, n65963 );
nand U137830 ( n65963, n76721, P2_P3_DATAO_REG_26_ );
nor U137831 ( n65962, n65964, n65965 );
nor U137832 ( n65964, n75389, n65911 );
nand U137833 ( n11636, n65970, n65971 );
nand U137834 ( n65971, n76721, P2_P3_DATAO_REG_24_ );
nor U137835 ( n65970, n65972, n65973 );
nor U137836 ( n65972, n75390, n65911 );
nor U137837 ( n24337, n76538, n75566 );
nor U137838 ( n24341, n76538, n75567 );
nor U137839 ( n24355, n76538, n75568 );
nor U137840 ( n24327, n76538, n75569 );
nor U137841 ( n24333, n76538, n75570 );
nor U137842 ( n24351, n76538, n75571 );
nor U137843 ( n24347, n76538, n75572 );
nand U137844 ( n7166, n24334, n24335 );
nand U137845 ( n24335, P1_P2_DATAO_REG_28_, n76771 );
nor U137846 ( n24334, n24336, n24337 );
nor U137847 ( n24336, n73394, n24329 );
nand U137848 ( n7161, n24338, n24339 );
nand U137849 ( n24339, P1_P2_DATAO_REG_27_, n76771 );
nor U137850 ( n24338, n24340, n24341 );
nor U137851 ( n24340, n75323, n24329 );
nand U137852 ( n7146, n24352, n24353 );
nand U137853 ( n24353, P1_P2_DATAO_REG_24_, n76771 );
nor U137854 ( n24352, n24354, n24355 );
nor U137855 ( n24354, n75344, n24329 );
nand U137856 ( n7176, n24324, n24325 );
nand U137857 ( n24325, P1_P2_DATAO_REG_30_, n76771 );
nor U137858 ( n24324, n24326, n24327 );
nor U137859 ( n24326, n75403, n24329 );
nand U137860 ( n7171, n24330, n24331 );
nand U137861 ( n24331, P1_P2_DATAO_REG_29_, n76771 );
nor U137862 ( n24330, n24332, n24333 );
nor U137863 ( n24332, n75205, n24329 );
nand U137864 ( n7151, n24348, n24349 );
nand U137865 ( n24349, P1_P2_DATAO_REG_25_, n76771 );
nor U137866 ( n24348, n24350, n24351 );
nor U137867 ( n24350, n75037, n24329 );
nand U137868 ( n7156, n24344, n24345 );
nand U137869 ( n24345, P1_P2_DATAO_REG_26_, n76771 );
nor U137870 ( n24344, n24346, n24347 );
nor U137871 ( n24346, n75345, n24329 );
nand U137872 ( n66830, n66831, P2_P3_PHYADDRPOINTER_REG_18_ );
nand U137873 ( n32184, n32185, P1_P3_PHYADDRPOINTER_REG_18_ );
nand U137874 ( n24954, n24955, P1_P2_PHYADDRPOINTER_REG_18_ );
nand U137875 ( n58089, n58090, P2_P2_PHYADDRPOINTER_REG_18_ );
nor U137876 ( n43308, P2_P1_PHYADDRPOINTER_REG_0_, n74467 );
nor U137877 ( n64054, P2_P3_PHYADDRPOINTER_REG_0_, n74469 );
nor U137878 ( n30037, P1_P3_PHYADDRPOINTER_REG_0_, n74470 );
nor U137879 ( n22714, P1_P2_PHYADDRPOINTER_REG_0_, n74471 );
nor U137880 ( n55830, P2_P2_PHYADDRPOINTER_REG_0_, n74472 );
and U137881 ( n68438, n68439, P2_P3_INSTADDRPOINTER_REG_5_ );
and U137882 ( n33682, n33683, P1_P3_INSTADDRPOINTER_REG_5_ );
and U137883 ( n47406, n47407, P2_P1_INSTADDRPOINTER_REG_5_ );
and U137884 ( n26437, n26438, P1_P2_INSTADDRPOINTER_REG_5_ );
and U137885 ( n59576, n59577, P2_P2_INSTADDRPOINTER_REG_5_ );
nor U137886 ( n57581, n76278, n75604 );
nor U137887 ( n66153, n76212, n75605 );
nor U137888 ( n57577, n76278, n75606 );
nor U137889 ( n66061, n76213, n75607 );
nor U137890 ( n66065, n76213, n75608 );
nor U137891 ( n66069, n76213, n75609 );
nor U137892 ( n66073, n76212, n75610 );
nor U137893 ( n66145, n76212, n75611 );
nor U137894 ( n57569, n76278, n75612 );
nor U137895 ( n66133, n76212, n75613 );
nor U137896 ( n57557, n76278, n75614 );
nor U137897 ( n66081, n76212, n75615 );
nor U137898 ( n57545, n76278, n75616 );
nor U137899 ( n57526, n76279, n75617 );
nor U137900 ( n66137, n76212, n75618 );
nor U137901 ( n57561, n76278, n75619 );
nor U137902 ( n57530, n76279, n75620 );
nor U137903 ( n57534, n76278, n75621 );
nor U137904 ( n66125, n76212, n75622 );
nor U137905 ( n57549, n76278, n75623 );
nor U137906 ( n57522, n76279, n75624 );
nor U137907 ( n66149, n76212, n75625 );
nor U137908 ( n57573, n76278, n75626 );
nor U137909 ( n66141, n76212, n75627 );
nor U137910 ( n57565, n76278, n75628 );
nor U137911 ( n66129, n76212, n75629 );
nor U137912 ( n57553, n76278, n75630 );
nor U137913 ( n57538, n76278, n75631 );
nor U137914 ( n57518, n76279, n75632 );
nor U137915 ( n66057, n76213, n75633 );
nor U137916 ( n66157, n76212, n75634 );
nor U137917 ( n66077, n76212, n75635 );
nand U137918 ( n13761, n57579, n57580 );
nand U137919 ( n57580, n76704, P2_P2_DATAO_REG_0_ );
nor U137920 ( n57579, n57581, n57582 );
nor U137921 ( n57582, n74490, n57515 );
nand U137922 ( n13766, n57575, n57576 );
nand U137923 ( n57576, n76704, P2_P2_DATAO_REG_1_ );
nor U137924 ( n57575, n57577, n57578 );
nor U137925 ( n57578, n73128, n57515 );
nand U137926 ( n13776, n57567, n57568 );
nand U137927 ( n57568, n76704, P2_P2_DATAO_REG_3_ );
nor U137928 ( n57567, n57569, n57570 );
nor U137929 ( n57570, n74509, n57515 );
nand U137930 ( n13791, n57555, n57556 );
nand U137931 ( n57556, n76704, P2_P2_DATAO_REG_6_ );
nor U137932 ( n57555, n57557, n57558 );
nor U137933 ( n57558, n75263, n57515 );
nand U137934 ( n13806, n57543, n57544 );
nand U137935 ( n57544, n76703, P2_P2_DATAO_REG_9_ );
nor U137936 ( n57543, n57545, n57546 );
nor U137937 ( n57546, n75249, n57515 );
nand U137938 ( n13826, n57524, n57525 );
nand U137939 ( n57525, n76703, P2_P2_DATAO_REG_13_ );
nor U137940 ( n57524, n57526, n57527 );
nor U137941 ( n57527, n74732, n57515 );
nand U137942 ( n13786, n57559, n57560 );
nand U137943 ( n57560, n76704, P2_P2_DATAO_REG_5_ );
nor U137944 ( n57559, n57561, n57562 );
nor U137945 ( n57562, n74542, n57515 );
nand U137946 ( n13821, n57528, n57529 );
nand U137947 ( n57529, n76703, P2_P2_DATAO_REG_12_ );
nor U137948 ( n57528, n57530, n57531 );
nor U137949 ( n57531, n75264, n57515 );
nand U137950 ( n13816, n57532, n57533 );
nand U137951 ( n57533, n76703, P2_P2_DATAO_REG_11_ );
nor U137952 ( n57532, n57534, n57535 );
nor U137953 ( n57535, n74678, n57515 );
nand U137954 ( n13801, n57547, n57548 );
nand U137955 ( n57548, n76703, P2_P2_DATAO_REG_8_ );
nor U137956 ( n57547, n57549, n57550 );
nor U137957 ( n57550, n75265, n57515 );
nand U137958 ( n13831, n57520, n57521 );
nand U137959 ( n57521, n76703, P2_P2_DATAO_REG_14_ );
nor U137960 ( n57520, n57522, n57523 );
nor U137961 ( n57523, n75266, n57515 );
nand U137962 ( n13771, n57571, n57572 );
nand U137963 ( n57572, n76704, P2_P2_DATAO_REG_2_ );
nor U137964 ( n57571, n57573, n57574 );
nor U137965 ( n57574, n75283, n57515 );
nand U137966 ( n13781, n57563, n57564 );
nand U137967 ( n57564, n76704, P2_P2_DATAO_REG_4_ );
nor U137968 ( n57563, n57565, n57566 );
nor U137969 ( n57566, n75267, n57515 );
nand U137970 ( n13796, n57551, n57552 );
nand U137971 ( n57552, n76703, P2_P2_DATAO_REG_7_ );
nor U137972 ( n57551, n57553, n57554 );
nor U137973 ( n57554, n74583, n57515 );
nand U137974 ( n13811, n57536, n57537 );
nand U137975 ( n57537, n76703, P2_P2_DATAO_REG_10_ );
nor U137976 ( n57536, n57538, n57539 );
nor U137977 ( n57539, n74632, n57515 );
nand U137978 ( n13836, n57516, n57517 );
nand U137979 ( n57517, n76703, P2_P2_DATAO_REG_15_ );
nor U137980 ( n57516, n57518, n57519 );
nor U137981 ( n57519, n74779, n57515 );
nand U137982 ( n11521, n66151, n66152 );
nand U137983 ( n66152, n76723, P2_P3_DATAO_REG_1_ );
nor U137984 ( n66151, n66153, n66154 );
nor U137985 ( n66154, n73127, n66054 );
nand U137986 ( n11586, n66059, n66060 );
nand U137987 ( n66060, n76722, P2_P3_DATAO_REG_14_ );
nor U137988 ( n66059, n66061, n66062 );
nor U137989 ( n66062, n75268, n66054 );
nand U137990 ( n11581, n66063, n66064 );
nand U137991 ( n66064, n76722, P2_P3_DATAO_REG_13_ );
nor U137992 ( n66063, n66065, n66066 );
nor U137993 ( n66066, n74730, n66054 );
nand U137994 ( n11576, n66067, n66068 );
nand U137995 ( n66068, n76722, P2_P3_DATAO_REG_12_ );
nor U137996 ( n66067, n66069, n66070 );
nor U137997 ( n66070, n75269, n66054 );
nand U137998 ( n11571, n66071, n66072 );
nand U137999 ( n66072, n76722, P2_P3_DATAO_REG_11_ );
nor U138000 ( n66071, n66073, n66074 );
nor U138001 ( n66074, n74675, n66054 );
nand U138002 ( n11531, n66143, n66144 );
nand U138003 ( n66144, n76723, P2_P3_DATAO_REG_3_ );
nor U138004 ( n66143, n66145, n66146 );
nor U138005 ( n66146, n74507, n66054 );
nand U138006 ( n11546, n66131, n66132 );
nand U138007 ( n66132, n76723, P2_P3_DATAO_REG_6_ );
nor U138008 ( n66131, n66133, n66134 );
nor U138009 ( n66134, n75270, n66054 );
nand U138010 ( n11561, n66079, n66080 );
nand U138011 ( n66080, n76722, P2_P3_DATAO_REG_9_ );
nor U138012 ( n66079, n66081, n66082 );
nor U138013 ( n66082, n75250, n66054 );
nand U138014 ( n11541, n66135, n66136 );
nand U138015 ( n66136, n76723, P2_P3_DATAO_REG_5_ );
nor U138016 ( n66135, n66137, n66138 );
nor U138017 ( n66138, n74539, n66054 );
nand U138018 ( n11556, n66123, n66124 );
nand U138019 ( n66124, n76722, P2_P3_DATAO_REG_8_ );
nor U138020 ( n66123, n66125, n66126 );
nor U138021 ( n66126, n75271, n66054 );
nand U138022 ( n11526, n66147, n66148 );
nand U138023 ( n66148, n76723, P2_P3_DATAO_REG_2_ );
nor U138024 ( n66147, n66149, n66150 );
nor U138025 ( n66150, n75284, n66054 );
nand U138026 ( n11536, n66139, n66140 );
nand U138027 ( n66140, n76723, P2_P3_DATAO_REG_4_ );
nor U138028 ( n66139, n66141, n66142 );
nor U138029 ( n66142, n75272, n66054 );
nand U138030 ( n11551, n66127, n66128 );
nand U138031 ( n66128, n76722, P2_P3_DATAO_REG_7_ );
nor U138032 ( n66127, n66129, n66130 );
nor U138033 ( n66130, n74581, n66054 );
nand U138034 ( n11591, n66055, n66056 );
nand U138035 ( n66056, n76722, P2_P3_DATAO_REG_15_ );
nor U138036 ( n66055, n66057, n66058 );
nor U138037 ( n66058, n74776, n66054 );
nand U138038 ( n11516, n66155, n66156 );
nand U138039 ( n66156, n76723, P2_P3_DATAO_REG_0_ );
nor U138040 ( n66155, n66157, n66158 );
nor U138041 ( n66158, n74487, n66054 );
nand U138042 ( n11566, n66075, n66076 );
nand U138043 ( n66076, n76722, P2_P3_DATAO_REG_10_ );
nor U138044 ( n66075, n66077, n66078 );
nor U138045 ( n66078, n74628, n66054 );
nand U138046 ( n63892, P2_P3_PHYADDRPOINTER_REG_6_, n5629 );
nand U138047 ( n29936, P1_P3_PHYADDRPOINTER_REG_6_, n3028 );
nand U138048 ( n29621, P1_P3_PHYADDRPOINTER_REG_18_, n3028 );
nand U138049 ( n22613, P1_P2_PHYADDRPOINTER_REG_6_, n3872 );
nand U138050 ( n55726, P2_P2_PHYADDRPOINTER_REG_6_, n6504 );
nor U138051 ( n24455, n76536, n75636 );
nor U138052 ( n24397, n76537, n75637 );
nor U138053 ( n24417, n76536, n75638 );
nor U138054 ( n24405, n76537, n75639 );
nor U138055 ( n24409, n76536, n75640 );
nor U138056 ( n24421, n76536, n75641 );
nor U138057 ( n24435, n76536, n75642 );
nor U138058 ( n24447, n76536, n75643 );
nor U138059 ( n24401, n76537, n75644 );
nor U138060 ( n24443, n76536, n75645 );
nor U138061 ( n24451, n76536, n75646 );
nor U138062 ( n24439, n76536, n75647 );
nor U138063 ( n24431, n76536, n75648 );
nor U138064 ( n24425, n76536, n75649 );
nor U138065 ( n24393, n76537, n75650 );
nor U138066 ( n24413, n76536, n75651 );
nand U138067 ( n7026, n24453, n24454 );
nand U138068 ( n24454, P1_P2_DATAO_REG_0_, n76769 );
nor U138069 ( n24453, n24455, n24456 );
nor U138070 ( n24456, n74491, n24390 );
nand U138071 ( n7096, n24395, n24396 );
nand U138072 ( n24396, P1_P2_DATAO_REG_14_, n76770 );
nor U138073 ( n24395, n24397, n24398 );
nor U138074 ( n24398, n75273, n24390 );
nand U138075 ( n7071, n24415, n24416 );
nand U138076 ( n24416, P1_P2_DATAO_REG_9_, n76769 );
nor U138077 ( n24415, n24417, n24418 );
nor U138078 ( n24418, n75251, n24390 );
nand U138079 ( n7086, n24403, n24404 );
nand U138080 ( n24404, P1_P2_DATAO_REG_12_, n76770 );
nor U138081 ( n24403, n24405, n24406 );
nor U138082 ( n24406, n75274, n24390 );
nand U138083 ( n7081, n24407, n24408 );
nand U138084 ( n24408, P1_P2_DATAO_REG_11_, n76769 );
nor U138085 ( n24407, n24409, n24410 );
nor U138086 ( n24410, n74679, n24390 );
nand U138087 ( n7066, n24419, n24420 );
nand U138088 ( n24420, P1_P2_DATAO_REG_8_, n76769 );
nor U138089 ( n24419, n24421, n24422 );
nor U138090 ( n24422, n75275, n24390 );
nand U138091 ( n7051, n24433, n24434 );
nand U138092 ( n24434, P1_P2_DATAO_REG_5_, n76769 );
nor U138093 ( n24433, n24435, n24436 );
nor U138094 ( n24436, n74543, n24390 );
nand U138095 ( n7036, n24445, n24446 );
nand U138096 ( n24446, P1_P2_DATAO_REG_2_, n76769 );
nor U138097 ( n24445, n24447, n24448 );
nor U138098 ( n24448, n75285, n24390 );
nand U138099 ( n7091, n24399, n24400 );
nand U138100 ( n24400, P1_P2_DATAO_REG_13_, n76770 );
nor U138101 ( n24399, n24401, n24402 );
nor U138102 ( n24402, n74733, n24390 );
nand U138103 ( n7041, n24441, n24442 );
nand U138104 ( n24442, P1_P2_DATAO_REG_3_, n76769 );
nor U138105 ( n24441, n24443, n24444 );
nor U138106 ( n24444, n74510, n24390 );
nand U138107 ( n7031, n24449, n24450 );
nand U138108 ( n24450, P1_P2_DATAO_REG_1_, n76769 );
nor U138109 ( n24449, n24451, n24452 );
nor U138110 ( n24452, n73129, n24390 );
nand U138111 ( n7046, n24437, n24438 );
nand U138112 ( n24438, P1_P2_DATAO_REG_4_, n76769 );
nor U138113 ( n24437, n24439, n24440 );
nor U138114 ( n24440, n75276, n24390 );
nand U138115 ( n7056, n24429, n24430 );
nand U138116 ( n24430, P1_P2_DATAO_REG_6_, n76769 );
nor U138117 ( n24429, n24431, n24432 );
nor U138118 ( n24432, n75277, n24390 );
nand U138119 ( n7061, n24423, n24424 );
nand U138120 ( n24424, P1_P2_DATAO_REG_7_, n76769 );
nor U138121 ( n24423, n24425, n24426 );
nor U138122 ( n24426, n74584, n24390 );
nand U138123 ( n7101, n24391, n24392 );
nand U138124 ( n24392, P1_P2_DATAO_REG_15_, n76770 );
nor U138125 ( n24391, n24393, n24394 );
nor U138126 ( n24394, n74780, n24390 );
nand U138127 ( n7076, n24411, n24412 );
nand U138128 ( n24412, P1_P2_DATAO_REG_10_, n76769 );
nor U138129 ( n24411, n24413, n24414 );
nor U138130 ( n24414, n74633, n24390 );
nand U138131 ( n63520, P2_P3_PHYADDRPOINTER_REG_18_, n5629 );
nand U138132 ( n22300, P1_P2_PHYADDRPOINTER_REG_18_, n3872 );
nand U138133 ( n55412, P2_P2_PHYADDRPOINTER_REG_18_, n6504 );
nor U138134 ( n8410, n8475, P1_P1_EBX_REG_29_ );
nand U138135 ( n8475, n8499, n5450 );
nor U138136 ( n8499, P1_P1_EBX_REG_28_, P1_P1_EBX_REG_27_ );
nand U138137 ( n9273, n9345, n73126 );
nor U138138 ( n9345, P1_P1_EBX_REG_2_, P1_P1_EBX_REG_1_ );
nand U138139 ( n43244, n43302, n73123 );
nor U138140 ( n43302, P2_P1_EBX_REG_2_, P2_P1_EBX_REG_1_ );
nand U138141 ( n63571, P2_P3_PHYADDRPOINTER_REG_16_, n5629 );
nand U138142 ( n63736, P2_P3_PHYADDRPOINTER_REG_12_, n5629 );
nand U138143 ( n63788, P2_P3_PHYADDRPOINTER_REG_10_, n5629 );
nand U138144 ( n29672, P1_P3_PHYADDRPOINTER_REG_16_, n3028 );
nand U138145 ( n29776, P1_P3_PHYADDRPOINTER_REG_12_, n3028 );
nand U138146 ( n29828, P1_P3_PHYADDRPOINTER_REG_10_, n3028 );
nand U138147 ( n22509, P1_P2_PHYADDRPOINTER_REG_10_, n3872 );
nand U138148 ( n22351, P1_P2_PHYADDRPOINTER_REG_16_, n3872 );
nand U138149 ( n22455, P1_P2_PHYADDRPOINTER_REG_12_, n3872 );
nand U138150 ( n55622, P2_P2_PHYADDRPOINTER_REG_10_, n6504 );
nand U138151 ( n55463, P2_P2_PHYADDRPOINTER_REG_16_, n6504 );
nand U138152 ( n55570, P2_P2_PHYADDRPOINTER_REG_12_, n6504 );
nand U138153 ( n43180, n43245, n8119 );
nor U138154 ( n43245, P2_P1_EBX_REG_4_, P2_P1_EBX_REG_3_ );
nand U138155 ( n9210, n9274, n5465 );
nor U138156 ( n9274, P1_P1_EBX_REG_4_, P1_P1_EBX_REG_3_ );
nand U138157 ( n8498, n8582, n5452 );
nor U138158 ( n8582, P1_P1_EBX_REG_26_, P1_P1_EBX_REG_25_ );
nand U138159 ( n8770, n8823, n5457 );
nor U138160 ( n8823, P1_P1_EBX_REG_18_, P1_P1_EBX_REG_17_ );
nand U138161 ( n8949, n9017, n5460 );
nor U138162 ( n9017, P1_P1_EBX_REG_12_, P1_P1_EBX_REG_11_ );
nand U138163 ( n9015, n9089, n5462 );
nor U138164 ( n9089, P1_P1_EBX_REG_9_, P1_P1_EBX_REG_10_ );
nand U138165 ( n9088, n9154, n5463 );
nor U138166 ( n9154, P1_P1_EBX_REG_8_, P1_P1_EBX_REG_7_ );
nand U138167 ( n9153, n9212, n5464 );
nor U138168 ( n9212, P1_P1_EBX_REG_6_, P1_P1_EBX_REG_5_ );
nand U138169 ( n42814, n42856, n8110 );
nor U138170 ( n42856, P2_P1_EBX_REG_18_, P2_P1_EBX_REG_17_ );
nand U138171 ( n42971, n43025, n8114 );
nor U138172 ( n43025, P2_P1_EBX_REG_12_, P2_P1_EBX_REG_11_ );
nand U138173 ( n43024, n43083, n8115 );
nor U138174 ( n43083, P2_P1_EBX_REG_9_, P2_P1_EBX_REG_10_ );
nand U138175 ( n43082, n43135, n8117 );
nor U138176 ( n43135, P2_P1_EBX_REG_8_, P2_P1_EBX_REG_7_ );
nand U138177 ( n43134, n43181, n8118 );
nor U138178 ( n43181, P2_P1_EBX_REG_6_, P2_P1_EBX_REG_5_ );
nand U138179 ( n42568, n42635, n8105 );
nor U138180 ( n42635, P2_P1_EBX_REG_26_, P2_P1_EBX_REG_25_ );
nand U138181 ( n42634, n42710, n8107 );
nor U138182 ( n42710, P2_P1_EBX_REG_24_, P2_P1_EBX_REG_23_ );
nand U138183 ( n42709, n42751, n8108 );
nor U138184 ( n42751, P2_P1_EBX_REG_22_, P2_P1_EBX_REG_21_ );
nand U138185 ( n42855, n42912, n8112 );
nor U138186 ( n42912, P2_P1_EBX_REG_16_, P2_P1_EBX_REG_15_ );
nand U138187 ( n43109, n7393, P2_P1_PHYADDRPOINTER_REG_9_ );
nand U138188 ( n43285, n7393, P2_P1_PHYADDRPOINTER_REG_3_ );
nand U138189 ( n42887, n7393, P2_P1_PHYADDRPOINTER_REG_17_ );
nand U138190 ( n63539, P2_P3_PHYADDRPOINTER_REG_17_, n5629 );
nand U138191 ( n63970, P2_P3_PHYADDRPOINTER_REG_3_, n5629 );
nand U138192 ( n29640, P1_P3_PHYADDRPOINTER_REG_17_, n3028 );
nand U138193 ( n30014, P1_P3_PHYADDRPOINTER_REG_3_, n3028 );
nand U138194 ( n22691, P1_P2_PHYADDRPOINTER_REG_3_, n3872 );
nand U138195 ( n22319, P1_P2_PHYADDRPOINTER_REG_17_, n3872 );
nand U138196 ( n55431, P2_P2_PHYADDRPOINTER_REG_17_, n6504 );
nand U138197 ( n8690, n8772, n5455 );
nor U138198 ( n8772, P1_P1_EBX_REG_20_, P1_P1_EBX_REG_19_ );
nand U138199 ( n8580, n8645, n5453 );
nor U138200 ( n8645, P1_P1_EBX_REG_24_, P1_P1_EBX_REG_23_ );
nand U138201 ( n8822, n8893, n5458 );
nor U138202 ( n8893, P1_P1_EBX_REG_16_, P1_P1_EBX_REG_15_ );
nand U138203 ( n8644, n8692, n5454 );
nor U138204 ( n8692, P1_P1_EBX_REG_22_, P1_P1_EBX_REG_21_ );
nand U138205 ( n8892, n8950, n5459 );
nor U138206 ( n8950, P1_P1_EBX_REG_14_, P1_P1_EBX_REG_13_ );
nand U138207 ( n42750, n42815, n8109 );
nor U138208 ( n42815, P2_P1_EBX_REG_20_, P2_P1_EBX_REG_19_ );
nand U138209 ( n42911, n42972, n8113 );
nor U138210 ( n42972, P2_P1_EBX_REG_14_, P2_P1_EBX_REG_13_ );
and U138211 ( n42550, n42569, n8104 );
nor U138212 ( n42569, P2_P1_EBX_REG_28_, P2_P1_EBX_REG_27_ );
nand U138213 ( n55807, P2_P2_PHYADDRPOINTER_REG_3_, n6504 );
nor U138214 ( n45157, n45159, n45160 );
nor U138215 ( n45160, n865, n74401 );
nor U138216 ( n45159, n45161, n45162 );
nand U138217 ( n45162, P3_REG2_REG_11_, n43559 );
nor U138218 ( n45062, n76357, n75488 );
nor U138219 ( n45094, n76357, n75489 );
nor U138220 ( n45090, n76357, n75490 );
nor U138221 ( n45102, n76357, n75491 );
nor U138222 ( n45058, n76357, n75492 );
nor U138223 ( n45110, n76357, n75493 );
nor U138224 ( n45106, n76357, n75494 );
nor U138225 ( n45054, n76357, n75495 );
nand U138226 ( n16111, n45059, n45060 );
nand U138227 ( n45060, n76679, P2_P1_DATAO_REG_21_ );
nor U138228 ( n45059, n45061, n45062 );
nor U138229 ( n45061, n73288, n45026 );
nand U138230 ( n16101, n45091, n45092 );
nand U138231 ( n45092, n76679, P2_P1_DATAO_REG_19_ );
nor U138232 ( n45091, n45093, n45094 );
nor U138233 ( n45093, n74953, n45026 );
nand U138234 ( n16106, n45087, n45088 );
nand U138235 ( n45088, n76679, P2_P1_DATAO_REG_20_ );
nor U138236 ( n45087, n45089, n45090 );
nor U138237 ( n45089, n74965, n45026 );
nand U138238 ( n16096, n45099, n45100 );
nand U138239 ( n45100, n76680, P2_P1_DATAO_REG_18_ );
nor U138240 ( n45099, n45101, n45102 );
nor U138241 ( n45101, n73265, n45026 );
nand U138242 ( n16116, n45055, n45056 );
nand U138243 ( n45056, n76679, P2_P1_DATAO_REG_22_ );
nor U138244 ( n45055, n45057, n45058 );
nor U138245 ( n45057, n75001, n45026 );
nand U138246 ( n16086, n45107, n45108 );
nand U138247 ( n45108, n76680, P2_P1_DATAO_REG_16_ );
nor U138248 ( n45107, n45109, n45110 );
nor U138249 ( n45109, n74902, n45026 );
nand U138250 ( n16091, n45103, n45104 );
nand U138251 ( n45104, n76680, P2_P1_DATAO_REG_17_ );
nor U138252 ( n45103, n45105, n45106 );
nor U138253 ( n45105, n74908, n45026 );
nand U138254 ( n16121, n45051, n45052 );
nand U138255 ( n45052, n76679, P2_P1_DATAO_REG_23_ );
nor U138256 ( n45051, n45053, n45054 );
nor U138257 ( n45053, n75012, n45026 );
nor U138258 ( n45222, n45224, n45225 );
nor U138259 ( n45225, n865, n74406 );
nor U138260 ( n45224, n45226, n45227 );
nand U138261 ( n45227, P3_REG1_REG_11_, n43559 );
nor U138262 ( n45024, n76358, n75573 );
nor U138263 ( n45034, n76358, n75574 );
nor U138264 ( n45038, n76358, n75575 );
nor U138265 ( n45042, n76358, n75576 );
nor U138266 ( n45030, n76358, n75577 );
nor U138267 ( n45050, n76358, n75578 );
nor U138268 ( n45046, n76358, n75579 );
nand U138269 ( n16156, n45021, n45022 );
nand U138270 ( n45022, n76679, P2_P1_DATAO_REG_30_ );
nor U138271 ( n45021, n45023, n45024 );
nor U138272 ( n45023, n75404, n45026 );
nand U138273 ( n16146, n45031, n45032 );
nand U138274 ( n45032, n76679, P2_P1_DATAO_REG_28_ );
nor U138275 ( n45031, n45033, n45034 );
nor U138276 ( n45033, n75324, n45026 );
nand U138277 ( n16141, n45035, n45036 );
nand U138278 ( n45036, n76679, P2_P1_DATAO_REG_27_ );
nor U138279 ( n45035, n45037, n45038 );
nor U138280 ( n45037, n73320, n45026 );
nand U138281 ( n16136, n45039, n45040 );
nand U138282 ( n45040, n76679, P2_P1_DATAO_REG_26_ );
nor U138283 ( n45039, n45041, n45042 );
nor U138284 ( n45041, n75084, n45026 );
nand U138285 ( n16151, n45027, n45028 );
nand U138286 ( n45028, n76679, P2_P1_DATAO_REG_29_ );
nor U138287 ( n45027, n45029, n45030 );
nor U138288 ( n45029, n75218, n45026 );
nand U138289 ( n16126, n45047, n45048 );
nand U138290 ( n45048, n76679, P2_P1_DATAO_REG_24_ );
nor U138291 ( n45047, n45049, n45050 );
nor U138292 ( n45049, n73306, n45026 );
nand U138293 ( n16131, n45043, n45044 );
nand U138294 ( n45044, n76679, P2_P1_DATAO_REG_25_ );
nor U138295 ( n45043, n45045, n45046 );
nor U138296 ( n45045, n75061, n45026 );
nand U138297 ( n9122, n4751, P1_P1_PHYADDRPOINTER_REG_9_ );
nand U138298 ( n9324, n4751, P1_P1_PHYADDRPOINTER_REG_3_ );
nand U138299 ( n8862, n4751, P1_P1_PHYADDRPOINTER_REG_17_ );
nand U138300 ( n13768, n13769, n74735 );
nand U138301 ( n13769, n13739, n13770 );
nand U138302 ( n13770, P1_P1_INSTADDRPOINTER_REG_9_, n13772 );
nand U138303 ( n13772, n4859, n13773 );
nor U138304 ( n45289, n76356, n75652 );
nor U138305 ( n45318, n76356, n75653 );
nor U138306 ( n45118, n76357, n75654 );
nor U138307 ( n45277, n76356, n75655 );
nor U138308 ( n45126, n76357, n75656 );
nor U138309 ( n45130, n76356, n75657 );
nor U138310 ( n45297, n76356, n75658 );
nor U138311 ( n45285, n76356, n75659 );
nor U138312 ( n45122, n76357, n75660 );
nor U138313 ( n45309, n76356, n75661 );
nor U138314 ( n45281, n76356, n75662 );
nor U138315 ( n45293, n76356, n75663 );
nor U138316 ( n45305, n76356, n75664 );
nor U138317 ( n45313, n76356, n75665 );
nor U138318 ( n45301, n76356, n75666 );
nor U138319 ( n45114, n76357, n75667 );
nand U138320 ( n16041, n45287, n45288 );
nand U138321 ( n45288, n76680, P2_P1_DATAO_REG_7_ );
nor U138322 ( n45287, n45289, n45290 );
nor U138323 ( n45290, n74738, n45111 );
nand U138324 ( n16006, n45315, n45316 );
nand U138325 ( n45316, n76681, P2_P1_DATAO_REG_0_ );
nor U138326 ( n45315, n45318, n45319 );
nor U138327 ( n45319, n73161, n45111 );
nand U138328 ( n16076, n45116, n45117 );
nand U138329 ( n45117, n76680, P2_P1_DATAO_REG_14_ );
nor U138330 ( n45116, n45118, n45119 );
nor U138331 ( n45119, n73251, n45111 );
nand U138332 ( n16056, n45275, n45276 );
nand U138333 ( n45276, n76680, P2_P1_DATAO_REG_10_ );
nor U138334 ( n45275, n45277, n45278 );
nor U138335 ( n45278, n74786, n45111 );
nand U138336 ( n16066, n45124, n45125 );
nand U138337 ( n45125, n76680, P2_P1_DATAO_REG_12_ );
nor U138338 ( n45124, n45126, n45127 );
nor U138339 ( n45127, n74803, n45111 );
nand U138340 ( n16061, n45128, n45129 );
nand U138341 ( n45129, n76680, P2_P1_DATAO_REG_11_ );
nor U138342 ( n45128, n45130, n45131 );
nor U138343 ( n45131, n73237, n45111 );
nand U138344 ( n16031, n45295, n45296 );
nand U138345 ( n45296, n76681, P2_P1_DATAO_REG_5_ );
nor U138346 ( n45295, n45297, n45298 );
nor U138347 ( n45298, n73195, n45111 );
nand U138348 ( n16046, n45283, n45284 );
nand U138349 ( n45284, n76680, P2_P1_DATAO_REG_8_ );
nor U138350 ( n45283, n45285, n45286 );
nor U138351 ( n45286, n73218, n45111 );
nand U138352 ( n16071, n45120, n45121 );
nand U138353 ( n45121, n76680, P2_P1_DATAO_REG_13_ );
nor U138354 ( n45120, n45122, n45123 );
nor U138355 ( n45123, n74842, n45111 );
nand U138356 ( n16016, n45307, n45308 );
nand U138357 ( n45308, n76681, P2_P1_DATAO_REG_2_ );
nor U138358 ( n45307, n45309, n45310 );
nor U138359 ( n45310, n73165, n45111 );
nand U138360 ( n16051, n45279, n45280 );
nand U138361 ( n45280, n76680, P2_P1_DATAO_REG_9_ );
nor U138362 ( n45279, n45281, n45282 );
nor U138363 ( n45282, n74757, n45111 );
nand U138364 ( n16036, n45291, n45292 );
nand U138365 ( n45292, n76680, P2_P1_DATAO_REG_6_ );
nor U138366 ( n45291, n45293, n45294 );
nor U138367 ( n45294, n74704, n45111 );
nand U138368 ( n16021, n45303, n45304 );
nand U138369 ( n45304, n76681, P2_P1_DATAO_REG_3_ );
nor U138370 ( n45303, n45305, n45306 );
nor U138371 ( n45306, n74631, n45111 );
nand U138372 ( n16011, n45311, n45312 );
nand U138373 ( n45312, n76681, P2_P1_DATAO_REG_1_ );
nor U138374 ( n45311, n45313, n45314 );
nor U138375 ( n45314, n74609, n45111 );
nand U138376 ( n16026, n45299, n45300 );
nand U138377 ( n45300, n76681, P2_P1_DATAO_REG_4_ );
nor U138378 ( n45299, n45301, n45302 );
nor U138379 ( n45302, n74681, n45111 );
nand U138380 ( n16081, n45112, n45113 );
nand U138381 ( n45113, n76680, P2_P1_DATAO_REG_15_ );
nor U138382 ( n45112, n45114, n45115 );
nor U138383 ( n45115, n74865, n45111 );
nor U138384 ( n11365, n76623, n75496 );
nor U138385 ( n11375, n76623, n75497 );
nor U138386 ( n11380, n76623, n75498 );
nor U138387 ( n11385, n76623, n75499 );
nor U138388 ( n11390, n76623, n75500 );
nor U138389 ( n11370, n76623, n75501 );
nor U138390 ( n11409, n76623, n75502 );
nor U138391 ( n11404, n76623, n75503 );
nand U138392 ( n9386, n11362, n11363 );
nand U138393 ( n11363, P1_P1_DATAO_REG_23_, n76747 );
nor U138394 ( n11362, n11364, n11365 );
nor U138395 ( n11364, n75013, n11325 );
nand U138396 ( n9376, n11372, n11373 );
nand U138397 ( n11373, P1_P1_DATAO_REG_21_, n76747 );
nor U138398 ( n11372, n11374, n11375 );
nor U138399 ( n11374, n73289, n11325 );
nand U138400 ( n9371, n11377, n11378 );
nand U138401 ( n11378, P1_P1_DATAO_REG_20_, n76747 );
nor U138402 ( n11377, n11379, n11380 );
nor U138403 ( n11379, n74966, n11325 );
nand U138404 ( n9366, n11382, n11383 );
nand U138405 ( n11383, P1_P1_DATAO_REG_19_, n76747 );
nor U138406 ( n11382, n11384, n11385 );
nor U138407 ( n11384, n74954, n11325 );
nand U138408 ( n9361, n11387, n11388 );
nand U138409 ( n11388, P1_P1_DATAO_REG_18_, n76747 );
nor U138410 ( n11387, n11389, n11390 );
nor U138411 ( n11389, n73266, n11325 );
nand U138412 ( n9381, n11367, n11368 );
nand U138413 ( n11368, P1_P1_DATAO_REG_22_, n76747 );
nor U138414 ( n11367, n11369, n11370 );
nor U138415 ( n11369, n75002, n11325 );
nand U138416 ( n9351, n11405, n11407 );
nand U138417 ( n11407, P1_P1_DATAO_REG_16_, n76747 );
nor U138418 ( n11405, n11408, n11409 );
nor U138419 ( n11408, n74903, n11325 );
nand U138420 ( n9356, n11400, n11402 );
nand U138421 ( n11402, P1_P1_DATAO_REG_17_, n76747 );
nor U138422 ( n11400, n11403, n11404 );
nor U138423 ( n11403, n74909, n11325 );
nor U138424 ( n11323, n76624, n75580 );
nor U138425 ( n11355, n76624, n75581 );
nor U138426 ( n11335, n76624, n75582 );
nor U138427 ( n11345, n76624, n75583 );
nor U138428 ( n11350, n76624, n75584 );
nor U138429 ( n11330, n76624, n75585 );
nor U138430 ( n11360, n76624, n75586 );
nand U138431 ( n9421, n11319, n11320 );
nand U138432 ( n11320, P1_P1_DATAO_REG_30_, n76748 );
nor U138433 ( n11319, n11322, n11323 );
nor U138434 ( n11322, n75405, n11325 );
nand U138435 ( n9396, n11352, n11353 );
nand U138436 ( n11353, P1_P1_DATAO_REG_25_, n76748 );
nor U138437 ( n11352, n11354, n11355 );
nor U138438 ( n11354, n75062, n11325 );
nand U138439 ( n9411, n11332, n11333 );
nand U138440 ( n11333, P1_P1_DATAO_REG_28_, n76748 );
nor U138441 ( n11332, n11334, n11335 );
nor U138442 ( n11334, n75325, n11325 );
nand U138443 ( n9406, n11342, n11343 );
nand U138444 ( n11343, P1_P1_DATAO_REG_27_, n76748 );
nor U138445 ( n11342, n11344, n11345 );
nor U138446 ( n11344, n73321, n11325 );
nand U138447 ( n9401, n11347, n11348 );
nand U138448 ( n11348, P1_P1_DATAO_REG_26_, n76748 );
nor U138449 ( n11347, n11349, n11350 );
nor U138450 ( n11349, n75085, n11325 );
nand U138451 ( n9416, n11327, n11328 );
nand U138452 ( n11328, P1_P1_DATAO_REG_29_, n76748 );
nor U138453 ( n11327, n11329, n11330 );
nor U138454 ( n11329, n75219, n11325 );
nand U138455 ( n9391, n11357, n11358 );
nand U138456 ( n11358, P1_P1_DATAO_REG_24_, n76748 );
nor U138457 ( n11357, n11359, n11360 );
nor U138458 ( n11359, n73307, n11325 );
nand U138459 ( n14705, P1_P1_INSTQUEUEWR_ADDR_REG_0_, P1_P1_INSTQUEUEWR_ADDR_REG_1_ );
nor U138460 ( n11414, n76623, n75668 );
nor U138461 ( n11495, n76622, n75669 );
nor U138462 ( n11419, n76623, n75670 );
nor U138463 ( n11444, n76622, n75671 );
nor U138464 ( n11439, n76622, n75672 );
nor U138465 ( n11429, n76623, n75673 );
nor U138466 ( n11434, n76622, n75674 );
nor U138467 ( n11449, n76622, n75675 );
nor U138468 ( n11469, n76622, n75676 );
nor U138469 ( n11424, n76623, n75677 );
nor U138470 ( n11484, n76622, n75678 );
nor U138471 ( n11479, n76622, n75679 );
nor U138472 ( n11489, n76622, n75680 );
nor U138473 ( n11464, n76622, n75681 );
nor U138474 ( n11474, n76622, n75682 );
nor U138475 ( n11459, n76622, n75683 );
nand U138476 ( n9346, n11412, n11413 );
nand U138477 ( n11413, P1_P1_DATAO_REG_15_, n76747 );
nor U138478 ( n11412, n11414, n11415 );
nor U138479 ( n11415, n74864, n11410 );
nand U138480 ( n9271, n11492, n11493 );
nand U138481 ( n11493, P1_P1_DATAO_REG_0_, n76746 );
nor U138482 ( n11492, n11495, n11497 );
nor U138483 ( n11497, n73162, n11410 );
nand U138484 ( n9341, n11417, n11418 );
nand U138485 ( n11418, P1_P1_DATAO_REG_14_, n76747 );
nor U138486 ( n11417, n11419, n11420 );
nor U138487 ( n11420, n73252, n11410 );
nand U138488 ( n9316, n11442, n11443 );
nand U138489 ( n11443, P1_P1_DATAO_REG_9_, n76746 );
nor U138490 ( n11442, n11444, n11445 );
nor U138491 ( n11445, n74756, n11410 );
nand U138492 ( n9321, n11437, n11438 );
nand U138493 ( n11438, P1_P1_DATAO_REG_10_, n76746 );
nor U138494 ( n11437, n11439, n11440 );
nor U138495 ( n11440, n74787, n11410 );
nand U138496 ( n9331, n11427, n11428 );
nand U138497 ( n11428, P1_P1_DATAO_REG_12_, n76747 );
nor U138498 ( n11427, n11429, n11430 );
nor U138499 ( n11430, n74802, n11410 );
nand U138500 ( n9326, n11432, n11433 );
nand U138501 ( n11433, P1_P1_DATAO_REG_11_, n76746 );
nor U138502 ( n11432, n11434, n11435 );
nor U138503 ( n11435, n73238, n11410 );
nand U138504 ( n9311, n11447, n11448 );
nand U138505 ( n11448, P1_P1_DATAO_REG_8_, n76746 );
nor U138506 ( n11447, n11449, n11450 );
nor U138507 ( n11450, n73219, n11410 );
nand U138508 ( n9296, n11467, n11468 );
nand U138509 ( n11468, P1_P1_DATAO_REG_5_, n76746 );
nor U138510 ( n11467, n11469, n11470 );
nor U138511 ( n11470, n73196, n11410 );
nand U138512 ( n9336, n11422, n11423 );
nand U138513 ( n11423, P1_P1_DATAO_REG_13_, n76747 );
nor U138514 ( n11422, n11424, n11425 );
nor U138515 ( n11425, n74843, n11410 );
nand U138516 ( n9281, n11482, n11483 );
nand U138517 ( n11483, P1_P1_DATAO_REG_2_, n76746 );
nor U138518 ( n11482, n11484, n11485 );
nor U138519 ( n11485, n73166, n11410 );
nand U138520 ( n9286, n11477, n11478 );
nand U138521 ( n11478, P1_P1_DATAO_REG_3_, n76746 );
nor U138522 ( n11477, n11479, n11480 );
nor U138523 ( n11480, n74630, n11410 );
nand U138524 ( n9276, n11487, n11488 );
nand U138525 ( n11488, P1_P1_DATAO_REG_1_, n76746 );
nor U138526 ( n11487, n11489, n11490 );
nor U138527 ( n11490, n74608, n11410 );
nand U138528 ( n9301, n11462, n11463 );
nand U138529 ( n11463, P1_P1_DATAO_REG_6_, n76746 );
nor U138530 ( n11462, n11464, n11465 );
nor U138531 ( n11465, n74705, n11410 );
nand U138532 ( n9291, n11472, n11473 );
nand U138533 ( n11473, P1_P1_DATAO_REG_4_, n76746 );
nor U138534 ( n11472, n11474, n11475 );
nor U138535 ( n11475, n74682, n11410 );
nand U138536 ( n9306, n11457, n11458 );
nand U138537 ( n11458, P1_P1_DATAO_REG_7_, n76746 );
nor U138538 ( n11457, n11459, n11460 );
nor U138539 ( n11460, n74739, n11410 );
nor U138540 ( n68114, P2_P3_INSTADDRPOINTER_REG_10_, n5714 );
nor U138541 ( n26111, P1_P2_INSTADDRPOINTER_REG_10_, n3957 );
nor U138542 ( n59252, P2_P2_INSTADDRPOINTER_REG_10_, n6589 );
nand U138543 ( n33442, n33443, n73115 );
nand U138544 ( n33443, n33420, n33444 );
nand U138545 ( n33444, P1_P3_INSTADDRPOINTER_REG_9_, n33445 );
nand U138546 ( n33445, n3118, n33446 );
nand U138547 ( n68800, n68803, n75054 );
nand U138548 ( n68803, n5689, n68804 );
nand U138549 ( n68804, P2_P3_INSTADDRPOINTER_REG_0_, n67826 );
nand U138550 ( n34044, n34047, n75055 );
nand U138551 ( n34047, n3088, n34048 );
nand U138552 ( n34048, P1_P3_INSTADDRPOINTER_REG_0_, n33070 );
nand U138553 ( n26801, n26804, n75056 );
nand U138554 ( n26804, n3932, n26805 );
nand U138555 ( n26805, P1_P2_INSTADDRPOINTER_REG_0_, n25823 );
nand U138556 ( n59941, n59944, n75057 );
nand U138557 ( n59944, n6564, n59945 );
nand U138558 ( n59945, P2_P2_INSTADDRPOINTER_REG_0_, n58961 );
nor U138559 ( n33357, P1_P3_INSTADDRPOINTER_REG_10_, n3113 );
nand U138560 ( n68193, n68194, n74758 );
nand U138561 ( n68194, n68170, n68195 );
nand U138562 ( n68195, P2_P3_INSTADDRPOINTER_REG_9_, n68196 );
nand U138563 ( n68196, n5719, n68197 );
nand U138564 ( n47162, n47163, n74734 );
nand U138565 ( n47163, n47139, n47164 );
nand U138566 ( n47164, P2_P1_INSTADDRPOINTER_REG_9_, n47165 );
nand U138567 ( n47165, n7505, n47166 );
nand U138568 ( n26192, n26193, n74759 );
nand U138569 ( n26193, n26169, n26194 );
nand U138570 ( n26194, P1_P2_INSTADDRPOINTER_REG_9_, n26195 );
nand U138571 ( n26195, n3962, n26196 );
nand U138572 ( n59331, n59332, n74760 );
nand U138573 ( n59332, n59308, n59333 );
nand U138574 ( n59333, P2_P2_INSTADDRPOINTER_REG_9_, n59334 );
nand U138575 ( n59334, n6594, n59335 );
nor U138576 ( n67771, P2_P3_INSTADDRPOINTER_REG_19_, n5714 );
nor U138577 ( n33015, P1_P3_INSTADDRPOINTER_REG_19_, n3113 );
nor U138578 ( n25768, P1_P2_INSTADDRPOINTER_REG_19_, n3957 );
nor U138579 ( n58906, P2_P2_INSTADDRPOINTER_REG_19_, n6589 );
nand U138580 ( n46818, P2_P1_INSTADDRPOINTER_REG_17_, P2_P1_INSTADDRPOINTER_REG_16_ );
nand U138581 ( n23148, n23149, n23150 );
nand U138582 ( n23149, P1_BUF2_REG_30_, n162 );
nand U138583 ( n23150, n163, P1_BUF1_REG_30_ );
nand U138584 ( n23293, n23294, n23295 );
nand U138585 ( n23294, P1_BUF2_REG_27_, n162 );
nand U138586 ( n23295, n163, P1_BUF1_REG_27_ );
nand U138587 ( n23438, n23439, n23440 );
nand U138588 ( n23439, P1_BUF2_REG_24_, n162 );
nand U138589 ( n23440, n163, P1_BUF1_REG_24_ );
nor U138590 ( n13755, P1_P1_INSTADDRPOINTER_REG_8_, n4832 );
nand U138591 ( n14523, n14527, n75059 );
nand U138592 ( n14527, n4832, n14528 );
nand U138593 ( n14528, P1_P1_INSTADDRPOINTER_REG_0_, n12828 );
nor U138594 ( n9353, P1_P1_PHYADDRPOINTER_REG_0_, n74477 );
nand U138595 ( n56269, n56270, n56271 );
nand U138596 ( n56270, n434, P2_BUF2_REG_30_ );
nand U138597 ( n56271, n435, P2_BUF1_REG_30_ );
nand U138598 ( n56417, n56418, n56419 );
nand U138599 ( n56418, n434, P2_BUF2_REG_27_ );
nand U138600 ( n56419, n435, P2_BUF1_REG_27_ );
nand U138601 ( n56560, n56561, n56562 );
nand U138602 ( n56561, n434, P2_BUF2_REG_24_ );
nand U138603 ( n56562, n435, P2_BUF1_REG_24_ );
nor U138604 ( n13669, P1_P1_INSTADDRPOINTER_REG_10_, n4855 );
nor U138605 ( n47083, P2_P1_INSTADDRPOINTER_REG_10_, n7500 );
nor U138606 ( n46724, P2_P1_INSTADDRPOINTER_REG_19_, n7500 );
nor U138607 ( n13235, P1_P1_INSTADDRPOINTER_REG_19_, n4855 );
nand U138608 ( n47779, n47782, n75058 );
nand U138609 ( n47782, n7474, n47783 );
nand U138610 ( n47783, P2_P1_INSTADDRPOINTER_REG_0_, n46779 );
xor U138611 ( n37828, n37829, n37830 );
xor U138612 ( n37830, n37827, P4_REG2_REG_7_ );
nor U138613 ( n13022, P1_P1_INSTADDRPOINTER_REG_23_, n4832 );
nand U138614 ( n67865, P2_P3_INSTADDRPOINTER_REG_17_, P2_P3_INSTADDRPOINTER_REG_16_ );
nand U138615 ( n25862, P1_P2_INSTADDRPOINTER_REG_17_, P1_P2_INSTADDRPOINTER_REG_16_ );
nand U138616 ( n59000, P2_P2_INSTADDRPOINTER_REG_17_, P2_P2_INSTADDRPOINTER_REG_16_ );
xnor U138617 ( n21337, n73141, P1_P1_INSTQUEUERD_ADDR_REG_1_ );
nor U138618 ( n13334, P1_P1_INSTADDRPOINTER_REG_17_, n4832 );
nand U138619 ( n46534, n46502, n46588 );
nand U138620 ( n46588, n46589, P2_P1_INSTADDRPOINTER_REG_24_ );
nand U138621 ( n46531, n46532, n74919 );
nand U138622 ( n46532, n46457, n46533 );
nand U138623 ( n46533, P2_P1_INSTADDRPOINTER_REG_25_, n46534 );
nand U138624 ( n21858, P1_READY21_REG, P1_READY12_REG );
nand U138625 ( n23309, n23310, n23311 );
nand U138626 ( n23311, P1_BUF2_REG_26_, n162 );
nand U138627 ( n23310, n164, n22830 );
nand U138628 ( n23453, n23454, n23455 );
nand U138629 ( n23455, P1_BUF2_REG_23_, n162 );
nand U138630 ( n23454, n164, n22859 );
nand U138631 ( n23642, n23643, n23644 );
nand U138632 ( n23644, P1_BUF2_REG_20_, n162 );
nand U138633 ( n23643, n164, n22889 );
nand U138634 ( n23686, n23687, n23688 );
nand U138635 ( n23688, P1_BUF2_REG_19_, n162 );
nand U138636 ( n23687, n164, n22899 );
nand U138637 ( n23731, n23732, n23733 );
nand U138638 ( n23733, P1_BUF2_REG_18_, n162 );
nand U138639 ( n23732, n164, n22908 );
nand U138640 ( n23597, n23598, n23599 );
nand U138641 ( n23599, P1_BUF2_REG_21_, n162 );
nand U138642 ( n23598, n164, n22880 );
nand U138643 ( n23553, n23554, n23555 );
nand U138644 ( n23555, P1_BUF2_REG_22_, n162 );
nand U138645 ( n23554, n164, n22870 );
nand U138646 ( n23164, n23165, n23166 );
nand U138647 ( n23166, P1_BUF2_REG_29_, n162 );
nand U138648 ( n23165, n164, n22804 );
nand U138649 ( n23356, n23357, n23358 );
nand U138650 ( n23358, P1_BUF2_REG_25_, n162 );
nand U138651 ( n23357, n164, n22840 );
nand U138652 ( n23775, n23776, n23777 );
nand U138653 ( n23777, P1_BUF2_REG_17_, n162 );
nand U138654 ( n23776, n164, n22918 );
nand U138655 ( n56719, n56720, n56721 );
nand U138656 ( n56721, n434, P2_BUF2_REG_21_ );
nand U138657 ( n56720, n437, n55995 );
nand U138658 ( n56764, n56765, n56766 );
nand U138659 ( n56766, n434, P2_BUF2_REG_20_ );
nand U138660 ( n56765, n437, n56004 );
nand U138661 ( n56285, n56286, n56287 );
nand U138662 ( n56287, n434, P2_BUF2_REG_29_ );
nand U138663 ( n56286, n437, n55918 );
nand U138664 ( n56433, n56434, n56435 );
nand U138665 ( n56435, n434, P2_BUF2_REG_26_ );
nand U138666 ( n56434, n437, n55944 );
nand U138667 ( n56480, n56481, n56482 );
nand U138668 ( n56482, n434, P2_BUF2_REG_25_ );
nand U138669 ( n56481, n437, n55957 );
nand U138670 ( n56575, n56576, n56577 );
nand U138671 ( n56577, n434, P2_BUF2_REG_23_ );
nand U138672 ( n56576, n437, n55976 );
nand U138673 ( n56675, n56676, n56677 );
nand U138674 ( n56677, n434, P2_BUF2_REG_22_ );
nand U138675 ( n56676, n437, n55985 );
nand U138676 ( n56808, n56809, n56810 );
nand U138677 ( n56810, n434, P2_BUF2_REG_19_ );
nand U138678 ( n56809, n437, n56014 );
nand U138679 ( n56853, n56854, n56855 );
nand U138680 ( n56855, n434, P2_BUF2_REG_18_ );
nand U138681 ( n56854, n437, n56023 );
nand U138682 ( n56900, n56901, n56902 );
nand U138683 ( n56902, n434, P2_BUF2_REG_17_ );
nand U138684 ( n56901, n437, n56033 );
nand U138685 ( n54949, P2_READY21_REG, P2_READY12_REG );
nand U138686 ( n67630, n67631, n73223 );
nand U138687 ( n67631, n5713, n67632 );
not U138688 ( n5713, n67596 );
nand U138689 ( n67632, P2_P3_INSTADDRPOINTER_REG_24_, n67633 );
nand U138690 ( n67857, n67858, n74574 );
nand U138691 ( n67858, n5710, n67859 );
not U138692 ( n5710, n67832 );
nand U138693 ( n67859, P2_P3_INSTADDRPOINTER_REG_18_, n67860 );
nand U138694 ( n46810, n46811, n74550 );
nand U138695 ( n46811, n7497, n46812 );
not U138696 ( n7497, n46785 );
nand U138697 ( n46812, P2_P1_INSTADDRPOINTER_REG_18_, n46813 );
nand U138698 ( n25854, n25855, n74575 );
nand U138699 ( n25855, n3953, n25856 );
not U138700 ( n3953, n25829 );
nand U138701 ( n25856, P1_P2_INSTADDRPOINTER_REG_18_, n25857 );
nand U138702 ( n58992, n58993, n74576 );
nand U138703 ( n58993, n6585, n58994 );
not U138704 ( n6585, n58967 );
nand U138705 ( n58994, P2_P2_INSTADDRPOINTER_REG_18_, n58995 );
nand U138706 ( n25625, n25626, n73224 );
nand U138707 ( n25626, n3955, n25627 );
not U138708 ( n3955, n25591 );
nand U138709 ( n25627, P1_P2_INSTADDRPOINTER_REG_24_, n25628 );
nand U138710 ( n58762, n58763, n73225 );
nand U138711 ( n58763, n6588, n58764 );
not U138712 ( n6588, n58728 );
nand U138713 ( n58764, P2_P2_INSTADDRPOINTER_REG_24_, n58765 );
nand U138714 ( n67860, n67836, n67861 );
nand U138715 ( n67861, n67862, P2_P3_INSTADDRPOINTER_REG_17_ );
nand U138716 ( n46813, n46789, n46814 );
nand U138717 ( n46814, n46815, P2_P1_INSTADDRPOINTER_REG_17_ );
nand U138718 ( n25857, n25833, n25858 );
nand U138719 ( n25858, n25859, P1_P2_INSTADDRPOINTER_REG_17_ );
nand U138720 ( n58995, n58971, n58996 );
nand U138721 ( n58996, n58997, P2_P2_INSTADDRPOINTER_REG_17_ );
nand U138722 ( n32872, n32873, n32874 );
nand U138723 ( n32874, n32875, P1_P3_INSTADDRPOINTER_REG_23_ );
nand U138724 ( n32869, n32870, n73232 );
nand U138725 ( n32870, n3112, n32871 );
not U138726 ( n3112, n32831 );
nand U138727 ( n32871, P1_P3_INSTADDRPOINTER_REG_24_, n32872 );
nand U138728 ( n67633, n67634, n67635 );
nand U138729 ( n67635, n67636, P2_P3_INSTADDRPOINTER_REG_23_ );
nand U138730 ( n25628, n25629, n25630 );
nand U138731 ( n25630, n25631, P1_P2_INSTADDRPOINTER_REG_23_ );
nand U138732 ( n58765, n58766, n58767 );
nand U138733 ( n58767, n58768, P2_P2_INSTADDRPOINTER_REG_23_ );
nand U138734 ( n33101, n33102, n74610 );
nand U138735 ( n33102, n3109, n33103 );
not U138736 ( n3109, n33076 );
nand U138737 ( n33103, P1_P3_INSTADDRPOINTER_REG_18_, n33104 );
nand U138738 ( n33104, n33080, n33105 );
nand U138739 ( n33105, n33106, P1_P3_INSTADDRPOINTER_REG_17_ );
nor U138740 ( n15385, n73134, P1_P1_INSTQUEUEWR_ADDR_REG_3_ );
nand U138741 ( n12840, n12764, n12894 );
nand U138742 ( n12894, P1_P1_INSTADDRPOINTER_REG_27_, n12895 );
and U138743 ( n12830, n12840, P1_P1_INSTADDRPOINTER_REG_28_ );
and U138744 ( n15793, n15710, P1_P1_INSTQUEUE_REG_8__7_ );
and U138745 ( n16209, n16129, P1_P1_INSTQUEUE_REG_12__7_ );
and U138746 ( n49238, n49179, P2_P1_INSTQUEUE_REG_12__7_ );
and U138747 ( n48869, n48810, P2_P1_INSTQUEUE_REG_8__7_ );
nor U138748 ( n71008, P1_P2_ADDRESS_REG_2_, n71009 );
nand U138749 ( n27125, n28391, n28392 );
nand U138750 ( n28391, P1_BUF1_REG_31_, n28287 );
nand U138751 ( n28392, P1_BUF2_REG_31_, n28286 );
nand U138752 ( n47315, P2_P1_INSTADDRPOINTER_REG_5_, n76100 );
nand U138753 ( n14739, P1_P1_INSTQUEUEWR_ADDR_REG_3_, n21113 );
nand U138754 ( n21113, n5204, P1_P1_INSTQUEUEWR_ADDR_REG_2_ );
nand U138755 ( n33343, P1_P3_INSTADDRPOINTER_REG_11_, n76127 );
nor U138756 ( n68345, n68299, n68347 );
nand U138757 ( n68347, P2_P3_INSTADDRPOINTER_REG_5_, n76057 );
nor U138758 ( n33589, n33543, n33591 );
nand U138759 ( n33591, P1_P3_INSTADDRPOINTER_REG_5_, n76127 );
nor U138760 ( n26344, n26298, n26346 );
nand U138761 ( n26346, P1_P2_INSTADDRPOINTER_REG_5_, n76155 );
nor U138762 ( n59483, n59437, n59485 );
nand U138763 ( n59485, P2_P2_INSTADDRPOINTER_REG_5_, n76083 );
nand U138764 ( n68100, P2_P3_INSTADDRPOINTER_REG_11_, n76057 );
nand U138765 ( n47069, P2_P1_INSTADDRPOINTER_REG_11_, n76100 );
nand U138766 ( n26097, P1_P2_INSTADDRPOINTER_REG_11_, n76155 );
nand U138767 ( n59238, P2_P2_INSTADDRPOINTER_REG_11_, n76083 );
nand U138768 ( n27062, n28320, n28321 );
nand U138769 ( n28320, n28287, P1_BUF1_REG_26_ );
nand U138770 ( n28321, n28286, P1_BUF2_REG_26_ );
nand U138771 ( n27095, n28363, n28364 );
nand U138772 ( n28363, n28287, P1_BUF1_REG_29_ );
nand U138773 ( n28364, n28286, P1_BUF2_REG_29_ );
nand U138774 ( n27073, n28334, n28335 );
nand U138775 ( n28334, n28287, P1_BUF1_REG_27_ );
nand U138776 ( n28335, n28286, P1_BUF2_REG_27_ );
nand U138777 ( n27051, n28306, n28307 );
nand U138778 ( n28306, n28287, P1_BUF1_REG_25_ );
nand U138779 ( n28307, n28286, P1_BUF2_REG_25_ );
nand U138780 ( n27084, n28349, n28350 );
nand U138781 ( n28349, n28287, P1_BUF1_REG_28_ );
nand U138782 ( n28350, n28286, P1_BUF2_REG_28_ );
nand U138783 ( n27037, n28284, n28285 );
nand U138784 ( n28284, n28287, P1_BUF1_REG_24_ );
nand U138785 ( n28285, n28286, P1_BUF2_REG_24_ );
nand U138786 ( n27106, n28377, n28378 );
nand U138787 ( n28377, n28287, P1_BUF1_REG_30_ );
nand U138788 ( n28378, n28286, P1_BUF2_REG_30_ );
nand U138789 ( n60239, n61640, n61641 );
nand U138790 ( n61640, n61509, P2_BUF1_REG_29_ );
nand U138791 ( n61641, n61508, P2_BUF2_REG_29_ );
nand U138792 ( n60214, n61556, n61557 );
nand U138793 ( n61556, n61509, P2_BUF1_REG_27_ );
nand U138794 ( n61557, n61508, P2_BUF2_REG_27_ );
nand U138795 ( n60203, n61542, n61543 );
nand U138796 ( n61542, n61509, P2_BUF1_REG_26_ );
nand U138797 ( n61543, n61508, P2_BUF2_REG_26_ );
nand U138798 ( n60192, n61528, n61529 );
nand U138799 ( n61528, n61509, P2_BUF1_REG_25_ );
nand U138800 ( n61529, n61508, P2_BUF2_REG_25_ );
nand U138801 ( n60225, n61571, n61572 );
nand U138802 ( n61571, n61509, P2_BUF1_REG_28_ );
nand U138803 ( n61572, n61508, P2_BUF2_REG_28_ );
nand U138804 ( n60250, n61654, n61655 );
nand U138805 ( n61654, n61509, P2_BUF1_REG_30_ );
nand U138806 ( n61655, n61508, P2_BUF2_REG_30_ );
nand U138807 ( n60269, n61672, n61673 );
nand U138808 ( n61672, n61509, P2_BUF1_REG_31_ );
nand U138809 ( n61673, n61508, P2_BUF2_REG_31_ );
nand U138810 ( n60178, n61506, n61507 );
nand U138811 ( n61506, n61509, P2_BUF1_REG_24_ );
nand U138812 ( n61507, n61508, P2_BUF2_REG_24_ );
nor U138813 ( n46515, P2_P1_INSTADDRPOINTER_REG_24_, n7509 );
nor U138814 ( n71016, P2_P2_ADDRESS_REG_2_, n71017 );
nand U138815 ( n9377, n9378, P1_P1_EBX_REG_0_ );
nor U138816 ( n9378, P1_P1_EBX_REG_1_, n8408 );
nor U138817 ( n67912, P2_P3_INSTADDRPOINTER_REG_15_, n5723 );
nor U138818 ( n32930, P1_P3_INSTADDRPOINTER_REG_21_, n3123 );
nor U138819 ( n46865, P2_P1_INSTADDRPOINTER_REG_15_, n7509 );
nor U138820 ( n25909, P1_P2_INSTADDRPOINTER_REG_15_, n3965 );
nor U138821 ( n59047, P2_P2_INSTADDRPOINTER_REG_15_, n6598 );
xnor U138822 ( n54320, n73052, P2_P1_INSTQUEUEWR_ADDR_REG_1_ );
nor U138823 ( n67576, P2_P3_INSTADDRPOINTER_REG_24_, n5723 );
nor U138824 ( n67691, P2_P3_INSTADDRPOINTER_REG_21_, n5723 );
nor U138825 ( n25686, P1_P2_INSTADDRPOINTER_REG_21_, n3965 );
nor U138826 ( n58826, P2_P2_INSTADDRPOINTER_REG_21_, n6598 );
nor U138827 ( n32811, P1_P3_INSTADDRPOINTER_REG_24_, n3123 );
nor U138828 ( n25571, P1_P2_INSTADDRPOINTER_REG_24_, n3965 );
nor U138829 ( n58708, P2_P2_INSTADDRPOINTER_REG_24_, n6598 );
nor U138830 ( n46644, P2_P1_INSTADDRPOINTER_REG_21_, n7509 );
nand U138831 ( n47926, P2_P1_INSTQUEUEWR_ADDR_REG_0_, P2_P1_INSTQUEUEWR_ADDR_REG_1_ );
nand U138832 ( n27497, n28322, n28323 );
nand U138833 ( n28322, n28287, P1_BUF1_REG_18_ );
nand U138834 ( n28323, n28286, P1_BUF2_REG_18_ );
nand U138835 ( n27524, n28365, n28366 );
nand U138836 ( n28365, n28287, P1_BUF1_REG_21_ );
nand U138837 ( n28366, n28286, P1_BUF2_REG_21_ );
nand U138838 ( n27506, n28337, n28338 );
nand U138839 ( n28337, n28287, P1_BUF1_REG_19_ );
nand U138840 ( n28338, n28286, P1_BUF2_REG_19_ );
nand U138841 ( n27488, n28308, n28309 );
nand U138842 ( n28308, n28287, P1_BUF1_REG_17_ );
nand U138843 ( n28309, n28286, P1_BUF2_REG_17_ );
nand U138844 ( n27515, n28351, n28352 );
nand U138845 ( n28351, n28287, P1_BUF1_REG_20_ );
nand U138846 ( n28352, n28286, P1_BUF2_REG_20_ );
nand U138847 ( n27475, n28292, n28293 );
nand U138848 ( n28292, n28287, P1_BUF1_REG_16_ );
nand U138849 ( n28293, n28286, P1_BUF2_REG_16_ );
nand U138850 ( n27533, n28379, n28380 );
nand U138851 ( n28379, n28287, P1_BUF1_REG_22_ );
nand U138852 ( n28380, n28286, P1_BUF2_REG_22_ );
nand U138853 ( n27542, n28393, n28394 );
nand U138854 ( n28393, n28287, P1_BUF1_REG_23_ );
nand U138855 ( n28394, n28286, P1_BUF2_REG_23_ );
nand U138856 ( n60676, n61642, n61643 );
nand U138857 ( n61642, n61509, P2_BUF1_REG_21_ );
nand U138858 ( n61643, n61508, P2_BUF2_REG_21_ );
nand U138859 ( n60655, n61559, n61560 );
nand U138860 ( n61559, n61509, P2_BUF1_REG_19_ );
nand U138861 ( n61560, n61508, P2_BUF2_REG_19_ );
nand U138862 ( n60646, n61544, n61545 );
nand U138863 ( n61544, n61509, P2_BUF1_REG_18_ );
nand U138864 ( n61545, n61508, P2_BUF2_REG_18_ );
nand U138865 ( n60637, n61530, n61531 );
nand U138866 ( n61530, n61509, P2_BUF1_REG_17_ );
nand U138867 ( n61531, n61508, P2_BUF2_REG_17_ );
nand U138868 ( n60664, n61573, n61574 );
nand U138869 ( n61573, n61509, P2_BUF1_REG_20_ );
nand U138870 ( n61574, n61508, P2_BUF2_REG_20_ );
nand U138871 ( n60685, n61656, n61657 );
nand U138872 ( n61656, n61509, P2_BUF1_REG_22_ );
nand U138873 ( n61657, n61508, P2_BUF2_REG_22_ );
nand U138874 ( n60694, n61674, n61675 );
nand U138875 ( n61674, n61509, P2_BUF1_REG_23_ );
nand U138876 ( n61675, n61508, P2_BUF2_REG_23_ );
nand U138877 ( n60624, n61514, n61515 );
nand U138878 ( n61514, n61509, P2_BUF1_REG_16_ );
nand U138879 ( n61515, n61508, P2_BUF2_REG_16_ );
nor U138880 ( n48711, P2_P1_INSTQUEUEWR_ADDR_REG_0_, n73140 );
nor U138881 ( n71019, P2_P3_ADDRESS_REG_2_, n71022 );
nand U138882 ( n43327, n43328, P2_P1_EBX_REG_0_ );
nor U138883 ( n43328, P2_P1_EBX_REG_1_, n42495 );
nand U138884 ( n45171, P3_REG2_REG_9_, n43230 );
nor U138885 ( n71010, P1_P3_ADDRESS_REG_2_, n71013 );
nand U138886 ( n47951, P2_P1_INSTQUEUEWR_ADDR_REG_3_, n54098 );
nand U138887 ( n54098, n7865, P2_P1_INSTQUEUEWR_ADDR_REG_2_ );
nand U138888 ( n45236, P3_REG1_REG_9_, n43230 );
nand U138889 ( n40369, n40370, n40371 );
nor U138890 ( n40370, P4_D_REG_4_, P4_D_REG_3_ );
nor U138891 ( n40371, P4_D_REG_6_, P4_D_REG_5_ );
nor U138892 ( n33156, P1_P3_INSTADDRPOINTER_REG_15_, n3123 );
nor U138893 ( n67450, P2_P3_INSTADDRPOINTER_REG_27_, n5723 );
nor U138894 ( n32685, P1_P3_INSTADDRPOINTER_REG_27_, n3123 );
nor U138895 ( n46386, P2_P1_INSTADDRPOINTER_REG_27_, n7509 );
nor U138896 ( n25445, P1_P2_INSTADDRPOINTER_REG_27_, n3965 );
nor U138897 ( n58582, P2_P2_INSTADDRPOINTER_REG_27_, n6598 );
nor U138898 ( n42518, P2_P1_EBX_REG_30_, n42497 );
nor U138899 ( n21976, P1_P2_EBX_REG_30_, n21952 );
nor U138900 ( n29291, P1_P3_EBX_REG_30_, n29269 );
nor U138901 ( n63058, P2_P3_EBX_REG_30_, n63036 );
nor U138902 ( n55086, P2_P2_EBX_REG_30_, n55064 );
nand U138903 ( n23823, P1_BUF2_REG_16_, n162 );
nor U138904 ( n40374, P4_D_REG_17_, P4_D_REG_16_ );
nand U138905 ( n40386, n40387, n40388 );
nor U138906 ( n40387, P4_D_REG_26_, P4_D_REG_25_ );
nor U138907 ( n40388, P4_D_REG_28_, P4_D_REG_27_ );
nand U138908 ( n68682, P2_P3_INSTADDRPOINTER_REG_0_, n67429 );
nand U138909 ( n33926, P1_P3_INSTADDRPOINTER_REG_0_, n32664 );
nand U138910 ( n26681, P1_P2_INSTADDRPOINTER_REG_0_, n25424 );
nand U138911 ( n59823, P2_P2_INSTADDRPOINTER_REG_0_, n58561 );
nand U138912 ( n47661, P2_P1_INSTADDRPOINTER_REG_0_, n46365 );
nand U138913 ( n14367, P1_P1_INSTADDRPOINTER_REG_0_, n12775 );
nand U138914 ( n7696, n21870, n21871 );
nand U138915 ( n21870, P1_P2_MORE_REG, n168 );
nand U138916 ( n21871, n21872, n21873 );
nand U138917 ( n14431, n54961, n54962 );
nand U138918 ( n54961, P2_P2_MORE_REG, n440 );
nand U138919 ( n54962, n54963, n54964 );
nand U138920 ( n16676, n42396, n42397 );
nand U138921 ( n42396, P2_P1_MORE_REG, n499 );
nand U138922 ( n42397, n42398, n42399 );
nand U138923 ( n5451, n29187, n29188 );
nand U138924 ( n29187, P1_P3_MORE_REG, n202 );
nand U138925 ( n29188, n29189, n29190 );
nand U138926 ( n12186, n62905, n62906 );
nand U138927 ( n62905, P2_P3_MORE_REG, n473 );
nand U138928 ( n62906, n62907, n62908 );
nor U138929 ( n40391, P4_D_REG_13_, P4_D_REG_12_ );
nor U138930 ( n40373, P4_D_REG_15_, P4_D_REG_14_ );
nor U138931 ( n13119, P1_P1_INSTADDRPOINTER_REG_21_, n4864 );
nand U138932 ( n46668, P2_P1_INSTADDRPOINTER_REG_21_, P2_P1_INSTADDRPOINTER_REG_20_ );
nand U138933 ( n46695, P2_P1_INSTADDRPOINTER_REG_19_, n7907 );
nand U138934 ( n40377, n40378, n40379 );
nor U138935 ( n40378, P4_D_REG_2_, P4_D_REG_29_ );
nor U138936 ( n40379, P4_D_REG_31_, P4_D_REG_30_ );
nor U138937 ( n40390, P4_D_REG_11_, P4_D_REG_10_ );
nor U138938 ( n48233, n7863, P2_P1_INSTQUEUEWR_ADDR_REG_0_ );
nand U138939 ( n56948, n434, P2_BUF2_REG_16_ );
nor U138940 ( n33436, P1_P3_INSTADDRPOINTER_REG_8_, n3088 );
nor U138941 ( n68183, P2_P3_INSTADDRPOINTER_REG_8_, n5689 );
nor U138942 ( n47152, P2_P1_INSTADDRPOINTER_REG_8_, n7474 );
nor U138943 ( n26182, P1_P2_INSTADDRPOINTER_REG_8_, n3932 );
nor U138944 ( n59321, P2_P2_INSTADDRPOINTER_REG_8_, n6564 );
nand U138945 ( n33375, n33376, n74458 );
nand U138946 ( n33376, n3119, n33377 );
nand U138947 ( n33377, P1_P3_INSTADDRPOINTER_REG_11_, n33378 );
nand U138948 ( n68127, n68128, n74438 );
nand U138949 ( n68128, n5720, n68129 );
nand U138950 ( n68129, P2_P3_INSTADDRPOINTER_REG_11_, n68130 );
nand U138951 ( n47096, n47097, n74427 );
nand U138952 ( n47097, n7507, n47098 );
nand U138953 ( n47098, P2_P1_INSTADDRPOINTER_REG_11_, n47099 );
nand U138954 ( n26124, n26125, n74439 );
nand U138955 ( n26125, n3963, n26126 );
nand U138956 ( n26126, P1_P2_INSTADDRPOINTER_REG_11_, n26127 );
nand U138957 ( n59265, n59266, n74440 );
nand U138958 ( n59266, n6595, n59267 );
nand U138959 ( n59267, P2_P2_INSTADDRPOINTER_REG_11_, n59268 );
nor U138960 ( n40381, P4_D_REG_9_, P4_D_REG_8_ );
nor U138961 ( n13409, P1_P1_INSTADDRPOINTER_REG_15_, n4864 );
nor U138962 ( n48515, n73133, P2_P1_INSTQUEUEWR_ADDR_REG_3_ );
nor U138963 ( n32853, P1_P3_INSTADDRPOINTER_REG_23_, n3088 );
nand U138964 ( n9941, n8312, n8313 );
nand U138965 ( n8312, P1_P1_MORE_REG, n228 );
nand U138966 ( n8313, n8314, n8315 );
nand U138967 ( n60086, P2_P2_INSTQUEUEWR_ADDR_REG_0_, P2_P2_INSTQUEUEWR_ADDR_REG_1_ );
nand U138968 ( n26946, P1_P2_INSTQUEUEWR_ADDR_REG_0_, P1_P2_INSTQUEUEWR_ADDR_REG_1_ );
nand U138969 ( n67715, P2_P3_INSTADDRPOINTER_REG_21_, P2_P3_INSTADDRPOINTER_REG_20_ );
nand U138970 ( n25710, P1_P2_INSTADDRPOINTER_REG_21_, P1_P2_INSTADDRPOINTER_REG_20_ );
nand U138971 ( n58850, P2_P2_INSTADDRPOINTER_REG_21_, P2_P2_INSTADDRPOINTER_REG_20_ );
nand U138972 ( n67742, P2_P3_INSTADDRPOINTER_REG_19_, n6118 );
nand U138973 ( n25737, P1_P2_INSTADDRPOINTER_REG_19_, n4340 );
nand U138974 ( n58877, P2_P2_INSTADDRPOINTER_REG_19_, n6973 );
nor U138975 ( n67618, P2_P3_INSTADDRPOINTER_REG_23_, n5689 );
nor U138976 ( n25613, P1_P2_INSTADDRPOINTER_REG_23_, n3932 );
nor U138977 ( n58750, P2_P2_INSTADDRPOINTER_REG_23_, n6564 );
nand U138978 ( n28265, n28266, n28267 );
nand U138979 ( n28267, n28203, n27542 );
nand U138980 ( n28266, P1_P2_INSTQUEUE_REG_14__7_, n28204 );
nand U138981 ( n61487, n61488, n61489 );
nand U138982 ( n61489, n61367, n60694 );
nand U138983 ( n61488, P2_P2_INSTQUEUE_REG_14__7_, n61368 );
nand U138984 ( n34191, P1_P3_INSTQUEUEWR_ADDR_REG_0_, P1_P3_INSTQUEUEWR_ADDR_REG_1_ );
nand U138985 ( n68945, P2_P3_INSTQUEUEWR_ADDR_REG_0_, P2_P3_INSTQUEUEWR_ADDR_REG_1_ );
nor U138986 ( n46805, P2_P1_INSTADDRPOINTER_REG_17_, n7474 );
nor U138987 ( n25849, P1_P2_INSTADDRPOINTER_REG_17_, n3932 );
nor U138988 ( n58987, P2_P2_INSTADDRPOINTER_REG_17_, n6564 );
nand U138989 ( n28245, n28246, n28247 );
nand U138990 ( n28247, n28203, n27524 );
nand U138991 ( n28246, P1_P2_INSTQUEUE_REG_14__5_, n28204 );
nand U138992 ( n61471, n61472, n61473 );
nand U138993 ( n61473, n61367, n60676 );
nand U138994 ( n61472, P2_P2_INSTQUEUE_REG_14__5_, n61368 );
nor U138995 ( n67852, P2_P3_INSTADDRPOINTER_REG_17_, n5689 );
nand U138996 ( n35433, n35434, n35435 );
nand U138997 ( n35435, n35436, n112 );
nand U138998 ( n35434, P1_P3_INSTQUEUE_REG_14__0_, n35437 );
nand U138999 ( n27940, n27941, n27942 );
nand U139000 ( n27942, n27882, n27542 );
nand U139001 ( n27941, P1_P2_INSTQUEUE_REG_10__7_, n27883 );
nand U139002 ( n27924, n27925, n27926 );
nand U139003 ( n27926, n27882, n27524 );
nand U139004 ( n27925, P1_P2_INSTQUEUE_REG_10__5_, n27883 );
nand U139005 ( n61077, n61078, n61079 );
nand U139006 ( n61079, n61029, n60676 );
nand U139007 ( n61078, P2_P2_INSTQUEUE_REG_10__5_, n61030 );
nand U139008 ( n61093, n61094, n61095 );
nand U139009 ( n61095, n61029, n60694 );
nand U139010 ( n61094, P2_P2_INSTQUEUE_REG_10__7_, n61030 );
nand U139011 ( n35118, n35119, n35120 );
nand U139012 ( n35120, n35121, n112 );
nand U139013 ( n35119, P1_P3_INSTQUEUE_REG_10__0_, n35122 );
nand U139014 ( n70163, n70164, n70165 );
nand U139015 ( n70165, n70166, n383 );
nand U139016 ( n70164, P2_P3_INSTQUEUE_REG_14__0_, n70167 );
nand U139017 ( n69854, n69855, n69856 );
nand U139018 ( n69856, n69857, n383 );
nand U139019 ( n69855, P2_P3_INSTQUEUE_REG_10__0_, n69858 );
nand U139020 ( n27932, n27933, n27934 );
nand U139021 ( n27934, n27882, n27533 );
nand U139022 ( n27933, P1_P2_INSTQUEUE_REG_10__6_, n27883 );
nand U139023 ( n28200, n28201, n28202 );
nand U139024 ( n28202, n28203, n27475 );
nand U139025 ( n28201, P1_P2_INSTQUEUE_REG_14__0_, n28204 );
nand U139026 ( n27879, n27880, n27881 );
nand U139027 ( n27881, n27882, n27475 );
nand U139028 ( n27880, P1_P2_INSTQUEUE_REG_10__0_, n27883 );
nand U139029 ( n61479, n61480, n61481 );
nand U139030 ( n61481, n61367, n60685 );
nand U139031 ( n61480, P2_P2_INSTQUEUE_REG_14__6_, n61368 );
nand U139032 ( n61085, n61086, n61087 );
nand U139033 ( n61087, n61029, n60685 );
nand U139034 ( n61086, P2_P2_INSTQUEUE_REG_10__6_, n61030 );
nand U139035 ( n61364, n61365, n61366 );
nand U139036 ( n61366, n61367, n60624 );
nand U139037 ( n61365, P2_P2_INSTQUEUE_REG_14__0_, n61368 );
nand U139038 ( n61026, n61027, n61028 );
nand U139039 ( n61028, n61029, n60624 );
nand U139040 ( n61027, P2_P2_INSTQUEUE_REG_10__0_, n61030 );
nand U139041 ( n28257, n28258, n28259 );
nand U139042 ( n28259, n28203, n27533 );
nand U139043 ( n28258, P1_P2_INSTQUEUE_REG_14__6_, n28204 );
nand U139044 ( n35446, n35447, n35448 );
nand U139045 ( n35448, n35436, n114 );
nand U139046 ( n35447, P1_P3_INSTQUEUE_REG_14__1_, n35437 );
nand U139047 ( n35163, n35164, n35165 );
nand U139048 ( n35165, n35121, n123 );
nand U139049 ( n35164, P1_P3_INSTQUEUE_REG_10__5_, n35122 );
nand U139050 ( n35478, n35479, n35480 );
nand U139051 ( n35480, n35436, n123 );
nand U139052 ( n35479, P1_P3_INSTQUEUE_REG_14__5_, n35437 );
nand U139053 ( n35171, n35172, n35173 );
nand U139054 ( n35173, n35121, n125 );
nand U139055 ( n35172, P1_P3_INSTQUEUE_REG_10__6_, n35122 );
nand U139056 ( n35486, n35487, n35488 );
nand U139057 ( n35488, n35436, n125 );
nand U139058 ( n35487, P1_P3_INSTQUEUE_REG_14__6_, n35437 );
nand U139059 ( n35496, n35497, n35498 );
nand U139060 ( n35498, n35436, n128 );
nand U139061 ( n35497, P1_P3_INSTQUEUE_REG_14__7_, n35437 );
nand U139062 ( n35179, n35180, n35181 );
nand U139063 ( n35181, n35121, n128 );
nand U139064 ( n35180, P1_P3_INSTQUEUE_REG_10__7_, n35122 );
nand U139065 ( n35462, n35463, n35464 );
nand U139066 ( n35464, n35436, n118 );
nand U139067 ( n35463, P1_P3_INSTQUEUE_REG_14__3_, n35437 );
nand U139068 ( n35147, n35148, n35149 );
nand U139069 ( n35149, n35121, n118 );
nand U139070 ( n35148, P1_P3_INSTQUEUE_REG_10__3_, n35122 );
nand U139071 ( n35470, n35471, n35472 );
nand U139072 ( n35472, n35436, n120 );
nand U139073 ( n35471, P1_P3_INSTQUEUE_REG_14__4_, n35437 );
nand U139074 ( n35155, n35156, n35157 );
nand U139075 ( n35157, n35121, n120 );
nand U139076 ( n35156, P1_P3_INSTQUEUE_REG_10__4_, n35122 );
nand U139077 ( n35139, n35140, n35141 );
nand U139078 ( n35141, n35121, n116 );
nand U139079 ( n35140, P1_P3_INSTQUEUE_REG_10__2_, n35122 );
nand U139080 ( n70176, n70177, n70178 );
nand U139081 ( n70178, n70166, n385 );
nand U139082 ( n70177, P2_P3_INSTQUEUE_REG_14__1_, n70167 );
nand U139083 ( n69867, n69868, n69869 );
nand U139084 ( n69869, n69857, n385 );
nand U139085 ( n69868, P2_P3_INSTQUEUE_REG_10__1_, n69858 );
nand U139086 ( n69875, n69876, n69877 );
nand U139087 ( n69877, n69857, n388 );
nand U139088 ( n69876, P2_P3_INSTQUEUE_REG_10__2_, n69858 );
nand U139089 ( n70192, n70193, n70194 );
nand U139090 ( n70194, n70166, n390 );
nand U139091 ( n70193, P2_P3_INSTQUEUE_REG_14__3_, n70167 );
nand U139092 ( n69907, n69908, n69909 );
nand U139093 ( n69909, n69857, n398 );
nand U139094 ( n69908, P2_P3_INSTQUEUE_REG_10__6_, n69858 );
nand U139095 ( n70216, n70217, n70218 );
nand U139096 ( n70218, n70166, n398 );
nand U139097 ( n70217, P2_P3_INSTQUEUE_REG_14__6_, n70167 );
nand U139098 ( n70224, n70225, n70226 );
nand U139099 ( n70226, n70166, n400 );
nand U139100 ( n70225, P2_P3_INSTQUEUE_REG_14__7_, n70167 );
nand U139101 ( n70200, n70201, n70202 );
nand U139102 ( n70202, n70166, n393 );
nand U139103 ( n70201, P2_P3_INSTQUEUE_REG_14__4_, n70167 );
nand U139104 ( n35454, n35455, n35456 );
nand U139105 ( n35456, n35436, n116 );
nand U139106 ( n35455, P1_P3_INSTQUEUE_REG_14__2_, n35437 );
nand U139107 ( n35131, n35132, n35133 );
nand U139108 ( n35133, n35121, n114 );
nand U139109 ( n35132, P1_P3_INSTQUEUE_REG_10__1_, n35122 );
nand U139110 ( n69883, n69884, n69885 );
nand U139111 ( n69885, n69857, n390 );
nand U139112 ( n69884, P2_P3_INSTQUEUE_REG_10__3_, n69858 );
nand U139113 ( n69915, n69916, n69917 );
nand U139114 ( n69917, n69857, n400 );
nand U139115 ( n69916, P2_P3_INSTQUEUE_REG_10__7_, n69858 );
nand U139116 ( n69899, n69900, n69901 );
nand U139117 ( n69901, n69857, n395 );
nand U139118 ( n69900, P2_P3_INSTQUEUE_REG_10__5_, n69858 );
nand U139119 ( n70208, n70209, n70210 );
nand U139120 ( n70210, n70166, n395 );
nand U139121 ( n70209, P2_P3_INSTQUEUE_REG_14__5_, n70167 );
nand U139122 ( n69891, n69892, n69893 );
nand U139123 ( n69893, n69857, n393 );
nand U139124 ( n69892, P2_P3_INSTQUEUE_REG_10__4_, n69858 );
nand U139125 ( n70184, n70185, n70186 );
nand U139126 ( n70186, n70166, n388 );
nand U139127 ( n70185, P2_P3_INSTQUEUE_REG_14__2_, n70167 );
nand U139128 ( n27892, n27893, n27894 );
nand U139129 ( n27894, n27882, n27488 );
nand U139130 ( n27893, P1_P2_INSTQUEUE_REG_10__1_, n27883 );
nand U139131 ( n28229, n28230, n28231 );
nand U139132 ( n28231, n28203, n27506 );
nand U139133 ( n28230, P1_P2_INSTQUEUE_REG_14__3_, n28204 );
nand U139134 ( n27908, n27909, n27910 );
nand U139135 ( n27910, n27882, n27506 );
nand U139136 ( n27909, P1_P2_INSTQUEUE_REG_10__3_, n27883 );
nand U139137 ( n28237, n28238, n28239 );
nand U139138 ( n28239, n28203, n27515 );
nand U139139 ( n28238, P1_P2_INSTQUEUE_REG_14__4_, n28204 );
nand U139140 ( n27916, n27917, n27918 );
nand U139141 ( n27918, n27882, n27515 );
nand U139142 ( n27917, P1_P2_INSTQUEUE_REG_10__4_, n27883 );
nand U139143 ( n28221, n28222, n28223 );
nand U139144 ( n28223, n28203, n27497 );
nand U139145 ( n28222, P1_P2_INSTQUEUE_REG_14__2_, n28204 );
nand U139146 ( n27900, n27901, n27902 );
nand U139147 ( n27902, n27882, n27497 );
nand U139148 ( n27901, P1_P2_INSTQUEUE_REG_10__2_, n27883 );
nand U139149 ( n61055, n61056, n61057 );
nand U139150 ( n61057, n61029, n60655 );
nand U139151 ( n61056, P2_P2_INSTQUEUE_REG_10__3_, n61030 );
nand U139152 ( n61377, n61378, n61379 );
nand U139153 ( n61379, n61367, n60637 );
nand U139154 ( n61378, P2_P2_INSTQUEUE_REG_14__1_, n61368 );
nand U139155 ( n61385, n61386, n61387 );
nand U139156 ( n61387, n61367, n60646 );
nand U139157 ( n61386, P2_P2_INSTQUEUE_REG_14__2_, n61368 );
nand U139158 ( n61047, n61048, n61049 );
nand U139159 ( n61049, n61029, n60646 );
nand U139160 ( n61048, P2_P2_INSTQUEUE_REG_10__2_, n61030 );
nand U139161 ( n61463, n61464, n61465 );
nand U139162 ( n61465, n61367, n60664 );
nand U139163 ( n61464, P2_P2_INSTQUEUE_REG_14__4_, n61368 );
nand U139164 ( n61063, n61064, n61065 );
nand U139165 ( n61065, n61029, n60664 );
nand U139166 ( n61064, P2_P2_INSTQUEUE_REG_10__4_, n61030 );
nand U139167 ( n61455, n61456, n61457 );
nand U139168 ( n61457, n61367, n60655 );
nand U139169 ( n61456, P2_P2_INSTQUEUE_REG_14__3_, n61368 );
nand U139170 ( n28213, n28214, n28215 );
nand U139171 ( n28215, n28203, n27488 );
nand U139172 ( n28214, P1_P2_INSTQUEUE_REG_14__1_, n28204 );
nand U139173 ( n61039, n61040, n61041 );
nand U139174 ( n61041, n61029, n60637 );
nand U139175 ( n61040, P2_P2_INSTQUEUE_REG_10__1_, n61030 );
and U139176 ( n14267, n14270, P1_P1_INSTADDRPOINTER_REG_3_ );
nor U139177 ( n33096, P1_P3_INSTADDRPOINTER_REG_17_, n3088 );
nor U139178 ( n46571, P2_P1_INSTADDRPOINTER_REG_23_, n7474 );
nand U139179 ( n69063, n70243, P2_BUF2_REG_18_ );
nand U139180 ( n69074, n70243, P2_BUF2_REG_19_ );
nand U139181 ( n69107, n70243, P2_BUF2_REG_22_ );
nand U139182 ( n69096, n70243, P2_BUF2_REG_21_ );
nand U139183 ( n69085, n70243, P2_BUF2_REG_20_ );
nand U139184 ( n69041, n70243, P2_BUF2_REG_16_ );
nand U139185 ( n69131, n70243, P2_BUF2_REG_23_ );
nand U139186 ( n69052, n70243, P2_BUF2_REG_17_ );
nand U139187 ( n34344, n35515, P1_BUF2_REG_21_ );
nand U139188 ( n34355, n35515, P1_BUF2_REG_22_ );
nand U139189 ( n34322, n35515, P1_BUF2_REG_19_ );
nand U139190 ( n34333, n35515, P1_BUF2_REG_20_ );
nand U139191 ( n34311, n35515, P1_BUF2_REG_18_ );
nand U139192 ( n34289, n35515, P1_BUF2_REG_16_ );
nand U139193 ( n34379, n35515, P1_BUF2_REG_23_ );
nand U139194 ( n34300, n35515, P1_BUF2_REG_17_ );
nand U139195 ( n35287, n35288, n35289 );
nand U139196 ( n35288, P1_P3_INSTQUEUE_REG_12__1_, n35278 );
nand U139197 ( n35289, n35277, n114 );
nand U139198 ( n34970, n34971, n34972 );
nand U139199 ( n34971, P1_P3_INSTQUEUE_REG_8__1_, n34961 );
nand U139200 ( n34972, n34960, n114 );
nand U139201 ( n35321, n35322, n35323 );
nand U139202 ( n35322, P1_P3_INSTQUEUE_REG_12__5_, n35278 );
nand U139203 ( n35323, n35277, n123 );
nand U139204 ( n35004, n35005, n35006 );
nand U139205 ( n35005, P1_P3_INSTQUEUE_REG_8__5_, n34961 );
nand U139206 ( n35006, n34960, n123 );
nand U139207 ( n35329, n35330, n35331 );
nand U139208 ( n35330, P1_P3_INSTQUEUE_REG_12__6_, n35278 );
nand U139209 ( n35331, n35277, n125 );
nand U139210 ( n35012, n35013, n35014 );
nand U139211 ( n35013, P1_P3_INSTQUEUE_REG_8__6_, n34961 );
nand U139212 ( n35014, n34960, n125 );
nand U139213 ( n35337, n35338, n35339 );
nand U139214 ( n35338, P1_P3_INSTQUEUE_REG_12__7_, n35278 );
nand U139215 ( n35339, n35277, n128 );
nand U139216 ( n35020, n35021, n35022 );
nand U139217 ( n35021, P1_P3_INSTQUEUE_REG_8__7_, n34961 );
nand U139218 ( n35022, n34960, n128 );
nand U139219 ( n35305, n35306, n35307 );
nand U139220 ( n35306, P1_P3_INSTQUEUE_REG_12__3_, n35278 );
nand U139221 ( n35307, n35277, n118 );
nand U139222 ( n34986, n34987, n34988 );
nand U139223 ( n34987, P1_P3_INSTQUEUE_REG_8__3_, n34961 );
nand U139224 ( n34988, n34960, n118 );
nand U139225 ( n35313, n35314, n35315 );
nand U139226 ( n35314, P1_P3_INSTQUEUE_REG_12__4_, n35278 );
nand U139227 ( n35315, n35277, n120 );
nand U139228 ( n34994, n34995, n34996 );
nand U139229 ( n34995, P1_P3_INSTQUEUE_REG_8__4_, n34961 );
nand U139230 ( n34996, n34960, n120 );
nand U139231 ( n35354, n35355, n35356 );
nand U139232 ( n35355, P1_P3_INSTQUEUE_REG_13__0_, n35358 );
nand U139233 ( n35356, n35357, n112 );
nand U139234 ( n35196, n35197, n35198 );
nand U139235 ( n35197, P1_P3_INSTQUEUE_REG_11__0_, n35200 );
nand U139236 ( n35198, n35199, n112 );
nand U139237 ( n35038, n35039, n35040 );
nand U139238 ( n35039, P1_P3_INSTQUEUE_REG_9__0_, n35042 );
nand U139239 ( n35040, n35041, n112 );
nand U139240 ( n34801, n34802, n34803 );
nand U139241 ( n34802, P1_P3_INSTQUEUE_REG_6__0_, n34805 );
nand U139242 ( n34803, n34804, n112 );
nand U139243 ( n34716, n34717, n34718 );
nand U139244 ( n34717, P1_P3_INSTQUEUE_REG_5__0_, n34720 );
nand U139245 ( n34718, n34719, n112 );
nand U139246 ( n35295, n35296, n35297 );
nand U139247 ( n35296, P1_P3_INSTQUEUE_REG_12__2_, n35278 );
nand U139248 ( n35297, n35277, n116 );
nand U139249 ( n34978, n34979, n34980 );
nand U139250 ( n34979, P1_P3_INSTQUEUE_REG_8__2_, n34961 );
nand U139251 ( n34980, n34960, n116 );
nand U139252 ( n70021, n70022, n70023 );
nand U139253 ( n70022, P2_P3_INSTQUEUE_REG_12__1_, n70012 );
nand U139254 ( n70023, n70011, n385 );
nand U139255 ( n69710, n69711, n69712 );
nand U139256 ( n69711, P2_P3_INSTQUEUE_REG_8__1_, n69701 );
nand U139257 ( n69712, n69700, n385 );
nand U139258 ( n70029, n70030, n70031 );
nand U139259 ( n70030, P2_P3_INSTQUEUE_REG_12__2_, n70012 );
nand U139260 ( n70031, n70011, n388 );
nand U139261 ( n69718, n69719, n69720 );
nand U139262 ( n69719, P2_P3_INSTQUEUE_REG_8__2_, n69701 );
nand U139263 ( n69720, n69700, n388 );
nand U139264 ( n70037, n70038, n70039 );
nand U139265 ( n70038, P2_P3_INSTQUEUE_REG_12__3_, n70012 );
nand U139266 ( n70039, n70011, n390 );
nand U139267 ( n69726, n69727, n69728 );
nand U139268 ( n69727, P2_P3_INSTQUEUE_REG_8__3_, n69701 );
nand U139269 ( n69728, n69700, n390 );
nand U139270 ( n70061, n70062, n70063 );
nand U139271 ( n70062, P2_P3_INSTQUEUE_REG_12__6_, n70012 );
nand U139272 ( n70063, n70011, n398 );
nand U139273 ( n69750, n69751, n69752 );
nand U139274 ( n69751, P2_P3_INSTQUEUE_REG_8__6_, n69701 );
nand U139275 ( n69752, n69700, n398 );
nand U139276 ( n70069, n70070, n70071 );
nand U139277 ( n70070, P2_P3_INSTQUEUE_REG_12__7_, n70012 );
nand U139278 ( n70071, n70011, n400 );
nand U139279 ( n69758, n69759, n69760 );
nand U139280 ( n69759, P2_P3_INSTQUEUE_REG_8__7_, n69701 );
nand U139281 ( n69760, n69700, n400 );
nand U139282 ( n70053, n70054, n70055 );
nand U139283 ( n70054, P2_P3_INSTQUEUE_REG_12__5_, n70012 );
nand U139284 ( n70055, n70011, n395 );
nand U139285 ( n69742, n69743, n69744 );
nand U139286 ( n69743, P2_P3_INSTQUEUE_REG_8__5_, n69701 );
nand U139287 ( n69744, n69700, n395 );
nand U139288 ( n70045, n70046, n70047 );
nand U139289 ( n70046, P2_P3_INSTQUEUE_REG_12__4_, n70012 );
nand U139290 ( n70047, n70011, n393 );
nand U139291 ( n69734, n69735, n69736 );
nand U139292 ( n69735, P2_P3_INSTQUEUE_REG_8__4_, n69701 );
nand U139293 ( n69736, n69700, n393 );
nand U139294 ( n70086, n70087, n70088 );
nand U139295 ( n70087, P2_P3_INSTQUEUE_REG_13__0_, n70090 );
nand U139296 ( n70088, n70089, n383 );
nand U139297 ( n69932, n69933, n69934 );
nand U139298 ( n69933, P2_P3_INSTQUEUE_REG_11__0_, n69936 );
nand U139299 ( n69934, n69935, n383 );
nand U139300 ( n69776, n69777, n69778 );
nand U139301 ( n69777, P2_P3_INSTQUEUE_REG_9__0_, n69780 );
nand U139302 ( n69778, n69779, n383 );
nand U139303 ( n69545, n69546, n69547 );
nand U139304 ( n69546, P2_P3_INSTQUEUE_REG_6__0_, n69549 );
nand U139305 ( n69547, n69548, n383 );
nand U139306 ( n69460, n69461, n69462 );
nand U139307 ( n69461, P2_P3_INSTQUEUE_REG_5__0_, n69464 );
nand U139308 ( n69462, n69463, n383 );
nand U139309 ( n35367, n35368, n35369 );
nand U139310 ( n35368, P1_P3_INSTQUEUE_REG_13__1_, n35358 );
nand U139311 ( n35369, n35357, n114 );
nand U139312 ( n35211, n35212, n35213 );
nand U139313 ( n35212, P1_P3_INSTQUEUE_REG_11__1_, n35200 );
nand U139314 ( n35213, n35199, n114 );
nand U139315 ( n35051, n35052, n35053 );
nand U139316 ( n35052, P1_P3_INSTQUEUE_REG_9__1_, n35042 );
nand U139317 ( n35053, n35041, n114 );
nand U139318 ( n34816, n34817, n34818 );
nand U139319 ( n34817, P1_P3_INSTQUEUE_REG_6__1_, n34805 );
nand U139320 ( n34818, n34804, n114 );
nand U139321 ( n34730, n34731, n34732 );
nand U139322 ( n34731, P1_P3_INSTQUEUE_REG_5__1_, n34720 );
nand U139323 ( n34732, n34719, n114 );
nand U139324 ( n35401, n35402, n35403 );
nand U139325 ( n35402, P1_P3_INSTQUEUE_REG_13__5_, n35358 );
nand U139326 ( n35403, n35357, n123 );
nand U139327 ( n35243, n35244, n35245 );
nand U139328 ( n35244, P1_P3_INSTQUEUE_REG_11__5_, n35200 );
nand U139329 ( n35245, n35199, n123 );
nand U139330 ( n35083, n35084, n35085 );
nand U139331 ( n35084, P1_P3_INSTQUEUE_REG_9__5_, n35042 );
nand U139332 ( n35085, n35041, n123 );
nand U139333 ( n34848, n34849, n34850 );
nand U139334 ( n34849, P1_P3_INSTQUEUE_REG_6__5_, n34805 );
nand U139335 ( n34850, n34804, n123 );
nand U139336 ( n34766, n34767, n34768 );
nand U139337 ( n34767, P1_P3_INSTQUEUE_REG_5__5_, n34720 );
nand U139338 ( n34768, n34719, n123 );
nand U139339 ( n35409, n35410, n35411 );
nand U139340 ( n35410, P1_P3_INSTQUEUE_REG_13__6_, n35358 );
nand U139341 ( n35411, n35357, n125 );
nand U139342 ( n35251, n35252, n35253 );
nand U139343 ( n35252, P1_P3_INSTQUEUE_REG_11__6_, n35200 );
nand U139344 ( n35253, n35199, n125 );
nand U139345 ( n35091, n35092, n35093 );
nand U139346 ( n35092, P1_P3_INSTQUEUE_REG_9__6_, n35042 );
nand U139347 ( n35093, n35041, n125 );
nand U139348 ( n34856, n34857, n34858 );
nand U139349 ( n34857, P1_P3_INSTQUEUE_REG_6__6_, n34805 );
nand U139350 ( n34858, n34804, n125 );
nand U139351 ( n34775, n34776, n34777 );
nand U139352 ( n34776, P1_P3_INSTQUEUE_REG_5__6_, n34720 );
nand U139353 ( n34777, n34719, n125 );
nand U139354 ( n35417, n35418, n35419 );
nand U139355 ( n35418, P1_P3_INSTQUEUE_REG_13__7_, n35358 );
nand U139356 ( n35419, n35357, n128 );
nand U139357 ( n35259, n35260, n35261 );
nand U139358 ( n35260, P1_P3_INSTQUEUE_REG_11__7_, n35200 );
nand U139359 ( n35261, n35199, n128 );
nand U139360 ( n35101, n35102, n35103 );
nand U139361 ( n35102, P1_P3_INSTQUEUE_REG_9__7_, n35042 );
nand U139362 ( n35103, n35041, n128 );
nand U139363 ( n34864, n34865, n34866 );
nand U139364 ( n34865, P1_P3_INSTQUEUE_REG_6__7_, n34805 );
nand U139365 ( n34866, n34804, n128 );
nand U139366 ( n34784, n34785, n34786 );
nand U139367 ( n34785, P1_P3_INSTQUEUE_REG_5__7_, n34720 );
nand U139368 ( n34786, n34719, n128 );
nand U139369 ( n35383, n35384, n35385 );
nand U139370 ( n35384, P1_P3_INSTQUEUE_REG_13__3_, n35358 );
nand U139371 ( n35385, n35357, n118 );
nand U139372 ( n35227, n35228, n35229 );
nand U139373 ( n35228, P1_P3_INSTQUEUE_REG_11__3_, n35200 );
nand U139374 ( n35229, n35199, n118 );
nand U139375 ( n35067, n35068, n35069 );
nand U139376 ( n35068, P1_P3_INSTQUEUE_REG_9__3_, n35042 );
nand U139377 ( n35069, n35041, n118 );
nand U139378 ( n34832, n34833, n34834 );
nand U139379 ( n34833, P1_P3_INSTQUEUE_REG_6__3_, n34805 );
nand U139380 ( n34834, n34804, n118 );
nand U139381 ( n34748, n34749, n34750 );
nand U139382 ( n34749, P1_P3_INSTQUEUE_REG_5__3_, n34720 );
nand U139383 ( n34750, n34719, n118 );
nand U139384 ( n35391, n35392, n35393 );
nand U139385 ( n35392, P1_P3_INSTQUEUE_REG_13__4_, n35358 );
nand U139386 ( n35393, n35357, n120 );
nand U139387 ( n35235, n35236, n35237 );
nand U139388 ( n35236, P1_P3_INSTQUEUE_REG_11__4_, n35200 );
nand U139389 ( n35237, n35199, n120 );
nand U139390 ( n35075, n35076, n35077 );
nand U139391 ( n35076, P1_P3_INSTQUEUE_REG_9__4_, n35042 );
nand U139392 ( n35077, n35041, n120 );
nand U139393 ( n34840, n34841, n34842 );
nand U139394 ( n34841, P1_P3_INSTQUEUE_REG_6__4_, n34805 );
nand U139395 ( n34842, n34804, n120 );
nand U139396 ( n34757, n34758, n34759 );
nand U139397 ( n34758, P1_P3_INSTQUEUE_REG_5__4_, n34720 );
nand U139398 ( n34759, n34719, n120 );
nand U139399 ( n35274, n35275, n35276 );
nand U139400 ( n35275, P1_P3_INSTQUEUE_REG_12__0_, n35278 );
nand U139401 ( n35276, n35277, n112 );
nand U139402 ( n34957, n34958, n34959 );
nand U139403 ( n34958, P1_P3_INSTQUEUE_REG_8__0_, n34961 );
nand U139404 ( n34959, n34960, n112 );
nand U139405 ( n35375, n35376, n35377 );
nand U139406 ( n35376, P1_P3_INSTQUEUE_REG_13__2_, n35358 );
nand U139407 ( n35377, n35357, n116 );
nand U139408 ( n35219, n35220, n35221 );
nand U139409 ( n35220, P1_P3_INSTQUEUE_REG_11__2_, n35200 );
nand U139410 ( n35221, n35199, n116 );
nand U139411 ( n35059, n35060, n35061 );
nand U139412 ( n35060, P1_P3_INSTQUEUE_REG_9__2_, n35042 );
nand U139413 ( n35061, n35041, n116 );
nand U139414 ( n34824, n34825, n34826 );
nand U139415 ( n34825, P1_P3_INSTQUEUE_REG_6__2_, n34805 );
nand U139416 ( n34826, n34804, n116 );
nand U139417 ( n34739, n34740, n34741 );
nand U139418 ( n34740, P1_P3_INSTQUEUE_REG_5__2_, n34720 );
nand U139419 ( n34741, n34719, n116 );
nand U139420 ( n70099, n70100, n70101 );
nand U139421 ( n70100, P2_P3_INSTQUEUE_REG_13__1_, n70090 );
nand U139422 ( n70101, n70089, n385 );
nand U139423 ( n69945, n69946, n69947 );
nand U139424 ( n69946, P2_P3_INSTQUEUE_REG_11__1_, n69936 );
nand U139425 ( n69947, n69935, n385 );
nand U139426 ( n69789, n69790, n69791 );
nand U139427 ( n69790, P2_P3_INSTQUEUE_REG_9__1_, n69780 );
nand U139428 ( n69791, n69779, n385 );
nand U139429 ( n69558, n69559, n69560 );
nand U139430 ( n69559, P2_P3_INSTQUEUE_REG_6__1_, n69549 );
nand U139431 ( n69560, n69548, n385 );
nand U139432 ( n69474, n69475, n69476 );
nand U139433 ( n69475, P2_P3_INSTQUEUE_REG_5__1_, n69464 );
nand U139434 ( n69476, n69463, n385 );
nand U139435 ( n70107, n70108, n70109 );
nand U139436 ( n70108, P2_P3_INSTQUEUE_REG_13__2_, n70090 );
nand U139437 ( n70109, n70089, n388 );
nand U139438 ( n69953, n69954, n69955 );
nand U139439 ( n69954, P2_P3_INSTQUEUE_REG_11__2_, n69936 );
nand U139440 ( n69955, n69935, n388 );
nand U139441 ( n69797, n69798, n69799 );
nand U139442 ( n69798, P2_P3_INSTQUEUE_REG_9__2_, n69780 );
nand U139443 ( n69799, n69779, n388 );
nand U139444 ( n69566, n69567, n69568 );
nand U139445 ( n69567, P2_P3_INSTQUEUE_REG_6__2_, n69549 );
nand U139446 ( n69568, n69548, n388 );
nand U139447 ( n69483, n69484, n69485 );
nand U139448 ( n69484, P2_P3_INSTQUEUE_REG_5__2_, n69464 );
nand U139449 ( n69485, n69463, n388 );
nand U139450 ( n70115, n70116, n70117 );
nand U139451 ( n70116, P2_P3_INSTQUEUE_REG_13__3_, n70090 );
nand U139452 ( n70117, n70089, n390 );
nand U139453 ( n69961, n69962, n69963 );
nand U139454 ( n69962, P2_P3_INSTQUEUE_REG_11__3_, n69936 );
nand U139455 ( n69963, n69935, n390 );
nand U139456 ( n69805, n69806, n69807 );
nand U139457 ( n69806, P2_P3_INSTQUEUE_REG_9__3_, n69780 );
nand U139458 ( n69807, n69779, n390 );
nand U139459 ( n69574, n69575, n69576 );
nand U139460 ( n69575, P2_P3_INSTQUEUE_REG_6__3_, n69549 );
nand U139461 ( n69576, n69548, n390 );
nand U139462 ( n69492, n69493, n69494 );
nand U139463 ( n69493, P2_P3_INSTQUEUE_REG_5__3_, n69464 );
nand U139464 ( n69494, n69463, n390 );
nand U139465 ( n70139, n70140, n70141 );
nand U139466 ( n70140, P2_P3_INSTQUEUE_REG_13__6_, n70090 );
nand U139467 ( n70141, n70089, n398 );
nand U139468 ( n69985, n69986, n69987 );
nand U139469 ( n69986, P2_P3_INSTQUEUE_REG_11__6_, n69936 );
nand U139470 ( n69987, n69935, n398 );
nand U139471 ( n69829, n69830, n69831 );
nand U139472 ( n69830, P2_P3_INSTQUEUE_REG_9__6_, n69780 );
nand U139473 ( n69831, n69779, n398 );
nand U139474 ( n69598, n69599, n69600 );
nand U139475 ( n69599, P2_P3_INSTQUEUE_REG_6__6_, n69549 );
nand U139476 ( n69600, n69548, n398 );
nand U139477 ( n69519, n69520, n69521 );
nand U139478 ( n69520, P2_P3_INSTQUEUE_REG_5__6_, n69464 );
nand U139479 ( n69521, n69463, n398 );
nand U139480 ( n70147, n70148, n70149 );
nand U139481 ( n70148, P2_P3_INSTQUEUE_REG_13__7_, n70090 );
nand U139482 ( n70149, n70089, n400 );
nand U139483 ( n69993, n69994, n69995 );
nand U139484 ( n69994, P2_P3_INSTQUEUE_REG_11__7_, n69936 );
nand U139485 ( n69995, n69935, n400 );
nand U139486 ( n69837, n69838, n69839 );
nand U139487 ( n69838, P2_P3_INSTQUEUE_REG_9__7_, n69780 );
nand U139488 ( n69839, n69779, n400 );
nand U139489 ( n69606, n69607, n69608 );
nand U139490 ( n69607, P2_P3_INSTQUEUE_REG_6__7_, n69549 );
nand U139491 ( n69608, n69548, n400 );
nand U139492 ( n69528, n69529, n69530 );
nand U139493 ( n69529, P2_P3_INSTQUEUE_REG_5__7_, n69464 );
nand U139494 ( n69530, n69463, n400 );
nand U139495 ( n70131, n70132, n70133 );
nand U139496 ( n70132, P2_P3_INSTQUEUE_REG_13__5_, n70090 );
nand U139497 ( n70133, n70089, n395 );
nand U139498 ( n69977, n69978, n69979 );
nand U139499 ( n69978, P2_P3_INSTQUEUE_REG_11__5_, n69936 );
nand U139500 ( n69979, n69935, n395 );
nand U139501 ( n69821, n69822, n69823 );
nand U139502 ( n69822, P2_P3_INSTQUEUE_REG_9__5_, n69780 );
nand U139503 ( n69823, n69779, n395 );
nand U139504 ( n69590, n69591, n69592 );
nand U139505 ( n69591, P2_P3_INSTQUEUE_REG_6__5_, n69549 );
nand U139506 ( n69592, n69548, n395 );
nand U139507 ( n69510, n69511, n69512 );
nand U139508 ( n69511, P2_P3_INSTQUEUE_REG_5__5_, n69464 );
nand U139509 ( n69512, n69463, n395 );
nand U139510 ( n70123, n70124, n70125 );
nand U139511 ( n70124, P2_P3_INSTQUEUE_REG_13__4_, n70090 );
nand U139512 ( n70125, n70089, n393 );
nand U139513 ( n69969, n69970, n69971 );
nand U139514 ( n69970, P2_P3_INSTQUEUE_REG_11__4_, n69936 );
nand U139515 ( n69971, n69935, n393 );
nand U139516 ( n69813, n69814, n69815 );
nand U139517 ( n69814, P2_P3_INSTQUEUE_REG_9__4_, n69780 );
nand U139518 ( n69815, n69779, n393 );
nand U139519 ( n69582, n69583, n69584 );
nand U139520 ( n69583, P2_P3_INSTQUEUE_REG_6__4_, n69549 );
nand U139521 ( n69584, n69548, n393 );
nand U139522 ( n69501, n69502, n69503 );
nand U139523 ( n69502, P2_P3_INSTQUEUE_REG_5__4_, n69464 );
nand U139524 ( n69503, n69463, n393 );
nand U139525 ( n70008, n70009, n70010 );
nand U139526 ( n70009, P2_P3_INSTQUEUE_REG_12__0_, n70012 );
nand U139527 ( n70010, n70011, n383 );
nand U139528 ( n69697, n69698, n69699 );
nand U139529 ( n69698, P2_P3_INSTQUEUE_REG_8__0_, n69701 );
nand U139530 ( n69699, n69700, n383 );
nand U139531 ( n28102, n28103, n28104 );
nand U139532 ( n28104, n28040, n27542 );
nand U139533 ( n28103, P1_P2_INSTQUEUE_REG_12__7_, n28041 );
nand U139534 ( n27779, n27780, n27781 );
nand U139535 ( n27781, n27715, n27542 );
nand U139536 ( n27780, P1_P2_INSTQUEUE_REG_8__7_, n27716 );
nand U139537 ( n28086, n28087, n28088 );
nand U139538 ( n28088, n28040, n27524 );
nand U139539 ( n28087, P1_P2_INSTQUEUE_REG_12__5_, n28041 );
nand U139540 ( n27763, n27764, n27765 );
nand U139541 ( n27765, n27715, n27524 );
nand U139542 ( n27764, P1_P2_INSTQUEUE_REG_8__5_, n27716 );
nand U139543 ( n61241, n61242, n61243 );
nand U139544 ( n61243, n61199, n60676 );
nand U139545 ( n61242, P2_P2_INSTQUEUE_REG_12__5_, n61200 );
nand U139546 ( n60911, n60912, n60913 );
nand U139547 ( n60913, n60866, n60676 );
nand U139548 ( n60912, P2_P2_INSTQUEUE_REG_8__5_, n60867 );
nand U139549 ( n61257, n61258, n61259 );
nand U139550 ( n61259, n61199, n60694 );
nand U139551 ( n61258, P2_P2_INSTQUEUE_REG_12__7_, n61200 );
nand U139552 ( n28050, n28051, n28052 );
nand U139553 ( n28052, n28040, n27488 );
nand U139554 ( n28051, P1_P2_INSTQUEUE_REG_12__1_, n28041 );
nand U139555 ( n27725, n27726, n27727 );
nand U139556 ( n27727, n27715, n27488 );
nand U139557 ( n27726, P1_P2_INSTQUEUE_REG_8__1_, n27716 );
nand U139558 ( n27741, n27742, n27743 );
nand U139559 ( n27743, n27715, n27506 );
nand U139560 ( n27742, P1_P2_INSTQUEUE_REG_8__3_, n27716 );
nand U139561 ( n28078, n28079, n28080 );
nand U139562 ( n28080, n28040, n27515 );
nand U139563 ( n28079, P1_P2_INSTQUEUE_REG_12__4_, n28041 );
nand U139564 ( n27755, n27756, n27757 );
nand U139565 ( n27757, n27715, n27515 );
nand U139566 ( n27756, P1_P2_INSTQUEUE_REG_8__4_, n27716 );
nand U139567 ( n28062, n28063, n28064 );
nand U139568 ( n28064, n28040, n27497 );
nand U139569 ( n28063, P1_P2_INSTQUEUE_REG_12__2_, n28041 );
nand U139570 ( n27733, n27734, n27735 );
nand U139571 ( n27735, n27715, n27497 );
nand U139572 ( n27734, P1_P2_INSTQUEUE_REG_8__2_, n27716 );
nand U139573 ( n61225, n61226, n61227 );
nand U139574 ( n61227, n61199, n60655 );
nand U139575 ( n61226, P2_P2_INSTQUEUE_REG_12__3_, n61200 );
nand U139576 ( n60927, n60928, n60929 );
nand U139577 ( n60929, n60866, n60694 );
nand U139578 ( n60928, P2_P2_INSTQUEUE_REG_8__7_, n60867 );
nand U139579 ( n28070, n28071, n28072 );
nand U139580 ( n28072, n28040, n27506 );
nand U139581 ( n28071, P1_P2_INSTQUEUE_REG_12__3_, n28041 );
nand U139582 ( n60895, n60896, n60897 );
nand U139583 ( n60897, n60866, n60655 );
nand U139584 ( n60896, P2_P2_INSTQUEUE_REG_8__3_, n60867 );
nand U139585 ( n61209, n61210, n61211 );
nand U139586 ( n61211, n61199, n60637 );
nand U139587 ( n61210, P2_P2_INSTQUEUE_REG_12__1_, n61200 );
nand U139588 ( n60879, n60880, n60881 );
nand U139589 ( n60881, n60866, n60637 );
nand U139590 ( n60880, P2_P2_INSTQUEUE_REG_8__1_, n60867 );
nand U139591 ( n61217, n61218, n61219 );
nand U139592 ( n61219, n61199, n60646 );
nand U139593 ( n61218, P2_P2_INSTQUEUE_REG_12__2_, n61200 );
nand U139594 ( n60887, n60888, n60889 );
nand U139595 ( n60889, n60866, n60646 );
nand U139596 ( n60888, P2_P2_INSTQUEUE_REG_8__2_, n60867 );
nand U139597 ( n61233, n61234, n61235 );
nand U139598 ( n61235, n61199, n60664 );
nand U139599 ( n61234, P2_P2_INSTQUEUE_REG_12__4_, n61200 );
nand U139600 ( n60903, n60904, n60905 );
nand U139601 ( n60905, n60866, n60664 );
nand U139602 ( n60904, P2_P2_INSTQUEUE_REG_8__4_, n60867 );
nand U139603 ( n28094, n28095, n28096 );
nand U139604 ( n28096, n28040, n27533 );
nand U139605 ( n28095, P1_P2_INSTQUEUE_REG_12__6_, n28041 );
nand U139606 ( n27771, n27772, n27773 );
nand U139607 ( n27773, n27715, n27533 );
nand U139608 ( n27772, P1_P2_INSTQUEUE_REG_8__6_, n27716 );
nand U139609 ( n28037, n28038, n28039 );
nand U139610 ( n28039, n28040, n27475 );
nand U139611 ( n28038, P1_P2_INSTQUEUE_REG_12__0_, n28041 );
nand U139612 ( n61249, n61250, n61251 );
nand U139613 ( n61251, n61199, n60685 );
nand U139614 ( n61250, P2_P2_INSTQUEUE_REG_12__6_, n61200 );
nand U139615 ( n27712, n27713, n27714 );
nand U139616 ( n27714, n27715, n27475 );
nand U139617 ( n27713, P1_P2_INSTQUEUE_REG_8__0_, n27716 );
nand U139618 ( n60919, n60920, n60921 );
nand U139619 ( n60921, n60866, n60685 );
nand U139620 ( n60920, P2_P2_INSTQUEUE_REG_8__6_, n60867 );
nand U139621 ( n61196, n61197, n61198 );
nand U139622 ( n61198, n61199, n60624 );
nand U139623 ( n61197, P2_P2_INSTQUEUE_REG_12__0_, n61200 );
nand U139624 ( n60863, n60864, n60865 );
nand U139625 ( n60865, n60866, n60624 );
nand U139626 ( n60864, P2_P2_INSTQUEUE_REG_8__0_, n60867 );
nand U139627 ( n13685, n13687, n74476 );
nand U139628 ( n13687, n4860, n13688 );
nand U139629 ( n13688, P1_P1_INSTADDRPOINTER_REG_11_, n13689 );
xor U139630 ( n42958, n42959, n42960 );
xor U139631 ( n42960, n42957, P3_REG1_REG_8_ );
nand U139632 ( n60993, n60994, n60995 );
nand U139633 ( n60995, n60948, n60676 );
nand U139634 ( n60994, P2_P2_INSTQUEUE_REG_9__5_, n60949 );
nand U139635 ( n61009, n61010, n61011 );
nand U139636 ( n61011, n60948, n60694 );
nand U139637 ( n61010, P2_P2_INSTQUEUE_REG_9__7_, n60949 );
nand U139638 ( n34646, n34647, n34648 );
nand U139639 ( n34648, P1_P3_INSTQUEUE_REG_4__1_, n34636 );
nand U139640 ( n34647, n34637, n133 );
nand U139641 ( n34686, n34687, n34688 );
nand U139642 ( n34688, P1_P3_INSTQUEUE_REG_4__6_, n34636 );
nand U139643 ( n34687, n34637, n145 );
nand U139644 ( n34654, n34655, n34656 );
nand U139645 ( n34656, P1_P3_INSTQUEUE_REG_4__2_, n34636 );
nand U139646 ( n34655, n34637, n135 );
nand U139647 ( n69392, n69393, n69394 );
nand U139648 ( n69394, P2_P3_INSTQUEUE_REG_4__1_, n69382 );
nand U139649 ( n69393, n69383, n405 );
nand U139650 ( n69400, n69401, n69402 );
nand U139651 ( n69402, P2_P3_INSTQUEUE_REG_4__2_, n69382 );
nand U139652 ( n69401, n69383, n408 );
nand U139653 ( n27862, n27863, n27864 );
nand U139654 ( n27864, n27800, n27542 );
nand U139655 ( n27863, P1_P2_INSTQUEUE_REG_9__7_, n27801 );
nand U139656 ( n27842, n27843, n27844 );
nand U139657 ( n27844, n27800, n27524 );
nand U139658 ( n27843, P1_P2_INSTQUEUE_REG_9__5_, n27801 );
nand U139659 ( n69408, n69409, n69410 );
nand U139660 ( n69410, P2_P3_INSTQUEUE_REG_4__3_, n69382 );
nand U139661 ( n69409, n69383, n410 );
nand U139662 ( n69432, n69433, n69434 );
nand U139663 ( n69434, P2_P3_INSTQUEUE_REG_4__6_, n69382 );
nand U139664 ( n69433, n69383, n418 );
nand U139665 ( n69440, n69441, n69442 );
nand U139666 ( n69442, P2_P3_INSTQUEUE_REG_4__7_, n69382 );
nand U139667 ( n69441, n69383, n419 );
nand U139668 ( n69424, n69425, n69426 );
nand U139669 ( n69426, P2_P3_INSTQUEUE_REG_4__5_, n69382 );
nand U139670 ( n69425, n69383, n415 );
nand U139671 ( n61155, n61156, n61157 );
nand U139672 ( n61157, n61113, n60676 );
nand U139673 ( n61156, P2_P2_INSTQUEUE_REG_11__5_, n61114 );
nand U139674 ( n61001, n61002, n61003 );
nand U139675 ( n61003, n60948, n60685 );
nand U139676 ( n61002, P2_P2_INSTQUEUE_REG_9__6_, n60949 );
nand U139677 ( n60945, n60946, n60947 );
nand U139678 ( n60947, n60948, n60624 );
nand U139679 ( n60946, P2_P2_INSTQUEUE_REG_9__0_, n60949 );
nand U139680 ( n61181, n61182, n61183 );
nand U139681 ( n61183, n61113, n60694 );
nand U139682 ( n61182, P2_P2_INSTQUEUE_REG_11__7_, n61114 );
nand U139683 ( n34678, n34679, n34680 );
nand U139684 ( n34680, P1_P3_INSTQUEUE_REG_4__5_, n34636 );
nand U139685 ( n34679, n34637, n143 );
nand U139686 ( n34662, n34663, n34664 );
nand U139687 ( n34664, P1_P3_INSTQUEUE_REG_4__3_, n34636 );
nand U139688 ( n34663, n34637, n138 );
nand U139689 ( n34670, n34671, n34672 );
nand U139690 ( n34672, P1_P3_INSTQUEUE_REG_4__4_, n34636 );
nand U139691 ( n34671, n34637, n140 );
nand U139692 ( n69416, n69417, n69418 );
nand U139693 ( n69418, P2_P3_INSTQUEUE_REG_4__4_, n69382 );
nand U139694 ( n69417, n69383, n413 );
nand U139695 ( n27854, n27855, n27856 );
nand U139696 ( n27856, n27800, n27533 );
nand U139697 ( n27855, P1_P2_INSTQUEUE_REG_9__6_, n27801 );
nand U139698 ( n27797, n27798, n27799 );
nand U139699 ( n27799, n27800, n27475 );
nand U139700 ( n27798, P1_P2_INSTQUEUE_REG_9__0_, n27801 );
nand U139701 ( n28006, n28007, n28008 );
nand U139702 ( n28008, n27964, n27524 );
nand U139703 ( n28007, P1_P2_INSTQUEUE_REG_11__5_, n27965 );
nand U139704 ( n34696, n34697, n34698 );
nand U139705 ( n34698, P1_P3_INSTQUEUE_REG_4__7_, n34636 );
nand U139706 ( n34697, n34637, n147 );
nand U139707 ( n28022, n28023, n28024 );
nand U139708 ( n28024, n27964, n27542 );
nand U139709 ( n28023, P1_P2_INSTQUEUE_REG_11__7_, n27965 );
nand U139710 ( n27810, n27811, n27812 );
nand U139711 ( n27812, n27800, n27488 );
nand U139712 ( n27811, P1_P2_INSTQUEUE_REG_9__1_, n27801 );
nand U139713 ( n28014, n28015, n28016 );
nand U139714 ( n28016, n27964, n27533 );
nand U139715 ( n28015, P1_P2_INSTQUEUE_REG_11__6_, n27965 );
nand U139716 ( n27961, n27962, n27963 );
nand U139717 ( n27963, n27964, n27475 );
nand U139718 ( n27962, P1_P2_INSTQUEUE_REG_11__0_, n27965 );
nand U139719 ( n28184, n28185, n28186 );
nand U139720 ( n28186, n28122, n27542 );
nand U139721 ( n28185, P1_P2_INSTQUEUE_REG_13__7_, n28123 );
nand U139722 ( n28168, n28169, n28170 );
nand U139723 ( n28170, n28122, n27524 );
nand U139724 ( n28169, P1_P2_INSTQUEUE_REG_13__5_, n28123 );
nand U139725 ( n27826, n27827, n27828 );
nand U139726 ( n27828, n27800, n27506 );
nand U139727 ( n27827, P1_P2_INSTQUEUE_REG_9__3_, n27801 );
nand U139728 ( n27834, n27835, n27836 );
nand U139729 ( n27836, n27800, n27515 );
nand U139730 ( n27835, P1_P2_INSTQUEUE_REG_9__4_, n27801 );
nand U139731 ( n27818, n27819, n27820 );
nand U139732 ( n27820, n27800, n27497 );
nand U139733 ( n27819, P1_P2_INSTQUEUE_REG_9__2_, n27801 );
nand U139734 ( n60977, n60978, n60979 );
nand U139735 ( n60979, n60948, n60655 );
nand U139736 ( n60978, P2_P2_INSTQUEUE_REG_9__3_, n60949 );
nand U139737 ( n61163, n61164, n61165 );
nand U139738 ( n61165, n61113, n60685 );
nand U139739 ( n61164, P2_P2_INSTQUEUE_REG_11__6_, n61114 );
nand U139740 ( n60958, n60959, n60960 );
nand U139741 ( n60960, n60948, n60637 );
nand U139742 ( n60959, P2_P2_INSTQUEUE_REG_9__1_, n60949 );
nand U139743 ( n61110, n61111, n61112 );
nand U139744 ( n61112, n61113, n60624 );
nand U139745 ( n61111, P2_P2_INSTQUEUE_REG_11__0_, n61114 );
nand U139746 ( n60966, n60967, n60968 );
nand U139747 ( n60968, n60948, n60646 );
nand U139748 ( n60967, P2_P2_INSTQUEUE_REG_9__2_, n60949 );
nand U139749 ( n60985, n60986, n60987 );
nand U139750 ( n60987, n60948, n60664 );
nand U139751 ( n60986, P2_P2_INSTQUEUE_REG_9__4_, n60949 );
nand U139752 ( n27974, n27975, n27976 );
nand U139753 ( n27976, n27964, n27488 );
nand U139754 ( n27975, P1_P2_INSTQUEUE_REG_11__1_, n27965 );
nand U139755 ( n28176, n28177, n28178 );
nand U139756 ( n28178, n28122, n27533 );
nand U139757 ( n28177, P1_P2_INSTQUEUE_REG_13__6_, n28123 );
nand U139758 ( n28119, n28120, n28121 );
nand U139759 ( n28121, n28122, n27475 );
nand U139760 ( n28120, P1_P2_INSTQUEUE_REG_13__0_, n28123 );
nand U139761 ( n27990, n27991, n27992 );
nand U139762 ( n27992, n27964, n27506 );
nand U139763 ( n27991, P1_P2_INSTQUEUE_REG_11__3_, n27965 );
nand U139764 ( n27998, n27999, n28000 );
nand U139765 ( n28000, n27964, n27515 );
nand U139766 ( n27999, P1_P2_INSTQUEUE_REG_11__4_, n27965 );
nand U139767 ( n27982, n27983, n27984 );
nand U139768 ( n27984, n27964, n27497 );
nand U139769 ( n27983, P1_P2_INSTQUEUE_REG_11__2_, n27965 );
nand U139770 ( n61332, n61333, n61334 );
nand U139771 ( n61334, n61277, n60676 );
nand U139772 ( n61333, P2_P2_INSTQUEUE_REG_13__5_, n61278 );
nand U139773 ( n61139, n61140, n61141 );
nand U139774 ( n61141, n61113, n60655 );
nand U139775 ( n61140, P2_P2_INSTQUEUE_REG_11__3_, n61114 );
nand U139776 ( n61340, n61341, n61342 );
nand U139777 ( n61342, n61277, n60685 );
nand U139778 ( n61341, P2_P2_INSTQUEUE_REG_13__6_, n61278 );
nand U139779 ( n61123, n61124, n61125 );
nand U139780 ( n61125, n61113, n60637 );
nand U139781 ( n61124, P2_P2_INSTQUEUE_REG_11__1_, n61114 );
nand U139782 ( n61131, n61132, n61133 );
nand U139783 ( n61133, n61113, n60646 );
nand U139784 ( n61132, P2_P2_INSTQUEUE_REG_11__2_, n61114 );
nand U139785 ( n61147, n61148, n61149 );
nand U139786 ( n61149, n61113, n60664 );
nand U139787 ( n61148, P2_P2_INSTQUEUE_REG_11__4_, n61114 );
nand U139788 ( n61348, n61349, n61350 );
nand U139789 ( n61350, n61277, n60694 );
nand U139790 ( n61349, P2_P2_INSTQUEUE_REG_13__7_, n61278 );
nand U139791 ( n34400, n34401, n34402 );
nand U139792 ( n34402, P1_P3_INSTQUEUE_REG_1__1_, n34388 );
nand U139793 ( n34401, n34389, n133 );
nand U139794 ( n34432, n34433, n34434 );
nand U139795 ( n34434, P1_P3_INSTQUEUE_REG_1__5_, n34388 );
nand U139796 ( n34433, n34389, n143 );
nand U139797 ( n34524, n34525, n34526 );
nand U139798 ( n34526, P1_P3_INSTQUEUE_REG_2__6_, n34472 );
nand U139799 ( n34525, n34473, n145 );
nand U139800 ( n34440, n34441, n34442 );
nand U139801 ( n34442, P1_P3_INSTQUEUE_REG_1__6_, n34388 );
nand U139802 ( n34441, n34389, n145 );
nand U139803 ( n69379, n69380, n69381 );
nand U139804 ( n69381, P2_P3_INSTQUEUE_REG_4__0_, n69382 );
nand U139805 ( n69380, n69383, n403 );
nand U139806 ( n61274, n61275, n61276 );
nand U139807 ( n61276, n61277, n60624 );
nand U139808 ( n61275, P2_P2_INSTQUEUE_REG_13__0_, n61278 );
nand U139809 ( n34482, n34483, n34484 );
nand U139810 ( n34484, P1_P3_INSTQUEUE_REG_2__1_, n34472 );
nand U139811 ( n34483, n34473, n133 );
nand U139812 ( n34516, n34517, n34518 );
nand U139813 ( n34518, P1_P3_INSTQUEUE_REG_2__5_, n34472 );
nand U139814 ( n34517, n34473, n143 );
nand U139815 ( n34614, n34615, n34616 );
nand U139816 ( n34616, P1_P3_INSTQUEUE_REG_3__7_, n34554 );
nand U139817 ( n34615, n34555, n147 );
nand U139818 ( n34448, n34449, n34450 );
nand U139819 ( n34450, P1_P3_INSTQUEUE_REG_1__7_, n34388 );
nand U139820 ( n34449, n34389, n147 );
nand U139821 ( n34500, n34501, n34502 );
nand U139822 ( n34502, P1_P3_INSTQUEUE_REG_2__3_, n34472 );
nand U139823 ( n34501, n34473, n138 );
nand U139824 ( n34416, n34417, n34418 );
nand U139825 ( n34418, P1_P3_INSTQUEUE_REG_1__3_, n34388 );
nand U139826 ( n34417, n34389, n138 );
nand U139827 ( n34588, n34589, n34590 );
nand U139828 ( n34590, P1_P3_INSTQUEUE_REG_3__4_, n34554 );
nand U139829 ( n34589, n34555, n140 );
nand U139830 ( n34508, n34509, n34510 );
nand U139831 ( n34510, P1_P3_INSTQUEUE_REG_2__4_, n34472 );
nand U139832 ( n34509, n34473, n140 );
nand U139833 ( n34424, n34425, n34426 );
nand U139834 ( n34426, P1_P3_INSTQUEUE_REG_1__4_, n34388 );
nand U139835 ( n34425, n34389, n140 );
nand U139836 ( n34469, n34470, n34471 );
nand U139837 ( n34471, P1_P3_INSTQUEUE_REG_2__0_, n34472 );
nand U139838 ( n34470, n34473, n130 );
nand U139839 ( n34385, n34386, n34387 );
nand U139840 ( n34387, P1_P3_INSTQUEUE_REG_1__0_, n34388 );
nand U139841 ( n34386, n34389, n130 );
nand U139842 ( n34490, n34491, n34492 );
nand U139843 ( n34492, P1_P3_INSTQUEUE_REG_2__2_, n34472 );
nand U139844 ( n34491, n34473, n135 );
nand U139845 ( n34408, n34409, n34410 );
nand U139846 ( n34410, P1_P3_INSTQUEUE_REG_1__2_, n34388 );
nand U139847 ( n34409, n34389, n135 );
nand U139848 ( n69312, n69313, n69314 );
nand U139849 ( n69314, P2_P3_INSTQUEUE_REG_3__1_, n69302 );
nand U139850 ( n69313, n69303, n405 );
nand U139851 ( n69232, n69233, n69234 );
nand U139852 ( n69234, P2_P3_INSTQUEUE_REG_2__1_, n69222 );
nand U139853 ( n69233, n69223, n405 );
nand U139854 ( n69150, n69151, n69152 );
nand U139855 ( n69152, P2_P3_INSTQUEUE_REG_1__1_, n69140 );
nand U139856 ( n69151, n69141, n405 );
nand U139857 ( n69320, n69321, n69322 );
nand U139858 ( n69322, P2_P3_INSTQUEUE_REG_3__2_, n69302 );
nand U139859 ( n69321, n69303, n408 );
nand U139860 ( n69240, n69241, n69242 );
nand U139861 ( n69242, P2_P3_INSTQUEUE_REG_2__2_, n69222 );
nand U139862 ( n69241, n69223, n408 );
nand U139863 ( n69158, n69159, n69160 );
nand U139864 ( n69160, P2_P3_INSTQUEUE_REG_1__2_, n69140 );
nand U139865 ( n69159, n69141, n408 );
nand U139866 ( n69328, n69329, n69330 );
nand U139867 ( n69330, P2_P3_INSTQUEUE_REG_3__3_, n69302 );
nand U139868 ( n69329, n69303, n410 );
nand U139869 ( n69248, n69249, n69250 );
nand U139870 ( n69250, P2_P3_INSTQUEUE_REG_2__3_, n69222 );
nand U139871 ( n69249, n69223, n410 );
nand U139872 ( n69166, n69167, n69168 );
nand U139873 ( n69168, P2_P3_INSTQUEUE_REG_1__3_, n69140 );
nand U139874 ( n69167, n69141, n410 );
nand U139875 ( n69352, n69353, n69354 );
nand U139876 ( n69354, P2_P3_INSTQUEUE_REG_3__6_, n69302 );
nand U139877 ( n69353, n69303, n418 );
nand U139878 ( n69272, n69273, n69274 );
nand U139879 ( n69274, P2_P3_INSTQUEUE_REG_2__6_, n69222 );
nand U139880 ( n69273, n69223, n418 );
nand U139881 ( n69190, n69191, n69192 );
nand U139882 ( n69192, P2_P3_INSTQUEUE_REG_1__6_, n69140 );
nand U139883 ( n69191, n69141, n418 );
nand U139884 ( n69344, n69345, n69346 );
nand U139885 ( n69346, P2_P3_INSTQUEUE_REG_3__5_, n69302 );
nand U139886 ( n69345, n69303, n415 );
nand U139887 ( n28132, n28133, n28134 );
nand U139888 ( n28134, n28122, n27488 );
nand U139889 ( n28133, P1_P2_INSTQUEUE_REG_13__1_, n28123 );
nand U139890 ( n28148, n28149, n28150 );
nand U139891 ( n28150, n28122, n27506 );
nand U139892 ( n28149, P1_P2_INSTQUEUE_REG_13__3_, n28123 );
nand U139893 ( n28160, n28161, n28162 );
nand U139894 ( n28162, n28122, n27515 );
nand U139895 ( n28161, P1_P2_INSTQUEUE_REG_13__4_, n28123 );
nand U139896 ( n28140, n28141, n28142 );
nand U139897 ( n28142, n28122, n27497 );
nand U139898 ( n28141, P1_P2_INSTQUEUE_REG_13__2_, n28123 );
nand U139899 ( n61316, n61317, n61318 );
nand U139900 ( n61318, n61277, n60655 );
nand U139901 ( n61317, P2_P2_INSTQUEUE_REG_13__3_, n61278 );
nand U139902 ( n61300, n61301, n61302 );
nand U139903 ( n61302, n61277, n60637 );
nand U139904 ( n61301, P2_P2_INSTQUEUE_REG_13__1_, n61278 );
nand U139905 ( n34580, n34581, n34582 );
nand U139906 ( n34582, P1_P3_INSTQUEUE_REG_3__3_, n34554 );
nand U139907 ( n34581, n34555, n138 );
nand U139908 ( n34633, n34634, n34635 );
nand U139909 ( n34635, P1_P3_INSTQUEUE_REG_4__0_, n34636 );
nand U139910 ( n34634, n34637, n130 );
nand U139911 ( n34572, n34573, n34574 );
nand U139912 ( n34574, P1_P3_INSTQUEUE_REG_3__2_, n34554 );
nand U139913 ( n34573, n34555, n135 );
nand U139914 ( n34532, n34533, n34534 );
nand U139915 ( n34534, P1_P3_INSTQUEUE_REG_2__7_, n34472 );
nand U139916 ( n34533, n34473, n147 );
nand U139917 ( n69360, n69361, n69362 );
nand U139918 ( n69362, P2_P3_INSTQUEUE_REG_3__7_, n69302 );
nand U139919 ( n69361, n69303, n419 );
nand U139920 ( n69280, n69281, n69282 );
nand U139921 ( n69282, P2_P3_INSTQUEUE_REG_2__7_, n69222 );
nand U139922 ( n69281, n69223, n419 );
nand U139923 ( n69198, n69199, n69200 );
nand U139924 ( n69200, P2_P3_INSTQUEUE_REG_1__7_, n69140 );
nand U139925 ( n69199, n69141, n419 );
nand U139926 ( n69264, n69265, n69266 );
nand U139927 ( n69266, P2_P3_INSTQUEUE_REG_2__5_, n69222 );
nand U139928 ( n69265, n69223, n415 );
nand U139929 ( n69182, n69183, n69184 );
nand U139930 ( n69184, P2_P3_INSTQUEUE_REG_1__5_, n69140 );
nand U139931 ( n69183, n69141, n415 );
nand U139932 ( n69336, n69337, n69338 );
nand U139933 ( n69338, P2_P3_INSTQUEUE_REG_3__4_, n69302 );
nand U139934 ( n69337, n69303, n413 );
nand U139935 ( n69256, n69257, n69258 );
nand U139936 ( n69258, P2_P3_INSTQUEUE_REG_2__4_, n69222 );
nand U139937 ( n69257, n69223, n413 );
nand U139938 ( n69174, n69175, n69176 );
nand U139939 ( n69176, P2_P3_INSTQUEUE_REG_1__4_, n69140 );
nand U139940 ( n69175, n69141, n413 );
nand U139941 ( n69299, n69300, n69301 );
nand U139942 ( n69301, P2_P3_INSTQUEUE_REG_3__0_, n69302 );
nand U139943 ( n69300, n69303, n403 );
nand U139944 ( n69219, n69220, n69221 );
nand U139945 ( n69221, P2_P3_INSTQUEUE_REG_2__0_, n69222 );
nand U139946 ( n69220, n69223, n403 );
nand U139947 ( n69137, n69138, n69139 );
nand U139948 ( n69139, P2_P3_INSTQUEUE_REG_1__0_, n69140 );
nand U139949 ( n69138, n69141, n403 );
nand U139950 ( n61308, n61309, n61310 );
nand U139951 ( n61310, n61277, n60646 );
nand U139952 ( n61309, P2_P2_INSTQUEUE_REG_13__2_, n61278 );
nand U139953 ( n61324, n61325, n61326 );
nand U139954 ( n61326, n61277, n60664 );
nand U139955 ( n61325, P2_P2_INSTQUEUE_REG_13__4_, n61278 );
nand U139956 ( n34564, n34565, n34566 );
nand U139957 ( n34566, P1_P3_INSTQUEUE_REG_3__1_, n34554 );
nand U139958 ( n34565, n34555, n133 );
nand U139959 ( n34598, n34599, n34600 );
nand U139960 ( n34600, P1_P3_INSTQUEUE_REG_3__5_, n34554 );
nand U139961 ( n34599, n34555, n143 );
nand U139962 ( n34606, n34607, n34608 );
nand U139963 ( n34608, P1_P3_INSTQUEUE_REG_3__6_, n34554 );
nand U139964 ( n34607, n34555, n145 );
nand U139965 ( n34551, n34552, n34553 );
nand U139966 ( n34553, P1_P3_INSTQUEUE_REG_3__0_, n34554 );
nand U139967 ( n34552, n34555, n130 );
and U139968 ( n16161, P2_P1_DATAO_REG_31_, n76679 );
nand U139969 ( n34359, n34360, n34361 );
nand U139970 ( n34361, P1_P3_INSTQUEUE_REG_0__7_, n34280 );
nand U139971 ( n34360, n147, n34281 );
nand U139972 ( n34326, n34327, n34328 );
nand U139973 ( n34328, P1_P3_INSTQUEUE_REG_0__4_, n34280 );
nand U139974 ( n34327, n140, n34281 );
nand U139975 ( n69045, n69046, n69047 );
nand U139976 ( n69047, P2_P3_INSTQUEUE_REG_0__1_, n69032 );
nand U139977 ( n69046, n405, n69033 );
nand U139978 ( n69056, n69057, n69058 );
nand U139979 ( n69058, P2_P3_INSTQUEUE_REG_0__2_, n69032 );
nand U139980 ( n69057, n408, n69033 );
nand U139981 ( n69067, n69068, n69069 );
nand U139982 ( n69069, P2_P3_INSTQUEUE_REG_0__3_, n69032 );
nand U139983 ( n69068, n410, n69033 );
nand U139984 ( n69100, n69101, n69102 );
nand U139985 ( n69102, P2_P3_INSTQUEUE_REG_0__6_, n69032 );
nand U139986 ( n69101, n418, n69033 );
nand U139987 ( n69111, n69112, n69113 );
nand U139988 ( n69113, P2_P3_INSTQUEUE_REG_0__7_, n69032 );
nand U139989 ( n69112, n419, n69033 );
nand U139990 ( n69089, n69090, n69091 );
nand U139991 ( n69091, P2_P3_INSTQUEUE_REG_0__5_, n69032 );
nand U139992 ( n69090, n415, n69033 );
nand U139993 ( n69078, n69079, n69080 );
nand U139994 ( n69080, P2_P3_INSTQUEUE_REG_0__4_, n69032 );
nand U139995 ( n69079, n413, n69033 );
nand U139996 ( n34293, n34294, n34295 );
nand U139997 ( n34295, P1_P3_INSTQUEUE_REG_0__1_, n34280 );
nand U139998 ( n34294, n133, n34281 );
nand U139999 ( n34337, n34338, n34339 );
nand U140000 ( n34339, P1_P3_INSTQUEUE_REG_0__5_, n34280 );
nand U140001 ( n34338, n143, n34281 );
nand U140002 ( n34348, n34349, n34350 );
nand U140003 ( n34350, P1_P3_INSTQUEUE_REG_0__6_, n34280 );
nand U140004 ( n34349, n145, n34281 );
nand U140005 ( n34315, n34316, n34317 );
nand U140006 ( n34317, P1_P3_INSTQUEUE_REG_0__3_, n34280 );
nand U140007 ( n34316, n138, n34281 );
nand U140008 ( n34304, n34305, n34306 );
nand U140009 ( n34306, P1_P3_INSTQUEUE_REG_0__2_, n34280 );
nand U140010 ( n34305, n135, n34281 );
nand U140011 ( n69029, n69030, n69031 );
nand U140012 ( n69031, P2_P3_INSTQUEUE_REG_0__0_, n69032 );
nand U140013 ( n69030, n403, n69033 );
nand U140014 ( n34277, n34278, n34279 );
nand U140015 ( n34279, P1_P3_INSTQUEUE_REG_0__0_, n34280 );
nand U140016 ( n34278, n130, n34281 );
nor U140017 ( n8494, n5449, n8495 );
nor U140018 ( n8495, n8497, n73384 );
not U140019 ( n5449, n8475 );
nor U140020 ( n8497, P1_P1_EBX_REG_27_, n8498 );
nand U140021 ( n60113, P2_P2_INSTQUEUEWR_ADDR_REG_3_, n61725 );
nand U140022 ( n61725, n6930, P2_P2_INSTQUEUEWR_ADDR_REG_2_ );
nand U140023 ( n26973, P1_P2_INSTQUEUEWR_ADDR_REG_3_, n28416 );
nand U140024 ( n28416, n4298, P1_P2_INSTQUEUEWR_ADDR_REG_2_ );
nand U140025 ( n34218, P1_P3_INSTQUEUEWR_ADDR_REG_3_, n35597 );
nand U140026 ( n35597, n3460, P1_P3_INSTQUEUEWR_ADDR_REG_2_ );
nand U140027 ( n68972, P2_P3_INSTQUEUEWR_ADDR_REG_3_, n70325 );
nand U140028 ( n70325, n6075, P2_P3_INSTQUEUEWR_ADDR_REG_2_ );
nand U140029 ( n66916, P2_P3_PHYADDRPOINTER_REG_13_, P2_P3_PHYADDRPOINTER_REG_12_ );
nand U140030 ( n32277, P1_P3_PHYADDRPOINTER_REG_13_, P1_P3_PHYADDRPOINTER_REG_12_ );
nand U140031 ( n25040, P1_P2_PHYADDRPOINTER_REG_13_, P1_P2_PHYADDRPOINTER_REG_12_ );
nand U140032 ( n58175, P2_P2_PHYADDRPOINTER_REG_13_, P2_P2_PHYADDRPOINTER_REG_12_ );
nor U140033 ( n48119, n48120, n48121 );
nor U140034 ( n48121, n48026, n48122 );
and U140035 ( n48120, n48024, P2_P1_INSTQUEUE_REG_0__7_ );
nand U140036 ( n15389, n14697, n21115 );
nand U140037 ( n21115, P1_P1_INSTQUEUEWR_ADDR_REG_1_, n74435 );
nor U140038 ( n48508, n48509, n48510 );
nor U140039 ( n48510, n48122, n48429 );
and U140040 ( n48509, n48426, P2_P1_INSTQUEUE_REG_4__7_ );
and U140041 ( n9426, n76748, P1_P1_DATAO_REG_31_ );
nand U140042 ( n27619, n27620, n27621 );
nand U140043 ( n27620, P1_P2_INSTQUEUE_REG_6__7_, n27562 );
nand U140044 ( n27621, n27561, n27542 );
nand U140045 ( n27539, n27540, n27541 );
nand U140046 ( n27540, P1_P2_INSTQUEUE_REG_5__7_, n27476 );
nand U140047 ( n27541, n27474, n27542 );
nand U140048 ( n27611, n27612, n27613 );
nand U140049 ( n27612, P1_P2_INSTQUEUE_REG_6__6_, n27562 );
nand U140050 ( n27613, n27561, n27533 );
nand U140051 ( n27530, n27531, n27532 );
nand U140052 ( n27531, P1_P2_INSTQUEUE_REG_5__6_, n27476 );
nand U140053 ( n27532, n27474, n27533 );
nand U140054 ( n27558, n27559, n27560 );
nand U140055 ( n27559, P1_P2_INSTQUEUE_REG_6__0_, n27562 );
nand U140056 ( n27560, n27561, n27475 );
nand U140057 ( n27471, n27472, n27473 );
nand U140058 ( n27472, P1_P2_INSTQUEUE_REG_5__0_, n27476 );
nand U140059 ( n27473, n27474, n27475 );
nand U140060 ( n27603, n27604, n27605 );
nand U140061 ( n27604, P1_P2_INSTQUEUE_REG_6__5_, n27562 );
nand U140062 ( n27605, n27561, n27524 );
nand U140063 ( n27521, n27522, n27523 );
nand U140064 ( n27522, P1_P2_INSTQUEUE_REG_5__5_, n27476 );
nand U140065 ( n27523, n27474, n27524 );
nand U140066 ( n60753, n60754, n60755 );
nand U140067 ( n60754, P2_P2_INSTQUEUE_REG_6__5_, n60712 );
nand U140068 ( n60755, n60711, n60676 );
nand U140069 ( n60673, n60674, n60675 );
nand U140070 ( n60674, P2_P2_INSTQUEUE_REG_5__5_, n60625 );
nand U140071 ( n60675, n60623, n60676 );
nand U140072 ( n60761, n60762, n60763 );
nand U140073 ( n60762, P2_P2_INSTQUEUE_REG_6__6_, n60712 );
nand U140074 ( n60763, n60711, n60685 );
nand U140075 ( n60682, n60683, n60684 );
nand U140076 ( n60683, P2_P2_INSTQUEUE_REG_5__6_, n60625 );
nand U140077 ( n60684, n60623, n60685 );
nand U140078 ( n60708, n60709, n60710 );
nand U140079 ( n60709, P2_P2_INSTQUEUE_REG_6__0_, n60712 );
nand U140080 ( n60710, n60711, n60624 );
nand U140081 ( n60620, n60621, n60622 );
nand U140082 ( n60621, P2_P2_INSTQUEUE_REG_5__0_, n60625 );
nand U140083 ( n60622, n60623, n60624 );
nand U140084 ( n60772, n60773, n60774 );
nand U140085 ( n60773, P2_P2_INSTQUEUE_REG_6__7_, n60712 );
nand U140086 ( n60774, n60711, n60694 );
nand U140087 ( n60691, n60692, n60693 );
nand U140088 ( n60692, P2_P2_INSTQUEUE_REG_5__7_, n60625 );
nand U140089 ( n60693, n60623, n60694 );
nand U140090 ( n27571, n27572, n27573 );
nand U140091 ( n27572, P1_P2_INSTQUEUE_REG_6__1_, n27562 );
nand U140092 ( n27573, n27561, n27488 );
nand U140093 ( n27485, n27486, n27487 );
nand U140094 ( n27486, P1_P2_INSTQUEUE_REG_5__1_, n27476 );
nand U140095 ( n27487, n27474, n27488 );
nand U140096 ( n27587, n27588, n27589 );
nand U140097 ( n27588, P1_P2_INSTQUEUE_REG_6__3_, n27562 );
nand U140098 ( n27589, n27561, n27506 );
nand U140099 ( n27503, n27504, n27505 );
nand U140100 ( n27504, P1_P2_INSTQUEUE_REG_5__3_, n27476 );
nand U140101 ( n27505, n27474, n27506 );
nand U140102 ( n27595, n27596, n27597 );
nand U140103 ( n27596, P1_P2_INSTQUEUE_REG_6__4_, n27562 );
nand U140104 ( n27597, n27561, n27515 );
nand U140105 ( n27512, n27513, n27514 );
nand U140106 ( n27513, P1_P2_INSTQUEUE_REG_5__4_, n27476 );
nand U140107 ( n27514, n27474, n27515 );
nand U140108 ( n27579, n27580, n27581 );
nand U140109 ( n27580, P1_P2_INSTQUEUE_REG_6__2_, n27562 );
nand U140110 ( n27581, n27561, n27497 );
nand U140111 ( n27494, n27495, n27496 );
nand U140112 ( n27495, P1_P2_INSTQUEUE_REG_5__2_, n27476 );
nand U140113 ( n27496, n27474, n27497 );
nand U140114 ( n60737, n60738, n60739 );
nand U140115 ( n60738, P2_P2_INSTQUEUE_REG_6__3_, n60712 );
nand U140116 ( n60739, n60711, n60655 );
nand U140117 ( n60652, n60653, n60654 );
nand U140118 ( n60653, P2_P2_INSTQUEUE_REG_5__3_, n60625 );
nand U140119 ( n60654, n60623, n60655 );
nand U140120 ( n60721, n60722, n60723 );
nand U140121 ( n60722, P2_P2_INSTQUEUE_REG_6__1_, n60712 );
nand U140122 ( n60723, n60711, n60637 );
nand U140123 ( n60634, n60635, n60636 );
nand U140124 ( n60635, P2_P2_INSTQUEUE_REG_5__1_, n60625 );
nand U140125 ( n60636, n60623, n60637 );
nand U140126 ( n60729, n60730, n60731 );
nand U140127 ( n60730, P2_P2_INSTQUEUE_REG_6__2_, n60712 );
nand U140128 ( n60731, n60711, n60646 );
nand U140129 ( n60643, n60644, n60645 );
nand U140130 ( n60644, P2_P2_INSTQUEUE_REG_5__2_, n60625 );
nand U140131 ( n60645, n60623, n60646 );
nand U140132 ( n60745, n60746, n60747 );
nand U140133 ( n60746, P2_P2_INSTQUEUE_REG_6__4_, n60712 );
nand U140134 ( n60747, n60711, n60664 );
nand U140135 ( n60661, n60662, n60663 );
nand U140136 ( n60662, P2_P2_INSTQUEUE_REG_5__4_, n60625 );
nand U140137 ( n60663, n60623, n60664 );
nor U140138 ( n29145, n34139, P1_P3_STATE2_REG_1_ );
nor U140139 ( n21830, n26894, P1_P2_STATE2_REG_1_ );
nor U140140 ( n62812, n68893, P2_P3_STATE2_REG_1_ );
nor U140141 ( n54906, n60034, P2_P2_STATE2_REG_1_ );
and U140142 ( n68602, n68605, P2_P3_INSTADDRPOINTER_REG_3_ );
and U140143 ( n33846, n33849, P1_P3_INSTADDRPOINTER_REG_3_ );
and U140144 ( n47581, n47584, P2_P1_INSTADDRPOINTER_REG_3_ );
and U140145 ( n26601, n26604, P1_P2_INSTADDRPOINTER_REG_3_ );
and U140146 ( n59743, n59746, P2_P2_INSTADDRPOINTER_REG_3_ );
nor U140147 ( n42565, n42550, n42566 );
nor U140148 ( n42566, n42567, n73385 );
nor U140149 ( n42567, P2_P1_EBX_REG_27_, n42568 );
nor U140150 ( n22024, n22009, n22025 );
nor U140151 ( n22025, n22026, n73386 );
nor U140152 ( n22026, P1_P2_EBX_REG_27_, n22027 );
nor U140153 ( n29343, n29328, n29344 );
nor U140154 ( n29344, n29345, n73387 );
nor U140155 ( n29345, P1_P3_EBX_REG_27_, n29346 );
nor U140156 ( n63106, n63091, n63107 );
nor U140157 ( n63107, n63108, n73388 );
nor U140158 ( n63108, P2_P3_EBX_REG_27_, n63109 );
nor U140159 ( n55134, n55119, n55135 );
nor U140160 ( n55135, n55136, n73389 );
nor U140161 ( n55136, P2_P2_EBX_REG_27_, n55137 );
nor U140162 ( n50341, n76927, n8243 );
not U140163 ( n8243, DIN_29_ );
and U140164 ( n49633, n50341, P3_DATAO_REG_0_ );
nor U140165 ( n31104, n75347, n30480 );
nor U140166 ( n30479, n75330, n30480 );
nor U140167 ( n30524, n75331, n30480 );
nor U140168 ( n30614, n75332, n30480 );
nor U140169 ( n30659, n75333, n30480 );
nor U140170 ( n30703, n75334, n30480 );
nor U140171 ( n30748, n75335, n30480 );
nor U140172 ( n30849, n75348, n30480 );
nor U140173 ( n30892, n75349, n30480 );
nor U140174 ( n30934, n75350, n30480 );
nor U140175 ( n30977, n75351, n30480 );
nor U140176 ( n64638, n75336, n64639 );
nor U140177 ( n64683, n75337, n64639 );
nor U140178 ( n64773, n75338, n64639 );
nor U140179 ( n64865, n75339, n64639 );
nor U140180 ( n64909, n75340, n64639 );
nor U140181 ( n64954, n75341, n64639 );
nor U140182 ( n65051, n75354, n64639 );
nor U140183 ( n65094, n75355, n64639 );
nor U140184 ( n65136, n75356, n64639 );
nor U140185 ( n65179, n75357, n64639 );
nor U140186 ( n65221, n75358, n64639 );
nor U140187 ( n65264, n75359, n64639 );
nor U140188 ( n31019, n75352, n30480 );
nor U140189 ( n31062, n75353, n30480 );
nor U140190 ( n65306, n75360, n64639 );
nand U140191 ( n27451, n27452, n27453 );
nand U140192 ( n27453, P1_P2_INSTQUEUE_REG_4__7_, n27391 );
nand U140193 ( n27452, n27392, n27125 );
nand U140194 ( n27114, n27115, n27116 );
nand U140195 ( n27116, P1_P2_INSTQUEUE_REG_0__7_, n27035 );
nand U140196 ( n27115, n27036, n27125 );
nand U140197 ( n27369, n27370, n27371 );
nand U140198 ( n27371, P1_P2_INSTQUEUE_REG_3__7_, n27309 );
nand U140199 ( n27370, n27310, n27125 );
nand U140200 ( n27287, n27288, n27289 );
nand U140201 ( n27289, P1_P2_INSTQUEUE_REG_2__7_, n27227 );
nand U140202 ( n27288, n27228, n27125 );
nand U140203 ( n27203, n27204, n27205 );
nand U140204 ( n27205, P1_P2_INSTQUEUE_REG_1__7_, n27145 );
nand U140205 ( n27204, n27146, n27125 );
nor U140206 ( n27464, n74516, P1_P2_INSTQUEUEWR_ADDR_REG_3_ );
nor U140207 ( n60613, n74517, P2_P2_INSTQUEUEWR_ADDR_REG_3_ );
nor U140208 ( n34709, n74513, P1_P3_INSTQUEUEWR_ADDR_REG_3_ );
nor U140209 ( n69453, n74514, P2_P3_INSTQUEUEWR_ADDR_REG_3_ );
nand U140210 ( n27401, n27402, n27403 );
nand U140211 ( n27403, P1_P2_INSTQUEUE_REG_4__1_, n27391 );
nand U140212 ( n27402, n27392, n27051 );
nand U140213 ( n27433, n27434, n27435 );
nand U140214 ( n27435, P1_P2_INSTQUEUE_REG_4__5_, n27391 );
nand U140215 ( n27434, n27392, n27095 );
nand U140216 ( n27417, n27418, n27419 );
nand U140217 ( n27419, P1_P2_INSTQUEUE_REG_4__3_, n27391 );
nand U140218 ( n27418, n27392, n27073 );
nand U140219 ( n27425, n27426, n27427 );
nand U140220 ( n27427, P1_P2_INSTQUEUE_REG_4__4_, n27391 );
nand U140221 ( n27426, n27392, n27084 );
nand U140222 ( n27409, n27410, n27411 );
nand U140223 ( n27411, P1_P2_INSTQUEUE_REG_4__2_, n27391 );
nand U140224 ( n27410, n27392, n27062 );
nand U140225 ( n27048, n27049, n27050 );
nand U140226 ( n27050, P1_P2_INSTQUEUE_REG_0__1_, n27035 );
nand U140227 ( n27049, n27036, n27051 );
nand U140228 ( n27092, n27093, n27094 );
nand U140229 ( n27094, P1_P2_INSTQUEUE_REG_0__5_, n27035 );
nand U140230 ( n27093, n27036, n27095 );
nand U140231 ( n27070, n27071, n27072 );
nand U140232 ( n27072, P1_P2_INSTQUEUE_REG_0__3_, n27035 );
nand U140233 ( n27071, n27036, n27073 );
nand U140234 ( n27081, n27082, n27083 );
nand U140235 ( n27083, P1_P2_INSTQUEUE_REG_0__4_, n27035 );
nand U140236 ( n27082, n27036, n27084 );
nand U140237 ( n27059, n27060, n27061 );
nand U140238 ( n27061, P1_P2_INSTQUEUE_REG_0__2_, n27035 );
nand U140239 ( n27060, n27036, n27062 );
nand U140240 ( n60584, n60585, n60586 );
nand U140241 ( n60586, P2_P2_INSTQUEUE_REG_4__5_, n60539 );
nand U140242 ( n60585, n60540, n60239 );
nand U140243 ( n60568, n60569, n60570 );
nand U140244 ( n60570, P2_P2_INSTQUEUE_REG_4__3_, n60539 );
nand U140245 ( n60569, n60540, n60214 );
nand U140246 ( n60557, n60558, n60559 );
nand U140247 ( n60559, P2_P2_INSTQUEUE_REG_4__2_, n60539 );
nand U140248 ( n60558, n60540, n60203 );
nand U140249 ( n60576, n60577, n60578 );
nand U140250 ( n60578, P2_P2_INSTQUEUE_REG_4__4_, n60539 );
nand U140251 ( n60577, n60540, n60225 );
nand U140252 ( n60549, n60550, n60551 );
nand U140253 ( n60551, P2_P2_INSTQUEUE_REG_4__1_, n60539 );
nand U140254 ( n60550, n60540, n60192 );
nand U140255 ( n60600, n60601, n60602 );
nand U140256 ( n60602, P2_P2_INSTQUEUE_REG_4__7_, n60539 );
nand U140257 ( n60601, n60540, n60269 );
nand U140258 ( n16179, P1_P1_INSTQUEUE_REG_12__4_, n16129 );
nand U140259 ( n15763, P1_P1_INSTQUEUE_REG_8__4_, n15710 );
nand U140260 ( n16169, P1_P1_INSTQUEUE_REG_12__3_, n16129 );
nand U140261 ( n15753, P1_P1_INSTQUEUE_REG_8__3_, n15710 );
nand U140262 ( n16159, P1_P1_INSTQUEUE_REG_12__2_, n16129 );
nand U140263 ( n15734, P1_P1_INSTQUEUE_REG_8__2_, n15710 );
nand U140264 ( n16189, P1_P1_INSTQUEUE_REG_12__5_, n16129 );
nand U140265 ( n15783, P1_P1_INSTQUEUE_REG_8__6_, n15710 );
nand U140266 ( n16149, P1_P1_INSTQUEUE_REG_12__1_, n16129 );
nand U140267 ( n15724, P1_P1_INSTQUEUE_REG_8__1_, n15710 );
nand U140268 ( n16199, P1_P1_INSTQUEUE_REG_12__6_, n16129 );
nand U140269 ( n15773, P1_P1_INSTQUEUE_REG_8__5_, n15710 );
nand U140270 ( n16128, P1_P1_INSTQUEUE_REG_12__0_, n16129 );
nand U140271 ( n15709, P1_P1_INSTQUEUE_REG_8__0_, n15710 );
nand U140272 ( n60236, n60237, n60238 );
nand U140273 ( n60238, P2_P2_INSTQUEUE_REG_0__5_, n60176 );
nand U140274 ( n60237, n60177, n60239 );
nand U140275 ( n60211, n60212, n60213 );
nand U140276 ( n60213, P2_P2_INSTQUEUE_REG_0__3_, n60176 );
nand U140277 ( n60212, n60177, n60214 );
nand U140278 ( n60189, n60190, n60191 );
nand U140279 ( n60191, P2_P2_INSTQUEUE_REG_0__1_, n60176 );
nand U140280 ( n60190, n60177, n60192 );
nand U140281 ( n60200, n60201, n60202 );
nand U140282 ( n60202, P2_P2_INSTQUEUE_REG_0__2_, n60176 );
nand U140283 ( n60201, n60177, n60203 );
nand U140284 ( n60222, n60223, n60224 );
nand U140285 ( n60224, P2_P2_INSTQUEUE_REG_0__4_, n60176 );
nand U140286 ( n60223, n60177, n60225 );
nand U140287 ( n60258, n60259, n60260 );
nand U140288 ( n60260, P2_P2_INSTQUEUE_REG_0__7_, n60176 );
nand U140289 ( n60259, n60177, n60269 );
nand U140290 ( n27388, n27389, n27390 );
nand U140291 ( n27390, P1_P2_INSTQUEUE_REG_4__0_, n27391 );
nand U140292 ( n27389, n27392, n27037 );
nand U140293 ( n27443, n27444, n27445 );
nand U140294 ( n27445, P1_P2_INSTQUEUE_REG_4__6_, n27391 );
nand U140295 ( n27444, n27392, n27106 );
nand U140296 ( n27103, n27104, n27105 );
nand U140297 ( n27105, P1_P2_INSTQUEUE_REG_0__6_, n27035 );
nand U140298 ( n27104, n27036, n27106 );
nand U140299 ( n27032, n27033, n27034 );
nand U140300 ( n27034, P1_P2_INSTQUEUE_REG_0__0_, n27035 );
nand U140301 ( n27033, n27036, n27037 );
nand U140302 ( n27319, n27320, n27321 );
nand U140303 ( n27321, P1_P2_INSTQUEUE_REG_3__1_, n27309 );
nand U140304 ( n27320, n27310, n27051 );
nand U140305 ( n27237, n27238, n27239 );
nand U140306 ( n27239, P1_P2_INSTQUEUE_REG_2__1_, n27227 );
nand U140307 ( n27238, n27228, n27051 );
nand U140308 ( n27155, n27156, n27157 );
nand U140309 ( n27157, P1_P2_INSTQUEUE_REG_1__1_, n27145 );
nand U140310 ( n27156, n27146, n27051 );
nand U140311 ( n27361, n27362, n27363 );
nand U140312 ( n27363, P1_P2_INSTQUEUE_REG_3__6_, n27309 );
nand U140313 ( n27362, n27310, n27106 );
nand U140314 ( n27279, n27280, n27281 );
nand U140315 ( n27281, P1_P2_INSTQUEUE_REG_2__6_, n27227 );
nand U140316 ( n27280, n27228, n27106 );
nand U140317 ( n27195, n27196, n27197 );
nand U140318 ( n27197, P1_P2_INSTQUEUE_REG_1__6_, n27145 );
nand U140319 ( n27196, n27146, n27106 );
nand U140320 ( n27306, n27307, n27308 );
nand U140321 ( n27308, P1_P2_INSTQUEUE_REG_3__0_, n27309 );
nand U140322 ( n27307, n27310, n27037 );
nand U140323 ( n27224, n27225, n27226 );
nand U140324 ( n27226, P1_P2_INSTQUEUE_REG_2__0_, n27227 );
nand U140325 ( n27225, n27228, n27037 );
nand U140326 ( n27142, n27143, n27144 );
nand U140327 ( n27144, P1_P2_INSTQUEUE_REG_1__0_, n27145 );
nand U140328 ( n27143, n27146, n27037 );
nand U140329 ( n27353, n27354, n27355 );
nand U140330 ( n27355, P1_P2_INSTQUEUE_REG_3__5_, n27309 );
nand U140331 ( n27354, n27310, n27095 );
nand U140332 ( n27271, n27272, n27273 );
nand U140333 ( n27273, P1_P2_INSTQUEUE_REG_2__5_, n27227 );
nand U140334 ( n27272, n27228, n27095 );
nand U140335 ( n27187, n27188, n27189 );
nand U140336 ( n27189, P1_P2_INSTQUEUE_REG_1__5_, n27145 );
nand U140337 ( n27188, n27146, n27095 );
nand U140338 ( n27335, n27336, n27337 );
nand U140339 ( n27337, P1_P2_INSTQUEUE_REG_3__3_, n27309 );
nand U140340 ( n27336, n27310, n27073 );
nand U140341 ( n27171, n27172, n27173 );
nand U140342 ( n27173, P1_P2_INSTQUEUE_REG_1__3_, n27145 );
nand U140343 ( n27172, n27146, n27073 );
nand U140344 ( n27345, n27346, n27347 );
nand U140345 ( n27347, P1_P2_INSTQUEUE_REG_3__4_, n27309 );
nand U140346 ( n27346, n27310, n27084 );
nand U140347 ( n27263, n27264, n27265 );
nand U140348 ( n27265, P1_P2_INSTQUEUE_REG_2__4_, n27227 );
nand U140349 ( n27264, n27228, n27084 );
nand U140350 ( n27179, n27180, n27181 );
nand U140351 ( n27181, P1_P2_INSTQUEUE_REG_1__4_, n27145 );
nand U140352 ( n27180, n27146, n27084 );
nand U140353 ( n27327, n27328, n27329 );
nand U140354 ( n27329, P1_P2_INSTQUEUE_REG_3__2_, n27309 );
nand U140355 ( n27328, n27310, n27062 );
nand U140356 ( n27247, n27248, n27249 );
nand U140357 ( n27249, P1_P2_INSTQUEUE_REG_2__2_, n27227 );
nand U140358 ( n27248, n27228, n27062 );
nand U140359 ( n27163, n27164, n27165 );
nand U140360 ( n27165, P1_P2_INSTQUEUE_REG_1__2_, n27145 );
nand U140361 ( n27164, n27146, n27062 );
nand U140362 ( n60536, n60537, n60538 );
nand U140363 ( n60538, P2_P2_INSTQUEUE_REG_4__0_, n60539 );
nand U140364 ( n60537, n60540, n60178 );
nand U140365 ( n60592, n60593, n60594 );
nand U140366 ( n60594, P2_P2_INSTQUEUE_REG_4__6_, n60539 );
nand U140367 ( n60593, n60540, n60250 );
nand U140368 ( n60247, n60248, n60249 );
nand U140369 ( n60249, P2_P2_INSTQUEUE_REG_0__6_, n60176 );
nand U140370 ( n60248, n60177, n60250 );
nand U140371 ( n27255, n27256, n27257 );
nand U140372 ( n27257, P1_P2_INSTQUEUE_REG_2__3_, n27227 );
nand U140373 ( n27256, n27228, n27073 );
nand U140374 ( n60173, n60174, n60175 );
nand U140375 ( n60175, P2_P2_INSTQUEUE_REG_0__0_, n60176 );
nand U140376 ( n60174, n60177, n60178 );
nand U140377 ( n60501, n60502, n60503 );
nand U140378 ( n60503, P2_P2_INSTQUEUE_REG_3__5_, n60452 );
nand U140379 ( n60502, n60453, n60239 );
nand U140380 ( n60414, n60415, n60416 );
nand U140381 ( n60416, P2_P2_INSTQUEUE_REG_2__5_, n60372 );
nand U140382 ( n60415, n60373, n60239 );
nand U140383 ( n60329, n60330, n60331 );
nand U140384 ( n60331, P2_P2_INSTQUEUE_REG_1__5_, n60287 );
nand U140385 ( n60330, n60288, n60239 );
nand U140386 ( n60485, n60486, n60487 );
nand U140387 ( n60487, P2_P2_INSTQUEUE_REG_3__3_, n60452 );
nand U140388 ( n60486, n60453, n60214 );
nand U140389 ( n60398, n60399, n60400 );
nand U140390 ( n60400, P2_P2_INSTQUEUE_REG_2__3_, n60372 );
nand U140391 ( n60399, n60373, n60214 );
nand U140392 ( n60313, n60314, n60315 );
nand U140393 ( n60315, P2_P2_INSTQUEUE_REG_1__3_, n60287 );
nand U140394 ( n60314, n60288, n60214 );
nand U140395 ( n60509, n60510, n60511 );
nand U140396 ( n60511, P2_P2_INSTQUEUE_REG_3__6_, n60452 );
nand U140397 ( n60510, n60453, n60250 );
nand U140398 ( n60422, n60423, n60424 );
nand U140399 ( n60424, P2_P2_INSTQUEUE_REG_2__6_, n60372 );
nand U140400 ( n60423, n60373, n60250 );
nand U140401 ( n60337, n60338, n60339 );
nand U140402 ( n60339, P2_P2_INSTQUEUE_REG_1__6_, n60287 );
nand U140403 ( n60338, n60288, n60250 );
nand U140404 ( n60465, n60466, n60467 );
nand U140405 ( n60467, P2_P2_INSTQUEUE_REG_3__1_, n60452 );
nand U140406 ( n60466, n60453, n60192 );
nand U140407 ( n60382, n60383, n60384 );
nand U140408 ( n60384, P2_P2_INSTQUEUE_REG_2__1_, n60372 );
nand U140409 ( n60383, n60373, n60192 );
nand U140410 ( n60297, n60298, n60299 );
nand U140411 ( n60299, P2_P2_INSTQUEUE_REG_1__1_, n60287 );
nand U140412 ( n60298, n60288, n60192 );
nand U140413 ( n60449, n60450, n60451 );
nand U140414 ( n60451, P2_P2_INSTQUEUE_REG_3__0_, n60452 );
nand U140415 ( n60450, n60453, n60178 );
nand U140416 ( n60369, n60370, n60371 );
nand U140417 ( n60371, P2_P2_INSTQUEUE_REG_2__0_, n60372 );
nand U140418 ( n60370, n60373, n60178 );
nand U140419 ( n60284, n60285, n60286 );
nand U140420 ( n60286, P2_P2_INSTQUEUE_REG_1__0_, n60287 );
nand U140421 ( n60285, n60288, n60178 );
nand U140422 ( n60473, n60474, n60475 );
nand U140423 ( n60475, P2_P2_INSTQUEUE_REG_3__2_, n60452 );
nand U140424 ( n60474, n60453, n60203 );
nand U140425 ( n60390, n60391, n60392 );
nand U140426 ( n60392, P2_P2_INSTQUEUE_REG_2__2_, n60372 );
nand U140427 ( n60391, n60373, n60203 );
nand U140428 ( n60305, n60306, n60307 );
nand U140429 ( n60307, P2_P2_INSTQUEUE_REG_1__2_, n60287 );
nand U140430 ( n60306, n60288, n60203 );
nand U140431 ( n60493, n60494, n60495 );
nand U140432 ( n60495, P2_P2_INSTQUEUE_REG_3__4_, n60452 );
nand U140433 ( n60494, n60453, n60225 );
nand U140434 ( n60406, n60407, n60408 );
nand U140435 ( n60408, P2_P2_INSTQUEUE_REG_2__4_, n60372 );
nand U140436 ( n60407, n60373, n60225 );
nand U140437 ( n60321, n60322, n60323 );
nand U140438 ( n60323, P2_P2_INSTQUEUE_REG_1__4_, n60287 );
nand U140439 ( n60322, n60288, n60225 );
nand U140440 ( n60517, n60518, n60519 );
nand U140441 ( n60519, P2_P2_INSTQUEUE_REG_3__7_, n60452 );
nand U140442 ( n60518, n60453, n60269 );
nand U140443 ( n60430, n60431, n60432 );
nand U140444 ( n60432, P2_P2_INSTQUEUE_REG_2__7_, n60372 );
nand U140445 ( n60431, n60373, n60269 );
nand U140446 ( n60348, n60349, n60350 );
nand U140447 ( n60350, P2_P2_INSTQUEUE_REG_1__7_, n60287 );
nand U140448 ( n60349, n60288, n60269 );
nand U140449 ( n49695, n50341, P3_DATAO_REG_1_ );
nor U140450 ( n14930, n14932, n14933 );
nor U140451 ( n14933, n14823, n14934 );
and U140452 ( n14932, n14820, P1_P1_INSTQUEUE_REG_0__7_ );
nand U140453 ( n48837, P2_P1_INSTQUEUE_REG_8__3_, n48810 );
nand U140454 ( n49214, P2_P1_INSTQUEUE_REG_12__4_, n49179 );
nand U140455 ( n48845, P2_P1_INSTQUEUE_REG_8__4_, n48810 );
nand U140456 ( n49198, P2_P1_INSTQUEUE_REG_12__2_, n49179 );
nand U140457 ( n48829, P2_P1_INSTQUEUE_REG_8__2_, n48810 );
nand U140458 ( n49222, P2_P1_INSTQUEUE_REG_12__5_, n49179 );
nand U140459 ( n48853, P2_P1_INSTQUEUE_REG_8__5_, n48810 );
nand U140460 ( n49178, P2_P1_INSTQUEUE_REG_12__0_, n49179 );
nand U140461 ( n48809, P2_P1_INSTQUEUE_REG_8__0_, n48810 );
nand U140462 ( n49190, P2_P1_INSTQUEUE_REG_12__1_, n49179 );
nand U140463 ( n48821, P2_P1_INSTQUEUE_REG_8__1_, n48810 );
nand U140464 ( n49230, P2_P1_INSTQUEUE_REG_12__6_, n49179 );
nand U140465 ( n48861, P2_P1_INSTQUEUE_REG_8__6_, n48810 );
nand U140466 ( n49206, P2_P1_INSTQUEUE_REG_12__3_, n49179 );
nor U140467 ( n15377, n15378, n15379 );
nor U140468 ( n15379, n14934, n15292 );
and U140469 ( n15378, n15288, P1_P1_INSTQUEUE_REG_4__7_ );
nand U140470 ( n4866, n31638, n31639 );
nand U140471 ( n31639, n2979, P1_P3_DATAO_REG_17_ );
nor U140472 ( n31638, n31640, n31641 );
nor U140473 ( n31641, n76147, n75599 );
nand U140474 ( n4876, n31630, n31631 );
nand U140475 ( n31631, n2979, P1_P3_DATAO_REG_19_ );
nor U140476 ( n31630, n31632, n31633 );
nor U140477 ( n31633, n76149, n75600 );
nand U140478 ( n4931, n31620, n31621 );
nand U140479 ( n31621, P1_P3_DATAO_REG_30_, n2979 );
nor U140480 ( n31620, n31622, n31623 );
nor U140481 ( n31623, n76150, n75601 );
nand U140482 ( n4861, n31642, n31643 );
nand U140483 ( n31643, n2979, P1_P3_DATAO_REG_16_ );
nor U140484 ( n31642, n31644, n31645 );
nor U140485 ( n31645, n76146, n75602 );
nand U140486 ( n4871, n31634, n31635 );
nand U140487 ( n31635, n2979, P1_P3_DATAO_REG_18_ );
nor U140488 ( n31634, n31636, n31637 );
nor U140489 ( n31637, n76148, n75603 );
nand U140490 ( n60062, n60114, n60115 );
nand U140491 ( n60115, n60116, n6554 );
nor U140492 ( n60114, n60118, n76259 );
and U140493 ( n60116, n60117, P2_P2_STATE2_REG_0_ );
nand U140494 ( n26922, n26974, n26975 );
nand U140495 ( n26975, n26976, n3922 );
nor U140496 ( n26974, n26978, n76517 );
and U140497 ( n26976, n26977, P1_P2_STATE2_REG_0_ );
nand U140498 ( n34167, n34219, n34220 );
nand U140499 ( n34220, n34221, n3078 );
nor U140500 ( n34219, n34223, n76461 );
and U140501 ( n34221, n34222, P1_P3_STATE2_REG_0_ );
nand U140502 ( n68921, n68973, n68974 );
nand U140503 ( n68974, n68975, n5679 );
nor U140504 ( n68973, n68977, n76193 );
and U140505 ( n68975, n68976, P2_P3_STATE2_REG_0_ );
nor U140506 ( n60077, n60080, n74556 );
nor U140507 ( n60080, n60081, n6513 );
nor U140508 ( n60081, P2_P2_INSTQUEUEWR_ADDR_REG_0_, n76912 );
nor U140509 ( n26937, n26940, n74555 );
nor U140510 ( n26940, n26941, n3880 );
nor U140511 ( n26941, P1_P2_INSTQUEUEWR_ADDR_REG_0_, n76916 );
nor U140512 ( n34182, n34185, n74561 );
nor U140513 ( n34185, n34186, n3037 );
nor U140514 ( n34186, P1_P3_INSTQUEUEWR_ADDR_REG_0_, n76918 );
nor U140515 ( n68936, n68939, n74562 );
nor U140516 ( n68939, n68940, n5638 );
nor U140517 ( n68940, P2_P3_INSTQUEUEWR_ADDR_REG_0_, n76914 );
nand U140518 ( n16742, n76928, n16748 );
xor U140519 ( n16748, n16749, n16750 );
nand U140520 ( n16750, DIN_30_, P4_DATAO_REG_1_ );
nand U140521 ( n16749, DIN_29_, P4_DATAO_REG_2_ );
nand U140522 ( n13281, n60059, n60060 );
nand U140523 ( n60060, n60061, n60062 );
nor U140524 ( n60059, n60063, n60064 );
nor U140525 ( n60064, P2_P2_INSTQUEUEWR_ADDR_REG_0_, n60065 );
nand U140526 ( n6546, n26919, n26920 );
nand U140527 ( n26920, n26921, n26922 );
nor U140528 ( n26919, n26923, n26924 );
nor U140529 ( n26924, P1_P2_INSTQUEUEWR_ADDR_REG_0_, n26925 );
nand U140530 ( n4301, n34164, n34165 );
nand U140531 ( n34165, n34166, n34167 );
nor U140532 ( n34164, n34168, n34169 );
nor U140533 ( n34169, P1_P3_INSTQUEUEWR_ADDR_REG_0_, n34170 );
nand U140534 ( n11036, n68918, n68919 );
nand U140535 ( n68919, n68920, n68921 );
nor U140536 ( n68918, n68922, n68923 );
nor U140537 ( n68923, P2_P3_INSTQUEUEWR_ADDR_REG_0_, n68924 );
nor U140538 ( n11312, P1_P1_EAX_REG_0_, n9908 );
nor U140539 ( n44991, P2_P1_EAX_REG_0_, n43808 );
nand U140540 ( n42402, n54123, P2_P1_STATE2_REG_2_ );
nor U140541 ( n54123, P2_P1_STATE2_REG_1_, n74648 );
nand U140542 ( n8319, n21140, P1_P1_STATE2_REG_2_ );
nor U140543 ( n21140, P1_P1_STATE2_REG_1_, n74649 );
nand U140544 ( n67467, n67420, n67510 );
nand U140545 ( n67510, P2_P3_INSTADDRPOINTER_REG_27_, n67511 );
nand U140546 ( n32702, n32655, n32745 );
nand U140547 ( n32745, P1_P3_INSTADDRPOINTER_REG_27_, n32746 );
nand U140548 ( n46403, n46356, n46446 );
nand U140549 ( n46446, P2_P1_INSTADDRPOINTER_REG_27_, n46447 );
nand U140550 ( n25462, n25415, n25505 );
nand U140551 ( n25505, P1_P2_INSTADDRPOINTER_REG_27_, n25506 );
nand U140552 ( n58599, n58552, n58642 );
nand U140553 ( n58642, P2_P2_INSTADDRPOINTER_REG_27_, n58643 );
nand U140554 ( n46400, n46401, n74986 );
nand U140555 ( n46401, n7485, n46402 );
not U140556 ( n7485, n46355 );
nand U140557 ( n46402, P2_P1_INSTADDRPOINTER_REG_28_, n46403 );
nand U140558 ( n25459, n25460, n75007 );
nand U140559 ( n25460, n3942, n25461 );
not U140560 ( n3942, n25414 );
nand U140561 ( n25461, P1_P2_INSTADDRPOINTER_REG_28_, n25462 );
nand U140562 ( n58596, n58597, n75008 );
nand U140563 ( n58597, n6574, n58598 );
not U140564 ( n6574, n58551 );
nand U140565 ( n58598, P2_P2_INSTADDRPOINTER_REG_28_, n58599 );
nand U140566 ( n67464, n67465, n75009 );
nand U140567 ( n67465, n5699, n67466 );
not U140568 ( n5699, n67419 );
nand U140569 ( n67466, P2_P3_INSTADDRPOINTER_REG_28_, n67467 );
nand U140570 ( n32699, n32700, n75010 );
nand U140571 ( n32700, n3098, n32701 );
not U140572 ( n3098, n32654 );
nand U140573 ( n32701, P1_P3_INSTADDRPOINTER_REG_28_, n32702 );
nor U140574 ( n9417, P1_P1_INSTQUEUERD_ADDR_REG_0_, n9383 );
nand U140575 ( n4266, n34245, n34246 );
nand U140576 ( n34246, n34247, n34228 );
nand U140577 ( n34245, n188, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U140578 ( n34247, n34248, n34249 );
nand U140579 ( n6511, n27000, n27001 );
nand U140580 ( n27001, n27002, n26983 );
nand U140581 ( n27000, n150, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U140582 ( n27002, n27003, n27004 );
nand U140583 ( n11001, n68999, n69000 );
nand U140584 ( n69000, n69001, n68982 );
nand U140585 ( n68999, n459, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U140586 ( n69001, n69002, n69003 );
nand U140587 ( n13246, n60143, n60144 );
nand U140588 ( n60144, n60145, n60126 );
nand U140589 ( n60143, n423, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U140590 ( n60145, n60146, n60147 );
nand U140591 ( n13256, n60123, n60124 );
nand U140592 ( n60124, n60125, n60126 );
nand U140593 ( n60123, n423, P2_P2_INSTQUEUERD_ADDR_REG_0_ );
nand U140594 ( n60125, n60127, n60128 );
nand U140595 ( n6521, n26980, n26981 );
nand U140596 ( n26981, n26982, n26983 );
nand U140597 ( n26980, n150, P1_P2_INSTQUEUERD_ADDR_REG_0_ );
nand U140598 ( n26982, n26984, n26985 );
nor U140599 ( n14157, n14163, n14164 );
nand U140600 ( n14164, P1_P1_INSTADDRPOINTER_REG_4_, P1_P1_INSTADDRPOINTER_REG_3_ );
nand U140601 ( n4276, n34225, n34226 );
nand U140602 ( n34226, n34227, n34228 );
nand U140603 ( n34225, n188, P1_P3_INSTQUEUERD_ADDR_REG_0_ );
nand U140604 ( n34227, n34229, n34230 );
nand U140605 ( n11011, n68979, n68980 );
nand U140606 ( n68980, n68981, n68982 );
nand U140607 ( n68979, n459, P2_P3_INSTQUEUERD_ADDR_REG_0_ );
nand U140608 ( n68981, n68983, n68984 );
nand U140609 ( n4256, n34264, n34265 );
nand U140610 ( n34265, n34266, n34267 );
nand U140611 ( n34264, n188, P1_P3_INSTQUEUERD_ADDR_REG_4_ );
nor U140612 ( n34266, n29169, n32707 );
nand U140613 ( n6501, n27019, n27020 );
nand U140614 ( n27020, n27021, n27022 );
nand U140615 ( n27019, n150, P1_P2_INSTQUEUERD_ADDR_REG_4_ );
nor U140616 ( n27021, n21856, n25467 );
nand U140617 ( n4261, n34254, n34255 );
nand U140618 ( n34255, n34256, n34228 );
nand U140619 ( n34254, n188, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U140620 ( n34256, n34257, n34258 );
nand U140621 ( n6506, n27011, n27012 );
nand U140622 ( n27012, n27013, n26983 );
nand U140623 ( n27011, n150, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U140624 ( n27013, n27014, n27015 );
nand U140625 ( n10996, n69008, n69009 );
nand U140626 ( n69009, n69010, n68982 );
nand U140627 ( n69008, n459, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U140628 ( n69010, n69011, n69012 );
nand U140629 ( n13241, n60152, n60153 );
nand U140630 ( n60153, n60154, n60126 );
nand U140631 ( n60152, n423, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U140632 ( n60154, n60155, n60156 );
nand U140633 ( n10991, n69016, n69017 );
nand U140634 ( n69017, n69018, n69019 );
nand U140635 ( n69016, n459, P2_P3_INSTQUEUERD_ADDR_REG_4_ );
nor U140636 ( n69018, n62891, n67472 );
nand U140637 ( n13236, n60160, n60161 );
nand U140638 ( n60161, n60162, n60163 );
nand U140639 ( n60160, n423, P2_P2_INSTQUEUERD_ADDR_REG_4_ );
nor U140640 ( n60162, n54947, n58604 );
nand U140641 ( n6516, n26990, n26991 );
nand U140642 ( n26991, n26992, n26983 );
nand U140643 ( n26990, n150, P1_P2_INSTQUEUERD_ADDR_REG_1_ );
nand U140644 ( n26992, n26993, n26994 );
nand U140645 ( n13251, n60133, n60134 );
nand U140646 ( n60134, n60135, n60126 );
nand U140647 ( n60133, n423, P2_P2_INSTQUEUERD_ADDR_REG_1_ );
nand U140648 ( n60135, n60136, n60137 );
nand U140649 ( n4271, n34235, n34236 );
nand U140650 ( n34236, n34237, n34228 );
nand U140651 ( n34235, n188, P1_P3_INSTQUEUERD_ADDR_REG_1_ );
nand U140652 ( n34237, n34238, n34239 );
nand U140653 ( n11006, n68989, n68990 );
nand U140654 ( n68990, n68991, n68982 );
nand U140655 ( n68989, n459, P2_P3_INSTQUEUERD_ADDR_REG_1_ );
nand U140656 ( n68991, n68992, n68993 );
nand U140657 ( n15491, n47991, n47992 );
nand U140658 ( n47992, n47993, n47974 );
nand U140659 ( n47991, n493, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U140660 ( n47993, n47994, n47995 );
nand U140661 ( n8756, n14779, n14780 );
nand U140662 ( n14780, n14782, n14752 );
nand U140663 ( n14779, n222, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U140664 ( n14782, n14783, n14784 );
nand U140665 ( n15501, n47971, n47972 );
nand U140666 ( n47972, n47973, n47974 );
nand U140667 ( n47971, n493, P2_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U140668 ( n47973, n47975, n47976 );
nand U140669 ( n8766, n14748, n14749 );
nand U140670 ( n14749, n14750, n14752 );
nand U140671 ( n14748, n222, P1_P1_INSTQUEUERD_ADDR_REG_0_ );
nand U140672 ( n14750, n14753, n14754 );
nand U140673 ( n15486, n48000, n48001 );
nand U140674 ( n48001, n48002, n47974 );
nand U140675 ( n48000, n493, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U140676 ( n48002, n48003, n48004 );
nand U140677 ( n8751, n14790, n14792 );
nand U140678 ( n14792, n14793, n14752 );
nand U140679 ( n14790, n222, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U140680 ( n14793, n14794, n14795 );
nand U140681 ( n8746, n14800, n14802 );
nand U140682 ( n14802, n14803, n14804 );
nand U140683 ( n14800, n222, P1_P1_INSTQUEUERD_ADDR_REG_4_ );
nor U140684 ( n14803, n8294, n12837 );
nand U140685 ( n15481, n48008, n48009 );
nand U140686 ( n48009, n48010, n48011 );
nand U140687 ( n48008, n493, P2_P1_INSTQUEUERD_ADDR_REG_4_ );
nor U140688 ( n48010, n42382, n46408 );
nand U140689 ( n8761, n14760, n14762 );
nand U140690 ( n14762, n14763, n14752 );
nand U140691 ( n14760, n222, P1_P1_INSTQUEUERD_ADDR_REG_1_ );
nand U140692 ( n14763, n14764, n14765 );
and U140693 ( n75982, P2_P2_STATE_REG_2_, n76301 );
nand U140694 ( n12316, n62619, n62620 );
nand U140695 ( n62620, P2_P2_ADDRESS_REG_16_, n76300 );
nor U140696 ( n62619, n62621, n62622 );
nor U140697 ( n62621, n74898, n76238 );
nand U140698 ( n12286, n62704, n62705 );
nand U140699 ( n62705, P2_P2_ADDRESS_REG_22_, n76300 );
nor U140700 ( n62704, n62706, n62707 );
nor U140701 ( n62706, n74990, n76237 );
nand U140702 ( n15496, n47981, n47982 );
nand U140703 ( n47982, n47983, n47974 );
nand U140704 ( n47981, n493, P2_P1_INSTQUEUERD_ADDR_REG_1_ );
nand U140705 ( n47983, n47984, n47985 );
nand U140706 ( n12301, n62692, n62693 );
nand U140707 ( n62693, P2_P2_ADDRESS_REG_19_, n76300 );
nor U140708 ( n62692, n62694, n62695 );
nor U140709 ( n62694, n74938, n76237 );
nand U140710 ( n12271, n62716, n62717 );
nand U140711 ( n62717, P2_P2_ADDRESS_REG_25_, n76300 );
nor U140712 ( n62716, n62718, n62719 );
nor U140713 ( n62718, n75000, n76237 );
nand U140714 ( n12331, n62607, n62608 );
nand U140715 ( n62608, P2_P2_ADDRESS_REG_13_, n76299 );
nor U140716 ( n62607, n62609, n62610 );
nor U140717 ( n62609, n74837, n76238 );
nand U140718 ( n12266, n62720, n62721 );
nand U140719 ( n62721, P2_P2_ADDRESS_REG_26_, n76300 );
nor U140720 ( n62720, n62722, n62723 );
nor U140721 ( n62722, n75300, n76237 );
nand U140722 ( n14697, P1_P1_INSTQUEUEWR_ADDR_REG_0_, n73141 );
nand U140723 ( n12296, n62696, n62697 );
nand U140724 ( n62697, P2_P2_ADDRESS_REG_20_, n76300 );
nor U140725 ( n62696, n62698, n62699 );
nor U140726 ( n62698, n73275, n76237 );
nand U140727 ( n12281, n62708, n62709 );
nand U140728 ( n62709, P2_P2_ADDRESS_REG_23_, n76300 );
nor U140729 ( n62708, n62710, n62711 );
nor U140730 ( n62710, n73290, n76237 );
nand U140731 ( n12256, n62787, n62788 );
nand U140732 ( n62788, P2_P2_ADDRESS_REG_28_, n76300 );
nor U140733 ( n62787, n62789, n62790 );
nor U140734 ( n62789, n75063, n76237 );
nand U140735 ( n12326, n62611, n62612 );
nand U140736 ( n62612, P2_P2_ADDRESS_REG_14_, n76300 );
nor U140737 ( n62611, n62613, n62614 );
nor U140738 ( n62613, n73247, n76238 );
nand U140739 ( n12311, n62623, n62624 );
nand U140740 ( n62624, P2_P2_ADDRESS_REG_17_, n76300 );
nor U140741 ( n62623, n62625, n62626 );
nor U140742 ( n62625, n73261, n76238 );
nand U140743 ( n12251, n62791, n62792 );
nand U140744 ( n62792, P2_P2_ADDRESS_REG_29_, n76300 );
nor U140745 ( n62791, n62793, n62794 );
nor U140746 ( n62793, n75177, n76237 );
nand U140747 ( n12346, n62595, n62596 );
nand U140748 ( n62596, P2_P2_ADDRESS_REG_10_, n76299 );
nor U140749 ( n62595, n62597, n62598 );
nor U140750 ( n62597, n74798, n76238 );
nand U140751 ( n12361, n62531, n62532 );
nand U140752 ( n62532, P2_P2_ADDRESS_REG_7_, n76299 );
nor U140753 ( n62531, n62533, n62534 );
nor U140754 ( n62533, n73214, n76238 );
nand U140755 ( n12291, n62700, n62701 );
nand U140756 ( n62701, P2_P2_ADDRESS_REG_21_, n76300 );
nor U140757 ( n62700, n62702, n62703 );
nor U140758 ( n62702, n74969, n76237 );
nand U140759 ( n12276, n62712, n62713 );
nand U140760 ( n62713, P2_P2_ADDRESS_REG_24_, n76300 );
nor U140761 ( n62712, n62714, n62715 );
nor U140762 ( n62714, n73295, n76237 );
nand U140763 ( n12321, n62615, n62616 );
nand U140764 ( n62616, P2_P2_ADDRESS_REG_15_, n76300 );
nor U140765 ( n62615, n62617, n62618 );
nor U140766 ( n62617, n74882, n76238 );
nand U140767 ( n12306, n62688, n62689 );
nand U140768 ( n62689, P2_P2_ADDRESS_REG_18_, n76300 );
nor U140769 ( n62688, n62690, n62691 );
nor U140770 ( n62690, n74925, n76237 );
nand U140771 ( n12366, n62527, n62528 );
nand U140772 ( n62528, P2_P2_ADDRESS_REG_6_, n76299 );
nor U140773 ( n62527, n62529, n62530 );
nor U140774 ( n62529, n74747, n76238 );
nand U140775 ( n12336, n62603, n62604 );
nand U140776 ( n62604, P2_P2_ADDRESS_REG_12_, n76299 );
nor U140777 ( n62603, n62605, n62606 );
nor U140778 ( n62605, n74827, n76238 );
nand U140779 ( n12351, n62591, n62592 );
nand U140780 ( n62592, P2_P2_ADDRESS_REG_9_, n76299 );
nor U140781 ( n62591, n62593, n62594 );
nor U140782 ( n62593, n74788, n76238 );
nand U140783 ( n12261, n62724, n62725 );
nand U140784 ( n62725, P2_P2_ADDRESS_REG_27_, n76300 );
nor U140785 ( n62724, n62726, n62727 );
nor U140786 ( n62726, n73316, n76237 );
nand U140787 ( n12341, n62599, n62600 );
nand U140788 ( n62600, P2_P2_ADDRESS_REG_11_, n76299 );
nor U140789 ( n62599, n62601, n62602 );
nor U140790 ( n62601, n73233, n76238 );
nand U140791 ( n12356, n62587, n62588 );
nand U140792 ( n62588, P2_P2_ADDRESS_REG_8_, n76299 );
nor U140793 ( n62587, n62589, n62590 );
nor U140794 ( n62589, n74743, n76238 );
nor U140795 ( n68514, n68519, n68520 );
nand U140796 ( n68520, P2_P3_INSTADDRPOINTER_REG_4_, P2_P3_INSTADDRPOINTER_REG_3_ );
nor U140797 ( n33758, n33763, n33764 );
nand U140798 ( n33764, P1_P3_INSTADDRPOINTER_REG_4_, P1_P3_INSTADDRPOINTER_REG_3_ );
nor U140799 ( n47493, n47498, n47499 );
nand U140800 ( n47499, P2_P1_INSTADDRPOINTER_REG_4_, P2_P1_INSTADDRPOINTER_REG_3_ );
nor U140801 ( n26513, n26518, n26519 );
nand U140802 ( n26519, P1_P2_INSTADDRPOINTER_REG_4_, P1_P2_INSTADDRPOINTER_REG_3_ );
nor U140803 ( n59652, n59657, n59658 );
nand U140804 ( n59658, P2_P2_INSTADDRPOINTER_REG_4_, P2_P2_INSTADDRPOINTER_REG_3_ );
nor U140805 ( n13883, n5214, n13892 );
nand U140806 ( n13892, P1_P1_INSTADDRPOINTER_REG_7_, n12732 );
and U140807 ( n75983, P1_P2_STATE_REG_2_, n76555 );
nand U140808 ( n5581, n29064, n29065 );
nand U140809 ( n29065, P1_P2_ADDRESS_REG_16_, n76554 );
nor U140810 ( n29064, n29066, n29067 );
nor U140811 ( n29066, n74899, n76507 );
nand U140812 ( n5551, n29092, n29093 );
nand U140813 ( n29093, P1_P2_ADDRESS_REG_22_, n76554 );
nor U140814 ( n29092, n29094, n29095 );
nor U140815 ( n29094, n74991, n76506 );
nand U140816 ( n5536, n29104, n29105 );
nand U140817 ( n29105, P1_P2_ADDRESS_REG_25_, n76554 );
nor U140818 ( n29104, n29106, n29107 );
nor U140819 ( n29106, n74999, n76506 );
nand U140820 ( n5566, n29076, n29077 );
nand U140821 ( n29077, P1_P2_ADDRESS_REG_19_, n76554 );
nor U140822 ( n29076, n29078, n29079 );
nor U140823 ( n29078, n74939, n76506 );
nand U140824 ( n5596, n29052, n29053 );
nand U140825 ( n29053, P1_P2_ADDRESS_REG_13_, n76553 );
nor U140826 ( n29052, n29054, n29055 );
nor U140827 ( n29054, n74838, n76507 );
nand U140828 ( n5531, n29108, n29109 );
nand U140829 ( n29109, P1_P2_ADDRESS_REG_26_, n76554 );
nor U140830 ( n29108, n29110, n29111 );
nor U140831 ( n29110, n75301, n76506 );
nand U140832 ( n5521, n29116, n29117 );
nand U140833 ( n29117, P1_P2_ADDRESS_REG_28_, n76554 );
nor U140834 ( n29116, n29118, n29119 );
nor U140835 ( n29118, n75064, n76506 );
nand U140836 ( n5546, n29096, n29097 );
nand U140837 ( n29097, P1_P2_ADDRESS_REG_23_, n76554 );
nor U140838 ( n29096, n29098, n29099 );
nor U140839 ( n29098, n73291, n76506 );
nand U140840 ( n5561, n29080, n29081 );
nand U140841 ( n29081, P1_P2_ADDRESS_REG_20_, n76554 );
nor U140842 ( n29080, n29082, n29083 );
nor U140843 ( n29082, n73276, n76506 );
nand U140844 ( n5576, n29068, n29069 );
nand U140845 ( n29069, P1_P2_ADDRESS_REG_17_, n76554 );
nor U140846 ( n29068, n29070, n29071 );
nor U140847 ( n29070, n73262, n76507 );
nand U140848 ( n5591, n29056, n29057 );
nand U140849 ( n29057, P1_P2_ADDRESS_REG_14_, n76554 );
nor U140850 ( n29056, n29058, n29059 );
nor U140851 ( n29058, n73248, n76507 );
nand U140852 ( n5516, n29120, n29121 );
nand U140853 ( n29121, P1_P2_ADDRESS_REG_29_, n76554 );
nor U140854 ( n29120, n29122, n29123 );
nor U140855 ( n29122, n75178, n76506 );
and U140856 ( n75984, P2_P1_STATE_REG_2_, n76373 );
nand U140857 ( n5586, n29060, n29061 );
nand U140858 ( n29061, P1_P2_ADDRESS_REG_15_, n76554 );
nor U140859 ( n29060, n29062, n29063 );
nor U140860 ( n29062, n74883, n76507 );
nand U140861 ( n5611, n29036, n29037 );
nand U140862 ( n29037, P1_P2_ADDRESS_REG_10_, n76553 );
nor U140863 ( n29036, n29038, n29039 );
nor U140864 ( n29038, n74799, n76507 );
nand U140865 ( n5626, n29024, n29025 );
nand U140866 ( n29025, P1_P2_ADDRESS_REG_7_, n76553 );
nor U140867 ( n29024, n29026, n29027 );
nor U140868 ( n29026, n73215, n76507 );
nand U140869 ( n14561, n54803, n54804 );
nand U140870 ( n54804, P2_P1_ADDRESS_REG_16_, n76372 );
nor U140871 ( n54803, n54805, n54806 );
nor U140872 ( n54805, n74914, n76307 );
nand U140873 ( n14531, n54842, n54843 );
nand U140874 ( n54843, P2_P1_ADDRESS_REG_22_, n76372 );
nor U140875 ( n54842, n54844, n54845 );
nor U140876 ( n54844, n75005, n76306 );
nand U140877 ( n5541, n29100, n29101 );
nand U140878 ( n29101, P1_P2_ADDRESS_REG_24_, n76554 );
nor U140879 ( n29100, n29102, n29103 );
nor U140880 ( n29102, n73294, n76506 );
nand U140881 ( n5556, n29088, n29089 );
nand U140882 ( n29089, P1_P2_ADDRESS_REG_21_, n76554 );
nor U140883 ( n29088, n29090, n29091 );
nor U140884 ( n29090, n74970, n76506 );
nand U140885 ( n14516, n54854, n54855 );
nand U140886 ( n54855, P2_P1_ADDRESS_REG_25_, n76372 );
nor U140887 ( n54854, n54856, n54857 );
nor U140888 ( n54856, n75014, n76306 );
nand U140889 ( n14546, n54830, n54831 );
nand U140890 ( n54831, P2_P1_ADDRESS_REG_19_, n76372 );
nor U140891 ( n54830, n54832, n54833 );
nor U140892 ( n54832, n74958, n76306 );
nand U140893 ( n5571, n29072, n29073 );
nand U140894 ( n29073, P1_P2_ADDRESS_REG_18_, n76554 );
nor U140895 ( n29072, n29074, n29075 );
nor U140896 ( n29074, n74926, n76506 );
nand U140897 ( n5601, n29048, n29049 );
nand U140898 ( n29049, P1_P2_ADDRESS_REG_12_, n76553 );
nor U140899 ( n29048, n29050, n29051 );
nor U140900 ( n29050, n74828, n76507 );
nand U140901 ( n5616, n29032, n29033 );
nand U140902 ( n29033, P1_P2_ADDRESS_REG_9_, n76553 );
nor U140903 ( n29032, n29034, n29035 );
nor U140904 ( n29034, n74789, n76507 );
nand U140905 ( n5631, n29020, n29021 );
nand U140906 ( n29021, P1_P2_ADDRESS_REG_6_, n76553 );
nor U140907 ( n29020, n29022, n29023 );
nor U140908 ( n29022, n74748, n76507 );
nand U140909 ( n14576, n54791, n54792 );
nand U140910 ( n54792, P2_P1_ADDRESS_REG_13_, n76371 );
nor U140911 ( n54791, n54793, n54794 );
nor U140912 ( n54793, n74868, n76307 );
nand U140913 ( n14511, n54858, n54859 );
nand U140914 ( n54859, P2_P1_ADDRESS_REG_26_, n76372 );
nor U140915 ( n54858, n54860, n54861 );
nor U140916 ( n54860, n75302, n76306 );
nand U140917 ( n5526, n29112, n29113 );
nand U140918 ( n29113, P1_P2_ADDRESS_REG_27_, n76554 );
nor U140919 ( n29112, n29114, n29115 );
nor U140920 ( n29114, n73317, n76506 );
nand U140921 ( n14541, n54834, n54835 );
nand U140922 ( n54835, P2_P1_ADDRESS_REG_20_, n76372 );
nor U140923 ( n54834, n54836, n54837 );
nor U140924 ( n54836, n73280, n76306 );
nand U140925 ( n14526, n54846, n54847 );
nand U140926 ( n54847, P2_P1_ADDRESS_REG_23_, n76372 );
nor U140927 ( n54846, n54848, n54849 );
nor U140928 ( n54848, n73304, n76306 );
nand U140929 ( n14501, n54881, n54882 );
nand U140930 ( n54882, P2_P1_ADDRESS_REG_28_, n76372 );
nor U140931 ( n54881, n54883, n54884 );
nor U140932 ( n54883, n75237, n76306 );
nand U140933 ( n5606, n29044, n29045 );
nand U140934 ( n29045, P1_P2_ADDRESS_REG_11_, n76553 );
nor U140935 ( n29044, n29046, n29047 );
nor U140936 ( n29046, n73234, n76507 );
nand U140937 ( n5621, n29028, n29029 );
nand U140938 ( n29029, P1_P2_ADDRESS_REG_8_, n76553 );
nor U140939 ( n29028, n29030, n29031 );
nor U140940 ( n29030, n74744, n76507 );
nand U140941 ( n14571, n54795, n54796 );
nand U140942 ( n54796, P2_P1_ADDRESS_REG_14_, n76372 );
nor U140943 ( n54795, n54797, n54798 );
nor U140944 ( n54797, n73253, n76307 );
nand U140945 ( n14556, n54822, n54823 );
nand U140946 ( n54823, P2_P1_ADDRESS_REG_17_, n76372 );
nor U140947 ( n54822, n54824, n54825 );
nor U140948 ( n54824, n73267, n76307 );
nand U140949 ( n14591, n54779, n54780 );
nand U140950 ( n54780, P2_P1_ADDRESS_REG_10_, n76371 );
nor U140951 ( n54779, n54781, n54782 );
nor U140952 ( n54781, n74815, n76307 );
nand U140953 ( n14606, n54763, n54764 );
nand U140954 ( n54764, P2_P1_ADDRESS_REG_7_, n76371 );
nor U140955 ( n54763, n54765, n54766 );
nor U140956 ( n54765, n73221, n76307 );
nand U140957 ( n14536, n54838, n54839 );
nand U140958 ( n54839, P2_P1_ADDRESS_REG_21_, n76372 );
nor U140959 ( n54838, n54840, n54841 );
nor U140960 ( n54840, n74995, n76306 );
nand U140961 ( n14521, n54850, n54851 );
nand U140962 ( n54851, P2_P1_ADDRESS_REG_24_, n76372 );
nor U140963 ( n54850, n54852, n54853 );
nor U140964 ( n54852, n73308, n76306 );
nand U140965 ( n14566, n54799, n54800 );
nand U140966 ( n54800, P2_P1_ADDRESS_REG_15_, n76372 );
nor U140967 ( n54799, n54801, n54802 );
nor U140968 ( n54801, n74904, n76307 );
nand U140969 ( n14551, n54826, n54827 );
nand U140970 ( n54827, P2_P1_ADDRESS_REG_18_, n76372 );
nor U140971 ( n54826, n54828, n54829 );
nor U140972 ( n54828, n74951, n76306 );
nand U140973 ( n14581, n54787, n54788 );
nand U140974 ( n54788, P2_P1_ADDRESS_REG_12_, n76371 );
nor U140975 ( n54787, n54789, n54790 );
nor U140976 ( n54789, n74860, n76307 );
nand U140977 ( n14596, n54775, n54776 );
nand U140978 ( n54776, P2_P1_ADDRESS_REG_9_, n76371 );
nor U140979 ( n54775, n54777, n54778 );
nor U140980 ( n54777, n74811, n76307 );
nand U140981 ( n14611, n54744, n54745 );
nand U140982 ( n54745, P2_P1_ADDRESS_REG_6_, n76371 );
nor U140983 ( n54744, n54746, n54747 );
nor U140984 ( n54746, n75965, n76307 );
nand U140985 ( n14496, n54885, n54886 );
nand U140986 ( n54886, P2_P1_ADDRESS_REG_29_, n76372 );
nor U140987 ( n54885, n54887, n54888 );
nor U140988 ( n54887, n75328, n76306 );
nand U140989 ( n14506, n54877, n54878 );
nand U140990 ( n54878, P2_P1_ADDRESS_REG_27_, n76372 );
nor U140991 ( n54877, n54879, n54880 );
nor U140992 ( n54879, n73391, n76306 );
nand U140993 ( n14586, n54783, n54784 );
nand U140994 ( n54784, P2_P1_ADDRESS_REG_11_, n76371 );
nor U140995 ( n54783, n54785, n54786 );
nor U140996 ( n54785, n73239, n76307 );
nand U140997 ( n14601, n54767, n54768 );
nand U140998 ( n54768, P2_P1_ADDRESS_REG_8_, n76371 );
nor U140999 ( n54767, n54769, n54770 );
nor U141000 ( n54769, n74769, n76307 );
nor U141001 ( n15053, n15389, P1_P1_INSTQUEUEWR_ADDR_REG_0_ );
nand U141002 ( n12386, n62511, n62512 );
nand U141003 ( n62512, P2_P2_ADDRESS_REG_2_, n76299 );
nor U141004 ( n62511, n62513, n62514 );
nor U141005 ( n62513, n74640, n76239 );
nand U141006 ( n12381, n62515, n62516 );
nand U141007 ( n62516, P2_P2_ADDRESS_REG_3_, n76299 );
nor U141008 ( n62515, n62517, n62518 );
nor U141009 ( n62517, n74693, n76239 );
nand U141010 ( n12376, n62519, n62520 );
nand U141011 ( n62520, P2_P2_ADDRESS_REG_4_, n76299 );
nor U141012 ( n62519, n62521, n62522 );
nor U141013 ( n62521, n74709, n76239 );
nand U141014 ( n12391, n62507, n62508 );
nand U141015 ( n62508, P2_P2_ADDRESS_REG_1_, n76299 );
nor U141016 ( n62507, n62509, n62510 );
nor U141017 ( n62509, n72960, n76239 );
nand U141018 ( n12396, n62503, n62504 );
nand U141019 ( n62504, P2_P2_ADDRESS_REG_0_, n76299 );
nor U141020 ( n62503, n62505, n62506 );
nor U141021 ( n62505, n74619, n76239 );
nand U141022 ( n12371, n62523, n62524 );
nand U141023 ( n62524, P2_P2_ADDRESS_REG_5_, n76299 );
nor U141024 ( n62523, n62525, n62526 );
nor U141025 ( n62525, n73198, n76239 );
nor U141026 ( n33537, n3463, n33544 );
nand U141027 ( n33544, P1_P3_INSTADDRPOINTER_REG_7_, n32630 );
nor U141028 ( n68293, n6078, n68300 );
nand U141029 ( n68300, P2_P3_INSTADDRPOINTER_REG_7_, n67395 );
nor U141030 ( n26292, n4300, n26299 );
nand U141031 ( n26299, P1_P2_INSTADDRPOINTER_REG_7_, n25390 );
nor U141032 ( n59431, n6933, n59438 );
nand U141033 ( n59438, P2_P2_INSTADDRPOINTER_REG_7_, n58527 );
nor U141034 ( n47262, n7868, n47269 );
nand U141035 ( n47269, P2_P1_INSTADDRPOINTER_REG_7_, n46331 );
nor U141036 ( n46451, n46457, n46458 );
nand U141037 ( n46458, P2_P1_INSTADDRPOINTER_REG_26_, P2_P1_INSTADDRPOINTER_REG_27_ );
nand U141038 ( n5651, n29004, n29005 );
nand U141039 ( n29005, P1_P2_ADDRESS_REG_2_, n76553 );
nor U141040 ( n29004, n29006, n29007 );
nor U141041 ( n29006, n74641, n76508 );
nand U141042 ( n5646, n29008, n29009 );
nand U141043 ( n29009, P1_P2_ADDRESS_REG_3_, n76553 );
nor U141044 ( n29008, n29010, n29011 );
nor U141045 ( n29010, n74694, n76508 );
nand U141046 ( n5641, n29012, n29013 );
nand U141047 ( n29013, P1_P2_ADDRESS_REG_4_, n76553 );
nor U141048 ( n29012, n29014, n29015 );
nor U141049 ( n29014, n74710, n76508 );
nand U141050 ( n5661, n28992, n28993 );
nand U141051 ( n28993, P1_P2_ADDRESS_REG_0_, n76553 );
nor U141052 ( n28992, n28994, n28995 );
nor U141053 ( n28994, n74620, n76508 );
nand U141054 ( n5656, n29000, n29001 );
nand U141055 ( n29001, P1_P2_ADDRESS_REG_1_, n76553 );
nor U141056 ( n29000, n29002, n29003 );
nor U141057 ( n29002, n72961, n76508 );
nand U141058 ( n14631, n54728, n54729 );
nand U141059 ( n54729, P2_P1_ADDRESS_REG_2_, n76371 );
nor U141060 ( n54728, n54730, n54731 );
nor U141061 ( n54730, n74672, n76308 );
nand U141062 ( n5636, n29016, n29017 );
nand U141063 ( n29017, P1_P2_ADDRESS_REG_5_, n76553 );
nor U141064 ( n29016, n29018, n29019 );
nor U141065 ( n29018, n73199, n76508 );
and U141066 ( n75985, P1_P1_STATE_REG_2_, n76645 );
nand U141067 ( n7841, n21740, n21741 );
nand U141068 ( n21741, P1_P1_ADDRESS_REG_13_, n76643 );
nor U141069 ( n21740, n21742, n21743 );
nor U141070 ( n21742, n74869, n76566 );
nand U141071 ( n7796, n21778, n21779 );
nand U141072 ( n21779, P1_P1_ADDRESS_REG_22_, n76644 );
nor U141073 ( n21778, n21780, n21781 );
nor U141074 ( n21780, n75006, n76565 );
nand U141075 ( n7826, n21752, n21753 );
nand U141076 ( n21753, P1_P1_ADDRESS_REG_16_, n76644 );
nor U141077 ( n21752, n21754, n21755 );
nor U141078 ( n21754, n74915, n76566 );
nand U141079 ( n7781, n21790, n21791 );
nand U141080 ( n21791, P1_P1_ADDRESS_REG_25_, n76644 );
nor U141081 ( n21790, n21792, n21793 );
nor U141082 ( n21792, n75015, n76565 );
xnor U141083 ( n37813, n37814, n37815 );
xor U141084 ( n37815, P4_REG2_REG_6_, n1930 );
nand U141085 ( n7811, n21764, n21765 );
nand U141086 ( n21765, P1_P1_ADDRESS_REG_19_, n76644 );
nor U141087 ( n21764, n21766, n21767 );
nor U141088 ( n21766, n74959, n76565 );
nand U141089 ( n7836, n21744, n21745 );
nand U141090 ( n21745, P1_P1_ADDRESS_REG_14_, n76644 );
nor U141091 ( n21744, n21746, n21747 );
nor U141092 ( n21746, n73254, n76566 );
nand U141093 ( n14626, n54732, n54733 );
nand U141094 ( n54733, P2_P1_ADDRESS_REG_3_, n76371 );
nor U141095 ( n54732, n54734, n54735 );
nor U141096 ( n54734, n74726, n76308 );
nand U141097 ( n7791, n21782, n21783 );
nand U141098 ( n21783, P1_P1_ADDRESS_REG_23_, n76644 );
nor U141099 ( n21782, n21784, n21785 );
nor U141100 ( n21784, n73305, n76565 );
nand U141101 ( n7776, n21794, n21795 );
nand U141102 ( n21795, P1_P1_ADDRESS_REG_26_, n76644 );
nor U141103 ( n21794, n21796, n21797 );
nor U141104 ( n21796, n75303, n76565 );
nand U141105 ( n7821, n21756, n21757 );
nand U141106 ( n21757, P1_P1_ADDRESS_REG_17_, n76644 );
nor U141107 ( n21756, n21758, n21759 );
nor U141108 ( n21758, n73268, n76566 );
nand U141109 ( n7856, n21728, n21729 );
nand U141110 ( n21729, P1_P1_ADDRESS_REG_10_, n76643 );
nor U141111 ( n21728, n21730, n21731 );
nor U141112 ( n21730, n74816, n76566 );
nand U141113 ( n7761, n21806, n21807 );
nand U141114 ( n21807, P1_P1_ADDRESS_REG_29_, n76644 );
nor U141115 ( n21806, n21808, n21809 );
nor U141116 ( n21808, n75329, n76565 );
nand U141117 ( n7806, n21770, n21771 );
nand U141118 ( n21771, P1_P1_ADDRESS_REG_20_, n76644 );
nor U141119 ( n21770, n21772, n21773 );
nor U141120 ( n21772, n73281, n76565 );
nand U141121 ( n7766, n21802, n21803 );
nand U141122 ( n21803, P1_P1_ADDRESS_REG_28_, n76644 );
nor U141123 ( n21802, n21804, n21805 );
nor U141124 ( n21804, n75238, n76565 );
nand U141125 ( n7771, n21798, n21799 );
nand U141126 ( n21799, P1_P1_ADDRESS_REG_27_, n76644 );
nor U141127 ( n21798, n21800, n21801 );
nor U141128 ( n21800, n73392, n76565 );
nand U141129 ( n14621, n54736, n54737 );
nand U141130 ( n54737, P2_P1_ADDRESS_REG_4_, n76371 );
nor U141131 ( n54736, n54738, n54739 );
nor U141132 ( n54738, n74728, n76308 );
nand U141133 ( n7786, n21786, n21787 );
nand U141134 ( n21787, P1_P1_ADDRESS_REG_24_, n76644 );
nor U141135 ( n21786, n21788, n21789 );
nor U141136 ( n21788, n73309, n76565 );
nand U141137 ( n7801, n21774, n21775 );
nand U141138 ( n21775, P1_P1_ADDRESS_REG_21_, n76644 );
nor U141139 ( n21774, n21776, n21777 );
nor U141140 ( n21776, n74996, n76565 );
nand U141141 ( n7831, n21748, n21749 );
nand U141142 ( n21749, P1_P1_ADDRESS_REG_15_, n76644 );
nor U141143 ( n21748, n21750, n21751 );
nor U141144 ( n21750, n74905, n76566 );
nand U141145 ( n7816, n21760, n21761 );
nand U141146 ( n21761, P1_P1_ADDRESS_REG_18_, n76644 );
nor U141147 ( n21760, n21762, n21763 );
nor U141148 ( n21762, n74952, n76565 );
nand U141149 ( n7846, n21736, n21737 );
nand U141150 ( n21737, P1_P1_ADDRESS_REG_12_, n76643 );
nor U141151 ( n21736, n21738, n21739 );
nor U141152 ( n21738, n74861, n76566 );
nand U141153 ( n7861, n21724, n21725 );
nand U141154 ( n21725, P1_P1_ADDRESS_REG_9_, n76643 );
nor U141155 ( n21724, n21726, n21727 );
nor U141156 ( n21726, n74812, n76566 );
nand U141157 ( n7871, n21716, n21717 );
nand U141158 ( n21717, P1_P1_ADDRESS_REG_7_, n76643 );
nor U141159 ( n21716, n21718, n21719 );
nor U141160 ( n21718, n73222, n76566 );
nand U141161 ( n7876, n21712, n21713 );
nand U141162 ( n21713, P1_P1_ADDRESS_REG_6_, n76643 );
nor U141163 ( n21712, n21714, n21715 );
nor U141164 ( n21714, n75967, n76566 );
nand U141165 ( n7851, n21732, n21733 );
nand U141166 ( n21733, P1_P1_ADDRESS_REG_11_, n76643 );
nor U141167 ( n21732, n21734, n21735 );
nor U141168 ( n21734, n73240, n76566 );
nand U141169 ( n7866, n21720, n21721 );
nand U141170 ( n21721, P1_P1_ADDRESS_REG_8_, n76643 );
nor U141171 ( n21720, n21722, n21723 );
nor U141172 ( n21722, n74770, n76566 );
nand U141173 ( n14641, n54720, n54721 );
nand U141174 ( n54721, P2_P1_ADDRESS_REG_0_, n76371 );
nor U141175 ( n54720, n54722, n54723 );
nor U141176 ( n54722, n74655, n76308 );
nand U141177 ( n14636, n54724, n54725 );
nand U141178 ( n54725, P2_P1_ADDRESS_REG_1_, n76371 );
nor U141179 ( n54724, n54726, n54727 );
nor U141180 ( n54726, n72964, n76308 );
nand U141181 ( n14616, n54740, n54741 );
nand U141182 ( n54741, P2_P1_ADDRESS_REG_5_, n76371 );
nor U141183 ( n54740, n54742, n54743 );
nor U141184 ( n54742, n73206, n76308 );
nor U141185 ( n67515, n67520, n67521 );
nand U141186 ( n67521, P2_P3_INSTADDRPOINTER_REG_26_, P2_P3_INSTADDRPOINTER_REG_27_ );
nor U141187 ( n32750, n32755, n32756 );
nand U141188 ( n32756, P1_P3_INSTADDRPOINTER_REG_26_, P1_P3_INSTADDRPOINTER_REG_27_ );
nor U141189 ( n25510, n25515, n25516 );
nand U141190 ( n25516, P1_P2_INSTADDRPOINTER_REG_26_, P1_P2_INSTADDRPOINTER_REG_27_ );
nor U141191 ( n58647, n58652, n58653 );
nand U141192 ( n58653, P2_P2_INSTADDRPOINTER_REG_26_, P2_P2_INSTADDRPOINTER_REG_27_ );
nand U141193 ( n7906, n21688, n21689 );
nand U141194 ( n21689, P1_P1_ADDRESS_REG_0_, n76643 );
nor U141195 ( n21688, n21690, n21691 );
nor U141196 ( n21690, n74656, n76567 );
nand U141197 ( n7896, n21696, n21697 );
nand U141198 ( n21697, P1_P1_ADDRESS_REG_2_, n76643 );
nor U141199 ( n21696, n21698, n21699 );
nor U141200 ( n21698, n74673, n76567 );
nand U141201 ( n7901, n21692, n21693 );
nand U141202 ( n21693, P1_P1_ADDRESS_REG_1_, n76643 );
nor U141203 ( n21692, n21694, n21695 );
nor U141204 ( n21694, n72965, n76567 );
nand U141205 ( n7886, n21704, n21705 );
nand U141206 ( n21705, P1_P1_ADDRESS_REG_4_, n76643 );
nor U141207 ( n21704, n21706, n21707 );
nor U141208 ( n21706, n74729, n76567 );
nand U141209 ( n7891, n21700, n21701 );
nand U141210 ( n21701, P1_P1_ADDRESS_REG_3_, n76643 );
nor U141211 ( n21700, n21702, n21703 );
nor U141212 ( n21702, n74727, n76567 );
nand U141213 ( n7881, n21708, n21709 );
nand U141214 ( n21709, P1_P1_ADDRESS_REG_5_, n76643 );
nor U141215 ( n21708, n21710, n21711 );
nor U141216 ( n21710, n73207, n76567 );
nor U141217 ( n63142, P2_P3_EBX_REG_27_, n6323 );
nor U141218 ( n29379, P1_P3_EBX_REG_27_, n3689 );
nor U141219 ( n42601, P2_P1_EBX_REG_27_, n8104 );
nor U141220 ( n22060, P1_P2_EBX_REG_27_, n4583 );
nor U141221 ( n55170, P2_P2_EBX_REG_27_, n7215 );
nor U141222 ( n8539, P1_P1_EBX_REG_27_, n5450 );
nor U141223 ( n63171, n6323, n63172 );
nor U141224 ( n63172, n63173, n75073 );
nor U141225 ( n63173, P2_P3_EBX_REG_25_, n63174 );
nor U141226 ( n29408, n3689, n29409 );
nor U141227 ( n29409, n29410, n75072 );
nor U141228 ( n29410, P1_P3_EBX_REG_25_, n29411 );
nor U141229 ( n22089, n4583, n22090 );
nor U141230 ( n22090, n22091, n75074 );
nor U141231 ( n22091, P1_P2_EBX_REG_25_, n22092 );
nor U141232 ( n55199, n7215, n55200 );
nor U141233 ( n55200, n55201, n75076 );
nor U141234 ( n55201, P2_P2_EBX_REG_25_, n55202 );
nand U141235 ( n27635, n27636, n27637 );
nand U141236 ( n27637, P1_P2_INSTQUEUE_REG_7__0_, n27638 );
nand U141237 ( n27636, n27639, n3 );
not U141238 ( n3, n27043 );
nand U141239 ( n60788, n60789, n60790 );
nand U141240 ( n60790, P2_P2_INSTQUEUE_REG_7__0_, n60791 );
nand U141241 ( n60789, n60792, n248 );
not U141242 ( n248, n60184 );
nand U141243 ( n806, n21625, n21626 );
nand U141244 ( n21626, P1_P3_DATAO_REG_1_, n76042 );
nor U141245 ( n21625, n21627, n21628 );
nor U141246 ( n21628, n13650, n73566 );
nand U141247 ( n12625, n14397, n14398 );
nand U141248 ( n14398, n14399, n4968 );
nand U141249 ( n14397, n14402, n14204 );
xor U141250 ( n14399, n14400, P1_P1_INSTADDRPOINTER_REG_2_ );
nand U141251 ( n4851, n31655, n31656 );
nand U141252 ( n31656, n2979, P1_P3_DATAO_REG_14_ );
nor U141253 ( n31655, n31657, n31658 );
nor U141254 ( n31657, n76153, n75684 );
nand U141255 ( n4846, n31659, n31660 );
nand U141256 ( n31660, n2979, P1_P3_DATAO_REG_13_ );
nor U141257 ( n31659, n31661, n31662 );
nor U141258 ( n31661, n76153, n75685 );
nand U141259 ( n4841, n31663, n31664 );
nand U141260 ( n31664, n2979, P1_P3_DATAO_REG_12_ );
nor U141261 ( n31663, n31665, n31666 );
nor U141262 ( n31665, n76153, n75686 );
nand U141263 ( n4836, n31667, n31668 );
nand U141264 ( n31668, n2979, P1_P3_DATAO_REG_11_ );
nor U141265 ( n31667, n31669, n31670 );
nor U141266 ( n31669, n76152, n75687 );
nand U141267 ( n4826, n31675, n31676 );
nand U141268 ( n31676, n2979, P1_P3_DATAO_REG_9_ );
nor U141269 ( n31675, n31677, n31678 );
nor U141270 ( n31677, n76151, n75688 );
nand U141271 ( n4821, n31679, n31680 );
nand U141272 ( n31680, n2979, P1_P3_DATAO_REG_8_ );
nor U141273 ( n31679, n31681, n31682 );
nor U141274 ( n31681, n76152, n75689 );
nand U141275 ( n4806, n31695, n31696 );
nand U141276 ( n31696, n2979, P1_P3_DATAO_REG_5_ );
nor U141277 ( n31695, n31697, n31698 );
nor U141278 ( n31697, n76150, n75690 );
nand U141279 ( n4791, n31707, n31708 );
nand U141280 ( n31708, n2979, P1_P3_DATAO_REG_2_ );
nor U141281 ( n31707, n31709, n31710 );
nor U141282 ( n31709, n76147, n75691 );
nand U141283 ( n4796, n31703, n31704 );
nand U141284 ( n31704, n2979, P1_P3_DATAO_REG_3_ );
nor U141285 ( n31703, n31705, n31706 );
nor U141286 ( n31705, n76148, n75692 );
nand U141287 ( n4786, n31711, n31712 );
nand U141288 ( n31712, n2979, P1_P3_DATAO_REG_1_ );
nor U141289 ( n31711, n31713, n31714 );
nor U141290 ( n31713, n76146, n75693 );
nand U141291 ( n4801, n31699, n31700 );
nand U141292 ( n31700, n2979, P1_P3_DATAO_REG_4_ );
nor U141293 ( n31699, n31701, n31702 );
nor U141294 ( n31701, n76149, n75694 );
nand U141295 ( n4811, n31687, n31688 );
nand U141296 ( n31688, n2979, P1_P3_DATAO_REG_6_ );
nor U141297 ( n31687, n31689, n31690 );
nor U141298 ( n31689, n76151, n75695 );
nand U141299 ( n4816, n31683, n31684 );
nand U141300 ( n31684, n2979, P1_P3_DATAO_REG_7_ );
nor U141301 ( n31683, n31685, n31686 );
nor U141302 ( n31685, n76152, n75696 );
nand U141303 ( n4856, n31651, n31652 );
nand U141304 ( n31652, n2979, P1_P3_DATAO_REG_15_ );
nor U141305 ( n31651, n31653, n31654 );
nor U141306 ( n31653, n76145, n75697 );
nand U141307 ( n4781, n31715, n31716 );
nand U141308 ( n31716, n2979, P1_P3_DATAO_REG_0_ );
nor U141309 ( n31715, n31717, n31718 );
nor U141310 ( n31717, n76145, n75698 );
nand U141311 ( n4831, n31671, n31672 );
nand U141312 ( n31672, n2979, P1_P3_DATAO_REG_10_ );
nor U141313 ( n31671, n31673, n31674 );
nor U141314 ( n31673, n76151, n75699 );
nand U141315 ( n27459, n26939, n28417 );
nand U141316 ( n28417, P1_P2_INSTQUEUEWR_ADDR_REG_1_, n74423 );
nand U141317 ( n60608, n60079, n61726 );
nand U141318 ( n61726, P2_P2_INSTQUEUEWR_ADDR_REG_1_, n74424 );
nand U141319 ( n69448, n68938, n70326 );
nand U141320 ( n70326, P2_P3_INSTQUEUEWR_ADDR_REG_1_, n74425 );
nand U141321 ( n34704, n34184, n35598 );
nand U141322 ( n35598, P1_P3_INSTQUEUEWR_ADDR_REG_1_, n74426 );
nand U141323 ( n4776, n31723, n31724 );
nand U141324 ( n31724, P1_P3_UWORD_REG_0_, n31725 );
nor U141325 ( n31723, n31726, n31727 );
nor U141326 ( n31726, n75421, n76138 );
nand U141327 ( n4696, n31757, n31758 );
nand U141328 ( n31758, P1_P3_LWORD_REG_1_, n31725 );
nor U141329 ( n31757, n31759, n31732 );
nor U141330 ( n31759, n72957, n76141 );
nand U141331 ( n4761, n31737, n31738 );
nand U141332 ( n31738, P1_P3_UWORD_REG_3_, n31725 );
nor U141333 ( n31737, n31739, n31740 );
nor U141334 ( n31739, n74876, n76136 );
nand U141335 ( n4771, n31729, n31730 );
nand U141336 ( n31730, P1_P3_UWORD_REG_1_, n76130 );
nor U141337 ( n31729, n31731, n31732 );
nor U141338 ( n31731, n74817, n76137 );
nand U141339 ( n4706, n31749, n31750 );
nand U141340 ( n31750, P1_P3_UWORD_REG_14_, n76130 );
nor U141341 ( n31749, n31751, n31752 );
nor U141342 ( n31751, n75447, n76135 );
nand U141343 ( n4631, n31810, n31811 );
nand U141344 ( n31811, P1_P3_LWORD_REG_14_, n76130 );
nor U141345 ( n31810, n31812, n31752 );
nor U141346 ( n31812, n75278, n76135 );
nand U141347 ( n4691, n31760, n31761 );
nand U141348 ( n31761, P1_P3_LWORD_REG_2_, n76130 );
nor U141349 ( n31760, n31762, n31736 );
nor U141350 ( n31762, n75286, n76141 );
nand U141351 ( n4766, n31733, n31734 );
nand U141352 ( n31734, P1_P3_UWORD_REG_2_, n76129 );
nor U141353 ( n31733, n31735, n31736 );
nor U141354 ( n31735, n75422, n76138 );
nand U141355 ( n4686, n31763, n31764 );
nand U141356 ( n31764, P1_P3_LWORD_REG_3_, n76129 );
nor U141357 ( n31763, n31765, n31740 );
nor U141358 ( n31765, n73135, n76141 );
nand U141359 ( n4701, n31753, n31754 );
nand U141360 ( n31754, P1_P3_LWORD_REG_0_, n76129 );
nor U141361 ( n31753, n31755, n31727 );
nor U141362 ( n31755, n74488, n76134 );
nand U141363 ( n66847, P2_P3_PHYADDRPOINTER_REG_16_, P2_P3_PHYADDRPOINTER_REG_15_ );
nand U141364 ( n24971, P1_P2_PHYADDRPOINTER_REG_16_, P1_P2_PHYADDRPOINTER_REG_15_ );
nand U141365 ( n58106, P2_P2_PHYADDRPOINTER_REG_16_, P2_P2_PHYADDRPOINTER_REG_15_ );
nand U141366 ( n32201, P1_P3_PHYADDRPOINTER_REG_16_, P1_P3_PHYADDRPOINTER_REG_15_ );
nand U141367 ( n27696, n27697, n27698 );
nand U141368 ( n27698, P1_P2_INSTQUEUE_REG_7__7_, n27638 );
nand U141369 ( n27697, n27639, n37 );
not U141370 ( n37, n27133 );
nand U141371 ( n27680, n27681, n27682 );
nand U141372 ( n27682, P1_P2_INSTQUEUE_REG_7__5_, n27638 );
nand U141373 ( n27681, n27639, n28 );
not U141374 ( n28, n27099 );
nand U141375 ( n60831, n60832, n60833 );
nand U141376 ( n60833, P2_P2_INSTQUEUE_REG_7__5_, n60791 );
nand U141377 ( n60832, n60792, n279 );
not U141378 ( n279, n60243 );
nand U141379 ( n60847, n60848, n60849 );
nand U141380 ( n60849, P2_P2_INSTQUEUE_REG_7__7_, n60791 );
nand U141381 ( n60848, n60792, n290 );
not U141382 ( n290, n60277 );
nand U141383 ( n27688, n27689, n27690 );
nand U141384 ( n27690, P1_P2_INSTQUEUE_REG_7__6_, n27638 );
nand U141385 ( n27689, n27639, n33 );
not U141386 ( n33, n27110 );
nand U141387 ( n60839, n60840, n60841 );
nand U141388 ( n60841, P2_P2_INSTQUEUE_REG_7__6_, n60791 );
nand U141389 ( n60840, n60792, n285 );
not U141390 ( n285, n60254 );
nand U141391 ( n45158, P3_REG2_REG_12_, n43666 );
nand U141392 ( n45223, P3_REG1_REG_12_, n43666 );
nand U141393 ( n4636, n31806, n31807 );
nand U141394 ( n31807, P1_P3_LWORD_REG_13_, n31725 );
nor U141395 ( n31806, n31808, n31809 );
nor U141396 ( n31808, n74731, n76136 );
nand U141397 ( n4681, n31766, n31767 );
nand U141398 ( n31767, P1_P3_LWORD_REG_4_, n31725 );
nor U141399 ( n31766, n31768, n31769 );
nor U141400 ( n31768, n75279, n76140 );
nand U141401 ( n4666, n31778, n31779 );
nand U141402 ( n31779, P1_P3_LWORD_REG_7_, n31725 );
nor U141403 ( n31778, n31780, n31781 );
nor U141404 ( n31780, n74582, n76140 );
nand U141405 ( n4651, n31794, n31795 );
nand U141406 ( n31795, P1_P3_LWORD_REG_10_, n31725 );
nor U141407 ( n31794, n31796, n31797 );
nor U141408 ( n31796, n74629, n76138 );
nand U141409 ( n4641, n31802, n31803 );
nand U141410 ( n31803, P1_P3_LWORD_REG_12_, n76129 );
nor U141411 ( n31802, n31804, n31805 );
nor U141412 ( n31804, n75280, n76137 );
nand U141413 ( n4646, n31798, n31799 );
nand U141414 ( n31799, P1_P3_LWORD_REG_11_, n76130 );
nor U141415 ( n31798, n31800, n31801 );
nor U141416 ( n31800, n74676, n76137 );
nand U141417 ( n4656, n31790, n31791 );
nand U141418 ( n31791, P1_P3_LWORD_REG_9_, n76129 );
nor U141419 ( n31790, n31792, n31793 );
nor U141420 ( n31792, n75252, n76139 );
nand U141421 ( n4661, n31782, n31783 );
nand U141422 ( n31783, P1_P3_LWORD_REG_8_, n76130 );
nor U141423 ( n31782, n31784, n31785 );
nor U141424 ( n31784, n75281, n76139 );
nand U141425 ( n4676, n31770, n31771 );
nand U141426 ( n31771, P1_P3_LWORD_REG_5_, n76130 );
nor U141427 ( n31770, n31772, n31773 );
nor U141428 ( n31772, n74540, n76139 );
nand U141429 ( n4671, n31774, n31775 );
nand U141430 ( n31775, P1_P3_LWORD_REG_6_, n76129 );
nor U141431 ( n31774, n31776, n31777 );
nor U141432 ( n31776, n75282, n76140 );
nand U141433 ( n4626, n31813, n31814 );
nand U141434 ( n31814, P1_P3_LWORD_REG_15_, n76129 );
nor U141435 ( n31813, n31815, n31816 );
nor U141436 ( n31815, n74778, n76134 );
nand U141437 ( n26939, P1_P2_INSTQUEUEWR_ADDR_REG_0_, n74555 );
nand U141438 ( n60079, P2_P2_INSTQUEUEWR_ADDR_REG_0_, n74556 );
nand U141439 ( n68938, P2_P3_INSTQUEUEWR_ADDR_REG_0_, n74562 );
nand U141440 ( n34184, P1_P3_INSTQUEUEWR_ADDR_REG_0_, n74561 );
nand U141441 ( n27646, n27647, n27648 );
nand U141442 ( n27648, P1_P2_INSTQUEUE_REG_7__1_, n27638 );
nand U141443 ( n27647, n27639, n8 );
not U141444 ( n8, n27055 );
nand U141445 ( n27664, n27665, n27666 );
nand U141446 ( n27666, P1_P2_INSTQUEUE_REG_7__3_, n27638 );
nand U141447 ( n27665, n27639, n18 );
not U141448 ( n18, n27077 );
nand U141449 ( n27672, n27673, n27674 );
nand U141450 ( n27674, P1_P2_INSTQUEUE_REG_7__4_, n27638 );
nand U141451 ( n27673, n27639, n23 );
not U141452 ( n23, n27088 );
nand U141453 ( n27656, n27657, n27658 );
nand U141454 ( n27658, P1_P2_INSTQUEUE_REG_7__2_, n27638 );
nand U141455 ( n27657, n27639, n13 );
not U141456 ( n13, n27066 );
nand U141457 ( n60815, n60816, n60817 );
nand U141458 ( n60817, P2_P2_INSTQUEUE_REG_7__3_, n60791 );
nand U141459 ( n60816, n60792, n267 );
not U141460 ( n267, n60218 );
nand U141461 ( n60799, n60800, n60801 );
nand U141462 ( n60801, P2_P2_INSTQUEUE_REG_7__1_, n60791 );
nand U141463 ( n60800, n60792, n254 );
not U141464 ( n254, n60196 );
nand U141465 ( n60807, n60808, n60809 );
nand U141466 ( n60809, P2_P2_INSTQUEUE_REG_7__2_, n60791 );
nand U141467 ( n60808, n60792, n260 );
not U141468 ( n260, n60207 );
nand U141469 ( n60823, n60824, n60825 );
nand U141470 ( n60825, P2_P2_INSTQUEUE_REG_7__4_, n60791 );
nand U141471 ( n60824, n60792, n273 );
not U141472 ( n273, n60229 );
nand U141473 ( n35789, P1_P3_STATE_REG_1_, n72928 );
nand U141474 ( n31722, n73192, n35787 );
nand U141475 ( n35787, n35788, n35789 );
nand U141476 ( n35788, P1_P3_STATE_REG_2_, n74654 );
nor U141477 ( n14717, P1_P1_INSTQUEUEWR_ADDR_REG_0_, n14692 );
nor U141478 ( n42632, n42633, n75071 );
nor U141479 ( n42633, P2_P1_EBX_REG_25_, n42634 );
nor U141480 ( n8578, n8579, n75075 );
nor U141481 ( n8579, P1_P1_EBX_REG_25_, n8580 );
nand U141482 ( n33109, P1_P3_INSTADDRPOINTER_REG_17_, P1_P3_INSTADDRPOINTER_REG_16_ );
nand U141483 ( n67270, n67271, n67272 );
nor U141484 ( n67271, P3_D_REG_4_, P3_D_REG_3_ );
nor U141485 ( n67272, P3_D_REG_6_, P3_D_REG_5_ );
nor U141486 ( n67275, P3_D_REG_17_, P3_D_REG_16_ );
nand U141487 ( n67287, n67288, n67289 );
nor U141488 ( n67288, P3_D_REG_26_, P3_D_REG_25_ );
nor U141489 ( n67289, P3_D_REG_28_, P3_D_REG_27_ );
nand U141490 ( n956, n10117, n10118 );
nand U141491 ( n10117, n10119, n76628 );
nor U141492 ( n10119, P3_IR_REG_30_, n10120 );
nand U141493 ( n24460, n74691, n28608 );
nand U141494 ( n28608, n28609, n28610 );
nand U141495 ( n28609, P1_P2_STATE_REG_2_, n73179 );
nand U141496 ( n28610, P1_P2_STATE_REG_1_, n74651 );
nor U141497 ( n67292, P3_D_REG_13_, P3_D_REG_12_ );
nor U141498 ( n67274, P3_D_REG_15_, P3_D_REG_14_ );
nor U141499 ( n27219, n27459, P1_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U141500 ( n60364, n60608, P2_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U141501 ( n23304, P1_P2_EAX_REG_26_, n23259 );
nor U141502 ( n56428, P2_P2_EAX_REG_26_, n56383 );
nor U141503 ( n34464, n34704, P1_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U141504 ( n69214, n69448, P2_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U141505 ( n64828, P2_P3_EAX_REG_26_, n64739 );
nand U141506 ( n67278, n67279, n67280 );
nor U141507 ( n67279, P3_D_REG_2_, P3_D_REG_29_ );
nor U141508 ( n67280, P3_D_REG_31_, P3_D_REG_30_ );
nor U141509 ( n30622, P1_P3_EAX_REG_26_, n30580 );
nand U141510 ( n67208, n68692, n68693 );
nand U141511 ( n68693, n68694, n5834 );
nand U141512 ( n68692, n68696, n68552 );
xor U141513 ( n68694, n68695, P2_P3_INSTADDRPOINTER_REG_2_ );
nand U141514 ( n46256, n47671, n47672 );
nand U141515 ( n47672, n47673, n7622 );
nand U141516 ( n47671, n47675, n47531 );
xor U141517 ( n47673, n47674, P2_P1_INSTADDRPOINTER_REG_2_ );
nand U141518 ( n25310, n26691, n26692 );
nand U141519 ( n26692, n26693, n4063 );
nand U141520 ( n26691, n26695, n26551 );
xor U141521 ( n26693, n26694, P1_P2_INSTADDRPOINTER_REG_2_ );
nand U141522 ( n58449, n59833, n59834 );
nand U141523 ( n59834, n59835, n6695 );
nand U141524 ( n59833, n59837, n59693 );
xor U141525 ( n59835, n59836, P2_P2_INSTADDRPOINTER_REG_2_ );
nor U141526 ( n67291, P3_D_REG_11_, P3_D_REG_10_ );
nand U141527 ( n32552, n33936, n33937 );
nand U141528 ( n33937, n33938, n3235 );
nand U141529 ( n33936, n33940, n33796 );
xor U141530 ( n33938, n33939, P1_P3_INSTADDRPOINTER_REG_2_ );
nand U141531 ( n32961, P1_P3_INSTADDRPOINTER_REG_21_, P1_P3_INSTADDRPOINTER_REG_20_ );
nand U141532 ( n32985, P1_P3_INSTADDRPOINTER_REG_19_, n3503 );
nor U141533 ( n67282, P3_D_REG_9_, P3_D_REG_8_ );
nand U141534 ( n66162, n73186, n70513 );
nand U141535 ( n70513, n70514, n70515 );
nand U141536 ( n70514, P2_P3_STATE_REG_2_, n74657 );
nand U141537 ( n70515, P2_P3_STATE_REG_1_, n72927 );
xor U141538 ( n68541, n68542, P2_P3_INSTADDRPOINTER_REG_4_ );
xor U141539 ( n47520, n47521, P2_P1_INSTADDRPOINTER_REG_4_ );
xor U141540 ( n26540, n26541, P1_P2_INSTADDRPOINTER_REG_4_ );
xor U141541 ( n59682, n59683, P2_P2_INSTADDRPOINTER_REG_4_ );
xor U141542 ( n33785, n33786, P1_P3_INSTADDRPOINTER_REG_4_ );
xor U141543 ( n14190, n14192, P1_P1_INSTADDRPOINTER_REG_4_ );
nand U141544 ( n57586, n74683, n61913 );
nand U141545 ( n61913, n61914, n61915 );
nand U141546 ( n61914, P2_P2_STATE_REG_2_, n73184 );
nand U141547 ( n61915, P2_P2_STATE_REG_1_, n74636 );
nand U141548 ( n13271, n60082, n60083 );
nand U141549 ( n60082, n60087, n60062 );
nand U141550 ( n60083, P2_P2_INSTQUEUEWR_ADDR_REG_2_, n60084 );
nand U141551 ( n60087, n60088, n60089 );
nand U141552 ( n6536, n26942, n26943 );
nand U141553 ( n26942, n26947, n26922 );
nand U141554 ( n26943, P1_P2_INSTQUEUEWR_ADDR_REG_2_, n26944 );
nand U141555 ( n26947, n26948, n26949 );
nand U141556 ( n4291, n34187, n34188 );
nand U141557 ( n34187, n34192, n34167 );
nand U141558 ( n34188, P1_P3_INSTQUEUEWR_ADDR_REG_2_, n34189 );
nand U141559 ( n34192, n34193, n34194 );
nand U141560 ( n11026, n68941, n68942 );
nand U141561 ( n68941, n68946, n68921 );
nand U141562 ( n68942, P2_P3_INSTQUEUEWR_ADDR_REG_2_, n68943 );
nand U141563 ( n68946, n68947, n68948 );
nand U141564 ( n34893, P1_P3_INSTQUEUE_REG_7__1_, n34883 );
nand U141565 ( n34927, P1_P3_INSTQUEUE_REG_7__5_, n34883 );
nand U141566 ( n34935, P1_P3_INSTQUEUE_REG_7__6_, n34883 );
nand U141567 ( n34943, P1_P3_INSTQUEUE_REG_7__7_, n34883 );
nand U141568 ( n34911, P1_P3_INSTQUEUE_REG_7__3_, n34883 );
nand U141569 ( n34919, P1_P3_INSTQUEUE_REG_7__4_, n34883 );
nand U141570 ( n34882, P1_P3_INSTQUEUE_REG_7__0_, n34883 );
nand U141571 ( n34901, P1_P3_INSTQUEUE_REG_7__2_, n34883 );
nand U141572 ( n69635, P2_P3_INSTQUEUE_REG_7__1_, n69625 );
nand U141573 ( n69643, P2_P3_INSTQUEUE_REG_7__2_, n69625 );
nand U141574 ( n69651, P2_P3_INSTQUEUE_REG_7__3_, n69625 );
nand U141575 ( n69675, P2_P3_INSTQUEUE_REG_7__6_, n69625 );
nand U141576 ( n69683, P2_P3_INSTQUEUE_REG_7__7_, n69625 );
nand U141577 ( n69667, P2_P3_INSTQUEUE_REG_7__5_, n69625 );
nand U141578 ( n69659, P2_P3_INSTQUEUE_REG_7__4_, n69625 );
nand U141579 ( n69624, P2_P3_INSTQUEUE_REG_7__0_, n69625 );
nand U141580 ( n30381, n30383, P1_P3_EBX_REG_1_ );
nor U141581 ( n30383, n74531, n73119 );
nand U141582 ( n23052, n23054, P1_P2_EBX_REG_1_ );
nor U141583 ( n23054, n74532, n73120 );
nand U141584 ( n64544, n64546, P2_P3_EBX_REG_1_ );
nor U141585 ( n64546, n74534, n73121 );
nand U141586 ( n56175, n56177, P2_P2_EBX_REG_1_ );
nor U141587 ( n56177, n74535, n73122 );
nand U141588 ( n43702, n43704, P2_P1_EBX_REG_1_ );
nor U141589 ( n43704, n74536, n73123 );
nor U141590 ( n46741, n46850, n46851 );
nand U141591 ( n46850, P2_P1_INSTADDRPOINTER_REG_15_, n7900 );
nand U141592 ( n9775, n9778, P1_P1_EBX_REG_1_ );
nor U141593 ( n9778, n74533, n73126 );
nor U141594 ( n13258, n13390, n13392 );
nand U141595 ( n13390, P1_P1_INSTADDRPOINTER_REG_15_, n5247 );
nand U141596 ( n16726, DIN_31_, n76928 );
xor U141597 ( n37796, n37797, n37798 );
xor U141598 ( n37798, n37799, P4_REG2_REG_5_ );
nor U141599 ( n12880, n12897, n12898 );
nand U141600 ( n12897, n12857, P1_P1_INSTADDRPOINTER_REG_25_ );
nand U141601 ( n42256, n42355, n42356 );
nand U141602 ( n42355, n42231, n42229 );
nand U141603 ( n42356, P3_REG1_REG_2_, n42357 );
or U141604 ( n42357, n42231, n42229 );
nor U141605 ( n63194, P2_P3_EBX_REG_25_, n6324 );
nor U141606 ( n29431, P1_P3_EBX_REG_25_, n3690 );
nor U141607 ( n42654, P2_P1_EBX_REG_25_, n8105 );
nor U141608 ( n22112, P1_P2_EBX_REG_25_, n4584 );
nor U141609 ( n8605, P1_P1_EBX_REG_25_, n5452 );
nor U141610 ( n55222, P2_P2_EBX_REG_25_, n7217 );
nor U141611 ( n63222, n6324, n63223 );
nor U141612 ( n63223, n63224, n75023 );
nor U141613 ( n63224, P2_P3_EBX_REG_23_, n63225 );
nor U141614 ( n29459, n3690, n29460 );
nor U141615 ( n29460, n29461, n75022 );
nor U141616 ( n29461, P1_P3_EBX_REG_23_, n29462 );
nor U141617 ( n22140, n4584, n22141 );
nor U141618 ( n22141, n22142, n75024 );
nor U141619 ( n22142, P1_P2_EBX_REG_23_, n22143 );
nor U141620 ( n55250, n7217, n55251 );
nor U141621 ( n55251, n55252, n75026 );
nor U141622 ( n55252, P2_P2_EBX_REG_23_, n55253 );
nor U141623 ( n14753, n14755, n14757 );
nor U141624 ( n14755, P1_P1_INSTQUEUERD_ADDR_REG_0_, n14759 );
nor U141625 ( n14757, n14758, n8294 );
nand U141626 ( n47577, P2_P1_INSTADDRPOINTER_REG_2_, P2_P1_INSTADDRPOINTER_REG_1_ );
nand U141627 ( n47660, n74580, n47734 );
nand U141628 ( n47734, P2_P1_INSTADDRPOINTER_REG_1_, P2_P1_INSTADDRPOINTER_REG_0_ );
nand U141629 ( n14365, n74579, n14467 );
nand U141630 ( n14467, P1_P1_INSTADDRPOINTER_REG_1_, P1_P1_INSTADDRPOINTER_REG_0_ );
nand U141631 ( n44508, n44545, n44546 );
nand U141632 ( n44546, n7817, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nor U141633 ( n44545, n44161, n44547 );
nor U141634 ( n44547, n7817, n44548 );
nand U141635 ( n10713, n10759, n10760 );
nand U141636 ( n10760, n5162, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nor U141637 ( n10759, n10297, n10762 );
nor U141638 ( n10762, n5162, n10763 );
nand U141639 ( n31129, n31166, n31167 );
nand U141640 ( n31167, n3414, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nor U141641 ( n31166, n30801, n31168 );
nor U141642 ( n31168, n3414, n31169 );
nand U141643 ( n65383, n65420, n65421 );
nand U141644 ( n65421, n6029, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nor U141645 ( n65420, n65003, n65422 );
nor U141646 ( n65422, n6029, n65423 );
nand U141647 ( n23837, n23874, n23875 );
nand U141648 ( n23875, n4252, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nor U141649 ( n23874, n23494, n23876 );
nor U141650 ( n23876, n4252, n23877 );
nand U141651 ( n56961, n56998, n56999 );
nand U141652 ( n56999, n6884, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nor U141653 ( n56998, n56616, n57000 );
nor U141654 ( n57000, n6884, n57001 );
nand U141655 ( n23824, P1_P2_ADDRESS_REG_29_, n63375 );
nand U141656 ( n63375, n63376, n63377 );
nor U141657 ( n63376, n63391, n63392 );
nor U141658 ( n63377, n63378, n63379 );
nand U141659 ( n47138, P2_P1_INSTADDRPOINTER_REG_9_, P2_P1_INSTADDRPOINTER_REG_10_ );
nand U141660 ( n5461, n29158, n29159 );
nand U141661 ( n29159, P1_P3_REQUESTPENDING_REG, n218 );
nor U141662 ( n29158, n29160, n29161 );
nor U141663 ( n29161, n218, n29162 );
nand U141664 ( n7706, n21845, n21846 );
nand U141665 ( n21846, P1_P2_REQUESTPENDING_REG, n184 );
nor U141666 ( n21845, n21847, n21848 );
nor U141667 ( n21848, n184, n21849 );
nand U141668 ( n12196, n62880, n62881 );
nand U141669 ( n62881, P2_P3_REQUESTPENDING_REG, n489 );
nor U141670 ( n62880, n62882, n62883 );
nor U141671 ( n62883, n489, n62884 );
nand U141672 ( n14441, n54936, n54937 );
nand U141673 ( n54937, P2_P2_REQUESTPENDING_REG, n455 );
nor U141674 ( n54936, n54938, n54939 );
nor U141675 ( n54939, n455, n54940 );
xor U141676 ( n68712, P2_P3_INSTADDRPOINTER_REG_2_, n68711 );
xor U141677 ( n47691, P2_P1_INSTADDRPOINTER_REG_2_, n47690 );
xor U141678 ( n26711, P1_P2_INSTADDRPOINTER_REG_2_, n26710 );
xor U141679 ( n59853, P2_P2_INSTADDRPOINTER_REG_2_, n59852 );
xor U141680 ( n33956, P1_P3_INSTADDRPOINTER_REG_2_, n33955 );
nand U141681 ( n13350, P1_P1_INSTADDRPOINTER_REG_17_, P1_P1_INSTADDRPOINTER_REG_16_ );
nand U141682 ( n16686, n42371, n42372 );
nand U141683 ( n42372, P2_P1_REQUESTPENDING_REG, n514 );
nor U141684 ( n42371, n42373, n42374 );
nor U141685 ( n42374, n514, n42375 );
nand U141686 ( n14547, P1_P1_INSTADDRPOINTER_REG_0_, n12999 );
nand U141687 ( n42246, n42341, n42342 );
nand U141688 ( n42341, n42227, n42229 );
nand U141689 ( n42342, P3_REG2_REG_2_, n42343 );
or U141690 ( n42343, n42227, n42229 );
nand U141691 ( n9951, n8280, n8282 );
nand U141692 ( n8282, P1_P1_REQUESTPENDING_REG, n243 );
nor U141693 ( n8280, n8283, n8284 );
nor U141694 ( n8284, n243, n8285 );
nor U141695 ( n60127, n60129, n60130 );
nor U141696 ( n60129, P2_P2_INSTQUEUERD_ADDR_REG_0_, n60132 );
and U141697 ( n60130, n60131, n6514 );
nor U141698 ( n26984, n26986, n26987 );
nor U141699 ( n26986, P1_P2_INSTQUEUERD_ADDR_REG_0_, n26989 );
and U141700 ( n26987, n26988, n3882 );
nor U141701 ( n34229, n34231, n34232 );
nor U141702 ( n34231, P1_P3_INSTQUEUERD_ADDR_REG_0_, n34234 );
and U141703 ( n34232, n34233, n3038 );
nor U141704 ( n68983, n68985, n68986 );
nor U141705 ( n68985, P2_P3_INSTQUEUERD_ADDR_REG_0_, n68988 );
and U141706 ( n68986, n68987, n5639 );
nor U141707 ( n47975, n47977, n47978 );
nor U141708 ( n47977, P2_P1_INSTQUEUERD_ADDR_REG_0_, n47980 );
and U141709 ( n47978, n47979, n7414 );
nand U141710 ( n63392, n63393, n63394 );
nor U141711 ( n63393, P1_P2_ADDRESS_REG_0_, n63397 );
nor U141712 ( n63394, n63395, n63396 );
nand U141713 ( n63397, n73450, n73029 );
nand U141714 ( n13158, P1_P1_INSTADDRPOINTER_REG_21_, P1_P1_INSTADDRPOINTER_REG_20_ );
nand U141715 ( n13197, P1_P1_INSTADDRPOINTER_REG_19_, n5253 );
nand U141716 ( n63391, n63398, n63399 );
nor U141717 ( n63399, n63400, n63401 );
nor U141718 ( n63398, P1_P2_ADDRESS_REG_16_, n63402 );
or U141719 ( n63400, P1_P2_ADDRESS_REG_20_, P1_P2_ADDRESS_REG_21_ );
or U141720 ( n63401, P1_P2_ADDRESS_REG_19_, P1_P2_ADDRESS_REG_1_ );
nand U141721 ( n26819, P1_P2_INSTADDRPOINTER_REG_0_, n76156 );
nand U141722 ( n59959, P2_P2_INSTADDRPOINTER_REG_0_, n76084 );
nand U141723 ( n47798, P2_P1_INSTADDRPOINTER_REG_0_, n76101 );
nand U141724 ( n34064, P1_P3_INSTADDRPOINTER_REG_0_, n76128 );
nand U141725 ( n68818, P2_P3_INSTADDRPOINTER_REG_0_, n76058 );
nor U141726 ( n67788, n67897, n67898 );
nand U141727 ( n67897, P2_P3_INSTADDRPOINTER_REG_15_, n6112 );
nor U141728 ( n25785, n25894, n25895 );
nand U141729 ( n25894, P1_P2_INSTADDRPOINTER_REG_15_, n4334 );
nor U141730 ( n58923, n59032, n59033 );
nand U141731 ( n59032, P2_P2_INSTADDRPOINTER_REG_15_, n6967 );
nor U141732 ( n33033, n33141, n33142 );
nand U141733 ( n33141, P1_P3_INSTADDRPOINTER_REG_15_, n3497 );
nand U141734 ( n63379, n63380, n63381 );
nor U141735 ( n63380, P1_P2_ADDRESS_REG_22_, n63384 );
nor U141736 ( n63381, n63382, n63383 );
or U141737 ( n63384, P1_P2_ADDRESS_REG_23_, P1_P2_ADDRESS_REG_24_ );
or U141738 ( n63383, P1_P2_ADDRESS_REG_25_, P1_P2_ADDRESS_REG_26_ );
nor U141739 ( n42707, n42708, n75021 );
nor U141740 ( n42708, P2_P1_EBX_REG_23_, n42709 );
nor U141741 ( n8642, n8643, n75025 );
nor U141742 ( n8643, P1_P1_EBX_REG_23_, n8644 );
or U141743 ( n63382, P1_P2_ADDRESS_REG_27_, P1_P2_ADDRESS_REG_28_ );
nand U141744 ( n45010, P3_REG2_REG_16_, n45007 );
nand U141745 ( n14262, P1_P1_INSTADDRPOINTER_REG_2_, P1_P1_INSTADDRPOINTER_REG_1_ );
nand U141746 ( n45018, P3_REG1_REG_16_, n45007 );
xor U141747 ( n14393, P1_P1_INSTADDRPOINTER_REG_2_, n14392 );
nand U141748 ( n33842, P1_P3_INSTADDRPOINTER_REG_2_, P1_P3_INSTADDRPOINTER_REG_1_ );
nand U141749 ( n68598, P2_P3_INSTADDRPOINTER_REG_2_, P2_P3_INSTADDRPOINTER_REG_1_ );
nand U141750 ( n26597, P1_P2_INSTADDRPOINTER_REG_2_, P1_P2_INSTADDRPOINTER_REG_1_ );
nand U141751 ( n59739, P2_P2_INSTADDRPOINTER_REG_2_, P2_P2_INSTADDRPOINTER_REG_1_ );
nor U141752 ( n32709, n32832, n32833 );
nand U141753 ( n32832, P1_P3_INSTADDRPOINTER_REG_23_, n3509 );
nor U141754 ( n67474, n67597, n67598 );
nand U141755 ( n67597, P2_P3_INSTADDRPOINTER_REG_23_, n6124 );
nor U141756 ( n25469, n25592, n25593 );
nand U141757 ( n25592, P1_P2_INSTADDRPOINTER_REG_23_, n4347 );
nor U141758 ( n58606, n58729, n58730 );
nand U141759 ( n58729, P2_P2_INSTADDRPOINTER_REG_23_, n6979 );
nand U141760 ( n68681, n74587, n68755 );
nand U141761 ( n68755, P2_P3_INSTADDRPOINTER_REG_1_, P2_P3_INSTADDRPOINTER_REG_0_ );
nand U141762 ( n33925, n74588, n33999 );
nand U141763 ( n33999, P1_P3_INSTADDRPOINTER_REG_1_, P1_P3_INSTADDRPOINTER_REG_0_ );
nand U141764 ( n26680, n74589, n26754 );
nand U141765 ( n26754, P1_P2_INSTADDRPOINTER_REG_1_, P1_P2_INSTADDRPOINTER_REG_0_ );
nand U141766 ( n59822, n74590, n59896 );
nand U141767 ( n59896, P2_P2_INSTADDRPOINTER_REG_1_, P2_P2_INSTADDRPOINTER_REG_0_ );
nor U141768 ( n56523, P2_P2_EAX_REG_24_, n56478 );
nor U141769 ( n23401, P1_P2_EAX_REG_24_, n23354 );
nor U141770 ( n64917, P2_P3_EAX_REG_24_, n64875 );
nor U141771 ( n30711, P1_P3_EAX_REG_24_, n30669 );
nor U141772 ( n45211, P3_REG1_REG_17_, n45077 );
nand U141773 ( n32878, P1_P3_INSTADDRPOINTER_REG_23_, P1_P3_INSTADDRPOINTER_REG_22_ );
nand U141774 ( n66784, P2_P3_PHYADDRPOINTER_REG_19_, P2_P3_PHYADDRPOINTER_REG_18_ );
nand U141775 ( n32138, P1_P3_PHYADDRPOINTER_REG_19_, P1_P3_PHYADDRPOINTER_REG_18_ );
nand U141776 ( n24906, P1_P2_PHYADDRPOINTER_REG_19_, P1_P2_PHYADDRPOINTER_REG_18_ );
nand U141777 ( n58043, P2_P2_PHYADDRPOINTER_REG_19_, P2_P2_PHYADDRPOINTER_REG_18_ );
nand U141778 ( n43348, n74684, n54285 );
nand U141779 ( n54285, n54286, n54287 );
nand U141780 ( n54286, P2_P1_STATE_REG_2_, n73177 );
nand U141781 ( n54287, P2_P1_STATE_REG_1_, n74650 );
nor U141782 ( n63325, n6325, n63326 );
nor U141783 ( n63326, n63327, n74980 );
nor U141784 ( n63327, P2_P3_EBX_REG_21_, n63328 );
nor U141785 ( n29496, n3692, n29497 );
nor U141786 ( n29497, n29498, n74979 );
nor U141787 ( n29498, P1_P3_EBX_REG_21_, n29499 );
nor U141788 ( n8687, n5453, n8688 );
nor U141789 ( n8688, n8689, n74981 );
nor U141790 ( n8689, P1_P1_EBX_REG_21_, n8690 );
nor U141791 ( n42747, n8107, n42748 );
nor U141792 ( n42748, n42749, n74978 );
nor U141793 ( n42749, P2_P1_EBX_REG_21_, n42750 );
nor U141794 ( n22177, n4585, n22178 );
nor U141795 ( n22178, n22179, n74982 );
nor U141796 ( n22179, P1_P2_EBX_REG_21_, n22180 );
nor U141797 ( n55291, n7218, n55292 );
nor U141798 ( n55292, n55293, n74983 );
nor U141799 ( n55293, P2_P2_EBX_REG_21_, n55294 );
nand U141800 ( n33419, P1_P3_INSTADDRPOINTER_REG_9_, P1_P3_INSTADDRPOINTER_REG_10_ );
nor U141801 ( n63243, P2_P3_EBX_REG_23_, n6325 );
nor U141802 ( n29480, P1_P3_EBX_REG_23_, n3692 );
nor U141803 ( n22161, P1_P2_EBX_REG_23_, n4585 );
nor U141804 ( n55275, P2_P2_EBX_REG_23_, n7218 );
nand U141805 ( n47011, P2_P1_INSTADDRPOINTER_REG_12_, P2_P1_INSTADDRPOINTER_REG_11_ );
nand U141806 ( n9402, n74713, n21302 );
nand U141807 ( n21302, n21303, n21304 );
nand U141808 ( n21303, P1_P1_STATE_REG_2_, n73185 );
nand U141809 ( n21304, P1_P1_STATE_REG_1_, n74670 );
nor U141810 ( n8264, n14640, P1_P1_STATE2_REG_1_ );
nand U141811 ( n14466, n54901, n54902 );
nand U141812 ( n54901, P2_P2_READREQUEST_REG, n54900 );
nand U141813 ( n54902, n54903, n6545 );
nand U141814 ( n54903, n54904, P2_P2_STATE2_REG_2_ );
nand U141815 ( n14471, n54897, n54898 );
nand U141816 ( n54897, P2_P2_MEMORYFETCH_REG, n54900 );
nand U141817 ( n54898, n54899, n6545 );
nand U141818 ( n54899, n6699, P2_P2_STATE2_REG_2_ );
nand U141819 ( n7731, n21825, n21826 );
nand U141820 ( n21825, P1_P2_READREQUEST_REG, n21824 );
nand U141821 ( n21826, n21827, n3913 );
nand U141822 ( n21827, n21828, P1_P2_STATE2_REG_2_ );
nand U141823 ( n7736, n21821, n21822 );
nand U141824 ( n21821, P1_P2_MEMORYFETCH_REG, n21824 );
nand U141825 ( n21822, n21823, n3913 );
nand U141826 ( n21823, n4067, P1_P2_STATE2_REG_2_ );
nand U141827 ( n5486, n29140, n29141 );
nand U141828 ( n29140, P1_P3_READREQUEST_REG, n29139 );
nand U141829 ( n29141, n29142, n3069 );
nand U141830 ( n29142, n29143, P1_P3_STATE2_REG_2_ );
nand U141831 ( n5491, n29136, n29137 );
nand U141832 ( n29136, P1_P3_MEMORYFETCH_REG, n29139 );
nand U141833 ( n29137, n29138, n3069 );
nand U141834 ( n29138, n3242, P1_P3_STATE2_REG_2_ );
nand U141835 ( n12221, n62807, n62808 );
nand U141836 ( n62807, P2_P3_READREQUEST_REG, n62806 );
nand U141837 ( n62808, n62809, n5670 );
nand U141838 ( n62809, n62810, P2_P3_STATE2_REG_2_ );
nand U141839 ( n12226, n62803, n62804 );
nand U141840 ( n62803, P2_P3_MEMORYFETCH_REG, n62806 );
nand U141841 ( n62804, n62805, n5670 );
nand U141842 ( n62805, n5842, P2_P3_STATE2_REG_2_ );
nand U141843 ( n26168, P1_P2_INSTADDRPOINTER_REG_9_, P1_P2_INSTADDRPOINTER_REG_10_ );
nand U141844 ( n59307, P2_P2_INSTADDRPOINTER_REG_9_, P2_P2_INSTADDRPOINTER_REG_10_ );
nand U141845 ( n46927, n46954, P2_P1_INSTADDRPOINTER_REG_15_ );
nand U141846 ( n68169, P2_P3_INSTADDRPOINTER_REG_9_, P2_P3_INSTADDRPOINTER_REG_10_ );
nor U141847 ( n26955, P1_P2_INSTQUEUEWR_ADDR_REG_0_, n26935 );
nor U141848 ( n34200, P1_P3_INSTQUEUEWR_ADDR_REG_0_, n34180 );
nor U141849 ( n60095, P2_P2_INSTQUEUEWR_ADDR_REG_0_, n60075 );
nor U141850 ( n68954, P2_P3_INSTQUEUEWR_ADDR_REG_0_, n68934 );
nand U141851 ( n16711, n42319, n42320 );
nand U141852 ( n42319, P2_P1_READREQUEST_REG, n42318 );
nand U141853 ( n42320, n42321, n7455 );
nand U141854 ( n42321, n42322, P2_P1_STATE2_REG_2_ );
nand U141855 ( n16716, n42315, n42316 );
nand U141856 ( n42315, P2_P1_MEMORYFETCH_REG, n42318 );
nand U141857 ( n42316, n42317, n7455 );
nand U141858 ( n42317, n7629, P2_P1_STATE2_REG_2_ );
nor U141859 ( n42324, n47873, P2_P1_STATE2_REG_1_ );
not U141860 ( n4813, P1_P1_STATE2_REG_3_ );
nand U141861 ( n9976, n8258, n8259 );
nand U141862 ( n8258, P1_P1_READREQUEST_REG, n8257 );
nand U141863 ( n8259, n8260, n4812 );
nand U141864 ( n8260, n8262, P1_P1_STATE2_REG_2_ );
nand U141865 ( n9981, n8253, n8254 );
nand U141866 ( n8253, P1_P1_MEMORYFETCH_REG, n8257 );
nand U141867 ( n8254, n8255, n4812 );
nand U141868 ( n8255, n4975, P1_P1_STATE2_REG_2_ );
nand U141869 ( n54249, n7799, P2_P1_INSTQUEUERD_ADDR_REG_1_ );
or U141870 ( n54250, n73497, n54197 );
nand U141871 ( n35751, n3397, P1_P3_INSTQUEUERD_ADDR_REG_1_ );
or U141872 ( n35752, n73524, n35699 );
nand U141873 ( n28572, n4234, P1_P2_INSTQUEUERD_ADDR_REG_1_ );
or U141874 ( n28573, n73503, n28520 );
nand U141875 ( n70477, n6012, P2_P3_INSTQUEUERD_ADDR_REG_1_ );
or U141876 ( n70478, n73502, n70425 );
nand U141877 ( n61877, n6867, P2_P2_INSTQUEUERD_ADDR_REG_1_ );
or U141878 ( n61878, n73504, n61825 );
nand U141879 ( n42297, n42298, n912 );
xor U141880 ( n42298, n42299, P3_REG2_REG_4_ );
nor U141881 ( n27297, P1_P2_INSTQUEUEWR_ADDR_REG_0_, n28413 );
nor U141882 ( n60440, P2_P2_INSTQUEUEWR_ADDR_REG_0_, n61722 );
nor U141883 ( n34542, P1_P3_INSTQUEUEWR_ADDR_REG_0_, n35594 );
nor U141884 ( n69290, P2_P3_INSTQUEUEWR_ADDR_REG_0_, n70322 );
and U141885 ( n9430, n21136, n21137 );
nor U141886 ( n21137, P1_P1_STATEBS16_REG, P1_P1_STATE2_REG_2_ );
nor U141887 ( n21136, P1_P1_STATE2_REG_0_, n74685 );
not U141888 ( n7457, P2_P1_STATE2_REG_3_ );
nand U141889 ( n31914, P2_P2_ADDRESS_REG_29_, n61682 );
nand U141890 ( n61682, n61683, n61684 );
nor U141891 ( n61683, n61698, n61699 );
nor U141892 ( n61684, n61685, n61686 );
xor U141893 ( n45074, n45077, P3_REG2_REG_17_ );
xor U141894 ( n45083, n45077, P3_REG1_REG_17_ );
and U141895 ( n43371, n54119, n54120 );
nor U141896 ( n54120, P2_P1_STATEBS16_REG, P2_P1_STATE2_REG_2_ );
nor U141897 ( n54119, P2_P1_STATE2_REG_0_, n74686 );
nand U141898 ( n61699, n61700, n61701 );
nor U141899 ( n61700, P2_P2_ADDRESS_REG_0_, n61704 );
nor U141900 ( n61701, n61702, n61703 );
nand U141901 ( n61704, n73063, n74266 );
nand U141902 ( n61698, n61705, n61706 );
nor U141903 ( n61706, n61707, n61708 );
nor U141904 ( n61705, P2_P2_ADDRESS_REG_16_, n61709 );
or U141905 ( n61707, P2_P2_ADDRESS_REG_20_, P2_P2_ADDRESS_REG_21_ );
nor U141906 ( n48137, n7860, P2_P1_INSTQUEUEWR_ADDR_REG_0_ );
nand U141907 ( n61686, n61687, n61688 );
nor U141908 ( n61687, P2_P2_ADDRESS_REG_22_, n61691 );
nor U141909 ( n61688, n61689, n61690 );
or U141910 ( n61691, P2_P2_ADDRESS_REG_23_, P2_P2_ADDRESS_REG_24_ );
or U141911 ( n61690, P2_P2_ADDRESS_REG_25_, P2_P2_ADDRESS_REG_26_ );
or U141912 ( n61708, P2_P2_ADDRESS_REG_19_, P2_P2_ADDRESS_REG_1_ );
nand U141913 ( n13738, P1_P1_INSTADDRPOINTER_REG_9_, P1_P1_INSTADDRPOINTER_REG_10_ );
nand U141914 ( n13052, P1_P1_INSTADDRPOINTER_REG_23_, P1_P1_INSTADDRPOINTER_REG_22_ );
or U141915 ( n61689, P2_P2_ADDRESS_REG_27_, P2_P2_ADDRESS_REG_28_ );
nand U141916 ( n42384, P2_READY11_REG, P1_P1_ADS_N_REG );
nand U141917 ( n8297, P2_P1_ADS_N_REG, P1_READY11_REG );
nand U141918 ( n9936, n8317, n8318 );
or U141919 ( n8317, n8322, n8319 );
nand U141920 ( n8318, P1_P1_FLUSH_REG, n228 );
xor U141921 ( n37968, n37969, P4_REG1_REG_17_ );
nand U141922 ( n5446, n29191, n29192 );
or U141923 ( n29191, n29195, n29193 );
nand U141924 ( n29192, P1_P3_FLUSH_REG, n202 );
nand U141925 ( n7691, n21874, n21875 );
or U141926 ( n21874, n21878, n21876 );
nand U141927 ( n21875, P1_P2_FLUSH_REG, n168 );
nand U141928 ( n12181, n62909, n62910 );
or U141929 ( n62909, n62913, n62911 );
nand U141930 ( n62910, P2_P3_FLUSH_REG, n473 );
nand U141931 ( n14426, n54965, n54966 );
or U141932 ( n54965, n54969, n54967 );
nand U141933 ( n54966, P2_P2_FLUSH_REG, n440 );
nand U141934 ( n21243, n5144, P1_P1_INSTQUEUERD_ADDR_REG_1_ );
or U141935 ( n21244, n73525, n21214 );
nor U141936 ( n23548, P1_P2_EAX_REG_22_, n23451 );
nor U141937 ( n56670, P2_P2_EAX_REG_22_, n56573 );
nor U141938 ( n65059, P2_P3_EAX_REG_22_, n64964 );
nor U141939 ( n30857, P1_P3_EAX_REG_22_, n30762 );
nand U141940 ( n16671, n42400, n42401 );
or U141941 ( n42400, n42404, n42402 );
nand U141942 ( n42401, P2_P1_FLUSH_REG, n499 );
nand U141943 ( n33287, P1_P3_INSTADDRPOINTER_REG_12_, P1_P3_INSTADDRPOINTER_REG_11_ );
nand U141944 ( n68046, P2_P3_INSTADDRPOINTER_REG_12_, P2_P3_INSTADDRPOINTER_REG_11_ );
nand U141945 ( n26043, P1_P2_INSTADDRPOINTER_REG_12_, P1_P2_INSTADDRPOINTER_REG_11_ );
nand U141946 ( n59184, P2_P2_INSTADDRPOINTER_REG_12_, P2_P2_INSTADDRPOINTER_REG_11_ );
nor U141947 ( n63361, P2_P3_EBX_REG_21_, n6327 );
nor U141948 ( n29532, P1_P3_EBX_REG_21_, n3693 );
nor U141949 ( n8732, P1_P1_EBX_REG_21_, n5454 );
nor U141950 ( n42783, P2_P1_EBX_REG_21_, n8108 );
nor U141951 ( n22213, P1_P2_EBX_REG_21_, n4587 );
nor U141952 ( n55327, P2_P2_EBX_REG_21_, n7219 );
and U141953 ( n55891, n61747, n61748 );
nor U141954 ( n61748, P2_P2_STATEBS16_REG, P2_P2_STATE2_REG_2_ );
nor U141955 ( n61747, P2_P2_STATE2_REG_0_, n73180 );
and U141956 ( n22777, n28442, n28443 );
nor U141957 ( n28443, P1_P2_STATEBS16_REG, P1_P2_STATE2_REG_2_ );
nor U141958 ( n28442, P1_P2_STATE2_REG_0_, n73181 );
and U141959 ( n30098, n35621, n35622 );
nor U141960 ( n35622, P1_P3_STATEBS16_REG, P1_P3_STATE2_REG_2_ );
nor U141961 ( n35621, P1_P3_STATE2_REG_0_, n73182 );
and U141962 ( n64115, n70347, n70348 );
nor U141963 ( n70348, P2_P3_STATEBS16_REG, P2_P3_STATE2_REG_2_ );
nor U141964 ( n70347, P2_P3_STATE2_REG_0_, n73183 );
nor U141965 ( n63463, n6327, n63464 );
nor U141966 ( n63464, n63465, n74934 );
nor U141967 ( n63465, P2_P3_EBX_REG_19_, n63466 );
nor U141968 ( n29560, n3693, n29561 );
nor U141969 ( n29561, n29562, n74933 );
nor U141970 ( n29562, P1_P3_EBX_REG_19_, n29563 );
nor U141971 ( n22243, n4587, n22244 );
nor U141972 ( n22244, n22245, n74936 );
nor U141973 ( n22245, P1_P2_EBX_REG_19_, n22246 );
nor U141974 ( n55355, n7219, n55356 );
nor U141975 ( n55356, n55357, n74937 );
nor U141976 ( n55357, P2_P2_EBX_REG_19_, n55358 );
nand U141977 ( n35728, n35729, n35730 );
nand U141978 ( n35729, n35731, n31509 );
nor U141979 ( n35731, P1_P3_INSTQUEUERD_ADDR_REG_3_, P1_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U141980 ( n28549, n28550, n28551 );
nand U141981 ( n28550, n28552, n24215 );
nor U141982 ( n28552, P1_P2_INSTQUEUERD_ADDR_REG_3_, P1_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U141983 ( n70454, n70455, n70456 );
nand U141984 ( n70455, n70457, n65759 );
nor U141985 ( n70457, P2_P3_INSTQUEUERD_ADDR_REG_3_, P2_P3_INSTQUEUERD_ADDR_REG_2_ );
nand U141986 ( n61854, n61855, n61856 );
nand U141987 ( n61855, n61857, n57337 );
nor U141988 ( n61857, P2_P2_INSTQUEUERD_ADDR_REG_3_, P2_P2_INSTQUEUERD_ADDR_REG_2_ );
nand U141989 ( n67974, n67989, P2_P3_INSTADDRPOINTER_REG_15_ );
nand U141990 ( n25971, n25986, P1_P2_INSTADDRPOINTER_REG_15_ );
nand U141991 ( n59109, n59124, P2_P2_INSTADDRPOINTER_REG_15_ );
nand U141992 ( n54226, n54227, n54228 );
nand U141993 ( n54227, n54229, n44894 );
nor U141994 ( n54229, P2_P1_INSTQUEUERD_ADDR_REG_3_, P2_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U141995 ( n33219, n33234, P1_P3_INSTADDRPOINTER_REG_15_ );
nor U141996 ( n14952, n5207, P1_P1_INSTQUEUEWR_ADDR_REG_0_ );
nand U141997 ( n66870, n66915, n6187 );
nor U141998 ( n66915, n66916, n74856 );
nand U141999 ( n24994, n25039, n4409 );
nor U142000 ( n25039, n25040, n74857 );
nand U142001 ( n58129, n58174, n7042 );
nor U142002 ( n58174, n58175, n74858 );
nand U142003 ( n32232, n32276, n3572 );
nor U142004 ( n32276, n32277, n74859 );
nand U142005 ( n70859, n70860, n76054 );
nand U142006 ( n70860, n70862, P2_P3_STATE_REG_0_ );
nor U142007 ( n70862, n70863, n74657 );
nor U142008 ( n70863, n472, n70864 );
nand U142009 ( n62478, n62479, n76239 );
nand U142010 ( n62479, n62481, P2_P2_STATE_REG_0_ );
nor U142011 ( n62481, n62482, n73184 );
nor U142012 ( n62482, n439, n62483 );
xor U142013 ( n37737, n37738, n37739 );
xor U142014 ( n37739, n37740, P4_REG2_REG_3_ );
nor U142015 ( n8768, n8769, n74935 );
nor U142016 ( n8769, P1_P1_EBX_REG_19_, n8770 );
nor U142017 ( n42812, n42813, n74932 );
nor U142018 ( n42813, P2_P1_EBX_REG_19_, n42814 );
nand U142019 ( n13578, P1_P1_INSTADDRPOINTER_REG_12_, P1_P1_INSTADDRPOINTER_REG_11_ );
nand U142020 ( n5666, n28976, n28977 );
nand U142021 ( n28977, P1_P2_STATE_REG_2_, n28978 );
nor U142022 ( n28976, n76504, n28981 );
nand U142023 ( n28978, n28979, n28980 );
xor U142024 ( n45015, n45007, P3_REG1_REG_16_ );
nand U142025 ( n14646, n54704, n54705 );
nand U142026 ( n54705, P2_P1_STATE_REG_2_, n54706 );
nor U142027 ( n54704, n76304, n54709 );
nand U142028 ( n54706, n54707, n54708 );
nand U142029 ( n13488, n13507, P1_P1_INSTADDRPOINTER_REG_15_ );
nor U142030 ( n54713, n54714, P2_P1_STATE_REG_2_ );
nor U142031 ( n54714, P2_P1_REQUESTPENDING_REG, n54715 );
nor U142032 ( n54715, n54716, n73177 );
nor U142033 ( n54716, NA, n42384 );
nor U142034 ( n21674, n21675, P1_P1_STATE_REG_2_ );
nor U142035 ( n21675, P1_P1_REQUESTPENDING_REG, n21676 );
nor U142036 ( n21676, n21677, n73185 );
nor U142037 ( n21677, NA, n8297 );
nand U142038 ( n7911, n21665, n21666 );
nand U142039 ( n21666, P1_P1_STATE_REG_2_, n21667 );
nor U142040 ( n21665, n76563, n21670 );
nand U142041 ( n21667, n21668, n21669 );
nor U142042 ( n36158, n36159, P1_P3_STATE_REG_2_ );
nor U142043 ( n36159, P1_P3_REQUESTPENDING_REG, n36160 );
nor U142044 ( n36160, n36161, n74654 );
nor U142045 ( n36161, NA, n29171 );
nand U142046 ( n3421, n36149, n36150 );
nand U142047 ( n36150, P1_P3_STATE_REG_2_, n36151 );
nor U142048 ( n36149, n2980, n36154 );
nand U142049 ( n36151, n36152, n36153 );
nor U142050 ( n28985, n28986, P1_P2_STATE_REG_2_ );
nor U142051 ( n28986, P1_P2_REQUESTPENDING_REG, n28987 );
nor U142052 ( n28987, n28988, n73179 );
nor U142053 ( n28988, NA, n21858 );
nand U142054 ( n9966, n8267, n8268 );
nand U142055 ( n8267, n8264, P1_P1_STATE2_REG_0_ );
nand U142056 ( n8268, P1_P1_CODEFETCH_REG, n8269 );
nand U142057 ( n8269, n8270, n4819 );
xor U142058 ( n44856, n44857, P3_REG2_REG_15_ );
nand U142059 ( n12228, n12283, n5320 );
nor U142060 ( n12283, n12284, n74870 );
nand U142061 ( n45919, n45964, n7975 );
nor U142062 ( n45964, n45965, n74871 );
nand U142063 ( n21228, n21229, n21230 );
nand U142064 ( n21229, n21231, n11184 );
nor U142065 ( n21231, P1_P1_INSTQUEUERD_ADDR_REG_3_, P1_P1_INSTQUEUERD_ADDR_REG_2_ );
nand U142066 ( n14446, n54932, n54933 );
nand U142067 ( n54933, P2_P2_D_C_N_REG, n76299 );
nor U142068 ( n54932, n54934, n54935 );
nor U142069 ( n54935, P2_P2_CODEFETCH_REG, n76299 );
nor U142070 ( n63478, P2_P3_EBX_REG_19_, n6328 );
nor U142071 ( n29579, P1_P3_EBX_REG_19_, n3694 );
nor U142072 ( n22258, P1_P2_EBX_REG_19_, n4588 );
nor U142073 ( n55370, P2_P2_EBX_REG_19_, n7220 );
nand U142074 ( n5476, n29147, n29148 );
nand U142075 ( n29147, n29145, P1_P3_STATE2_REG_0_ );
nand U142076 ( n29148, P1_P3_CODEFETCH_REG, n29149 );
nand U142077 ( n29149, n29150, n3077 );
nand U142078 ( n7721, n21832, n21833 );
nand U142079 ( n21832, n21830, P1_P2_STATE2_REG_0_ );
nand U142080 ( n21833, P1_P2_CODEFETCH_REG, n21834 );
nand U142081 ( n21834, n21835, n3920 );
nand U142082 ( n14456, n54925, n54926 );
nand U142083 ( n54925, n54906, P2_P2_STATE2_REG_0_ );
nand U142084 ( n54926, P2_P2_CODEFETCH_REG, n54927 );
nand U142085 ( n54927, n54928, n6553 );
nand U142086 ( n12211, n62814, n62815 );
nand U142087 ( n62814, n62812, P2_P3_STATE2_REG_0_ );
nand U142088 ( n62815, P2_P3_CODEFETCH_REG, n62816 );
nand U142089 ( n62816, n62817, n5678 );
xor U142090 ( n37944, n37941, P4_REG1_REG_15_ );
nand U142091 ( n54687, n54688, n54689 );
or U142092 ( n54689, n54690, P2_P1_STATE_REG_1_ );
nand U142093 ( n54688, n76372, n75253 );
nand U142094 ( n16691, n42367, n42368 );
nand U142095 ( n42368, P2_P1_D_C_N_REG, n76371 );
nor U142096 ( n42367, n42369, n42370 );
nor U142097 ( n42370, P2_P1_CODEFETCH_REG, n76371 );
nand U142098 ( n28959, n28960, n28961 );
or U142099 ( n28961, n28962, P1_P2_STATE_REG_1_ );
nand U142100 ( n28960, n76554, n75254 );
nand U142101 ( n5456, n29182, n29183 );
nand U142102 ( n29183, BS, n76497 );
nor U142103 ( n29182, n29156, n29185 );
nor U142104 ( n29185, n76496, n74887 );
nand U142105 ( n7711, n21839, n21840 );
nand U142106 ( n21840, P1_P2_D_C_N_REG, n76553 );
nor U142107 ( n21839, n21841, n21842 );
nor U142108 ( n21842, P1_P2_CODEFETCH_REG, n76553 );
nor U142109 ( n63504, n6328, n63505 );
nor U142110 ( n63505, n63506, n74894 );
nor U142111 ( n63506, P2_P3_EBX_REG_17_, n63507 );
nor U142112 ( n29605, n3694, n29606 );
nor U142113 ( n29606, n29607, n74893 );
nor U142114 ( n29607, P1_P3_EBX_REG_17_, n29608 );
nor U142115 ( n42852, n8109, n42853 );
nor U142116 ( n42853, n42854, n74892 );
nor U142117 ( n42854, P2_P1_EBX_REG_17_, n42855 );
nor U142118 ( n22284, n4588, n22285 );
nor U142119 ( n22285, n22286, n74896 );
nor U142120 ( n22286, P1_P2_EBX_REG_17_, n22287 );
nor U142121 ( n8818, n5455, n8819 );
nor U142122 ( n8819, n8820, n74895 );
nor U142123 ( n8820, P1_P1_EBX_REG_17_, n8822 );
nor U142124 ( n55396, n7220, n55397 );
nor U142125 ( n55397, n55398, n74897 );
nor U142126 ( n55398, P2_P2_EBX_REG_17_, n55399 );
nand U142127 ( n16701, n42360, n42361 );
nand U142128 ( n42360, n42324, P2_P1_STATE2_REG_0_ );
nand U142129 ( n42361, P2_P1_CODEFETCH_REG, n42362 );
nand U142130 ( n42362, n42363, n7463 );
nand U142131 ( n21649, n21650, n21651 );
or U142132 ( n21651, n21652, P1_P1_STATE_REG_1_ );
nand U142133 ( n21650, n76644, n75255 );
nand U142134 ( n9956, n8275, n8277 );
nand U142135 ( n8277, P1_P1_D_C_N_REG, n76643 );
nor U142136 ( n8275, n8278, n8279 );
nor U142137 ( n8279, P1_P1_CODEFETCH_REG, n76643 );
nor U142138 ( n23637, P1_P2_EAX_REG_20_, n23595 );
nor U142139 ( n56759, P2_P2_EAX_REG_20_, n56717 );
nor U142140 ( n30942, P1_P3_EAX_REG_20_, n30902 );
nor U142141 ( n65144, P2_P3_EAX_REG_20_, n65104 );
nand U142142 ( n9946, n8305, n8307 );
nand U142143 ( n8307, BS, n76640 );
nor U142144 ( n8305, n8278, n8309 );
nor U142145 ( n8309, n76639, n74906 );
nand U142146 ( n16681, n42391, n42392 );
nand U142147 ( n42392, BS, n76368 );
nor U142148 ( n42391, n42369, n42394 );
nor U142149 ( n42394, n76367, n74907 );
nand U142150 ( n7701, n21865, n21866 );
nand U142151 ( n21866, BS, n76550 );
nor U142152 ( n21865, n21841, n21868 );
nor U142153 ( n21868, n76549, n74888 );
nand U142154 ( n12191, n62900, n62901 );
nand U142155 ( n62901, BS, n76230 );
nor U142156 ( n62900, n62878, n62903 );
nor U142157 ( n62903, n76229, n74889 );
nand U142158 ( n14436, n54956, n54957 );
nand U142159 ( n54957, BS, n76296 );
nor U142160 ( n54956, n54934, n54959 );
nor U142161 ( n54959, n76295, n74890 );
nand U142162 ( n38139, n63403, n63404 );
nor U142163 ( n63403, n63407, n63408 );
nor U142164 ( n63404, n63405, n63406 );
nand U142165 ( n63408, P1_P2_W_R_N_REG, P1_P2_M_IO_N_REG );
or U142166 ( n63406, P1_P2_BE_N_REG_1_, P1_P2_BE_N_REG_2_ );
nand U142167 ( n21769, n31915, n31916 );
nor U142168 ( n31915, n31919, n31920 );
nor U142169 ( n31916, n31917, n31918 );
nand U142170 ( n31920, P2_P2_W_R_N_REG, P2_P2_M_IO_N_REG );
or U142171 ( n31918, P2_P2_BE_N_REG_1_, P2_P2_BE_N_REG_2_ );
not U142172 ( n8209, NA );
nor U142173 ( n34380, n3455, P1_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U142174 ( n27135, n4293, P1_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U142175 ( n69132, n6070, P2_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U142176 ( n60279, n6925, P2_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U142177 ( n70870, n73186, n70871 );
nand U142178 ( n70871, HOLD, n70872 );
nand U142179 ( n70872, n72927, n70873 );
nand U142180 ( n70873, n70874, n75227 );
nand U142181 ( n70874, P2_P3_STATE_REG_1_, n70875 );
nand U142182 ( n70875, n472, n8209 );
nand U142183 ( n62493, P2_P2_STATE_REG_1_, n62494 );
nand U142184 ( n62494, n439, n8209 );
nor U142185 ( n62489, n74683, n62490 );
nand U142186 ( n62490, HOLD, n62491 );
nand U142187 ( n62491, n74636, n62492 );
nand U142188 ( n62492, n62493, n75228 );
nand U142189 ( n15516, n47922, n47923 );
nand U142190 ( n47923, P2_P1_INSTQUEUEWR_ADDR_REG_2_, n47924 );
nand U142191 ( n47922, n47927, n47901 );
nand U142192 ( n47924, n47901, n47925 );
xor U142193 ( n37929, P4_REG1_REG_14_, n1972 );
or U142194 ( n63405, P1_P2_BE_N_REG_3_, P1_P2_D_C_N_REG );
or U142195 ( n31917, P2_P2_BE_N_REG_3_, P2_P2_D_C_N_REG );
xor U142196 ( n42675, n42678, P3_REG2_REG_7_ );
xor U142197 ( n42336, n42344, P3_REG2_REG_5_ );
or U142198 ( n63407, P1_P2_ADS_N_REG, P1_P2_BE_N_REG_0_ );
or U142199 ( n31919, P2_P2_ADS_N_REG, P2_P2_BE_N_REG_0_ );
xor U142200 ( n42684, n42678, P3_REG1_REG_7_ );
xor U142201 ( n42350, n42344, P3_REG1_REG_5_ );
nand U142202 ( n26954, P1_P2_STATEBS16_REG, n3912 );
nand U142203 ( n60094, P2_P2_STATEBS16_REG, n6544 );
not U142204 ( n76647, n8247 );
nand U142205 ( n8247, P2_P3_STATE_REG_1_, n73186 );
nand U142206 ( n12201, n62876, n62877 );
nand U142207 ( n62877, P2_P3_D_C_N_REG, n76646 );
nor U142208 ( n62876, n62878, n62879 );
nor U142209 ( n62879, P2_P3_CODEFETCH_REG, n76646 );
nor U142210 ( n34248, n34251, n34252 );
nor U142211 ( n34251, n73077, n34253 );
nor U142212 ( n34252, n34115, n34234 );
nand U142213 ( n34253, P1_P3_STATE2_REG_1_, n34243 );
nor U142214 ( n27003, n27006, n27007 );
nor U142215 ( n27006, n73075, n27008 );
nor U142216 ( n27007, n26870, n26989 );
nand U142217 ( n27008, P1_P2_STATE2_REG_1_, n26998 );
nor U142218 ( n69002, n69005, n69006 );
nor U142219 ( n69005, n73076, n69007 );
nor U142220 ( n69006, n68869, n68988 );
nand U142221 ( n69007, P2_P3_STATE2_REG_1_, n68997 );
nor U142222 ( n60146, n60149, n60150 );
nor U142223 ( n60149, n73074, n60151 );
nor U142224 ( n60150, n60010, n60132 );
nand U142225 ( n60151, P2_P2_STATE2_REG_1_, n60141 );
nor U142226 ( n26993, n26996, n26997 );
nor U142227 ( n26996, n26998, n26999 );
nor U142228 ( n26997, n26885, n26989 );
nand U142229 ( n26999, P1_P2_INSTADDRPOINTER_REG_0_, P1_P2_STATE2_REG_1_ );
nor U142230 ( n60136, n60139, n60140 );
nor U142231 ( n60139, n60141, n60142 );
nor U142232 ( n60140, n60025, n60132 );
nand U142233 ( n60142, P2_P2_INSTADDRPOINTER_REG_0_, P2_P2_STATE2_REG_1_ );
nor U142234 ( n34238, n34241, n34242 );
nor U142235 ( n34241, n34243, n34244 );
nor U142236 ( n34242, n34130, n34234 );
nand U142237 ( n34244, P1_P3_INSTADDRPOINTER_REG_0_, P1_P3_STATE2_REG_1_ );
nor U142238 ( n68992, n68995, n68996 );
nor U142239 ( n68995, n68997, n68998 );
nor U142240 ( n68996, n68884, n68988 );
nand U142241 ( n68998, P2_P3_INSTADDRPOINTER_REG_0_, P2_P3_STATE2_REG_1_ );
not U142242 ( n76501, n29153 );
nand U142243 ( n29153, P1_P3_STATE_REG_1_, n73192 );
nand U142244 ( n5466, n29154, n29155 );
nand U142245 ( n29155, P1_P3_D_C_N_REG, n76500 );
nor U142246 ( n29154, n29156, n29157 );
nor U142247 ( n29157, P1_P3_CODEFETCH_REG, n76500 );
nand U142248 ( n3441, n36116, n36117 );
nand U142249 ( n36116, P1_P3_DATAWIDTH_REG_1_, n76499 );
nand U142250 ( n36117, n36118, n76497 );
nand U142251 ( n36118, n8210, n29186 );
or U142252 ( n63411, n75986, P1_P1_BE_N_REG_2_ );
or U142253 ( n75986, P1_P1_D_C_N_REG, P1_P1_BE_N_REG_3_ );
or U142254 ( n31923, n75987, P2_P1_BE_N_REG_2_ );
or U142255 ( n75987, P2_P1_D_C_N_REG, P2_P1_BE_N_REG_3_ );
nand U142256 ( n14421, n54970, n54971 );
nand U142257 ( n54970, P2_P2_W_R_N_REG, n76299 );
or U142258 ( n54971, n76300, P2_P2_READREQUEST_REG );
xnor U142259 ( n43856, n43866, P3_REG2_REG_13_ );
xnor U142260 ( n43870, n43866, P3_REG1_REG_13_ );
nand U142261 ( n36162, P1_P3_STATE_REG_1_, n8209 );
nand U142262 ( n54717, P2_P1_STATE_REG_1_, n8209 );
nand U142263 ( n21678, P1_P1_STATE_REG_1_, n8209 );
nand U142264 ( n28989, P1_P2_STATE_REG_1_, n8209 );
nand U142265 ( n7931, n21633, n21634 );
nand U142266 ( n21633, P1_P1_DATAWIDTH_REG_1_, n76642 );
nand U142267 ( n21634, n21635, n76640 );
nand U142268 ( n21635, n8210, n8310 );
nand U142269 ( n36132, n36133, n36134 );
or U142270 ( n36134, n36135, P1_P3_STATE_REG_1_ );
nand U142271 ( n36133, n76500, n75256 );
nand U142272 ( n16666, n42405, n42406 );
nand U142273 ( n42405, P2_P1_W_R_N_REG, n76371 );
or U142274 ( n42406, n76372, P2_P1_READREQUEST_REG );
nand U142275 ( n14666, n54655, n54656 );
nand U142276 ( n54655, P2_P1_DATAWIDTH_REG_1_, n76370 );
nand U142277 ( n54656, n54657, n76368 );
nand U142278 ( n54657, n8210, n42395 );
nand U142279 ( n5686, n28943, n28944 );
nand U142280 ( n28943, P1_P2_DATAWIDTH_REG_1_, n76552 );
nand U142281 ( n28944, n28945, n76550 );
nand U142282 ( n28945, n8210, n21869 );
nand U142283 ( n7686, n21879, n21880 );
nand U142284 ( n21879, P1_P2_W_R_N_REG, n76553 );
or U142285 ( n21880, n76554, P1_P2_READREQUEST_REG );
nand U142286 ( n12236, n62799, n62800 );
nand U142287 ( n62800, P2_P2_BYTEENABLE_REG_2_, n76301 );
nand U142288 ( n62799, P2_P2_BE_N_REG_2_, n76300 );
nand U142289 ( n12241, n62797, n62798 );
nand U142290 ( n62798, P2_P2_BYTEENABLE_REG_1_, n76301 );
nand U142291 ( n62797, P2_P2_BE_N_REG_1_, n76300 );
nand U142292 ( n12246, n62795, n62796 );
nand U142293 ( n62796, P2_P2_BYTEENABLE_REG_0_, n76301 );
nand U142294 ( n62795, P2_P2_BE_N_REG_0_, n76300 );
nand U142295 ( n12231, n62801, n62802 );
nand U142296 ( n62802, P2_P2_BYTEENABLE_REG_3_, n76301 );
nand U142297 ( n62801, P2_P2_BE_N_REG_3_, n76299 );
nand U142298 ( n14451, n54929, n54930 );
nand U142299 ( n54930, n76301, P2_P2_MEMORYFETCH_REG );
nand U142300 ( n54929, P2_P2_M_IO_N_REG, n76299 );
nand U142301 ( n9931, n8323, n8324 );
nand U142302 ( n8323, P1_P1_W_R_N_REG, n76643 );
or U142303 ( n8324, n76644, P1_P1_READREQUEST_REG );
nor U142304 ( n29176, P1_P3_STATEBS16_REG, n29177 );
nor U142305 ( n21863, P1_P2_STATEBS16_REG, n21864 );
nor U142306 ( n62898, P2_P3_STATEBS16_REG, n62899 );
nor U142307 ( n54954, P2_P2_STATEBS16_REG, n54955 );
nor U142308 ( n42389, P2_P1_STATEBS16_REG, n42390 );
nor U142309 ( n8303, P1_P1_STATEBS16_REG, n8304 );
xor U142310 ( n37916, n37913, P4_REG1_REG_13_ );
nand U142311 ( n14481, n54893, n54894 );
nand U142312 ( n54894, P2_P1_BYTEENABLE_REG_2_, n76373 );
nand U142313 ( n54893, P2_P1_BE_N_REG_2_, n76372 );
nand U142314 ( n14486, n54891, n54892 );
nand U142315 ( n54892, P2_P1_BYTEENABLE_REG_1_, n76373 );
nand U142316 ( n54891, P2_P1_BE_N_REG_1_, n76372 );
nand U142317 ( n14491, n54889, n54890 );
nand U142318 ( n54890, P2_P1_BYTEENABLE_REG_0_, n76373 );
nand U142319 ( n54889, P2_P1_BE_N_REG_0_, n76372 );
nand U142320 ( n5501, n29132, n29133 );
nand U142321 ( n29133, P1_P2_BYTEENABLE_REG_2_, n76555 );
nand U142322 ( n29132, P1_P2_BE_N_REG_2_, n76554 );
nand U142323 ( n14476, n54895, n54896 );
nand U142324 ( n54896, P2_P1_BYTEENABLE_REG_3_, n76373 );
nand U142325 ( n54895, P2_P1_BE_N_REG_3_, n76371 );
nand U142326 ( n5506, n29130, n29131 );
nand U142327 ( n29131, P1_P2_BYTEENABLE_REG_1_, n76555 );
nand U142328 ( n29130, P1_P2_BE_N_REG_1_, n76554 );
nand U142329 ( n5511, n29124, n29125 );
nand U142330 ( n29125, P1_P2_BYTEENABLE_REG_0_, n76555 );
nand U142331 ( n29124, P1_P2_BE_N_REG_0_, n76554 );
nand U142332 ( n16696, n42364, n42365 );
nand U142333 ( n42365, n76373, P2_P1_MEMORYFETCH_REG );
nand U142334 ( n42364, P2_P1_M_IO_N_REG, n76371 );
nand U142335 ( n5496, n29134, n29135 );
nand U142336 ( n29135, P1_P2_BYTEENABLE_REG_3_, n76555 );
nand U142337 ( n29134, P1_P2_BE_N_REG_3_, n76553 );
nand U142338 ( n7716, n21836, n21837 );
nand U142339 ( n21837, n76555, P1_P2_MEMORYFETCH_REG );
nand U142340 ( n21836, P1_P2_M_IO_N_REG, n76553 );
nand U142341 ( n10176, n70836, n70837 );
nand U142342 ( n70836, P2_P3_DATAWIDTH_REG_1_, n76232 );
nand U142343 ( n70837, n70838, n76230 );
nand U142344 ( n70838, n8210, n62904 );
or U142345 ( n63414, n75988, P1_P1_ADS_N_REG );
nand U142346 ( n12421, n62399, n62400 );
nand U142347 ( n62399, P2_P2_DATAWIDTH_REG_1_, n76298 );
nand U142348 ( n62400, n62401, n76296 );
nand U142349 ( n62401, n8210, n54960 );
nand U142350 ( n7746, n21817, n21818 );
nand U142351 ( n21818, P1_P1_BYTEENABLE_REG_2_, n76645 );
nand U142352 ( n21817, P1_P1_BE_N_REG_2_, n76644 );
nand U142353 ( n7751, n21815, n21816 );
nand U142354 ( n21816, P1_P1_BYTEENABLE_REG_1_, n76645 );
nand U142355 ( n21815, P1_P1_BE_N_REG_1_, n76644 );
nand U142356 ( n7756, n21813, n21814 );
nand U142357 ( n21814, P1_P1_BYTEENABLE_REG_0_, n76645 );
nand U142358 ( n21813, P1_P1_BE_N_REG_0_, n76644 );
nand U142359 ( n7741, n21819, n21820 );
nand U142360 ( n21820, P1_P1_BYTEENABLE_REG_3_, n76645 );
nand U142361 ( n21819, P1_P1_BE_N_REG_3_, n76643 );
nand U142362 ( n9961, n8272, n8273 );
nand U142363 ( n8273, n76645, P1_P1_MEMORYFETCH_REG );
nand U142364 ( n8272, P1_P1_M_IO_N_REG, n76643 );
xor U142365 ( n37812, P4_REG1_REG_6_, n1930 );
nand U142366 ( n34199, P1_P3_STATEBS16_REG, n3068 );
nand U142367 ( n68953, P2_P3_STATEBS16_REG, n5669 );
nor U142368 ( n63560, n6329, n63561 );
nor U142369 ( n63561, n63562, n74833 );
nor U142370 ( n63562, P2_P3_EBX_REG_15_, n63563 );
nor U142371 ( n29661, n3695, n29662 );
nor U142372 ( n29662, n29663, n74832 );
nor U142373 ( n29663, P1_P3_EBX_REG_15_, n29664 );
nor U142374 ( n22340, n4589, n22341 );
nor U142375 ( n22341, n22342, n74835 );
nor U142376 ( n22342, P1_P2_EBX_REG_15_, n22343 );
nor U142377 ( n55452, n7222, n55453 );
nor U142378 ( n55453, n55454, n74836 );
nor U142379 ( n55454, P2_P2_EBX_REG_15_, n55455 );
nand U142380 ( n31927, P2_P1_W_R_N_REG, P2_P1_M_IO_N_REG );
nand U142381 ( n46788, P2_P1_INSTADDRPOINTER_REG_19_, P2_P1_INSTADDRPOINTER_REG_18_ );
xor U142382 ( n37871, P4_REG1_REG_10_, n1950 );
nand U142383 ( n70847, n70848, n70849 );
or U142384 ( n70848, n70842, n8209 );
nand U142385 ( n70849, n70850, P2_P3_STATE_REG_0_ );
nor U142386 ( n70850, n74657, n8208 );
xor U142387 ( n37882, n37883, P4_REG1_REG_11_ );
xor U142388 ( n37854, n37855, P4_REG1_REG_9_ );
xor U142389 ( n37826, n37827, P4_REG1_REG_7_ );
nand U142390 ( n62410, n62411, n62412 );
or U142391 ( n62411, n62405, n8209 );
nand U142392 ( n62412, n62413, P2_P2_STATE_REG_0_ );
nor U142393 ( n62413, n8208, n73184 );
nand U142394 ( n28954, n28955, n28956 );
or U142395 ( n28955, n28949, n8209 );
nand U142396 ( n28956, n28957, P1_P2_STATE_REG_0_ );
nor U142397 ( n28957, n8208, n73179 );
nand U142398 ( n36127, n36128, n36129 );
or U142399 ( n36128, n36122, n8209 );
nand U142400 ( n36129, n36130, P1_P3_STATE_REG_0_ );
nor U142401 ( n36130, n8208, n74654 );
nand U142402 ( n54682, n54683, n54684 );
or U142403 ( n54683, n54661, n8209 );
nand U142404 ( n54684, n54685, P2_P1_STATE_REG_0_ );
nor U142405 ( n54685, n8208, n73177 );
xor U142406 ( n43665, n43666, P3_REG2_REG_12_ );
xor U142407 ( n43558, n43559, P3_REG2_REG_11_ );
xor U142408 ( n37802, n37799, P4_REG1_REG_5_ );
xor U142409 ( n37743, n37740, P4_REG1_REG_3_ );
xor U142410 ( n43229, n43230, P3_REG2_REG_9_ );
nand U142411 ( n54690, P2_P1_STATE_REG_2_, HOLD );
nand U142412 ( n28962, P1_P2_STATE_REG_2_, HOLD );
nand U142413 ( n36135, P1_P3_STATE_REG_2_, HOLD );
xor U142414 ( n42213, n42214, n42215 );
nand U142415 ( n42215, P3_REG1_REG_0_, P3_IR_REG_0_ );
nand U142416 ( n42214, n42216, n42217 );
nand U142417 ( n42217, n917, n73825 );
nor U142418 ( n23726, P1_P2_EAX_REG_18_, n23684 );
nor U142419 ( n56848, P2_P2_EAX_REG_18_, n56806 );
nor U142420 ( n65229, P2_P3_EAX_REG_18_, n65189 );
nor U142421 ( n31027, P1_P3_EAX_REG_18_, n30987 );
nand U142422 ( n21652, HOLD, P1_P1_STATE_REG_2_ );
nand U142423 ( n8781, n14700, n14702 );
nand U142424 ( n14702, P1_P1_INSTQUEUEWR_ADDR_REG_2_, n14703 );
nand U142425 ( n14700, n14707, n14675 );
nand U142426 ( n14703, n14675, n14704 );
nand U142427 ( n10141, n70895, n70896 );
nor U142428 ( n70895, n70897, n70898 );
nand U142429 ( n70896, P2_P3_ADDRESS_REG_2_, n76646 );
nor U142430 ( n70897, n74642, n76056 );
nand U142431 ( n10101, n70927, n70928 );
nor U142432 ( n70927, n70929, n70930 );
nand U142433 ( n70928, P2_P3_ADDRESS_REG_10_, n76646 );
nor U142434 ( n70929, n74800, n76051 );
nand U142435 ( n10106, n70923, n70924 );
nor U142436 ( n70923, n70925, n70926 );
nand U142437 ( n70924, P2_P3_ADDRESS_REG_9_, n76646 );
nor U142438 ( n70925, n74790, n76052 );
nand U142439 ( n10111, n70919, n70920 );
nor U142440 ( n70919, n70921, n70922 );
nand U142441 ( n70920, P2_P3_ADDRESS_REG_8_, n76646 );
nor U142442 ( n70921, n74745, n76053 );
nand U142443 ( n10116, n70915, n70916 );
nor U142444 ( n70915, n70917, n70918 );
nand U142445 ( n70916, P2_P3_ADDRESS_REG_7_, n76646 );
nor U142446 ( n70917, n73216, n76049 );
nand U142447 ( n10121, n70911, n70912 );
nor U142448 ( n70911, n70913, n70914 );
nand U142449 ( n70912, P2_P3_ADDRESS_REG_6_, n76646 );
nor U142450 ( n70913, n74749, n76054 );
nand U142451 ( n10126, n70907, n70908 );
nor U142452 ( n70907, n70909, n70910 );
nand U142453 ( n70908, P2_P3_ADDRESS_REG_5_, n8247 );
nor U142454 ( n70909, n72966, n76056 );
nand U142455 ( n10131, n70903, n70904 );
nor U142456 ( n70903, n70905, n70906 );
nand U142457 ( n70904, P2_P3_ADDRESS_REG_4_, n76646 );
nor U142458 ( n70905, n74711, n76055 );
nand U142459 ( n10136, n70899, n70900 );
nor U142460 ( n70899, n70901, n70902 );
nand U142461 ( n70900, P2_P3_ADDRESS_REG_3_, n8247 );
nor U142462 ( n70901, n73193, n76055 );
nand U142463 ( n10146, n70891, n70892 );
nor U142464 ( n70891, n70893, n70894 );
nand U142465 ( n70892, P2_P3_ADDRESS_REG_1_, n76646 );
nor U142466 ( n70893, n73168, n76047 );
nand U142467 ( n10151, n70887, n70888 );
nor U142468 ( n70887, n70889, n70890 );
nand U142469 ( n70888, P2_P3_ADDRESS_REG_0_, n8247 );
nor U142470 ( n70889, n74621, n76048 );
xor U142471 ( n42956, n42957, P3_REG2_REG_8_ );
nand U142472 ( n9991, n8248, n8249 );
nand U142473 ( n8249, P2_P3_BYTEENABLE_REG_2_, n76647 );
nand U142474 ( n8248, P2_P3_BE_N_REG_2_, n8247 );
nand U142475 ( n10001, n70995, n70996 );
nand U142476 ( n70996, P2_P3_BYTEENABLE_REG_0_, n76647 );
nand U142477 ( n70995, P2_P3_BE_N_REG_0_, n8247 );
nand U142478 ( n12206, n62874, n62875 );
nand U142479 ( n62875, P2_P3_MEMORYFETCH_REG, n76647 );
nand U142480 ( n62874, P2_P3_M_IO_N_REG, n8247 );
nand U142481 ( n9996, n8244, n8245 );
nand U142482 ( n8245, P2_P3_BYTEENABLE_REG_1_, n76647 );
nand U142483 ( n8244, P2_P3_BE_N_REG_1_, n8247 );
nand U142484 ( n9986, n8250, n8252 );
nand U142485 ( n8252, P2_P3_BYTEENABLE_REG_3_, n76647 );
nand U142486 ( n8250, P2_P3_BE_N_REG_3_, n8247 );
nand U142487 ( n12176, n62914, n62915 );
or U142488 ( n62915, n76646, P2_P3_READREQUEST_REG );
nand U142489 ( n62914, P2_P3_W_R_N_REG, n8247 );
nand U142490 ( n3406, n36178, n36179 );
nor U142491 ( n36178, n36180, n36181 );
nand U142492 ( n36179, P1_P3_ADDRESS_REG_2_, n76500 );
nor U142493 ( n36180, n74643, n76126 );
nand U142494 ( n3351, n36224, n36225 );
nor U142495 ( n36224, n36226, n36227 );
nand U142496 ( n36225, P1_P3_ADDRESS_REG_13_, n76500 );
nor U142497 ( n36226, n74839, n76122 );
nand U142498 ( n3356, n36220, n36221 );
nor U142499 ( n36220, n36222, n36223 );
nand U142500 ( n36221, P1_P3_ADDRESS_REG_12_, n76500 );
nor U142501 ( n36222, n74829, n76123 );
nand U142502 ( n3361, n36214, n36215 );
nor U142503 ( n36214, n36216, n36217 );
nand U142504 ( n36215, P1_P3_ADDRESS_REG_11_, n76500 );
nor U142505 ( n36216, n73235, n76120 );
nand U142506 ( n3366, n36210, n36211 );
nor U142507 ( n36210, n36212, n36213 );
nand U142508 ( n36211, P1_P3_ADDRESS_REG_10_, n76500 );
nor U142509 ( n36212, n74801, n76121 );
nand U142510 ( n3371, n36206, n36207 );
nor U142511 ( n36206, n36208, n36209 );
nand U142512 ( n36207, P1_P3_ADDRESS_REG_9_, n29153 );
nor U142513 ( n36208, n74791, n76122 );
nand U142514 ( n3376, n36202, n36203 );
nor U142515 ( n36202, n36204, n36205 );
nand U142516 ( n36203, P1_P3_ADDRESS_REG_8_, n29153 );
nor U142517 ( n36204, n74746, n76123 );
nand U142518 ( n3381, n36198, n36199 );
nor U142519 ( n36198, n36200, n36201 );
nand U142520 ( n36199, P1_P3_ADDRESS_REG_7_, n76500 );
nor U142521 ( n36200, n73217, n76119 );
nand U142522 ( n3386, n36194, n36195 );
nor U142523 ( n36194, n36196, n36197 );
nand U142524 ( n36195, P1_P3_ADDRESS_REG_6_, n29153 );
nor U142525 ( n36196, n74750, n76124 );
nand U142526 ( n3391, n36190, n36191 );
nor U142527 ( n36190, n36192, n36193 );
nand U142528 ( n36191, P1_P3_ADDRESS_REG_5_, n29153 );
nor U142529 ( n36192, n72967, n76126 );
nand U142530 ( n3396, n36186, n36187 );
nor U142531 ( n36186, n36188, n36189 );
nand U142532 ( n36187, P1_P3_ADDRESS_REG_4_, n76500 );
nor U142533 ( n36188, n74712, n76125 );
nand U142534 ( n3401, n36182, n36183 );
nor U142535 ( n36182, n36184, n36185 );
nand U142536 ( n36183, P1_P3_ADDRESS_REG_3_, n29153 );
nor U142537 ( n36184, n73194, n76125 );
nand U142538 ( n3411, n36172, n36173 );
nor U142539 ( n36172, n36174, n36175 );
nand U142540 ( n36173, P1_P3_ADDRESS_REG_1_, n76500 );
nor U142541 ( n36174, n73169, n76117 );
nand U142542 ( n3416, n36168, n36169 );
nor U142543 ( n36168, n36170, n36171 );
nand U142544 ( n36169, P1_P3_ADDRESS_REG_0_, n29153 );
nor U142545 ( n36170, n74622, n76118 );
nand U142546 ( n3251, n36258, n36259 );
nand U142547 ( n36259, P1_P3_BYTEENABLE_REG_3_, n76501 );
nand U142548 ( n36258, P1_P3_BE_N_REG_3_, n29153 );
nand U142549 ( n5471, n29151, n29152 );
nand U142550 ( n29152, n76501, P1_P3_MEMORYFETCH_REG );
nand U142551 ( n29151, P1_P3_M_IO_N_REG, n29153 );
nand U142552 ( n5441, n29196, n29197 );
or U142553 ( n29197, n76500, P1_P3_READREQUEST_REG );
nand U142554 ( n29196, P1_P3_W_R_N_REG, n29153 );
nand U142555 ( n10061, n70959, n70960 );
nor U142556 ( n70959, n70961, n70962 );
nand U142557 ( n70960, P2_P3_ADDRESS_REG_18_, n76646 );
nor U142558 ( n70961, n74928, n76047 );
nand U142559 ( n10066, n70955, n70956 );
nor U142560 ( n70955, n70957, n70958 );
nand U142561 ( n70956, P2_P3_ADDRESS_REG_17_, n76646 );
nor U142562 ( n70957, n73263, n76048 );
nand U142563 ( n10071, n70951, n70952 );
nor U142564 ( n70951, n70953, n70954 );
nand U142565 ( n70952, P2_P3_ADDRESS_REG_16_, n76646 );
nor U142566 ( n70953, n74900, n76049 );
nand U142567 ( n10076, n70947, n70948 );
nor U142568 ( n70947, n70949, n70950 );
nand U142569 ( n70948, P2_P3_ADDRESS_REG_15_, n76646 );
nor U142570 ( n70949, n74884, n76050 );
nand U142571 ( n10081, n70943, n70944 );
nor U142572 ( n70943, n70945, n70946 );
nand U142573 ( n70944, P2_P3_ADDRESS_REG_14_, n76646 );
nor U142574 ( n70945, n73249, n76051 );
nand U142575 ( n10086, n70939, n70940 );
nor U142576 ( n70939, n70941, n70942 );
nand U142577 ( n70940, P2_P3_ADDRESS_REG_13_, n76646 );
nor U142578 ( n70941, n74840, n76052 );
nand U142579 ( n10091, n70935, n70936 );
nor U142580 ( n70935, n70937, n70938 );
nand U142581 ( n70936, P2_P3_ADDRESS_REG_12_, n76646 );
nor U142582 ( n70937, n74830, n76053 );
nand U142583 ( n10096, n70931, n70932 );
nor U142584 ( n70931, n70933, n70934 );
nand U142585 ( n70932, P2_P3_ADDRESS_REG_11_, n76646 );
nor U142586 ( n70933, n73236, n76050 );
nor U142587 ( n70878, n62893, n70879 );
nand U142588 ( n70879, P2_P3_STATE_REG_1_, n70880 );
nand U142589 ( n70880, n72927, n70881 );
nand U142590 ( n70881, n70882, P2_P3_REQUESTPENDING_REG );
nor U142591 ( n70882, NA, n73186 );
nor U142592 ( n62497, n54949, n62498 );
nand U142593 ( n62498, P2_P2_STATE_REG_1_, n62499 );
nand U142594 ( n62499, n74636, n62500 );
nand U142595 ( n62500, n62501, P2_P2_REQUESTPENDING_REG );
nor U142596 ( n62501, NA, n74683 );
nand U142597 ( n3326, n36244, n36245 );
nor U142598 ( n36244, n36246, n36247 );
nand U142599 ( n36245, P1_P3_ADDRESS_REG_18_, n76500 );
nor U142600 ( n36246, n74929, n76117 );
nand U142601 ( n3331, n36240, n36241 );
nor U142602 ( n36240, n36242, n36243 );
nand U142603 ( n36241, P1_P3_ADDRESS_REG_17_, n76500 );
nor U142604 ( n36242, n73264, n76118 );
nand U142605 ( n3336, n36236, n36237 );
nor U142606 ( n36236, n36238, n36239 );
nand U142607 ( n36237, P1_P3_ADDRESS_REG_16_, n76500 );
nor U142608 ( n36238, n74901, n76119 );
nand U142609 ( n3341, n36232, n36233 );
nor U142610 ( n36232, n36234, n36235 );
nand U142611 ( n36233, P1_P3_ADDRESS_REG_15_, n76500 );
nor U142612 ( n36234, n74885, n76120 );
nand U142613 ( n3346, n36228, n36229 );
nor U142614 ( n36228, n36230, n36231 );
nand U142615 ( n36229, P1_P3_ADDRESS_REG_14_, n76500 );
nor U142616 ( n36230, n73250, n76121 );
nand U142617 ( n3256, n36256, n36257 );
nand U142618 ( n36257, P1_P3_BYTEENABLE_REG_2_, n76501 );
nand U142619 ( n36256, P1_P3_BE_N_REG_2_, n76500 );
nand U142620 ( n3261, n36252, n36253 );
nand U142621 ( n36253, P1_P3_BYTEENABLE_REG_1_, n76501 );
nand U142622 ( n36252, P1_P3_BE_N_REG_1_, n76500 );
nand U142623 ( n3266, n36250, n36251 );
nand U142624 ( n36251, P1_P3_BYTEENABLE_REG_0_, n76501 );
nand U142625 ( n36250, P1_P3_BE_N_REG_0_, n76500 );
nor U142626 ( n42909, n42910, n74831 );
nor U142627 ( n42910, P2_P1_EBX_REG_15_, n42911 );
nor U142628 ( n8889, n8890, n74834 );
nor U142629 ( n8890, P1_P1_EBX_REG_15_, n8892 );
nand U142630 ( n21644, n21645, n21646 );
nand U142631 ( n21646, n21647, HOLD );
or U142632 ( n21645, n8209, n21639 );
nor U142633 ( n54699, HOLD, n498 );
nor U142634 ( n21660, HOLD, n227 );
nor U142635 ( n28971, HOLD, n167 );
nor U142636 ( n36144, HOLD, n200 );
nand U142637 ( n791, n21681, n21682 );
nor U142638 ( n21682, n21683, n21684 );
nor U142639 ( n21681, n21685, n21686 );
or U142640 ( n21683, P2_P3_D_C_N_REG, P2_P3_W_R_N_REG );
buf U142641 ( n76556, n21812 );
nor U142642 ( n21812, n21769, P2_P2_ADDRESS_REG_29_ );
nand U142643 ( n451, n32416, n32417 );
nor U142644 ( n32417, n32418, n32419 );
nor U142645 ( n32416, n32420, n32421 );
or U142646 ( n32418, P1_P3_D_C_N_REG, P1_P3_W_R_N_REG );
buf U142647 ( n76463, n33423 );
nor U142648 ( n33423, n38139, P1_P2_ADDRESS_REG_29_ );
nand U142649 ( n13313, P1_P1_INSTADDRPOINTER_REG_19_, P1_P1_INSTADDRPOINTER_REG_18_ );
nor U142650 ( n63584, P2_P3_EBX_REG_15_, n6330 );
nor U142651 ( n29685, P1_P3_EBX_REG_15_, n3697 );
nor U142652 ( n22364, P1_P2_EBX_REG_15_, n4590 );
nor U142653 ( n55476, P2_P2_EBX_REG_15_, n7223 );
nand U142654 ( n67835, P2_P3_INSTADDRPOINTER_REG_19_, P2_P3_INSTADDRPOINTER_REG_18_ );
nand U142655 ( n33079, P1_P3_INSTADDRPOINTER_REG_19_, P1_P3_INSTADDRPOINTER_REG_18_ );
nand U142656 ( n25832, P1_P2_INSTADDRPOINTER_REG_19_, P1_P2_INSTADDRPOINTER_REG_18_ );
nand U142657 ( n58970, P2_P2_INSTADDRPOINTER_REG_19_, P2_P2_INSTADDRPOINTER_REG_18_ );
nand U142658 ( n46592, P2_P1_INSTADDRPOINTER_REG_23_, P2_P1_INSTADDRPOINTER_REG_22_ );
nand U142659 ( n46734, P2_P1_INSTADDRPOINTER_REG_19_, P2_P1_INSTADDRPOINTER_REG_20_ );
nand U142660 ( n28973, P1_P2_STATE_REG_0_, n28962 );
nand U142661 ( n36146, P1_P3_STATE_REG_0_, n36135 );
nand U142662 ( n54701, P2_P1_STATE_REG_0_, n54690 );
nand U142663 ( n736, n23055, n23056 );
nand U142664 ( n23056, P2_P2_DATAO_REG_23_, n76032 );
nand U142665 ( n23055, P2_BUF2_REG_23_, n76557 );
nand U142666 ( n726, n23936, n23937 );
nand U142667 ( n23937, P2_P2_DATAO_REG_21_, n76032 );
nand U142668 ( n23936, P2_BUF2_REG_21_, n76557 );
nand U142669 ( n731, n23392, n23393 );
nand U142670 ( n23393, P2_P2_DATAO_REG_22_, n76032 );
nand U142671 ( n23392, P2_BUF2_REG_22_, n76557 );
nand U142672 ( n756, n22484, n22485 );
nand U142673 ( n22485, P2_P2_DATAO_REG_27_, n76033 );
nand U142674 ( n22484, P2_BUF2_REG_27_, n76557 );
nand U142675 ( n741, n22963, n22964 );
nand U142676 ( n22964, P2_P2_DATAO_REG_24_, n76033 );
nand U142677 ( n22963, P2_BUF2_REG_24_, n76557 );
nand U142678 ( n721, n24270, n24271 );
nand U142679 ( n24271, P2_P2_DATAO_REG_20_, n76032 );
nand U142680 ( n24270, P2_BUF2_REG_20_, n76558 );
nand U142681 ( n766, n21960, n21961 );
nand U142682 ( n21961, P2_P2_DATAO_REG_29_, n76033 );
nand U142683 ( n21960, P2_BUF2_REG_29_, n76557 );
nand U142684 ( n746, n22866, n22867 );
nand U142685 ( n22867, P2_P2_DATAO_REG_25_, n76033 );
nand U142686 ( n22866, P2_BUF2_REG_25_, n76557 );
nand U142687 ( n771, n21843, n21844 );
nand U142688 ( n21844, P2_P2_DATAO_REG_30_, n76033 );
nand U142689 ( n21843, P2_BUF2_REG_30_, n76557 );
nand U142690 ( n716, n24342, n24343 );
nand U142691 ( n24343, P2_P2_DATAO_REG_19_, n76032 );
nand U142692 ( n24342, P2_BUF2_REG_19_, n76558 );
nand U142693 ( n711, n24384, n24385 );
nand U142694 ( n24385, P2_P2_DATAO_REG_18_, n76032 );
nand U142695 ( n24384, P2_BUF2_REG_18_, n76558 );
nand U142696 ( n701, n24475, n24476 );
nand U142697 ( n24476, P2_P2_DATAO_REG_16_, n76032 );
nand U142698 ( n24475, P2_BUF2_REG_16_, n76558 );
nand U142699 ( n751, n22744, n22745 );
nand U142700 ( n22745, P2_P2_DATAO_REG_26_, n76033 );
nand U142701 ( n22744, P2_BUF2_REG_26_, n76557 );
nand U142702 ( n706, n24427, n24428 );
nand U142703 ( n24428, P2_P2_DATAO_REG_17_, n76032 );
nand U142704 ( n24427, P2_BUF2_REG_17_, n76558 );
nand U142705 ( n761, n22222, n22223 );
nand U142706 ( n22223, P2_P2_DATAO_REG_28_, n76033 );
nand U142707 ( n22222, P2_BUF2_REG_28_, n76557 );
nand U142708 ( n776, n21810, n21811 );
nand U142709 ( n21811, P2_P2_DATAO_REG_31_, n76033 );
nand U142710 ( n21810, P2_BUF2_REG_31_, n76557 );
nand U142711 ( n666, n25754, n25755 );
nand U142712 ( n25755, P2_P2_DATAO_REG_9_, n76031 );
nand U142713 ( n25754, P2_BUF2_REG_9_, n76558 );
nand U142714 ( n686, n24664, n24665 );
nand U142715 ( n24665, P2_P2_DATAO_REG_13_, n76032 );
nand U142716 ( n24664, P2_BUF2_REG_13_, n76558 );
nand U142717 ( n681, n24930, n24931 );
nand U142718 ( n24931, P2_P2_DATAO_REG_12_, n76032 );
nand U142719 ( n24930, P2_BUF2_REG_12_, n76558 );
nand U142720 ( n676, n25158, n25159 );
nand U142721 ( n25159, P2_P2_DATAO_REG_11_, n76031 );
nand U142722 ( n25158, P2_BUF2_REG_11_, n76558 );
nand U142723 ( n691, n24560, n24561 );
nand U142724 ( n24561, P2_P2_DATAO_REG_14_, n76032 );
nand U142725 ( n24560, P2_BUF2_REG_14_, n76558 );
nand U142726 ( n671, n25348, n25349 );
nand U142727 ( n25349, P2_P2_DATAO_REG_10_, n76031 );
nand U142728 ( n25348, P2_BUF2_REG_10_, n76558 );
nand U142729 ( n696, n24517, n24518 );
nand U142730 ( n24518, P2_P2_DATAO_REG_15_, n76032 );
nand U142731 ( n24517, P2_BUF2_REG_15_, n76558 );
nand U142732 ( n626, n27553, n27554 );
nand U142733 ( n27554, P2_P2_DATAO_REG_1_, n76031 );
nand U142734 ( n27553, P2_BUF2_REG_1_, n76558 );
nand U142735 ( n636, n27340, n27341 );
nand U142736 ( n27341, P2_P2_DATAO_REG_3_, n76031 );
nand U142737 ( n27340, P2_BUF2_REG_3_, n76558 );
nand U142738 ( n651, n27009, n27010 );
nand U142739 ( n27010, P2_P2_DATAO_REG_6_, n76031 );
nand U142740 ( n27009, P2_BUF2_REG_6_, n76558 );
nand U142741 ( n646, n27137, n27138 );
nand U142742 ( n27138, P2_P2_DATAO_REG_5_, n76031 );
nand U142743 ( n27137, P2_BUF2_REG_5_, n76558 );
nand U142744 ( n631, n27438, n27439 );
nand U142745 ( n27439, P2_P2_DATAO_REG_2_, n76031 );
nand U142746 ( n27438, P2_BUF2_REG_2_, n76558 );
nand U142747 ( n641, n27242, n27243 );
nand U142748 ( n27243, P2_P2_DATAO_REG_4_, n76031 );
nand U142749 ( n27242, P2_BUF2_REG_4_, n76558 );
nand U142750 ( n656, n26757, n26758 );
nand U142751 ( n26758, P2_P2_DATAO_REG_7_, n76031 );
nand U142752 ( n26757, P2_BUF2_REG_7_, n76558 );
nand U142753 ( n621, n27651, n27652 );
nand U142754 ( n27652, P2_P2_DATAO_REG_0_, n76031 );
nand U142755 ( n27651, P2_BUF2_REG_0_, n76557 );
nand U142756 ( n13247, P1_P1_INSTADDRPOINTER_REG_19_, P1_P1_INSTADDRPOINTER_REG_20_ );
nand U142757 ( n21662, P1_P1_STATE_REG_0_, n21652 );
nand U142758 ( n661, n26137, n26138 );
nand U142759 ( n26138, P2_P2_DATAO_REG_8_, n76031 );
nand U142760 ( n26137, P2_BUF2_REG_8_, n76558 );
nand U142761 ( n406, n34691, n34692 );
nand U142762 ( n34692, P1_P2_DATAO_REG_25_, n76020 );
nand U142763 ( n34691, P1_BUF2_REG_25_, n76464 );
nand U142764 ( n396, n34904, n34905 );
nand U142765 ( n34905, P1_P2_DATAO_REG_23_, n76019 );
nand U142766 ( n34904, P1_BUF2_REG_23_, n76464 );
nand U142767 ( n391, n34999, n35000 );
nand U142768 ( n35000, P1_P2_DATAO_REG_22_, n76019 );
nand U142769 ( n34999, P1_BUF2_REG_22_, n76464 );
nand U142770 ( n386, n35096, n35097 );
nand U142771 ( n35097, P1_P2_DATAO_REG_21_, n76019 );
nand U142772 ( n35096, P1_BUF2_REG_21_, n76464 );
nand U142773 ( n376, n35300, n35301 );
nand U142774 ( n35301, P1_P2_DATAO_REG_19_, n76019 );
nand U142775 ( n35300, P1_BUF2_REG_19_, n76465 );
nand U142776 ( n381, n35206, n35207 );
nand U142777 ( n35207, P1_P2_DATAO_REG_20_, n76019 );
nand U142778 ( n35206, P1_BUF2_REG_20_, n76465 );
nand U142779 ( n416, n34495, n34496 );
nand U142780 ( n34496, P1_P2_DATAO_REG_27_, n76020 );
nand U142781 ( n34495, P1_BUF2_REG_27_, n76464 );
nand U142782 ( n401, n34811, n34812 );
nand U142783 ( n34812, P1_P2_DATAO_REG_24_, n76020 );
nand U142784 ( n34811, P1_BUF2_REG_24_, n76464 );
nand U142785 ( n371, n35396, n35397 );
nand U142786 ( n35397, P1_P2_DATAO_REG_18_, n76019 );
nand U142787 ( n35396, P1_BUF2_REG_18_, n76465 );
nand U142788 ( n431, n34049, n34050 );
nand U142789 ( n34050, P1_P2_DATAO_REG_30_, n76020 );
nand U142790 ( n34049, P1_BUF2_REG_30_, n76464 );
nand U142791 ( n426, n34262, n34263 );
nand U142792 ( n34263, P1_P2_DATAO_REG_29_, n76020 );
nand U142793 ( n34262, P1_BUF2_REG_29_, n76464 );
nand U142794 ( n361, n35614, n35615 );
nand U142795 ( n35615, P1_P2_DATAO_REG_16_, n76019 );
nand U142796 ( n35614, P1_BUF2_REG_16_, n76465 );
nand U142797 ( n411, n34593, n34594 );
nand U142798 ( n34594, P1_P2_DATAO_REG_26_, n76020 );
nand U142799 ( n34593, P1_BUF2_REG_26_, n76464 );
nand U142800 ( n366, n35491, n35492 );
nand U142801 ( n35492, P1_P2_DATAO_REG_17_, n76019 );
nand U142802 ( n35491, P1_BUF2_REG_17_, n76465 );
nand U142803 ( n421, n34395, n34396 );
nand U142804 ( n34396, P1_P2_DATAO_REG_28_, n76020 );
nand U142805 ( n34395, P1_BUF2_REG_28_, n76464 );
nand U142806 ( n436, n33421, n33422 );
nand U142807 ( n33422, P1_P2_DATAO_REG_31_, n76020 );
nand U142808 ( n33421, P1_BUF2_REG_31_, n76464 );
nand U142809 ( n356, n36110, n36111 );
nand U142810 ( n36111, P1_P2_DATAO_REG_15_, n76019 );
nand U142811 ( n36110, P1_BUF2_REG_15_, n76465 );
nand U142812 ( n351, n36112, n36113 );
nand U142813 ( n36113, P1_P2_DATAO_REG_14_, n76019 );
nand U142814 ( n36112, P1_BUF2_REG_14_, n76465 );
nand U142815 ( n326, n36254, n36255 );
nand U142816 ( n36255, P1_P2_DATAO_REG_9_, n76018 );
nand U142817 ( n36254, P1_BUF2_REG_9_, n76465 );
nand U142818 ( n341, n36176, n36177 );
nand U142819 ( n36177, P1_P2_DATAO_REG_12_, n76019 );
nand U142820 ( n36176, P1_BUF2_REG_12_, n76465 );
nand U142821 ( n336, n36218, n36219 );
nand U142822 ( n36219, P1_P2_DATAO_REG_11_, n76018 );
nand U142823 ( n36218, P1_BUF2_REG_11_, n76465 );
nand U142824 ( n346, n36114, n36115 );
nand U142825 ( n36115, P1_P2_DATAO_REG_13_, n76019 );
nand U142826 ( n36114, P1_BUF2_REG_13_, n76465 );
nand U142827 ( n331, n36248, n36249 );
nand U142828 ( n36249, P1_P2_DATAO_REG_10_, n76018 );
nand U142829 ( n36248, P1_BUF2_REG_10_, n76465 );
nand U142830 ( n306, n37621, n37622 );
nand U142831 ( n37622, P1_P2_DATAO_REG_5_, n76018 );
nand U142832 ( n37621, P1_BUF2_REG_5_, n76465 );
nand U142833 ( n291, n37729, n37730 );
nand U142834 ( n37730, P1_P2_DATAO_REG_2_, n76018 );
nand U142835 ( n37729, P1_BUF2_REG_2_, n76465 );
nand U142836 ( n296, n37665, n37666 );
nand U142837 ( n37666, P1_P2_DATAO_REG_3_, n76018 );
nand U142838 ( n37665, P1_BUF2_REG_3_, n76465 );
nand U142839 ( n286, n37902, n37903 );
nand U142840 ( n37903, P1_P2_DATAO_REG_1_, n76018 );
nand U142841 ( n37902, P1_BUF2_REG_1_, n76465 );
nand U142842 ( n301, n37643, n37644 );
nand U142843 ( n37644, P1_P2_DATAO_REG_4_, n76018 );
nand U142844 ( n37643, P1_BUF2_REG_4_, n76465 );
nand U142845 ( n311, n36784, n36785 );
nand U142846 ( n36785, P1_P2_DATAO_REG_6_, n76018 );
nand U142847 ( n36784, P1_BUF2_REG_6_, n76465 );
nand U142848 ( n316, n36595, n36596 );
nand U142849 ( n36596, P1_P2_DATAO_REG_7_, n76018 );
nand U142850 ( n36595, P1_BUF2_REG_7_, n76465 );
nand U142851 ( n281, n38137, n38138 );
nand U142852 ( n38138, P1_P2_DATAO_REG_0_, n76018 );
nand U142853 ( n38137, P1_BUF2_REG_0_, n76464 );
nand U142854 ( n321, n36361, n36362 );
nand U142855 ( n36362, P1_P2_DATAO_REG_8_, n76018 );
nand U142856 ( n36361, P1_BUF2_REG_8_, n76465 );
nor U142857 ( n23815, P1_P2_EAX_REG_16_, n23773 );
nor U142858 ( n56940, P2_P2_EAX_REG_16_, n56898 );
nor U142859 ( n31112, P1_P3_EAX_REG_16_, n31072 );
nor U142860 ( n65366, P2_P3_EAX_REG_16_, n65274 );
nand U142861 ( n10118, LOGIC0, n76041 );
nand U142862 ( n47901, n47965, n47966 );
nand U142863 ( n47966, n47967, n7464 );
nor U142864 ( n47965, n47969, n76325 );
and U142865 ( n47967, n47968, P2_P1_STATE2_REG_0_ );
nor U142866 ( n47910, n47911, n73140 );
nor U142867 ( n47911, n47912, n7413 );
nor U142868 ( n47912, P2_P1_INSTQUEUEWR_ADDR_REG_0_, n7457 );
nand U142869 ( n46369, P2_P1_INSTADDRPOINTER_REG_28_, P2_P1_INSTADDRPOINTER_REG_27_ );
nand U142870 ( n48017, P2_P1_STATE2_REG_1_, P2_P1_STATE2_REG_2_ );
nand U142871 ( n14812, P1_P1_STATE2_REG_1_, P1_P1_STATE2_REG_2_ );
nand U142872 ( n15526, n47898, n47899 );
nand U142873 ( n47899, n47900, n47901 );
nor U142874 ( n47898, n47902, n47903 );
nor U142875 ( n47903, P2_P1_INSTQUEUEWR_ADDR_REG_0_, n47904 );
nand U142876 ( n14675, n14740, n14742 );
nand U142877 ( n14742, n14743, n4820 );
nor U142878 ( n14740, n14745, n76591 );
and U142879 ( n14743, n14744, P1_P1_STATE2_REG_0_ );
nor U142880 ( n14694, n14698, n73141 );
nor U142881 ( n14698, n14699, n4769 );
nor U142882 ( n14699, P1_P1_INSTQUEUEWR_ADDR_REG_0_, n4813 );
nor U142883 ( n63607, n63608, n74793 );
nor U142884 ( n63608, P2_P3_EBX_REG_13_, n63609 );
nor U142885 ( n29708, n29709, n74792 );
nor U142886 ( n29709, P1_P3_EBX_REG_13_, n29710 );
nor U142887 ( n8947, n8948, n74794 );
nor U142888 ( n8948, P1_P1_EBX_REG_13_, n8949 );
nor U142889 ( n42969, n42970, n74795 );
nor U142890 ( n42970, P2_P1_EBX_REG_13_, n42971 );
nor U142891 ( n22387, n22388, n74796 );
nor U142892 ( n22388, P1_P2_EBX_REG_13_, n22389 );
nor U142893 ( n55499, n55500, n74797 );
nor U142894 ( n55500, P2_P2_EBX_REG_13_, n55501 );
nand U142895 ( n8791, n14672, n14673 );
nand U142896 ( n14673, n14674, n14675 );
nor U142897 ( n14672, n14677, n14678 );
nor U142898 ( n14678, P1_P1_INSTQUEUEWR_ADDR_REG_0_, n14679 );
nand U142899 ( n32668, P1_P3_INSTADDRPOINTER_REG_28_, P1_P3_INSTADDRPOINTER_REG_27_ );
nand U142900 ( n25428, P1_P2_INSTADDRPOINTER_REG_28_, P1_P2_INSTADDRPOINTER_REG_27_ );
nand U142901 ( n58565, P2_P2_INSTADDRPOINTER_REG_28_, P2_P2_INSTADDRPOINTER_REG_27_ );
nand U142902 ( n67433, P2_P3_INSTADDRPOINTER_REG_28_, P2_P3_INSTADDRPOINTER_REG_27_ );
nor U142903 ( n30082, P1_P3_EBX_REG_31_, n205 );
nand U142904 ( n67781, P2_P3_INSTADDRPOINTER_REG_19_, P2_P3_INSTADDRPOINTER_REG_20_ );
nand U142905 ( n25778, P1_P2_INSTADDRPOINTER_REG_19_, P1_P2_INSTADDRPOINTER_REG_20_ );
nand U142906 ( n58916, P2_P2_INSTADDRPOINTER_REG_19_, P2_P2_INSTADDRPOINTER_REG_20_ );
nor U142907 ( n64099, P2_P3_EBX_REG_31_, n477 );
nand U142908 ( n33024, P1_P3_INSTADDRPOINTER_REG_19_, P1_P3_INSTADDRPOINTER_REG_20_ );
and U142909 ( n12839, P1_P1_INSTADDRPOINTER_REG_28_, n12857 );
not U142910 ( n8210, BS );
nand U142911 ( n67639, P2_P3_INSTADDRPOINTER_REG_23_, P2_P3_INSTADDRPOINTER_REG_22_ );
nand U142912 ( n25634, P1_P2_INSTADDRPOINTER_REG_23_, P1_P2_INSTADDRPOINTER_REG_22_ );
nand U142913 ( n58771, P2_P2_INSTADDRPOINTER_REG_23_, P2_P2_INSTADDRPOINTER_REG_22_ );
nand U142914 ( n27028, P1_P2_STATE2_REG_1_, P1_P2_STATE2_REG_2_ );
nor U142915 ( n34708, P1_P3_INSTQUEUEWR_ADDR_REG_1_, P1_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U142916 ( n27463, P1_P2_INSTQUEUEWR_ADDR_REG_1_, P1_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U142917 ( n69452, P2_P3_INSTQUEUEWR_ADDR_REG_1_, P2_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U142918 ( n60612, P2_P2_INSTQUEUEWR_ADDR_REG_1_, P2_P2_INSTQUEUEWR_ADDR_REG_0_ );
nand U142919 ( n60169, P2_P2_STATE2_REG_1_, P2_P2_STATE2_REG_2_ );
nand U142920 ( n34268, n35698, n74611 );
nand U142921 ( n35698, n35699, P1_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U142922 ( n27023, n28519, n74612 );
nand U142923 ( n28519, n28520, P1_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U142924 ( n69020, n70424, n74613 );
nand U142925 ( n70424, n70425, P2_P3_INSTQUEUERD_ADDR_REG_3_ );
nand U142926 ( n60164, n61824, n74614 );
nand U142927 ( n61824, n61825, P2_P2_INSTQUEUERD_ADDR_REG_3_ );
nand U142928 ( n48012, n54196, n74626 );
nand U142929 ( n54196, n54197, P2_P1_INSTQUEUERD_ADDR_REG_3_ );
nand U142930 ( n14805, n21213, n74646 );
nand U142931 ( n21213, n21214, P1_P1_INSTQUEUERD_ADDR_REG_3_ );
nor U142932 ( n63635, P2_P3_EBX_REG_13_, n6332 );
nor U142933 ( n29736, P1_P3_EBX_REG_13_, n3698 );
nor U142934 ( n22415, P1_P2_EBX_REG_13_, n4592 );
nor U142935 ( n55530, P2_P2_EBX_REG_13_, n7224 );
nor U142936 ( n48514, P2_P1_INSTQUEUEWR_ADDR_REG_1_, P2_P1_INSTQUEUEWR_ADDR_REG_0_ );
nand U142937 ( n10171, n70839, n70840 );
nand U142938 ( n70839, P2_P3_DATAWIDTH_REG_0_, n76232 );
nand U142939 ( n70840, n70841, n62904 );
nor U142940 ( n70841, BS, n76232 );
nand U142941 ( n12416, n62402, n62403 );
nand U142942 ( n62402, P2_P2_DATAWIDTH_REG_0_, n76298 );
nand U142943 ( n62403, n62404, n54960 );
nor U142944 ( n62404, BS, n76298 );
nand U142945 ( n14661, n54658, n54659 );
nand U142946 ( n54658, P2_P1_DATAWIDTH_REG_0_, n76370 );
nand U142947 ( n54659, n54660, n42395 );
nor U142948 ( n54660, BS, n76370 );
nand U142949 ( n7926, n21636, n21637 );
nand U142950 ( n21636, P1_P1_DATAWIDTH_REG_0_, n76642 );
nand U142951 ( n21637, n21638, n8310 );
nor U142952 ( n21638, BS, n76642 );
nand U142953 ( n5681, n28946, n28947 );
nand U142954 ( n28946, P1_P2_DATAWIDTH_REG_0_, n76552 );
nand U142955 ( n28947, n28948, n21869 );
nor U142956 ( n28948, BS, n76552 );
nand U142957 ( n3436, n36119, n36120 );
nand U142958 ( n36119, P1_P3_DATAWIDTH_REG_0_, n76499 );
nand U142959 ( n36120, n36121, n29186 );
nor U142960 ( n36121, BS, n76499 );
nand U142961 ( n46499, P2_P1_INSTADDRPOINTER_REG_25_, P2_P1_INSTADDRPOINTER_REG_24_ );
nand U142962 ( n57682, n61646, n61647 );
nand U142963 ( n61647, P2_BUF2_REG_5_, n31914 );
nand U142964 ( n61646, P2_BUF1_REG_5_, n6429 );
nand U142965 ( n57686, n61660, n61661 );
nand U142966 ( n61661, P2_BUF2_REG_6_, n31914 );
nand U142967 ( n61660, P2_BUF1_REG_6_, n6429 );
nand U142968 ( n57690, n61680, n61681 );
nand U142969 ( n61681, P2_BUF2_REG_7_, n31914 );
nand U142970 ( n61680, P2_BUF1_REG_7_, n6429 );
nand U142971 ( n57659, n61520, n61521 );
nand U142972 ( n61521, P2_BUF2_REG_0_, n31914 );
nand U142973 ( n61520, P2_BUF1_REG_0_, n6429 );
nand U142974 ( n12952, P1_P1_INSTADDRPOINTER_REG_25_, P1_P1_INSTADDRPOINTER_REG_24_ );
nand U142975 ( n24551, n28369, n28370 );
nand U142976 ( n28370, P1_BUF2_REG_5_, n23824 );
nand U142977 ( n28369, n3797, P1_BUF1_REG_5_ );
nand U142978 ( n24555, n28383, n28384 );
nand U142979 ( n28384, P1_BUF2_REG_6_, n23824 );
nand U142980 ( n28383, n3797, P1_BUF1_REG_6_ );
nand U142981 ( n24559, n28399, n28400 );
nand U142982 ( n28400, P1_BUF2_REG_7_, n23824 );
nand U142983 ( n28399, n3797, P1_BUF1_REG_7_ );
nand U142984 ( n24531, n28298, n28299 );
nand U142985 ( n28299, P1_BUF2_REG_0_, n23824 );
nand U142986 ( n28298, n3797, P1_BUF1_REG_0_ );
nand U142987 ( n12003, P1_P1_PHYADDRPOINTER_REG_22_, P1_P1_PHYADDRPOINTER_REG_21_ );
nand U142988 ( n45735, P2_P1_PHYADDRPOINTER_REG_22_, P2_P1_PHYADDRPOINTER_REG_21_ );
nand U142989 ( n66661, P2_P3_PHYADDRPOINTER_REG_22_, P2_P3_PHYADDRPOINTER_REG_21_ );
nand U142990 ( n32058, P1_P3_PHYADDRPOINTER_REG_22_, P1_P3_PHYADDRPOINTER_REG_21_ );
nand U142991 ( n24826, P1_P2_PHYADDRPOINTER_REG_22_, P1_P2_PHYADDRPOINTER_REG_21_ );
nand U142992 ( n57960, P2_P2_PHYADDRPOINTER_REG_22_, P2_P2_PHYADDRPOINTER_REG_21_ );
nand U142993 ( n47918, P2_P1_STATEBS16_REG, n7454 );
nand U142994 ( n34273, P1_P3_STATE2_REG_1_, P1_P3_STATE2_REG_2_ );
nand U142995 ( n69025, P2_P3_STATE2_REG_1_, P2_P3_STATE2_REG_2_ );
nand U142996 ( n57671, n61563, n61564 );
nand U142997 ( n61564, P2_BUF2_REG_3_, n31914 );
nand U142998 ( n61563, P2_BUF1_REG_3_, n6429 );
nand U142999 ( n57667, n61548, n61549 );
nand U143000 ( n61549, P2_BUF2_REG_2_, n31914 );
nand U143001 ( n61548, P2_BUF1_REG_2_, n6429 );
nand U143002 ( n57675, n61577, n61578 );
nand U143003 ( n61578, P2_BUF2_REG_4_, n31914 );
nand U143004 ( n61577, P2_BUF1_REG_4_, n6429 );
nand U143005 ( n57663, n61534, n61535 );
nand U143006 ( n61535, P2_BUF2_REG_1_, n31914 );
nand U143007 ( n61534, P2_BUF1_REG_1_, n6429 );
nand U143008 ( n14715, P1_P1_STATEBS16_REG, n4810 );
nor U143009 ( n63721, n63722, n74763 );
nor U143010 ( n63722, P2_P3_EBX_REG_11_, n63723 );
nor U143011 ( n29761, n29762, n74762 );
nor U143012 ( n29762, P1_P3_EBX_REG_11_, n29763 );
nor U143013 ( n9013, n9014, n74764 );
nor U143014 ( n9014, P1_P1_EBX_REG_11_, n9015 );
nor U143015 ( n43022, n43023, n74765 );
nor U143016 ( n43023, P2_P1_EBX_REG_11_, n43024 );
nor U143017 ( n22440, n22441, n74766 );
nor U143018 ( n22441, P1_P2_EBX_REG_11_, n22442 );
nor U143019 ( n55555, n55556, n74767 );
nor U143020 ( n55556, P2_P2_EBX_REG_11_, n55557 );
nand U143021 ( n24543, n28341, n28342 );
nand U143022 ( n28342, P1_BUF2_REG_3_, n23824 );
nand U143023 ( n28341, n3797, P1_BUF1_REG_3_ );
nand U143024 ( n24539, n28326, n28327 );
nand U143025 ( n28327, P1_BUF2_REG_2_, n23824 );
nand U143026 ( n28326, n3797, P1_BUF1_REG_2_ );
nand U143027 ( n24547, n28355, n28356 );
nand U143028 ( n28356, P1_BUF2_REG_4_, n23824 );
nand U143029 ( n28355, n3797, P1_BUF1_REG_4_ );
nand U143030 ( n24535, n28312, n28313 );
nand U143031 ( n28313, P1_BUF2_REG_1_, n23824 );
nand U143032 ( n28312, n3797, P1_BUF1_REG_1_ );
and U143033 ( n12778, n12782, P1_P1_INSTADDRPOINTER_REG_28_ );
nor U143034 ( n12782, n73279, n72970 );
nand U143035 ( n25557, P1_P2_INSTADDRPOINTER_REG_25_, P1_P2_INSTADDRPOINTER_REG_24_ );
nand U143036 ( n58694, P2_P2_INSTADDRPOINTER_REG_25_, P2_P2_INSTADDRPOINTER_REG_24_ );
nand U143037 ( n67562, P2_P3_INSTADDRPOINTER_REG_25_, P2_P3_INSTADDRPOINTER_REG_24_ );
nor U143038 ( n22761, P1_P2_EBX_REG_31_, n172 );
nor U143039 ( n55875, P2_P2_EBX_REG_31_, n444 );
nand U143040 ( n32797, P1_P3_INSTADDRPOINTER_REG_25_, P1_P3_INSTADDRPOINTER_REG_24_ );
nor U143041 ( n63748, P2_P3_EBX_REG_11_, n6333 );
nor U143042 ( n29788, P1_P3_EBX_REG_11_, n3699 );
nor U143043 ( n22467, P1_P2_EBX_REG_11_, n4593 );
nor U143044 ( n55582, P2_P2_EBX_REG_11_, n7225 );
nor U143045 ( n48982, P2_P1_INSTQUEUEWR_ADDR_REG_2_, n74525 );
nor U143046 ( n63778, n6333, n63779 );
nor U143047 ( n63779, n63780, n74720 );
nor U143048 ( n63780, P2_P3_EBX_REG_9_, n63781 );
nor U143049 ( n29818, n3699, n29819 );
nor U143050 ( n29819, n29820, n74719 );
nor U143051 ( n29820, P1_P3_EBX_REG_9_, n29821 );
nor U143052 ( n22499, n4593, n22500 );
nor U143053 ( n22500, n22501, n74723 );
nor U143054 ( n22501, P1_P2_EBX_REG_9_, n22502 );
nor U143055 ( n55612, n7225, n55613 );
nor U143056 ( n55613, n55614, n74724 );
nor U143057 ( n55614, P2_P2_EBX_REG_9_, n55615 );
nor U143058 ( n15915, P1_P1_INSTQUEUEWR_ADDR_REG_2_, n74538 );
nand U143059 ( n48871, n48875, n48127 );
nor U143060 ( n48875, P2_P1_INSTQUEUEWR_ADDR_REG_1_, n74525 );
nand U143061 ( n15795, n15800, n14940 );
nor U143062 ( n15800, P1_P1_INSTQUEUEWR_ADDR_REG_1_, n74538 );
nor U143063 ( n15600, P1_P1_INSTQUEUEWR_ADDR_REG_0_, n73141 );
nor U143064 ( n48320, P2_P1_INSTQUEUEWR_ADDR_REG_3_, n73140 );
nand U143065 ( n5481, n76499, n29146 );
nand U143066 ( n29146, P1_P3_ADS_N_REG, P1_P3_STATE_REG_0_ );
nor U143067 ( n15168, P1_P1_INSTQUEUEWR_ADDR_REG_3_, n73141 );
nand U143068 ( n12216, n76232, n62813 );
nand U143069 ( n62813, P2_P3_ADS_N_REG, P2_P3_STATE_REG_0_ );
nand U143070 ( n9971, n76642, n8265 );
nand U143071 ( n8265, P1_P1_ADS_N_REG, P1_P1_STATE_REG_0_ );
nand U143072 ( n16706, n76370, n42359 );
nand U143073 ( n42359, P2_P1_STATE_REG_0_, P2_P1_ADS_N_REG );
nand U143074 ( n7726, n76552, n21831 );
nand U143075 ( n21831, P1_P2_ADS_N_REG, P1_P2_STATE_REG_0_ );
nand U143076 ( n24747, P1_P2_PHYADDRPOINTER_REG_25_, P1_P2_PHYADDRPOINTER_REG_24_ );
nand U143077 ( n57881, P2_P2_PHYADDRPOINTER_REG_25_, P2_P2_PHYADDRPOINTER_REG_24_ );
nand U143078 ( n14461, n76298, n54907 );
nand U143079 ( n54907, P2_P2_ADS_N_REG, P2_P2_STATE_REG_0_ );
nand U143080 ( n66582, P2_P3_PHYADDRPOINTER_REG_25_, P2_P3_PHYADDRPOINTER_REG_24_ );
nand U143081 ( n31979, P1_P3_PHYADDRPOINTER_REG_25_, P1_P3_PHYADDRPOINTER_REG_24_ );
nor U143082 ( n43355, P2_P1_EBX_REG_31_, n503 );
nor U143083 ( n9410, P1_P1_EBX_REG_31_, n232 );
nor U143084 ( n9085, n9087, n74721 );
nor U143085 ( n9087, P1_P1_EBX_REG_9_, n9088 );
nor U143086 ( n43080, n43081, n74722 );
nor U143087 ( n43081, P2_P1_EBX_REG_9_, n43082 );
nor U143088 ( n14940, P1_P1_INSTQUEUEWR_ADDR_REG_2_, P1_P1_INSTQUEUEWR_ADDR_REG_0_ );
nand U143089 ( n45658, P2_P1_PHYADDRPOINTER_REG_25_, P2_P1_PHYADDRPOINTER_REG_24_ );
nand U143090 ( n11912, P1_P1_PHYADDRPOINTER_REG_25_, P1_P1_PHYADDRPOINTER_REG_24_ );
and U143091 ( n56272, n57724, n57725 );
nand U143092 ( n57725, P2_BUF2_REG_14_, n31914 );
nand U143093 ( n57724, P2_BUF1_REG_14_, n6429 );
and U143094 ( n56320, n57719, n57720 );
nand U143095 ( n57720, P2_BUF2_REG_13_, n31914 );
nand U143096 ( n57719, P2_BUF1_REG_13_, n6429 );
and U143097 ( n56369, n57714, n57715 );
nand U143098 ( n57715, P2_BUF2_REG_12_, n31914 );
nand U143099 ( n57714, P2_BUF1_REG_12_, n6429 );
and U143100 ( n56420, n57709, n57710 );
nand U143101 ( n57710, P2_BUF2_REG_11_, n31914 );
nand U143102 ( n57709, P2_BUF1_REG_11_, n6429 );
and U143103 ( n56468, n57704, n57705 );
nand U143104 ( n57705, P2_BUF2_REG_10_, n31914 );
nand U143105 ( n57704, P2_BUF1_REG_10_, n6429 );
and U143106 ( n56515, n57699, n57700 );
nand U143107 ( n57700, P2_BUF2_REG_9_, n31914 );
nand U143108 ( n57699, P2_BUF1_REG_9_, n6429 );
and U143109 ( n56563, n57694, n57695 );
nand U143110 ( n57695, P2_BUF2_REG_8_, n31914 );
nand U143111 ( n57694, P2_BUF1_REG_8_, n6429 );
nor U143112 ( n27875, P1_P2_INSTQUEUEWR_ADDR_REG_2_, n73136 );
nor U143113 ( n61022, P2_P2_INSTQUEUEWR_ADDR_REG_2_, n73137 );
nor U143114 ( n35114, P1_P3_INSTQUEUEWR_ADDR_REG_2_, n73138 );
nor U143115 ( n69850, P2_P3_INSTQUEUEWR_ADDR_REG_2_, n73139 );
nor U143116 ( n48127, P2_P1_INSTQUEUEWR_ADDR_REG_2_, P2_P1_INSTQUEUEWR_ADDR_REG_0_ );
and U143117 ( n23199, n24590, n24591 );
nand U143118 ( n24591, P1_BUF2_REG_13_, n23824 );
nand U143119 ( n24590, n3797, P1_BUF1_REG_13_ );
and U143120 ( n23248, n24585, n24586 );
nand U143121 ( n24586, P1_BUF2_REG_12_, n23824 );
nand U143122 ( n24585, n3797, P1_BUF1_REG_12_ );
and U143123 ( n23296, n24580, n24581 );
nand U143124 ( n24581, P1_BUF2_REG_11_, n23824 );
nand U143125 ( n24580, n3797, P1_BUF1_REG_11_ );
and U143126 ( n23151, n24595, n24596 );
nand U143127 ( n24596, P1_BUF2_REG_14_, n23824 );
nand U143128 ( n24595, n3797, P1_BUF1_REG_14_ );
and U143129 ( n23344, n24575, n24576 );
nand U143130 ( n24576, P1_BUF2_REG_10_, n23824 );
nand U143131 ( n24575, n3797, P1_BUF1_REG_10_ );
and U143132 ( n23391, n24570, n24571 );
nand U143133 ( n24571, P1_BUF2_REG_9_, n23824 );
nand U143134 ( n24570, n3797, P1_BUF1_REG_9_ );
and U143135 ( n23441, n24565, n24566 );
nand U143136 ( n24566, P1_BUF2_REG_8_, n23824 );
nand U143137 ( n24565, n3797, P1_BUF1_REG_8_ );
nor U143138 ( n63830, n6334, n63831 );
nor U143139 ( n63831, n63832, n74666 );
nor U143140 ( n63832, P2_P3_EBX_REG_7_, n63833 );
nor U143141 ( n29874, n3700, n29875 );
nor U143142 ( n29875, n29876, n74664 );
nor U143143 ( n29876, P1_P3_EBX_REG_7_, n29877 );
nor U143144 ( n22551, n4594, n22552 );
nor U143145 ( n22552, n22553, n74668 );
nor U143146 ( n22553, P1_P2_EBX_REG_7_, n22554 );
nor U143147 ( n55664, n7227, n55665 );
nor U143148 ( n55665, n55666, n74669 );
nor U143149 ( n55666, P2_P2_EBX_REG_7_, n55667 );
nor U143150 ( n60784, P2_P2_INSTQUEUEWR_ADDR_REG_0_, n74556 );
nor U143151 ( n27631, P1_P2_INSTQUEUEWR_ADDR_REG_0_, n74555 );
nor U143152 ( n69618, P2_P3_INSTQUEUEWR_ADDR_REG_0_, n74562 );
nor U143153 ( n34876, P1_P3_INSTQUEUEWR_ADDR_REG_0_, n74561 );
and U143154 ( n57006, n57740, n57741 );
nand U143155 ( n57741, P2_BUF2_REG_15_, n31914 );
nand U143156 ( n57740, P2_BUF1_REG_15_, n6429 );
or U143157 ( n10899, n10852, P1_P1_EAX_REG_13_ );
or U143158 ( n44652, n44614, P2_P1_EAX_REG_13_ );
and U143159 ( n23882, n24608, n24609 );
nand U143160 ( n24609, P1_BUF2_REG_15_, n23824 );
nand U143161 ( n24608, n3797, P1_BUF1_REG_15_ );
nor U143162 ( n27302, P1_P2_INSTQUEUEWR_ADDR_REG_3_, n74555 );
nor U143163 ( n34547, P1_P3_INSTQUEUEWR_ADDR_REG_3_, n74561 );
nor U143164 ( n69295, P2_P3_INSTQUEUEWR_ADDR_REG_3_, n74562 );
nor U143165 ( n60445, P2_P2_INSTQUEUEWR_ADDR_REG_3_, n74556 );
nor U143166 ( n15384, P1_P1_INSTQUEUEWR_ADDR_REG_1_, P1_P1_INSTQUEUEWR_ADDR_REG_0_ );
nor U143167 ( n14939, P1_P1_INSTQUEUEWR_ADDR_REG_3_, P1_P1_INSTQUEUEWR_ADDR_REG_1_ );
nor U143168 ( n15059, P1_P1_INSTQUEUEWR_ADDR_REG_3_, P1_P1_INSTQUEUEWR_ADDR_REG_2_ );
nor U143169 ( n48238, P2_P1_INSTQUEUEWR_ADDR_REG_3_, P2_P1_INSTQUEUEWR_ADDR_REG_2_ );
nand U143170 ( n12915, P1_P1_INSTADDRPOINTER_REG_26_, n72970 );
and U143171 ( n47969, n48016, P2_P1_FLUSH_REG );
nor U143172 ( n48016, n74648, n48017 );
and U143173 ( n34223, n34272, P1_P3_FLUSH_REG );
nor U143174 ( n34272, n74591, n34273 );
and U143175 ( n26978, n27027, P1_P2_FLUSH_REG );
nor U143176 ( n27027, n74592, n27028 );
and U143177 ( n14745, n14810, P1_P1_FLUSH_REG );
nor U143178 ( n14810, n74649, n14812 );
and U143179 ( n68977, n69024, P2_P3_FLUSH_REG );
nor U143180 ( n69024, n74593, n69025 );
and U143181 ( n60118, n60168, P2_P2_FLUSH_REG );
nor U143182 ( n60168, n74594, n60169 );
nor U143183 ( n27789, P1_P2_INSTQUEUEWR_ADDR_REG_1_, n73136 );
nor U143184 ( n60937, P2_P2_INSTQUEUEWR_ADDR_REG_1_, n73137 );
nor U143185 ( n35030, P1_P3_INSTQUEUEWR_ADDR_REG_1_, n73138 );
nor U143186 ( n69768, P2_P3_INSTQUEUEWR_ADDR_REG_1_, n73139 );
and U143187 ( n22001, n22004, P1_P2_REIP_REG_28_ );
nor U143188 ( n22004, n73294, n74999 );
and U143189 ( n55111, n55114, P2_P2_REIP_REG_28_ );
nor U143190 ( n55114, n73295, n75000 );
nor U143191 ( n34374, P1_P3_INSTQUEUEWR_ADDR_REG_2_, P1_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U143192 ( n69126, P2_P3_INSTQUEUEWR_ADDR_REG_2_, P2_P3_INSTQUEUEWR_ADDR_REG_0_ );
nor U143193 ( n27130, P1_P2_INSTQUEUEWR_ADDR_REG_2_, P1_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U143194 ( n60274, P2_P2_INSTQUEUEWR_ADDR_REG_2_, P2_P2_INSTQUEUEWR_ADDR_REG_0_ );
nor U143195 ( n48126, P2_P1_INSTQUEUEWR_ADDR_REG_3_, P2_P1_INSTQUEUEWR_ADDR_REG_1_ );
nor U143196 ( n9150, n9152, n74665 );
nor U143197 ( n9152, P1_P1_EBX_REG_7_, n9153 );
nor U143198 ( n43132, n43133, n74667 );
nor U143199 ( n43133, P2_P1_EBX_REG_7_, n43134 );
nand U143200 ( n68030, P2_P3_INSTADDRPOINTER_REG_13_, n74431 );
nand U143201 ( n46995, P2_P1_INSTADDRPOINTER_REG_13_, n74417 );
nand U143202 ( n26027, P1_P2_INSTADDRPOINTER_REG_13_, n74432 );
nand U143203 ( n59168, P2_P2_INSTADDRPOINTER_REG_13_, n74433 );
nand U143204 ( n33271, P1_P3_INSTADDRPOINTER_REG_13_, n73160 );
and U143205 ( n42543, n42545, P2_P1_REIP_REG_28_ );
nor U143206 ( n42545, n73308, n75014 );
and U143207 ( n8468, n8470, P1_P1_REIP_REG_28_ );
nor U143208 ( n8470, n73309, n75015 );
nand U143209 ( n13558, P1_P1_INSTADDRPOINTER_REG_13_, n73117 );
and U143210 ( n63083, n63086, P2_P3_REIP_REG_28_ );
nor U143211 ( n63086, n73296, n75003 );
and U143212 ( n29320, n29323, P1_P3_REIP_REG_28_ );
nor U143213 ( n29323, n73297, n75004 );
nand U143214 ( n11813, P1_P1_PHYADDRPOINTER_REG_28_, P1_P1_PHYADDRPOINTER_REG_27_ );
nand U143215 ( n45569, P2_P1_PHYADDRPOINTER_REG_28_, P2_P1_PHYADDRPOINTER_REG_27_ );
nor U143216 ( n12913, n72970, P1_P1_INSTADDRPOINTER_REG_26_ );
nand U143217 ( n46314, P2_P1_INSTADDRPOINTER_REG_31_, n75016 );
nand U143218 ( n66494, P2_P3_PHYADDRPOINTER_REG_28_, P2_P3_PHYADDRPOINTER_REG_27_ );
nand U143219 ( n31871, P1_P3_PHYADDRPOINTER_REG_28_, P1_P3_PHYADDRPOINTER_REG_27_ );
nand U143220 ( n24657, P1_P2_PHYADDRPOINTER_REG_28_, P1_P2_PHYADDRPOINTER_REG_27_ );
nand U143221 ( n57793, P2_P2_PHYADDRPOINTER_REG_28_, P2_P2_PHYADDRPOINTER_REG_27_ );
nor U143222 ( n63852, P2_P3_EBX_REG_7_, n6335 );
nor U143223 ( n29896, P1_P3_EBX_REG_7_, n3702 );
nor U143224 ( n22573, P1_P2_EBX_REG_7_, n4595 );
nor U143225 ( n55686, P2_P2_EBX_REG_7_, n7228 );
nor U143226 ( n47994, n47997, n47998 );
nor U143227 ( n47997, n73071, n47999 );
nor U143228 ( n47998, n47849, n47980 );
nand U143229 ( n47999, P2_P1_STATE2_REG_1_, n47989 );
nor U143230 ( n14783, n14787, n14788 );
nor U143231 ( n14787, n73079, n14789 );
nor U143232 ( n14788, n14610, n14759 );
nand U143233 ( n14789, P1_P1_STATE2_REG_1_, n14770 );
nor U143234 ( n34465, P1_P3_INSTQUEUEWR_ADDR_REG_3_, P1_P3_INSTQUEUEWR_ADDR_REG_2_ );
nor U143235 ( n69215, P2_P3_INSTQUEUEWR_ADDR_REG_3_, P2_P3_INSTQUEUEWR_ADDR_REG_2_ );
nor U143236 ( n27220, P1_P2_INSTQUEUEWR_ADDR_REG_3_, P1_P2_INSTQUEUEWR_ADDR_REG_2_ );
nor U143237 ( n60365, P2_P2_INSTQUEUEWR_ADDR_REG_3_, P2_P2_INSTQUEUEWR_ADDR_REG_2_ );
nor U143238 ( n13555, n73117, P1_P1_INSTADDRPOINTER_REG_13_ );
nor U143239 ( n27129, P1_P2_INSTQUEUEWR_ADDR_REG_3_, P1_P2_INSTQUEUEWR_ADDR_REG_1_ );
nor U143240 ( n34373, P1_P3_INSTQUEUEWR_ADDR_REG_3_, P1_P3_INSTQUEUEWR_ADDR_REG_1_ );
nor U143241 ( n69125, P2_P3_INSTQUEUEWR_ADDR_REG_3_, P2_P3_INSTQUEUEWR_ADDR_REG_1_ );
nor U143242 ( n60273, P2_P2_INSTQUEUEWR_ADDR_REG_3_, P2_P2_INSTQUEUEWR_ADDR_REG_1_ );
nand U143243 ( n32614, P1_P3_INSTADDRPOINTER_REG_31_, n75042 );
nand U143244 ( n25374, P1_P2_INSTADDRPOINTER_REG_31_, n75038 );
nand U143245 ( n67379, P2_P3_INSTADDRPOINTER_REG_31_, n75039 );
nand U143246 ( n58511, P2_P2_INSTADDRPOINTER_REG_31_, n75040 );
nor U143247 ( n33269, n73160, P1_P3_INSTADDRPOINTER_REG_13_ );
or U143248 ( n11049, n11002, P1_P1_EAX_REG_10_ );
or U143249 ( n44772, n44734, P2_P1_EAX_REG_10_ );
nor U143250 ( n68028, n74431, P2_P3_INSTADDRPOINTER_REG_13_ );
nor U143251 ( n46993, n74417, P2_P1_INSTADDRPOINTER_REG_13_ );
nor U143252 ( n26025, n74432, P1_P2_INSTADDRPOINTER_REG_13_ );
nor U143253 ( n59166, n74433, P2_P2_INSTADDRPOINTER_REG_13_ );
nand U143254 ( n36163, n200, P1_P3_REQUESTPENDING_REG );
nor U143255 ( n63877, n63878, n74603 );
nor U143256 ( n63878, P2_P3_EBX_REG_5_, n63879 );
nor U143257 ( n29921, n29922, n74601 );
nor U143258 ( n29922, P1_P3_EBX_REG_5_, n29923 );
nor U143259 ( n22598, n22599, n74605 );
nor U143260 ( n22599, P1_P2_EBX_REG_5_, n22600 );
nor U143261 ( n55711, n55712, n74606 );
nor U143262 ( n55712, P2_P2_EBX_REG_5_, n55713 );
nor U143263 ( n9208, n9209, n74602 );
nor U143264 ( n9209, P1_P1_EBX_REG_5_, n9210 );
nor U143265 ( n43178, n43179, n74604 );
nor U143266 ( n43179, P2_P1_EBX_REG_5_, n43180 );
and U143267 ( n47900, n7464, n54112 );
nand U143268 ( n54112, n47968, n75229 );
and U143269 ( n34166, n3078, n35612 );
nand U143270 ( n35612, n34222, n75230 );
and U143271 ( n26921, n3922, n28435 );
nand U143272 ( n28435, n26977, n75231 );
and U143273 ( n14674, n4820, n21129 );
nand U143274 ( n21129, n14744, n75232 );
and U143275 ( n68920, n5679, n70340 );
nand U143276 ( n70340, n68976, n75233 );
and U143277 ( n60061, n6554, n61740 );
nand U143278 ( n61740, n60117, n75234 );
nand U143279 ( n35603, n35627, n200 );
nor U143280 ( n35627, P1_P3_STATE2_REG_2_, n74591 );
nand U143281 ( n42442, n42449, n7354 );
nor U143282 ( n42449, P2_P1_REIP_REG_1_, P2_P1_DATAWIDTH_REG_1_ );
nand U143283 ( n21893, n21900, n3833 );
nor U143284 ( n21900, P1_P2_REIP_REG_1_, P1_P2_DATAWIDTH_REG_1_ );
nand U143285 ( n8340, n8349, n4720 );
nor U143286 ( n8349, P1_P1_REIP_REG_1_, P1_P1_DATAWIDTH_REG_1_ );
nand U143287 ( n55005, n55012, n6465 );
nor U143288 ( n55012, P2_P2_REIP_REG_1_, P2_P2_DATAWIDTH_REG_1_ );
nand U143289 ( n29210, n29217, n2989 );
nor U143290 ( n29217, P1_P3_REIP_REG_1_, P1_P3_DATAWIDTH_REG_1_ );
nand U143291 ( n62928, n62984, n5590 );
nor U143292 ( n62984, P2_P3_REIP_REG_1_, P2_P3_DATAWIDTH_REG_1_ );
nor U143293 ( n62927, P2_P3_DATAWIDTH_REG_0_, n62928 );
nor U143294 ( n29209, P1_P3_DATAWIDTH_REG_0_, n29210 );
nor U143295 ( n42441, P2_P1_DATAWIDTH_REG_0_, n42442 );
nor U143296 ( n21892, P1_P2_DATAWIDTH_REG_0_, n21893 );
nor U143297 ( n55004, P2_P2_DATAWIDTH_REG_0_, n55005 );
nor U143298 ( n8339, P1_P1_DATAWIDTH_REG_0_, n8340 );
and U143299 ( n63009, P2_P3_DATAWIDTH_REG_0_, P2_P3_DATAWIDTH_REG_1_ );
and U143300 ( n29242, P1_P3_DATAWIDTH_REG_0_, P1_P3_DATAWIDTH_REG_1_ );
and U143301 ( n42474, P2_P1_DATAWIDTH_REG_0_, P2_P1_DATAWIDTH_REG_1_ );
and U143302 ( n21925, P1_P2_DATAWIDTH_REG_0_, P1_P2_DATAWIDTH_REG_1_ );
and U143303 ( n55037, P2_P2_DATAWIDTH_REG_0_, P2_P2_DATAWIDTH_REG_1_ );
and U143304 ( n8380, P1_P1_DATAWIDTH_REG_0_, P1_P1_DATAWIDTH_REG_1_ );
nand U143305 ( n12161, n62924, n62925 );
nor U143306 ( n62924, n62931, n62932 );
nor U143307 ( n62925, n62926, n62927 );
and U143308 ( n62932, n62918, P2_P3_BYTEENABLE_REG_2_ );
nand U143309 ( n5426, n29206, n29207 );
nor U143310 ( n29206, n29213, n29214 );
nor U143311 ( n29207, n29208, n29209 );
and U143312 ( n29214, n29200, P1_P3_BYTEENABLE_REG_2_ );
nand U143313 ( n16651, n42438, n42439 );
nor U143314 ( n42438, n42445, n42446 );
nor U143315 ( n42439, n42440, n42441 );
and U143316 ( n42446, n42409, P2_P1_BYTEENABLE_REG_2_ );
nand U143317 ( n7671, n21889, n21890 );
nor U143318 ( n21889, n21896, n21897 );
nor U143319 ( n21890, n21891, n21892 );
and U143320 ( n21897, n21883, P1_P2_BYTEENABLE_REG_2_ );
nand U143321 ( n14406, n55001, n55002 );
nor U143322 ( n55001, n55008, n55009 );
nor U143323 ( n55002, n55003, n55004 );
and U143324 ( n55009, n54974, P2_P2_BYTEENABLE_REG_2_ );
nand U143325 ( n9916, n8335, n8337 );
nor U143326 ( n8335, n8344, n8345 );
nor U143327 ( n8337, n8338, n8339 );
and U143328 ( n8345, n8328, P1_P1_BYTEENABLE_REG_2_ );
nand U143329 ( n70331, n70353, n472 );
nor U143330 ( n70353, P2_P3_STATE2_REG_2_, n74593 );
nor U143331 ( n63905, P2_P3_EBX_REG_5_, n6337 );
nor U143332 ( n29949, P1_P3_EBX_REG_5_, n3703 );
nor U143333 ( n22626, P1_P2_EBX_REG_5_, n4597 );
nor U143334 ( n55739, P2_P2_EBX_REG_5_, n7229 );
nand U143335 ( n35632, n35633, P1_P3_STATE2_REG_0_ );
nor U143336 ( n35633, P1_P3_STATE2_REG_2_, n200 );
nor U143337 ( n63926, n6337, n63927 );
nor U143338 ( n63927, n63928, n74570 );
nor U143339 ( n63928, P2_P3_EBX_REG_3_, n63929 );
nor U143340 ( n29970, n3703, n29971 );
nor U143341 ( n29971, n29972, n74568 );
nor U143342 ( n29972, P1_P3_EBX_REG_3_, n29973 );
nor U143343 ( n9269, n5464, n9270 );
nor U143344 ( n9270, n9272, n74569 );
nor U143345 ( n9272, P1_P1_EBX_REG_3_, n9273 );
nor U143346 ( n43241, n8118, n43242 );
nor U143347 ( n43242, n43243, n74571 );
nor U143348 ( n43243, P2_P1_EBX_REG_3_, n43244 );
nor U143349 ( n22647, n4597, n22648 );
nor U143350 ( n22648, n22649, n74572 );
nor U143351 ( n22649, P1_P2_EBX_REG_3_, n22650 );
nor U143352 ( n55760, n7229, n55761 );
nor U143353 ( n55761, n55762, n74573 );
nor U143354 ( n55762, P2_P2_EBX_REG_3_, n55763 );
and U143355 ( n62931, P2_P3_REIP_REG_0_, n62919 );
and U143356 ( n29213, P1_P3_REIP_REG_0_, n29201 );
and U143357 ( n42445, P2_P1_REIP_REG_0_, n42410 );
and U143358 ( n21896, P1_P2_REIP_REG_0_, n21884 );
and U143359 ( n55008, P2_P2_REIP_REG_0_, n54975 );
and U143360 ( n8344, P1_P1_REIP_REG_0_, n8329 );
nand U143361 ( n33180, P1_P3_INSTADDRPOINTER_REG_15_, P1_P3_INSTADDRPOINTER_REG_16_ );
nand U143362 ( n13439, P1_P1_INSTADDRPOINTER_REG_15_, P1_P1_INSTADDRPOINTER_REG_16_ );
nor U143363 ( n62926, n62929, n62930 );
nand U143364 ( n62929, n75257, n73163 );
nand U143365 ( n62930, n5590, P2_P3_DATAWIDTH_REG_0_ );
nor U143366 ( n29208, n29211, n29212 );
nand U143367 ( n29211, n75258, n73164 );
nand U143368 ( n29212, n2989, P1_P3_DATAWIDTH_REG_0_ );
nor U143369 ( n42440, n42443, n42444 );
nand U143370 ( n42443, n75259, n72962 );
nand U143371 ( n42444, n7354, P2_P1_DATAWIDTH_REG_0_ );
nor U143372 ( n21891, n21894, n21895 );
nand U143373 ( n21894, n75260, n72958 );
nand U143374 ( n21895, n3833, P1_P2_DATAWIDTH_REG_0_ );
nor U143375 ( n55003, n55006, n55007 );
nand U143376 ( n55006, n75261, n72959 );
nand U143377 ( n55007, n6465, P2_P2_DATAWIDTH_REG_0_ );
nor U143378 ( n8338, n8342, n8343 );
nand U143379 ( n8342, n75262, n72963 );
nand U143380 ( n8343, n4720, P1_P1_DATAWIDTH_REG_0_ );
nand U143381 ( n70358, n70359, P2_P3_STATE2_REG_0_ );
nor U143382 ( n70359, P2_P3_STATE2_REG_2_, n472 );
nand U143383 ( n16646, n42447, n42448 );
nand U143384 ( n42448, P2_P1_BYTEENABLE_REG_3_, n42409 );
nor U143385 ( n42447, n42437, n7353 );
not U143386 ( n7353, n42442 );
nand U143387 ( n7666, n21898, n21899 );
nand U143388 ( n21899, P1_P2_BYTEENABLE_REG_3_, n21883 );
nor U143389 ( n21898, n21888, n3832 );
not U143390 ( n3832, n21893 );
nand U143391 ( n9911, n8347, n8348 );
nand U143392 ( n8348, P1_P1_BYTEENABLE_REG_3_, n8328 );
nor U143393 ( n8347, n8334, n4719 );
not U143394 ( n4719, n8340 );
nand U143395 ( n14401, n55010, n55011 );
nand U143396 ( n55011, P2_P2_BYTEENABLE_REG_3_, n54974 );
nor U143397 ( n55010, n54979, n6464 );
not U143398 ( n6464, n55005 );
nand U143399 ( n5421, n29215, n29216 );
nand U143400 ( n29216, P1_P3_BYTEENABLE_REG_3_, n29200 );
nor U143401 ( n29215, n29205, n2988 );
not U143402 ( n2988, n29210 );
nand U143403 ( n12156, n62982, n62983 );
nand U143404 ( n62983, P2_P3_BYTEENABLE_REG_3_, n62918 );
nor U143405 ( n62982, n62923, n5589 );
not U143406 ( n5589, n62928 );
nor U143407 ( n47984, n47987, n47988 );
nor U143408 ( n47987, n47989, n47990 );
nor U143409 ( n47988, n47864, n47980 );
nand U143410 ( n47990, P2_P1_INSTADDRPOINTER_REG_0_, P2_P1_STATE2_REG_1_ );
nor U143411 ( n14764, n14768, n14769 );
nor U143412 ( n14768, n14770, n14772 );
nor U143413 ( n14769, n14629, n14759 );
nand U143414 ( n14772, P1_P1_INSTADDRPOINTER_REG_0_, P1_P1_STATE2_REG_1_ );
and U143415 ( n42437, n42450, n42451 );
nor U143416 ( n42451, P2_P1_REIP_REG_0_, P2_P1_DATAWIDTH_REG_1_ );
nor U143417 ( n42450, P2_P1_DATAWIDTH_REG_0_, n42409 );
and U143418 ( n21888, n21901, n21902 );
nor U143419 ( n21902, P1_P2_REIP_REG_0_, P1_P2_DATAWIDTH_REG_1_ );
nor U143420 ( n21901, P1_P2_DATAWIDTH_REG_0_, n21883 );
and U143421 ( n8334, n8350, n8352 );
nor U143422 ( n8352, P1_P1_REIP_REG_0_, P1_P1_DATAWIDTH_REG_1_ );
nor U143423 ( n8350, P1_P1_DATAWIDTH_REG_0_, n8328 );
and U143424 ( n54979, n55013, n55014 );
nor U143425 ( n55014, P2_P2_REIP_REG_0_, P2_P2_DATAWIDTH_REG_1_ );
nor U143426 ( n55013, P2_P2_DATAWIDTH_REG_0_, n54974 );
and U143427 ( n29205, n29218, n29219 );
nor U143428 ( n29219, P1_P3_REIP_REG_0_, P1_P3_DATAWIDTH_REG_1_ );
nor U143429 ( n29218, P1_P3_DATAWIDTH_REG_0_, n29200 );
and U143430 ( n62923, n62985, n62986 );
nor U143431 ( n62986, P2_P3_REIP_REG_0_, P2_P3_DATAWIDTH_REG_1_ );
nor U143432 ( n62985, P2_P3_DATAWIDTH_REG_0_, n62918 );
nand U143433 ( n12166, n62921, n62922 );
nand U143434 ( n62922, P2_P3_BYTEENABLE_REG_1_, n62918 );
nor U143435 ( n62921, n62923, n62919 );
nand U143436 ( n5431, n29203, n29204 );
nand U143437 ( n29204, P1_P3_BYTEENABLE_REG_1_, n29200 );
nor U143438 ( n29203, n29205, n29201 );
nand U143439 ( n16656, n42435, n42436 );
nand U143440 ( n42436, P2_P1_BYTEENABLE_REG_1_, n42409 );
nor U143441 ( n42435, n42437, n42410 );
nand U143442 ( n7676, n21886, n21887 );
nand U143443 ( n21887, P1_P2_BYTEENABLE_REG_1_, n21883 );
nor U143444 ( n21886, n21888, n21884 );
nand U143445 ( n14411, n54977, n54978 );
nand U143446 ( n54978, P2_P2_BYTEENABLE_REG_1_, n54974 );
nor U143447 ( n54977, n54979, n54975 );
nand U143448 ( n9921, n8332, n8333 );
nand U143449 ( n8333, P1_P1_BYTEENABLE_REG_1_, n8328 );
nor U143450 ( n8332, n8334, n8329 );
or U143451 ( n11220, n11152, P1_P1_EAX_REG_7_ );
or U143452 ( n44923, n44868, P2_P1_EAX_REG_7_ );
nand U143453 ( n54718, n498, P2_P1_REQUESTPENDING_REG );
nand U143454 ( n21679, n227, P1_P1_REQUESTPENDING_REG );
nand U143455 ( n54103, n54125, n498 );
nor U143456 ( n54125, P2_P1_STATE2_REG_2_, n74648 );
nand U143457 ( n21120, n21142, n227 );
nor U143458 ( n21142, P1_P1_STATE2_REG_2_, n74649 );
nand U143459 ( n28426, n28448, n167 );
nor U143460 ( n28448, P1_P2_STATE2_REG_2_, n74592 );
nand U143461 ( n61731, n61753, n439 );
nor U143462 ( n61753, P2_P2_STATE2_REG_2_, n74594 );
nand U143463 ( n12171, n62916, n62917 );
nand U143464 ( n62917, P2_P3_BYTEENABLE_REG_0_, n62918 );
nor U143465 ( n62916, n62919, n62920 );
nor U143466 ( n62920, n62918, n75257 );
nand U143467 ( n5436, n29198, n29199 );
nand U143468 ( n29199, P1_P3_BYTEENABLE_REG_0_, n29200 );
nor U143469 ( n29198, n29201, n29202 );
nor U143470 ( n29202, n29200, n75258 );
nand U143471 ( n16661, n42407, n42408 );
nand U143472 ( n42408, P2_P1_BYTEENABLE_REG_0_, n42409 );
nor U143473 ( n42407, n42410, n42411 );
nor U143474 ( n42411, n42409, n75259 );
nand U143475 ( n7681, n21881, n21882 );
nand U143476 ( n21882, P1_P2_BYTEENABLE_REG_0_, n21883 );
nor U143477 ( n21881, n21884, n21885 );
nor U143478 ( n21885, n21883, n75260 );
nand U143479 ( n14416, n54972, n54973 );
nand U143480 ( n54973, P2_P2_BYTEENABLE_REG_0_, n54974 );
nor U143481 ( n54972, n54975, n54976 );
nor U143482 ( n54976, n54974, n75261 );
nand U143483 ( n9926, n8325, n8327 );
nand U143484 ( n8327, P1_P1_BYTEENABLE_REG_0_, n8328 );
nor U143485 ( n8325, n8329, n8330 );
nor U143486 ( n8330, n8328, n75262 );
nand U143487 ( n28990, n167, P1_P2_REQUESTPENDING_REG );
nor U143488 ( n63966, P2_P3_EBX_REG_3_, n6338 );
nor U143489 ( n30010, P1_P3_EBX_REG_3_, n3704 );
nor U143490 ( n22687, P1_P2_EBX_REG_3_, n4598 );
nor U143491 ( n55803, P2_P2_EBX_REG_3_, n7230 );
xor U143492 ( n26998, P1_P2_INSTADDRPOINTER_REG_31_, P1_P2_INSTADDRPOINTER_REG_1_ );
xor U143493 ( n60141, P2_P2_INSTADDRPOINTER_REG_31_, P2_P2_INSTADDRPOINTER_REG_1_ );
xor U143494 ( n47989, P2_P1_INSTADDRPOINTER_REG_31_, P2_P1_INSTADDRPOINTER_REG_1_ );
xor U143495 ( n34243, P1_P3_INSTADDRPOINTER_REG_31_, P1_P3_INSTADDRPOINTER_REG_1_ );
xor U143496 ( n14770, P1_P1_INSTADDRPOINTER_REG_31_, P1_P1_INSTADDRPOINTER_REG_1_ );
xor U143497 ( n68997, P2_P3_INSTADDRPOINTER_REG_31_, P2_P3_INSTADDRPOINTER_REG_1_ );
nand U143498 ( n54130, n54131, P2_P1_STATE2_REG_0_ );
nor U143499 ( n54131, P2_P1_STATE2_REG_2_, n498 );
nand U143500 ( n21147, n21148, P1_P1_STATE2_REG_0_ );
nor U143501 ( n21148, P1_P1_STATE2_REG_2_, n227 );
nor U143502 ( n64046, n64047, n74534 );
nor U143503 ( n64047, P2_P3_EBX_REG_1_, P2_P3_EBX_REG_0_ );
nor U143504 ( n30029, n30030, n74531 );
nor U143505 ( n30030, P1_P3_EBX_REG_1_, P1_P3_EBX_REG_0_ );
nor U143506 ( n9343, n9344, n74533 );
nor U143507 ( n9344, P1_P1_EBX_REG_1_, P1_P1_EBX_REG_0_ );
nor U143508 ( n43300, n43301, n74536 );
nor U143509 ( n43301, P2_P1_EBX_REG_1_, P2_P1_EBX_REG_0_ );
nor U143510 ( n22706, n22707, n74532 );
nor U143511 ( n22707, P1_P2_EBX_REG_1_, P1_P2_EBX_REG_0_ );
nor U143512 ( n55822, n55823, n74535 );
nor U143513 ( n55823, P2_P2_EBX_REG_1_, P2_P2_EBX_REG_0_ );
or U143514 ( n44953, n44945, P2_P1_EAX_REG_4_ );
or U143515 ( n11264, n11254, P1_P1_EAX_REG_4_ );
nand U143516 ( n28453, n28454, P1_P2_STATE2_REG_0_ );
nor U143517 ( n28454, P1_P2_STATE2_REG_2_, n167 );
nand U143518 ( n61758, n61759, P2_P2_STATE2_REG_0_ );
nor U143519 ( n61759, P2_P2_STATE2_REG_2_, n439 );
nand U143520 ( n54129, P2_P1_STATEBS16_REG, n74648 );
nand U143521 ( n35631, P1_P3_STATEBS16_REG, n74591 );
nand U143522 ( n28452, P1_P2_STATEBS16_REG, n74592 );
nand U143523 ( n21146, P1_P1_STATEBS16_REG, n74649 );
nand U143524 ( n70357, P2_P3_STATEBS16_REG, n74593 );
nand U143525 ( n61757, P2_P2_STATEBS16_REG, n74594 );
nor U143526 ( n29156, n29186, P1_P3_STATE_REG_0_ );
nor U143527 ( n21841, P1_P2_STATE_REG_0_, n21869 );
nor U143528 ( n8278, n8310, P1_P1_STATE_REG_0_ );
nor U143529 ( n42369, n42395, P2_P1_STATE_REG_0_ );
nor U143530 ( n54934, P2_P2_STATE_REG_0_, n54960 );
nor U143531 ( n62878, n62904, P2_P3_STATE_REG_0_ );
nand U143532 ( n60128, P2_P2_STATE2_REG_1_, n73074 );
nand U143533 ( n26985, P1_P2_STATE2_REG_1_, n73075 );
nand U143534 ( n34230, P1_P3_STATE2_REG_1_, n73077 );
nand U143535 ( n68984, P2_P3_STATE2_REG_1_, n73076 );
nand U143536 ( n47976, P2_P1_STATE2_REG_1_, n73071 );
nand U143537 ( n14754, P1_P1_STATE2_REG_1_, n73079 );
nand U143538 ( n30321, P1_P3_EBX_REG_9_, n74719 );
nand U143539 ( n64440, P2_P3_EBX_REG_9_, n74720 );
nand U143540 ( n9697, P1_P1_EBX_REG_9_, n74721 );
nand U143541 ( n43628, P2_P1_EBX_REG_9_, n74722 );
nand U143542 ( n43501, P2_P1_EBX_REG_21_, n74978 );
nand U143543 ( n43520, P2_P1_EBX_REG_19_, n74932 );
nand U143544 ( n43539, P2_P1_EBX_REG_17_, n74892 );
nand U143545 ( n43571, P2_P1_EBX_REG_15_, n74831 );
nand U143546 ( n30199, P1_P3_EBX_REG_21_, n74979 );
nand U143547 ( n30222, P1_P3_EBX_REG_19_, n74933 );
nand U143548 ( n30241, P1_P3_EBX_REG_17_, n74893 );
nand U143549 ( n30260, P1_P3_EBX_REG_15_, n74832 );
nand U143550 ( n30279, P1_P3_EBX_REG_13_, n74792 );
nand U143551 ( n30298, P1_P3_EBX_REG_11_, n74762 );
nand U143552 ( n64265, P2_P3_EBX_REG_21_, n74980 );
nand U143553 ( n64284, P2_P3_EBX_REG_19_, n74934 );
nand U143554 ( n64303, P2_P3_EBX_REG_17_, n74894 );
nand U143555 ( n64322, P2_P3_EBX_REG_15_, n74833 );
nand U143556 ( n64402, P2_P3_EBX_REG_13_, n74793 );
nand U143557 ( n64421, P2_P3_EBX_REG_11_, n74763 );
nand U143558 ( n30340, P1_P3_EBX_REG_7_, n74664 );
nand U143559 ( n30357, P1_P3_EBX_REG_5_, n74601 );
nand U143560 ( n30374, P1_P3_EBX_REG_3_, n74568 );
nand U143561 ( n9552, P1_P1_EBX_REG_21_, n74981 );
nand U143562 ( n9575, P1_P1_EBX_REG_19_, n74935 );
nand U143563 ( n9598, P1_P1_EBX_REG_17_, n74895 );
nand U143564 ( n9645, P1_P1_EBX_REG_13_, n74794 );
nand U143565 ( n9673, P1_P1_EBX_REG_11_, n74764 );
nand U143566 ( n9720, P1_P1_EBX_REG_7_, n74665 );
nand U143567 ( n9742, P1_P1_EBX_REG_5_, n74602 );
nand U143568 ( n9763, P1_P1_EBX_REG_3_, n74569 );
nand U143569 ( n64459, P2_P3_EBX_REG_7_, n74666 );
nand U143570 ( n64476, P2_P3_EBX_REG_5_, n74603 );
nand U143571 ( n64537, P2_P3_EBX_REG_3_, n74570 );
nand U143572 ( n43590, P2_P1_EBX_REG_13_, n74795 );
nand U143573 ( n43609, P2_P1_EBX_REG_11_, n74765 );
nand U143574 ( n43647, P2_P1_EBX_REG_7_, n74667 );
nand U143575 ( n43678, P2_P1_EBX_REG_5_, n74604 );
nand U143576 ( n43695, P2_P1_EBX_REG_3_, n74571 );
nand U143577 ( n9622, P1_P1_EBX_REG_15_, n74834 );
nand U143578 ( n22992, P1_P2_EBX_REG_9_, n74723 );
nand U143579 ( n56108, P2_P2_EBX_REG_9_, n74724 );
nand U143580 ( n43463, P2_P1_EBX_REG_25_, n75071 );
nand U143581 ( n43482, P2_P1_EBX_REG_23_, n75021 );
nand U143582 ( n30161, P1_P3_EBX_REG_25_, n75072 );
nand U143583 ( n30180, P1_P3_EBX_REG_23_, n75022 );
nand U143584 ( n64174, P2_P3_EBX_REG_25_, n75073 );
nand U143585 ( n64246, P2_P3_EBX_REG_23_, n75023 );
nand U143586 ( n22836, P1_P2_EBX_REG_25_, n75074 );
nand U143587 ( n22855, P1_P2_EBX_REG_23_, n75024 );
nand U143588 ( n22876, P1_P2_EBX_REG_21_, n74982 );
nand U143589 ( n22895, P1_P2_EBX_REG_19_, n74936 );
nand U143590 ( n22914, P1_P2_EBX_REG_17_, n74896 );
nand U143591 ( n22933, P1_P2_EBX_REG_15_, n74835 );
nand U143592 ( n22952, P1_P2_EBX_REG_13_, n74796 );
nand U143593 ( n22973, P1_P2_EBX_REG_11_, n74766 );
nand U143594 ( n23011, P1_P2_EBX_REG_7_, n74668 );
nand U143595 ( n23028, P1_P2_EBX_REG_5_, n74605 );
nand U143596 ( n23045, P1_P2_EBX_REG_3_, n74572 );
nand U143597 ( n9504, P1_P1_EBX_REG_25_, n75075 );
nand U143598 ( n9528, P1_P1_EBX_REG_23_, n75025 );
nand U143599 ( n55950, P2_P2_EBX_REG_25_, n75076 );
nand U143600 ( n55972, P2_P2_EBX_REG_23_, n75026 );
nand U143601 ( n55991, P2_P2_EBX_REG_21_, n74983 );
nand U143602 ( n56010, P2_P2_EBX_REG_19_, n74937 );
nand U143603 ( n56029, P2_P2_EBX_REG_17_, n74897 );
nand U143604 ( n56048, P2_P2_EBX_REG_15_, n74836 );
nand U143605 ( n56070, P2_P2_EBX_REG_13_, n74797 );
nand U143606 ( n56089, P2_P2_EBX_REG_11_, n74767 );
nand U143607 ( n56127, P2_P2_EBX_REG_7_, n74669 );
nand U143608 ( n56144, P2_P2_EBX_REG_5_, n74606 );
nand U143609 ( n56164, P2_P2_EBX_REG_3_, n74573 );
nand U143610 ( n43405, P2_P1_EBX_REG_28_, n75190 );
nand U143611 ( n30136, P1_P3_EBX_REG_28_, n75181 );
nand U143612 ( n64149, P2_P3_EBX_REG_28_, n75182 );
nand U143613 ( n22811, P1_P2_EBX_REG_28_, n75183 );
nand U143614 ( n9473, P1_P1_EBX_REG_28_, n75189 );
nand U143615 ( n55925, P2_P2_EBX_REG_28_, n75184 );
nand U143616 ( n30391, P1_P3_EBX_REG_0_, n74531 );
nand U143617 ( n23064, P1_P2_EBX_REG_0_, n74532 );
nand U143618 ( n9788, P1_P1_EBX_REG_0_, n74533 );
nand U143619 ( n64554, P2_P3_EBX_REG_0_, n74534 );
nand U143620 ( n56185, P2_P2_EBX_REG_0_, n74535 );
nand U143621 ( n43712, P2_P1_EBX_REG_0_, n74536 );
nand U143622 ( n11300, P1_P1_EAX_REG_0_, n74608 );
nand U143623 ( n44982, P2_P1_EAX_REG_0_, n74609 );
nand U143624 ( n10953, P1_P1_EAX_REG_11_, n74802 );
nand U143625 ( n11103, P1_P1_EAX_REG_8_, n74756 );
nand U143626 ( n11280, P1_P1_EAX_REG_2_, n74630 );
nand U143627 ( n44695, P2_P1_EAX_REG_11_, n74803 );
nand U143628 ( n44815, P2_P1_EAX_REG_8_, n74757 );
nand U143629 ( n44936, P2_P1_EAX_REG_5_, n74704 );
nand U143630 ( n44966, P2_P1_EAX_REG_2_, n74631 );
nand U143631 ( n10780, P1_P1_EAX_REG_14_, n74864 );
nand U143632 ( n11237, P1_P1_EAX_REG_5_, n74705 );
nand U143633 ( n44557, P2_P1_EAX_REG_14_, n74865 );
nor U143634 ( n30111, P1_P3_EBX_REG_31_, n75213 );
nor U143635 ( n64124, P2_P3_EBX_REG_31_, n75214 );
nor U143636 ( n22786, P1_P2_EBX_REG_31_, n75215 );
nor U143637 ( n55900, P2_P2_EBX_REG_31_, n75216 );
nor U143638 ( n43380, P2_P1_EBX_REG_31_, n75220 );
nor U143639 ( n21648, P1_P1_STATE_REG_2_, P1_P1_STATE_REG_0_ );
nor U143640 ( n54686, P2_P1_STATE_REG_2_, P2_P1_STATE_REG_0_ );
nor U143641 ( n28958, P1_P2_STATE_REG_2_, P1_P2_STATE_REG_0_ );
nor U143642 ( n36131, P1_P3_STATE_REG_2_, P1_P3_STATE_REG_0_ );
nor U143643 ( n9442, P1_P1_EBX_REG_31_, n75217 );
nor U143644 ( n62414, P2_P2_STATE_REG_2_, P2_P2_STATE_REG_0_ );
nor U143645 ( n70851, P2_P3_STATE_REG_2_, P2_P3_STATE_REG_0_ );
or U143646 ( n32419, P1_P3_BE_N_REG_2_, P1_P3_BE_N_REG_3_ );
or U143647 ( n21684, P2_P3_BE_N_REG_2_, P2_P3_BE_N_REG_3_ );
or U143648 ( n32420, P1_P3_BE_N_REG_0_, P1_P3_BE_N_REG_1_ );
or U143649 ( n21685, P2_P3_BE_N_REG_0_, P2_P3_BE_N_REG_1_ );
nor U143650 ( n49656, n48501, n49462 );
nor U143651 ( n48862, n48501, n48815 );
nor U143652 ( n49231, n48501, n49184 );
nor U143653 ( n48599, n48501, n48535 );
nor U143654 ( n48693, n48501, n48629 );
nor U143655 ( n48964, n48501, n48896 );
nor U143656 ( n49059, n48501, n48995 );
nor U143657 ( n49153, n48501, n7834 );
nor U143658 ( n49328, n48501, n49280 );
nor U143659 ( n49421, n48501, n49358 );
nor U143660 ( n48765, n48501, n48719 );
nand U143661 ( n48107, n347, n48025 );
nand U143662 ( n48215, n48150, n347 );
nand U143663 ( n48298, n48248, n347 );
nand U143664 ( n48395, n48345, n347 );
nand U143665 ( n48499, n48427, n347 );
not U143666 ( n347, n48501 );
xnor U143667 ( n49630, n49631, n49632 );
xor U143668 ( n49604, n49605, n1213 );
nand U143669 ( n50354, n49631, n49634 );
or U143670 ( n50356, n49634, n49631 );
nand U143671 ( n50594, n1213, n49603 );
nor U143672 ( n50598, n50602, n50603 );
nand U143673 ( n50636, n50863, n8240 );
nor U143674 ( n50864, n50868, n50869 );
nand U143675 ( n50865, n50866, n50867 );
and U143676 ( n51109, n51110, n50867 );
nor U143677 ( n50868, n50867, n50872 );
xor U143678 ( n50870, n50871, n50867 );
nor U143679 ( n51116, n51123, n1328 );
nand U143680 ( n51152, n1328, n51123 );
nor U143681 ( n51161, n51162, n51163 );
nor U143682 ( n51863, n51864, n51861 );
nand U143683 ( n51518, n51859, n51861 );
nor U143684 ( n52367, n51880, n1402 );
nand U143685 ( n52792, n52793, n1433 );
nor U143686 ( n52794, n1433, n52802 );
nor U143687 ( n52799, n1422, n1433 );
not U143688 ( n1433, n52801 );
nand U143689 ( n53182, n1489, n53068 );
nor U143690 ( n53069, n1477, n1489 );
nor U143691 ( n53270, n53272, n53273 );
nor U143692 ( n53311, n53273, n53267 );
nor U143693 ( n53378, n53379, n53380 );
nand U143694 ( n53443, n53380, n53385 );
nor U143695 ( n53550, n53553, n53554 );
nor U143696 ( n53663, n53619, n53612 );
nand U143697 ( n53611, n53612, n53613 );
nor U143698 ( n53614, n53613, n53620 );
nor U143699 ( n53616, n53618, n53619 );
nor U143700 ( n53619, n53621, n53613 );
not U143701 ( n1602, n53613 );
nor U143702 ( n8426, n15683, n15684 );
nor U143703 ( n14925, n14927, n14928 );
nor U143704 ( n15037, n14927, n15038 );
nor U143705 ( n15147, n14927, n15148 );
nor U143706 ( n15257, n14927, n15258 );
nor U143707 ( n15373, n14927, n15374 );
nor U143708 ( n15484, n14927, n15485 );
nor U143709 ( n15582, n14927, n15583 );
nor U143710 ( n15788, n14927, n15789 );
nor U143711 ( n15897, n14927, n15898 );
nor U143712 ( n16004, n14927, n16005 );
nor U143713 ( n16103, n14927, n16104 );
nor U143714 ( n16204, n14927, n16205 );
nor U143715 ( n16314, n14927, n16315 );
nor U143716 ( n16417, n14927, n16418 );
nor U143717 ( n16705, n14927, n16707 );
nor U143718 ( n15684, n14927, n15685 );
xor U143719 ( n16619, n16622, n16623 );
nor U143720 ( n17388, n16659, n17389 );
not U143721 ( n2354, n17389 );
nand U143722 ( n17393, n16620, n16622 );
or U143723 ( n17639, n16622, n16620 );
nand U143724 ( n17644, n17632, n17631 );
nor U143725 ( n17645, n17631, n17649 );
nor U143726 ( n17646, n2392, n17647 );
not U143727 ( n2364, n17631 );
nand U143728 ( n17903, n17904, n17631 );
xor U143729 ( n17647, n17631, n17648 );
nor U143730 ( n17908, n17912, n17913 );
nor U143731 ( n17913, n2400, n17914 );
nor U143732 ( n18161, n18162, n18163 );
nand U143733 ( n18165, n18163, n18164 );
not U143734 ( n2447, n18163 );
nor U143735 ( n18200, n18204, n18205 );
nor U143736 ( n18205, n18206, n18207 );
nor U143737 ( n19248, n19251, n19252 );
nor U143738 ( n18922, n18926, n18927 );
not U143739 ( n2522, n18927 );
nor U143740 ( n19842, n19844, n19845 );
nand U143741 ( n19968, n19845, n19841 );
nand U143742 ( n20106, n20107, n20108 );
nand U143743 ( n16982, n16981, n16983 );
nor U143744 ( n20109, n20108, n20115 );
nand U143745 ( n20328, n2613, n20112 );
nor U143746 ( n20114, n20116, n20108 );
not U143747 ( n2613, n20108 );
nor U143748 ( n20418, n20420, n20421 );
nand U143749 ( n20454, n20421, n20417 );
nor U143750 ( n20520, n20521, n20522 );
nand U143751 ( n20755, n20522, n20527 );
not U143752 ( n2667, n20522 );
nor U143753 ( n20702, n20706, n20707 );
nand U143754 ( n20703, n20704, n20705 );
nand U143755 ( n20764, n2693, n20705 );
nor U143756 ( n20762, n20763, n20705 );
nor U143757 ( n18660, n16983, n73417 );
not U143758 ( n2689, n20705 );
xnor U143759 ( n20802, n20884, n20770 );
or U143760 ( n20765, n20770, n20769 );
nand U143761 ( n20767, n20769, n20770 );
nor U143762 ( n18517, n16983, n75916 );
nand U143763 ( n20886, n20799, n20887 );
nor U143764 ( n20888, n20887, n20893 );
nor U143765 ( n20305, n16983, n73407 );
nor U143766 ( n19938, n16983, n73006 );
nor U143767 ( n20600, n16983, n73011 );
nor U143768 ( n19046, n73000, n16983 );
nor U143769 ( n20798, n20892, n20887 );
nor U143770 ( n19368, n73398, n16983 );
not U143771 ( n2723, n20887 );
nor U143772 ( n18104, n16983, n73409 );
nor U143773 ( n20672, n16983, n73007 );
nor U143774 ( n17853, n16983, n73004 );
nor U143775 ( n17583, n16983, n73399 );
nor U143776 ( n17367, n73396, n16983 );
nand U143777 ( n16488, n8222, n16983 );
not U143778 ( n8224, n16983 );
nor U143779 ( n48115, n48116, n48117 );
nor U143780 ( n48220, n48116, n48221 );
nor U143781 ( n48303, n48116, n48304 );
nor U143782 ( n48400, n48116, n48401 );
nor U143783 ( n48505, n48116, n48506 );
nor U143784 ( n48602, n48116, n48603 );
nor U143785 ( n48696, n48116, n48697 );
nor U143786 ( n48773, n48116, n48774 );
nor U143787 ( n48865, n48116, n48866 );
nor U143788 ( n48967, n48116, n48968 );
nor U143789 ( n49062, n48116, n49063 );
nor U143790 ( n49156, n48116, n49157 );
nor U143791 ( n49234, n48116, n49235 );
nor U143792 ( n49331, n48116, n49332 );
nor U143793 ( n49424, n48116, n49425 );
nor U143794 ( n49664, n48116, n49665 );
nor U143795 ( n50343, n49634, n50344 );
not U143796 ( n1212, n50344 );
nand U143797 ( n50348, n1247, n50351 );
not U143798 ( n1213, n50351 );
nand U143799 ( n50599, n1270, n50600 );
nor U143800 ( n50602, n50600, n50606 );
nor U143801 ( n50603, n1277, n50604 );
nand U143802 ( n50858, n50859, n50600 );
not U143803 ( n1248, n50600 );
nor U143804 ( n50869, n1284, n50870 );
nand U143805 ( n51143, n50921, n51144 );
not U143806 ( n1324, n51144 );
and U143807 ( n51149, n51145, n51144 );
nor U143808 ( n51118, n51119, n51120 );
nand U143809 ( n51122, n51120, n51121 );
not U143810 ( n1328, n51120 );
and U143811 ( n51515, n51516, n51159 );
nand U143812 ( n51157, n51158, n51159 );
or U143813 ( n51165, n1400, n51159 );
xor U143814 ( n51163, n51159, n51164 );
nor U143815 ( n51878, n51882, n51883 );
not U143816 ( n1402, n51883 );
nor U143817 ( n52796, n52798, n52799 );
nor U143818 ( n52798, n52800, n52801 );
nor U143819 ( n52923, n52799, n52793 );
nand U143820 ( n52924, n52801, n52797 );
xor U143821 ( n52801, n52921, n53054 );
nand U143822 ( n49939, n49938, n49940 );
nand U143823 ( n53062, n53063, n53064 );
nor U143824 ( n53065, n53064, n53071 );
not U143825 ( n1489, n53064 );
xnor U143826 ( n53064, n53277, n53278 );
nand U143827 ( n53419, n1515, n53307 );
nor U143828 ( n53272, n53274, n53275 );
and U143829 ( n53306, n53307, n1515 );
nand U143830 ( n53312, n53275, n53271 );
nor U143831 ( n53305, n1515, n53307 );
nand U143832 ( n53510, n53439, n53436 );
xor U143833 ( n53275, n53307, n53386 );
nor U143834 ( n53437, n1550, n53439 );
not U143835 ( n1564, n53439 );
nor U143836 ( n53554, n53555, n53556 );
nand U143837 ( n53586, n53556, n53561 );
nor U143838 ( n51620, n73016, n49940 );
not U143839 ( n1587, n53556 );
nor U143840 ( n51481, n73415, n49940 );
nand U143841 ( n53679, n53680, n53681 );
nand U143842 ( n53723, n1615, n53685 );
nor U143843 ( n53682, n53681, n53688 );
nor U143844 ( n53836, n73401, n49940 );
nor U143845 ( n52891, n73001, n49940 );
nor U143846 ( n53883, n73005, n49940 );
nor U143847 ( n51058, n73010, n49940 );
not U143848 ( n1615, n53681 );
nor U143849 ( n50798, n73405, n49940 );
nor U143850 ( n53871, n73403, n49940 );
nor U143851 ( n50542, n73402, n49940 );
nand U143852 ( n49482, n76649, n49940 );
not U143853 ( n76173, P2_P1_STATE2_REG_3_ );
not U143854 ( n76174, P2_P1_STATE2_REG_3_ );
not U143855 ( n76175, n76173 );
not U143856 ( n76176, n76173 );
not U143857 ( n76177, n76173 );
not U143858 ( n76178, n76173 );
not U143859 ( n76179, n76174 );
not U143860 ( n76180, n76174 );
not U143861 ( n76181, n76174 );
not U143862 ( n76182, n76174 );
not U143863 ( n76183, P1_P1_STATE2_REG_3_ );
not U143864 ( n76184, P1_P1_STATE2_REG_3_ );
not U143865 ( n76185, n76183 );
not U143866 ( n76186, n76183 );
not U143867 ( n76187, n76183 );
not U143868 ( n76188, n76183 );
not U143869 ( n76189, n76184 );
not U143870 ( n76190, n76184 );
not U143871 ( n76191, n76184 );
not U143872 ( n76192, n76184 );
endmodule

