
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule

module s9234_ori ( clk, reset, g89, g102, g557, g558, g559, g560, g561, g562, g563, g564, g705, g2584, g3222,
g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282,
g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728
);
input clk, reset, g89, g102, g557, g558, g559, g560, g561, g562, g563, g564, g705;
output g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728;
wire ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, g564, g705, g567, g571, g598, g606, g634, g642, g646, g650, g654, g22,
g41, g47, g663, g665, g667, g666, g664, g699, g702, g684, g4321,
g4307, g18, g24, g1, g28, g2, g6, g10, g40, g14, g32, g36, g37, g42,
g38, g39, g45, g3600, g46, new_g2670_, new_g2859_, new_g2861_,
new_g3454_, new_g3599_, new_g3814_, new_g3910_, new_g3768_,
new_g3828_, new_g3844_, new_g4157_, new_g4219_, new_g4430_,
new_g4433_, new_g4434_, new_g4436_, new_g4438_, new_g4440_,
new_g4441_, new_g4443_, new_g4444_, new_g4446_, new_g4447_,
new_g4450_, new_g4451_, new_g4454_, new_g4455_, new_g4458_,
new_g4460_, new_g4501_, new_g4687_, new_g4761_, new_g5019_,
new_g4872_, new_g5017_, new_g5149_, new_g5167_, new_g5231_,
new_g5386_, new_g5531_, new_g5532_, new_g5533_, new_g5535_,
new_g5622_, new_g5624_, new_g5625_, new_g5626_, new_g5627_,
new_g5628_, new_g5629_, new_g5630_, new_g6142_, new_g6287_,
new_g6286_, new_g6290_, new_g6289_, new_g6294_, new_g6292_,
new_g6293_, new_g6298_, new_g6296_, new_g6297_, new_g6300_,
new_g6301_, new_g6303_, new_g6307_, new_g6309_, new_g6310_,
new_g6291_, new_g6295_, new_g6299_, new_g6304_, new_g6485_,
new_g6482_, new_g6479_, new_g6426_, new_g6480_, new_g6481_,
new_g6483_, new_g6437_, new_g6684_, new_g6685_, new_g6686_,
new_g6687_, new_g6688_, new_g6689_, new_g6690_, new_g6691_,
new_g6658_, new_g6704_, new_g6702_, new_g6774_, new_g6778_,
new_g6791_, new_g6792_, new_g6793_, new_g6794_, new_g6787_,
new_g6788_, new_g6789_, new_g6790_, new_g6844_, new_g6845_, g212,
g224, g230, g236, g242, g248, g254, g676, n9, n53, n71, n72, n699,
n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
n1517, n1518, n1519, n1520, n1521, n1522;
assign g4422 = g564;
assign g3222 = g705;
assign g5469 = g4321;
assign g5468 = g4307;
assign g5137 = g3600;
assign g6728 = 1'b0;
assign g5692 = 1'b0;

dff g46_reg ( clk, reset, g46, g46 );
dff g45_reg ( clk, reset, g45, g45 );
not U_inv0 ( n1476, g45 );
dff g42_reg ( clk, reset, g42, g42 );
dff g40_reg ( clk, reset, g40, g40 );
not U_inv1 ( n1444, g40 );
dff g39_reg ( clk, reset, g39, g39 );
not U_inv2 ( n1443, g39 );
dff g38_reg ( clk, reset, g38, g38 );
not U_inv3 ( n1442, g38 );
dff g37_reg ( clk, reset, g37, g37 );
not U_inv4 ( n1455, g37 );
dff g36_reg ( clk, reset, g36, g36 );
not U_inv5 ( n1454, g36 );
dff g32_reg ( clk, reset, g32, g32 );
not U_inv6 ( n1446, g32 );
dff g47_reg ( clk, reset, g47, g47 );
not U_inv7 ( n9, g47 );
dff g41_reg ( clk, reset, g41, g41 );
not U_inv8 ( n1477, g41 );
dff g22_reg ( clk, reset, g22, g22 );
not U_inv9 ( n1440, g22 );
dff g266_reg ( clk, reset, n774, new_g3910_ );
not U_inv10 ( n53, n774 );
dff g658_reg ( clk, reset, n764, new_g3814_ );
dff g667_reg ( clk, reset, g667, g45 );
dff g666_reg ( clk, reset, g666, g46 );
dff g662_reg ( clk, reset, ex_wire0, n53 );
not U_inv11 ( n1498, ex_wire0 );
dff g663_reg ( clk, reset, g663, g42 );
dff g664_reg ( clk, reset, g664, g663 );
dff g471_reg ( clk, reset, n728, g664 );
not U_inv12 ( n1464, n728 );
dff g665_reg ( clk, reset, g665, g42 );
dff g478_reg ( clk, reset, n729, g665 );
not U_inv13 ( n1465, n729 );
dff g638_reg ( clk, reset, ex_wire1, g667 );
not U_inv14 ( n1499, ex_wire1 );
dff g567_reg ( clk, reset, g567, new_g3599_ );
not U_inv15 ( n1473, g567 );
dff g212_reg ( clk, reset, g212, g567 );
dff g598_reg ( clk, reset, g598, new_g2859_ );
not U_inv16 ( n1472, g598 );
dff g218_reg ( clk, reset, ex_wire2, g598 );
not U_inv17 ( n1469, ex_wire2 );
dff g634_reg ( clk, reset, g634, new_g3454_ );
not U_inv18 ( n1488, g634 );
dff g224_reg ( clk, reset, g224, g634 );
dff g642_reg ( clk, reset, g642, new_g3844_ );
not U_inv19 ( n1489, g642 );
dff g230_reg ( clk, reset, g230, g642 );
dff g606_reg ( clk, reset, g606, new_g4219_ );
not U_inv20 ( n1490, g606 );
dff g236_reg ( clk, reset, g236, g606 );
dff g646_reg ( clk, reset, g646, new_g4501_ );
not U_inv21 ( n1459, g646 );
dff g242_reg ( clk, reset, g242, g646 );
dff g650_reg ( clk, reset, g650, new_g4761_ );
dff g248_reg ( clk, reset, g248, g650 );
dff g654_reg ( clk, reset, g654, new_g5017_ );
not U_inv22 ( n1456, g654 );
dff g254_reg ( clk, reset, g254, g654 );
dff g571_reg ( clk, reset, g571, new_g5149_ );
not U_inv23 ( n1441, g571 );
dff g260_reg ( clk, reset, ex_wire3, g571 );
not U_inv24 ( n1468, ex_wire3 );
dff g639_reg ( clk, reset, n714, g666 );
not U_inv25 ( n1500, n714 );
dff g602_reg ( clk, reset, ex_wire4, new_g2861_ );
not U_inv26 ( n1475, ex_wire4 );
dff g610_reg ( clk, reset, ex_wire5, new_g2670_ );
not U_inv27 ( n1474, ex_wire5 );
dff g613_reg ( clk, reset, ex_wire6, new_g3828_ );
not U_inv28 ( n1471, ex_wire6 );
dff g616_reg ( clk, reset, n772, new_g3768_ );
not U_inv29 ( n1495, n772 );
dff g619_reg ( clk, reset, ex_wire7, new_g4157_ );
not U_inv30 ( n1496, ex_wire7 );
dff g622_reg ( clk, reset, ex_wire8, new_g4460_ );
not U_inv31 ( n1460, ex_wire8 );
dff g625_reg ( clk, reset, ex_wire9, new_g4687_ );
not U_inv32 ( n1458, ex_wire9 );
dff g628_reg ( clk, reset, ex_wire10, new_g4872_ );
not U_inv33 ( n1457, ex_wire10 );
dff g631_reg ( clk, reset, ex_wire11, new_g5167_ );
not U_inv34 ( n1497, ex_wire11 );
dff g578_reg ( clk, reset, n719, new_g6291_ );
not U_inv35 ( n1491, n719 );
dff g590_reg ( clk, reset, ex_wire12, new_g6437_ );
not U_inv36 ( n1432, ex_wire12 );
dff g594_reg ( clk, reset, n744, new_g6304_ );
not U_inv37 ( n1431, n744 );
dff g586_reg ( clk, reset, n727, new_g6299_ );
not U_inv38 ( n1493, n727 );
dff g574_reg ( clk, reset, n771, new_g6426_ );
not U_inv39 ( n1494, n771 );
dff g582_reg ( clk, reset, n743, new_g6295_ );
not U_inv40 ( n1492, n743 );
dff g699_reg ( clk, reset, g699, n9 );
not U_inv41 ( n1501, g699 );
dff g702_reg ( clk, reset, g702, g699 );
not U_inv42 ( n1502, g702 );
dff g675_reg ( clk, reset, ex_wire13, g702 );
not U_inv43 ( n1439, ex_wire13 );
dff g685_reg ( clk, reset, n767, g32 );
dff g687_reg ( clk, reset, ex_wire14, g37 );
not U_inv44 ( n1513, ex_wire14 );
dff g688_reg ( clk, reset, ex_wire15, g38 );
not U_inv45 ( n1430, ex_wire15 );
dff g689_reg ( clk, reset, n749, g39 );
not U_inv46 ( n1514, n749 );
dff g698_reg ( clk, reset, n704, g40 );
not U_inv47 ( n1515, n704 );
dff g492_reg ( clk, reset, ex_wire16, new_g6704_ );
not U_inv48 ( n1522, ex_wire16 );
dff g7_reg ( clk, reset, new_g6688_, new_g6480_ );
not U_inv49 ( n778, new_g6688_ );
dff g2_reg ( clk, reset, g2, new_g6688_ );
not U_inv50 ( n1447, g2 );
dff g678_reg ( clk, reset, n705, g2 );
not U_inv51 ( n1511, n705 );
dff g691_reg ( clk, reset, n711, g2 );
not U_inv52 ( n72, n711 );
dff g489_reg ( clk, reset, n763, n72 );
dff g48_reg ( clk, reset, ex_wire17, new_g6658_ );
not U_inv53 ( n1445, ex_wire17 );
dff g676_reg ( clk, reset, g676, new_g5019_ );
dff g669_reg ( clk, reset, ex_wire18, new_g5386_ );
not U_inv54 ( n1503, ex_wire18 );
dff g3_reg ( clk, reset, new_g6686_, new_g6479_ );
not U_inv55 ( n779, new_g6686_ );
dff g1_reg ( clk, reset, g1, new_g6686_ );
not U_inv56 ( n1453, g1 );
dff g677_reg ( clk, reset, n748, g1 );
not U_inv57 ( n1510, n748 );
dff g690_reg ( clk, reset, n712, g1 );
not U_inv58 ( n71, n712 );
dff g486_reg ( clk, reset, n762, n71 );
dff g532_reg ( clk, reset, n723, new_g6301_ );
dff g465_reg ( clk, reset, n700, new_g6297_ );
not U_inv59 ( n1518, n700 );
dff g504_reg ( clk, reset, ex_wire19, new_g6296_ );
not U_inv60 ( n1470, ex_wire19 );
dff g500_reg ( clk, reset, ex_wire20, new_g6292_ );
not U_inv61 ( n1467, ex_wire20 );
dff g528_reg ( clk, reset, n725, new_g6286_ );
dff g536_reg ( clk, reset, n756, new_g6293_ );
not U_inv62 ( n1519, n756 );
dff g402_reg ( clk, reset, n755, new_g4438_ );
not U_inv63 ( n1466, n755 );
dff g406_reg ( clk, reset, n754, new_g4441_ );
not U_inv64 ( n1463, n754 );
dff g410_reg ( clk, reset, n733, new_g4444_ );
dff g414_reg ( clk, reset, n732, new_g4447_ );
dff g418_reg ( clk, reset, n731, new_g4451_ );
dff g422_reg ( clk, reset, n730, new_g4455_ );
dff g426_reg ( clk, reset, n736, new_g4458_ );
dff g430_reg ( clk, reset, n737, new_g4434_ );
dff g461_reg ( clk, reset, n735, new_g4440_ );
dff g457_reg ( clk, reset, n734, new_g4443_ );
dff g453_reg ( clk, reset, n753, new_g4446_ );
not U_inv65 ( n1462, n753 );
dff g449_reg ( clk, reset, n752, new_g4450_ );
not U_inv66 ( n1461, n752 );
dff g445_reg ( clk, reset, n739, new_g4454_ );
dff g441_reg ( clk, reset, n740, new_g4430_ );
dff g437_reg ( clk, reset, n738, new_g4433_ );
dff g434_reg ( clk, reset, n761, new_g4436_ );
dff g33_reg ( clk, reset, new_g6687_, new_g6845_ );
not U_inv67 ( n747, new_g6687_ );
dff g28_reg ( clk, reset, g28, new_g6687_ );
not U_inv68 ( n1449, g28 );
dff g684_reg ( clk, reset, g684, g28 );
dff g697_reg ( clk, reset, n706, g28 );
dff g211_reg ( clk, reset, n718, new_g6792_ );
not U_inv69 ( n1438, n718 );
dff g210_reg ( clk, reset, n703, new_g6791_ );
not U_inv70 ( n1487, n703 );
dff g29_reg ( clk, reset, new_g6685_, new_g6844_ );
not U_inv71 ( n776, new_g6685_ );
dff g24_reg ( clk, reset, g24, new_g6685_ );
not U_inv72 ( n1448, g24 );
dff g696_reg ( clk, reset, n699, g24 );
not U_inv73 ( n1509, n699 );
dff g524_reg ( clk, reset, n726, new_g6310_ );
dff g683_reg ( clk, reset, ex_wire21, g24 );
not U_inv74 ( n1512, ex_wire21 );
dff g269_reg ( clk, reset, n707, new_g6290_ );
not U_inv75 ( n1517, n707 );
dff g197_reg ( clk, reset, n708, new_g6287_ );
not U_inv76 ( n1516, n708 );
dff g208_reg ( clk, reset, n742, new_g5533_ );
not U_inv77 ( n1486, n742 );
dff g19_reg ( clk, reset, new_g6691_, new_g6483_ );
not U_inv78 ( n746, new_g6691_ );
dff g14_reg ( clk, reset, g14, new_g6691_ );
not U_inv79 ( n1451, g14 );
dff g694_reg ( clk, reset, n713, g14 );
not U_inv80 ( n1507, n713 );
dff g516_reg ( clk, reset, n720, new_g6307_ );
dff g681_reg ( clk, reset, ex_wire22, g14 );
not U_inv81 ( n1428, ex_wire22 );
dff g25_reg ( clk, reset, new_g6684_, new_g6485_ );
not U_inv82 ( n780, new_g6684_ );
dff g18_reg ( clk, reset, g18, new_g6684_ );
not U_inv83 ( n1452, g18 );
dff g695_reg ( clk, reset, n701, g18 );
not U_inv84 ( n1508, n701 );
dff g520_reg ( clk, reset, n722, new_g6309_ );
dff g682_reg ( clk, reset, ex_wire23, g18 );
not U_inv85 ( n1429, ex_wire23 );
dff g11_reg ( clk, reset, new_g6689_, new_g6481_ );
not U_inv86 ( n745, new_g6689_ );
dff g6_reg ( clk, reset, g6, new_g6689_ );
not U_inv87 ( n1450, g6 );
dff g679_reg ( clk, reset, n775, g6 );
not U_inv88 ( n1426, n775 );
dff g692_reg ( clk, reset, n710, g6 );
not U_inv89 ( n1505, n710 );
dff g508_reg ( clk, reset, n724, new_g6300_ );
dff g293_reg ( clk, reset, n760, new_g6294_ );
dff g206_reg ( clk, reset, n751, new_g5624_ );
not U_inv90 ( n1485, n751 );
dff g209_reg ( clk, reset, n766, new_g5629_ );
not U_inv91 ( n1437, n766 );
dff g204_reg ( clk, reset, n716, new_g5531_ );
not U_inv92 ( n1483, n716 );
dff g205_reg ( clk, reset, n769, new_g5622_ );
not U_inv93 ( n1484, n769 );
dff g207_reg ( clk, reset, ex_wire24, new_g5626_ );
not U_inv94 ( n1436, ex_wire24 );
dff g15_reg ( clk, reset, new_g6690_, new_g6482_ );
not U_inv95 ( n777, new_g6690_ );
dff g10_reg ( clk, reset, g10, new_g6690_ );
dff g680_reg ( clk, reset, n770, g10 );
not U_inv96 ( n1427, n770 );
dff g693_reg ( clk, reset, n709, g10 );
not U_inv97 ( n1506, n709 );
dff g512_reg ( clk, reset, n721, new_g6303_ );
dff g297_reg ( clk, reset, n759, new_g6298_ );
dff g279_reg ( clk, reset, ex_wire25, new_g5628_ );
not U_inv98 ( n1433, ex_wire25 );
dff g283_reg ( clk, reset, n717, new_g6794_ );
not U_inv99 ( n1435, n717 );
dff g276_reg ( clk, reset, n715, new_g5532_ );
not U_inv100 ( n1478, n715 );
dff g277_reg ( clk, reset, n768, new_g5625_ );
not U_inv101 ( n1479, n768 );
dff g278_reg ( clk, reset, n750, new_g5627_ );
not U_inv102 ( n1480, n750 );
dff g280_reg ( clk, reset, n741, new_g5535_ );
not U_inv103 ( n1481, n741 );
dff g281_reg ( clk, reset, n765, new_g5630_ );
not U_inv104 ( n1434, n765 );
dff g541_reg ( clk, reset, n773, new_g6289_ );
not U_inv105 ( n1520, n773 );
dff g282_reg ( clk, reset, n702, new_g6793_ );
not U_inv106 ( n1482, n702 );
dff g551_reg ( clk, reset, ex_wire26, new_g6789_ );
not U_inv107 ( n1425, ex_wire26 );
dff g554_reg ( clk, reset, ex_wire27, new_g6790_ );
not U_inv108 ( n1424, ex_wire27 );
dff g485_reg ( clk, reset, g4307, new_g6778_ );
dff g496_reg ( clk, reset, ex_wire28, new_g6702_ );
not U_inv109 ( n1521, ex_wire28 );
dff g545_reg ( clk, reset, n758, new_g6787_ );
dff g548_reg ( clk, reset, n757, new_g6788_ );
dff g668_reg ( clk, reset, g4321, new_g6774_ );
dff g43_reg ( clk, reset, g3600, new_g6142_ );
dff g672_reg ( clk, reset, ex_wire29, new_g5231_ );
not U_inv110 ( n1504, ex_wire29 );
nand U808 ( new_g6845_, n781, n782 );
nor U809 ( n782, n783, n784 );
nand U810 ( n784, n785, n786 );
nand U811 ( n786, n787, new_g6794_ );
nand U812 ( n785, n788, n706 );
nand U813 ( n783, n789, n790 );
nand U814 ( n789, n791, new_g6792_ );
nor U815 ( n781, n792, n793 );
nand U816 ( n793, n794, n795 );
nand U817 ( n795, g557, n796 );
nand U818 ( n794, n797, n725 );
nand U819 ( n792, n798, n799 );
nand U820 ( n799, n800, n761 );
nand U821 ( n798, n801, n737 );
nand U822 ( new_g6844_, n802, n803 );
nor U823 ( n803, n804, n805 );
nand U824 ( n805, n806, n807 );
nand U825 ( n807, n787, new_g6793_ );
nand U826 ( n806, n788, n699 );
nand U827 ( n804, n808, n790 );
nand U828 ( n808, n791, new_g6791_ );
nor U829 ( n802, n809, n810 );
nand U830 ( n810, n811, n812 );
nand U831 ( n812, g558, n796 );
nand U832 ( n811, n797, n726 );
nand U833 ( n809, n813, n814 );
nand U834 ( n814, n800, n738 );
nand U835 ( n813, n801, n736 );
nand U836 ( new_g6794_, n815, n816 );
nand U837 ( n816, n1517, n706 );
nand U838 ( n815, n817, n707 );
nand U839 ( new_g6793_, n818, n819 );
nand U840 ( n819, n1517, n699 );
nand U841 ( n818, n820, n707 );
nand U842 ( new_g6792_, n821, n822 );
nand U843 ( n822, n1516, n706 );
nand U844 ( n821, n823, n708 );
nand U845 ( new_g6791_, n824, n825 );
nand U846 ( n825, n1516, n699 );
nand U847 ( n824, n826, n708 );
nand U848 ( new_g6790_, n827, n828 );
nand U849 ( n828, n829, n817 );
or U850 ( n827, n829, n1424 );
nand U851 ( new_g6789_, n830, n831 );
nand U852 ( n831, n829, n820 );
or U853 ( n830, n829, n1425 );
nand U854 ( new_g6788_, n832, n833 );
nand U855 ( n833, n829, n823 );
nand U856 ( n832, n834, n757 );
nand U857 ( new_g6787_, n835, n836 );
nand U858 ( n836, n829, n826 );
not U859 ( n829, n834 );
nand U860 ( n835, n834, n758 );
nand U861 ( new_g6778_, n817, n820 );
nand U862 ( n820, n837, n838 );
nand U863 ( n838, n839, n717 );
nor U864 ( n837, n840, n841 );
nor U865 ( n841, n842, n843 );
nand U866 ( n843, n844, n702 );
nand U867 ( n817, n845, n846 );
not U868 ( n846, n842 );
nor U869 ( n842, n847, n839 );
nor U870 ( n845, n848, n849 );
nor U871 ( n849, n850, n851 );
nand U872 ( n851, n847, n702 );
nor U873 ( n848, n1435, n839 );
nand U874 ( new_g6774_, n823, n826 );
nand U875 ( n826, n852, n853 );
nand U876 ( n853, n854, n718 );
nor U877 ( n852, n855, n856 );
nor U878 ( n856, n857, n858 );
nand U879 ( n858, n859, n703 );
nand U880 ( n823, n860, n861 );
not U881 ( n861, n857 );
nor U882 ( n857, n862, n854 );
nor U883 ( n860, n863, n864 );
nor U884 ( n864, n865, n866 );
nand U885 ( n866, n862, n703 );
nor U886 ( n863, n1438, n854 );
nand U887 ( new_g6704_, n1522, n867 );
nand U888 ( n867, n868, n717 );
nand U889 ( n868, n847, n869 );
or U890 ( n869, n844, n1482 );
nand U891 ( n844, n870, n871 );
xnor U892 ( n870, n1465, n872 );
nand U893 ( n847, n873, n874 );
xnor U894 ( n874, n1465, n875 );
nand U895 ( n875, n876, n877 );
nand U896 ( n877, n878, n750 );
nor U897 ( n878, n879, n880 );
nand U898 ( n880, n881, n882 );
nand U899 ( n882, n883, n1479 );
nor U900 ( n883, n884, n885 );
nor U901 ( n885, n1506, n715 );
nor U902 ( n884, n1478, n1505 );
nand U903 ( n881, n886, n72 );
and U904 ( n879, n71, n887 );
nand U905 ( n876, n888, n1480 );
nor U906 ( n888, n889, n890 );
nand U907 ( n890, n891, n892 );
nand U908 ( n892, n886, n1508 );
nand U909 ( n891, n887, n1507 );
nor U910 ( n889, n768, n893 );
nand U911 ( n893, n894, n895 );
nand U912 ( n895, n699, n715 );
nand U913 ( n894, n1478, n706 );
nor U914 ( n873, n1482, n871 );
nand U915 ( new_g6702_, n1521, n896 );
nand U916 ( n896, n897, n718 );
nand U917 ( n897, n862, n898 );
or U918 ( n898, n859, n1487 );
nand U919 ( n859, n899, n900 );
xnor U920 ( n899, n1464, n901 );
nand U921 ( n862, n902, n903 );
xnor U922 ( n903, n1464, n904 );
nand U923 ( n904, n905, n906 );
nand U924 ( n906, n907, n751 );
nor U925 ( n907, n908, n909 );
nand U926 ( n909, n910, n911 );
nand U927 ( n911, n912, n1484 );
nor U928 ( n912, n913, n914 );
nor U929 ( n914, n1506, n716 );
nor U930 ( n913, n1483, n1505 );
nand U931 ( n910, n72, n915 );
and U932 ( n908, n916, n71 );
nand U933 ( n905, n917, n1485 );
nor U934 ( n917, n918, n919 );
nand U935 ( n919, n920, n921 );
nand U936 ( n921, n1508, n915 );
nand U937 ( n920, n1507, n916 );
nor U938 ( n918, n769, n922 );
nand U939 ( n922, n923, n924 );
nand U940 ( n924, n699, n716 );
nand U941 ( n923, n1483, n706 );
nor U942 ( n902, n1487, n900 );
not U943 ( new_g6658_, n925 );
nand U944 ( new_g6485_, n926, n927 );
nor U945 ( n927, n928, n929 );
nand U946 ( n929, n930, n931 );
nand U947 ( n931, n787, new_g5630_ );
nand U948 ( n930, n788, n701 );
nand U949 ( n928, n932, n790 );
nand U950 ( n932, n791, new_g5629_ );
nor U951 ( n926, n933, n934 );
nand U952 ( n934, n935, n936 );
nand U953 ( n936, g559, n796 );
nand U954 ( n935, n797, n722 );
nand U955 ( n933, n937, n938 );
nand U956 ( n938, n800, n740 );
nand U957 ( n937, n801, n730 );
nand U958 ( new_g6483_, n939, n940 );
nor U959 ( n940, n941, n942 );
nand U960 ( n942, n943, n944 );
nand U961 ( n944, n787, new_g5535_ );
nand U962 ( n943, n788, n713 );
nand U963 ( n941, n945, n790 );
nand U964 ( n945, n791, new_g5533_ );
nor U965 ( n939, n946, n947 );
nand U966 ( n947, n948, n949 );
nand U967 ( n949, g560, n796 );
nand U968 ( n948, n797, n720 );
nand U969 ( n946, n950, n951 );
nand U970 ( n951, n800, n739 );
nand U971 ( n950, n801, n731 );
nand U972 ( new_g6482_, n952, n953 );
nor U973 ( n953, n954, n955 );
nand U974 ( n955, n956, n957 );
nand U975 ( n957, n801, n732 );
nor U976 ( n956, n958, n959 );
nor U977 ( n959, n1461, n960 );
nor U978 ( n958, n1506, n961 );
nand U979 ( n954, n962, n963 );
nand U980 ( n963, n787, new_g5628_ );
nor U981 ( n962, n964, n965 );
and U982 ( n965, new_g5626_, n791 );
nor U983 ( n952, n966, n967 );
nand U984 ( n967, n968, n969 );
nand U985 ( n969, n970, n759 );
nand U986 ( n968, n971, n773 );
nand U987 ( n966, n972, n973 );
nand U988 ( n973, n797, n721 );
nor U989 ( n972, n974, n975 );
nor U990 ( n975, n1424, n976 );
and U991 ( n974, g561, n796 );
nand U992 ( new_g6481_, n977, n978 );
nor U993 ( n978, n979, n980 );
nand U994 ( n980, n981, n982 );
nand U995 ( n982, n801, n733 );
nor U996 ( n981, n983, n984 );
nor U997 ( n984, n1462, n960 );
nor U998 ( n983, n1505, n961 );
nand U999 ( n979, n985, n986 );
nand U1000 ( n986, n787, new_g5627_ );
nor U1001 ( n985, n964, n987 );
and U1002 ( n987, new_g5624_, n791 );
nor U1003 ( n977, n988, n989 );
nand U1004 ( n989, n990, n991 );
nand U1005 ( n991, n970, n760 );
not U1006 ( n970, n992 );
nand U1007 ( n990, n971, n756 );
nand U1008 ( n988, n993, n994 );
nand U1009 ( n994, n797, n724 );
nor U1010 ( n993, n995, n996 );
nor U1011 ( n996, n1425, n976 );
and U1012 ( n995, g562, n796 );
nand U1013 ( new_g6480_, n997, n998 );
nor U1014 ( n998, n999, n1000 );
nand U1015 ( n1000, n1001, n1002 );
nand U1016 ( n1002, n800, n734 );
nor U1017 ( n1001, n1003, n1004 );
nor U1018 ( n1004, n72, n961 );
and U1019 ( n1003, new_g5625_, n787 );
nand U1020 ( n999, n1005, n1006 );
nor U1021 ( n1006, n964, n1007 );
nor U1022 ( n1007, n1008, n1009 );
or U1023 ( n1009, n1504, n1427 );
nor U1024 ( n1005, n1010, n1011 );
and U1025 ( n1011, new_g5622_, n791 );
nor U1026 ( n1010, n1012, n1013 );
nand U1027 ( n1013, n1014, n1015 );
nand U1028 ( n1015, n705, n763 );
nand U1029 ( n1014, n1522, n1511 );
nor U1030 ( n997, n1016, n1017 );
nand U1031 ( n1017, n1018, n1019 );
nand U1032 ( n1019, n971, n700 );
nor U1033 ( n1018, n1020, n1021 );
nor U1034 ( n1021, n1517, n992 );
nor U1035 ( n1020, n1470, n1022 );
nand U1036 ( n1016, n1023, n1024 );
nand U1037 ( n1024, n1025, n757 );
nor U1038 ( n1023, n1026, n1027 );
and U1039 ( n1027, g563, n796 );
nor U1040 ( n1026, n1463, n1028 );
nand U1041 ( new_g6479_, n1029, n1030 );
nor U1042 ( n1030, n1031, n1032 );
nand U1043 ( n1032, n1033, n1034 );
nand U1044 ( n1034, n800, n735 );
nor U1045 ( n1033, n1035, n1036 );
nor U1046 ( n1036, n71, n961 );
and U1047 ( n1035, new_g5532_, n787 );
not U1048 ( n787, n1037 );
nand U1049 ( n1031, n1038, n1039 );
nor U1050 ( n1039, n964, n1040 );
nor U1051 ( n1040, n1008, n1041 );
or U1052 ( n1041, n1503, n1427 );
not U1053 ( n964, n790 );
nand U1054 ( n790, n1042, n1043 );
nor U1055 ( n1043, n1044, n1045 );
nand U1056 ( n1045, n1046, n1037 );
nand U1057 ( n1037, n1047, n1048 );
nor U1058 ( n1048, n1513, n1049 );
nor U1059 ( n1047, n704, n749 );
nor U1060 ( n1046, n800, n788 );
not U1061 ( n788, n961 );
nand U1062 ( n961, n1050, n749 );
nand U1063 ( n1050, n1051, n1052 );
or U1064 ( n1052, n767, n1049 );
nand U1065 ( n1051, n1515, n1053 );
not U1066 ( n800, n960 );
nand U1067 ( n960, n1054, n1510 );
nor U1068 ( n1054, n1429, n1055 );
nand U1069 ( n1044, n1056, n1028 );
nor U1070 ( n1056, n1025, n796 );
nor U1071 ( n1042, n1057, n1058 );
nand U1072 ( n1058, n1059, n992 );
nor U1073 ( n1059, n797, n971 );
not U1074 ( n797, n1022 );
nand U1075 ( n1057, n1060, n1008 );
nand U1076 ( n1008, n1511, n1061 );
and U1077 ( n1060, n1062, n1012 );
nor U1078 ( n1038, n1063, n1064 );
and U1079 ( n1064, new_g5531_, n791 );
not U1080 ( n791, n1062 );
nand U1081 ( n1062, n1065, n1066 );
nor U1082 ( n1066, n1049, n704 );
nand U1083 ( n1049, n1053, n1430 );
nor U1084 ( n1053, n1067, n1068 );
or U1085 ( n1067, n1498, n1069 );
and U1086 ( n1065, n1514, n1513 );
nor U1087 ( n1063, n1012, n1070 );
nand U1088 ( n1070, n1071, n1072 );
nand U1089 ( n1072, n705, n762 );
nand U1090 ( n1071, n1521, n1511 );
nand U1091 ( n1012, n1061, n1427 );
nor U1092 ( n1061, n775, n1073 );
nor U1093 ( n1029, n1074, n1075 );
nand U1094 ( n1075, n1076, n1077 );
nand U1095 ( n1077, n971, n723 );
and U1096 ( n971, n1078, n1079 );
nor U1097 ( n1078, n1055, n748 );
nor U1098 ( n1076, n1080, n1081 );
nor U1099 ( n1081, n1516, n992 );
nand U1100 ( n992, n1082, n1512 );
nor U1101 ( n1082, n1083, n1084 );
nor U1102 ( n1080, n1467, n1022 );
nand U1103 ( n1022, n1085, n1079 );
not U1104 ( n1079, n1086 );
nor U1105 ( n1085, n1510, n1055 );
nand U1106 ( n1074, n1087, n1088 );
nand U1107 ( n1088, n1025, n758 );
not U1108 ( n1025, n976 );
nand U1109 ( n976, n1089, n1429 );
nor U1110 ( n1089, n1428, n1055 );
nor U1111 ( n1087, n1090, n1091 );
and U1112 ( n1091, g564, n796 );
and U1113 ( n796, n1092, n1093 );
nor U1114 ( n1093, n1426, n1511 );
nor U1115 ( n1092, n1073, n770 );
nand U1116 ( n1073, n1094, n1095 );
nor U1117 ( n1095, n1430, n1514 );
nor U1118 ( n1094, n1515, n1084 );
not U1119 ( n1084, n1096 );
nor U1120 ( n1090, n1466, n1028 );
not U1121 ( n1028, n801 );
nor U1122 ( n801, n1097, n1055 );
nand U1123 ( n1055, n1098, n1096 );
nor U1124 ( n1096, n1069, n1099 );
and U1125 ( n1099, n53, n1498 );
nand U1126 ( n1069, n1100, n1101 );
nor U1127 ( n1101, n1477, n1501 );
nor U1128 ( n1100, n1502, n764 );
nor U1129 ( n1098, n1512, n1083 );
or U1130 ( n1097, n1429, n1510 );
nand U1131 ( new_g6437_, n1102, n1103 );
xnor U1132 ( n1103, n1432, n1104 );
nand U1133 ( new_g6426_, n1102, n1105 );
xnor U1134 ( n1105, n1494, n1106 );
nand U1135 ( n1106, n1107, n727 );
not U1136 ( n1102, n1108 );
nand U1137 ( new_g6310_, n1109, n1110 );
nand U1138 ( n1110, n1111, n699 );
nand U1139 ( n1109, n1112, n726 );
nand U1140 ( new_g6309_, n1113, n1114 );
nand U1141 ( n1114, n1111, n701 );
nand U1142 ( n1113, n1112, n722 );
nand U1143 ( new_g6307_, n1115, n1116 );
nand U1144 ( n1116, n1111, n713 );
nand U1145 ( n1115, n1112, n720 );
nor U1146 ( new_g6304_, n1117, n1108 );
nor U1147 ( n1117, n1118, n744 );
nor U1148 ( n1118, n1432, n1104 );
nand U1149 ( new_g6303_, n1119, n1120 );
nand U1150 ( n1120, n1111, n709 );
nand U1151 ( n1119, n1112, n721 );
nand U1152 ( new_g6301_, n1121, n1122 );
nand U1153 ( n1122, n1123, n712 );
nand U1154 ( n1121, n1124, n723 );
nand U1155 ( new_g6300_, n1125, n1126 );
nand U1156 ( n1126, n1111, n710 );
nand U1157 ( n1125, n1112, n724 );
nor U1158 ( new_g6299_, n1108, n1127 );
xnor U1159 ( n1127, n727, n1107 );
nand U1160 ( new_g6298_, n1128, n1129 );
nand U1161 ( n1129, n1130, n709 );
nand U1162 ( n1128, n1131, n759 );
nand U1163 ( new_g6297_, n1132, n1133 );
nand U1164 ( n1133, n1123, n711 );
nand U1165 ( n1132, n1124, n700 );
nand U1166 ( new_g6296_, n1134, n1135 );
nand U1167 ( n1135, n1111, n711 );
or U1168 ( n1134, n1111, n1470 );
nor U1169 ( new_g6295_, n1108, n1136 );
xnor U1170 ( n1136, n1492, n1137 );
nand U1171 ( new_g6294_, n1138, n1139 );
nand U1172 ( n1139, n1130, n710 );
nand U1173 ( n1138, n1131, n760 );
nand U1174 ( new_g6293_, n1140, n1141 );
nand U1175 ( n1141, n1123, n710 );
nand U1176 ( n1140, n1142, n1124 );
nor U1177 ( n1142, n1519, n1143 );
nor U1178 ( n1143, n834, n1144 );
nand U1179 ( n1144, n1145, n1146 );
nand U1180 ( n1146, n1147, n700 );
nand U1181 ( n1145, n1518, n1148 );
nand U1182 ( new_g6292_, n1149, n1150 );
nand U1183 ( n1150, n1111, n712 );
or U1184 ( n1149, n1111, n1467 );
nor U1185 ( new_g6291_, n1108, n1151 );
xnor U1186 ( n1151, n719, n1152 );
nand U1187 ( n1108, n714, n1153 );
nand U1188 ( n1153, n1154, n1155 );
not U1189 ( n1155, n1104 );
nand U1190 ( n1104, n1156, n1107 );
nor U1191 ( n1107, n1137, n1492 );
nand U1192 ( n1137, n1152, n719 );
nor U1193 ( n1152, n1157, n1497 );
nor U1194 ( n1156, n1493, n1494 );
nor U1195 ( n1154, n1431, n1432 );
nand U1196 ( new_g6290_, n1158, n1159 );
nand U1197 ( n1159, n1130, n711 );
nand U1198 ( n1158, n1131, n707 );
nand U1199 ( new_g6289_, n1160, n1161 );
nand U1200 ( n1161, n1123, n709 );
not U1201 ( n1123, n1124 );
nand U1202 ( n1160, n1162, n1124 );
nand U1203 ( n1124, n1163, n1510 );
nand U1204 ( n1162, n1520, n1164 );
nand U1205 ( n1164, n1165, n1166 );
nor U1206 ( n1166, n1167, n1168 );
nor U1207 ( n1168, n854, n700 );
not U1208 ( n854, n865 );
nor U1209 ( n1167, n1518, n839 );
not U1210 ( n839, n850 );
nand U1211 ( new_g6287_, n1169, n1170 );
nand U1212 ( n1170, n1130, n712 );
not U1213 ( n1130, n1131 );
nand U1214 ( n1169, n1131, n708 );
nand U1215 ( n1131, n1171, n1512 );
nand U1216 ( new_g6286_, n1172, n1173 );
nand U1217 ( n1173, n1111, n706 );
not U1218 ( n1111, n1112 );
nand U1219 ( n1172, n1112, n725 );
nand U1220 ( n1112, n1163, n748 );
and U1221 ( n1163, n1174, n1171 );
and U1222 ( n1171, n1175, n1176 );
nor U1223 ( n1176, n1083, n1177 );
or U1224 ( n1177, n1502, n1501 );
nand U1225 ( n1083, n1178, n1179 );
nor U1226 ( n1179, n1514, n1180 );
nand U1227 ( n1180, n767, g684 );
and U1228 ( n1178, n704, n1430 );
nor U1229 ( n1175, g41, n1068 );
nor U1230 ( n1174, n1512, n1086 );
nand U1231 ( n1086, n1428, n1429 );
nand U1232 ( g6366, n1181, n747 );
nand U1233 ( g6362, n1181, n776 );
nand U1234 ( g6360, n1181, n780 );
nand U1235 ( g6374, n1181, n746 );
nand U1236 ( g6372, n1181, n777 );
nand U1237 ( g6370, n1181, n745 );
nand U1238 ( g6368, n1181, n778 );
nand U1239 ( g6364, n1181, n779 );
nor U1240 ( new_g6142_, n1182, n1183 );
nor U1241 ( n1183, n1184, n1185 );
nand U1242 ( n1185, n1186, n1187 );
nand U1243 ( n1187, n1188, n727 );
nor U1244 ( n1188, n1189, n1190 );
nand U1245 ( n1190, n1191, n1192 );
nand U1246 ( n1192, n1491, n1193 );
nand U1247 ( n1193, n1194, n1195 );
nand U1248 ( n1195, n72, n743 );
nand U1249 ( n1191, n1196, n71 );
nor U1250 ( n1189, n1194, n710 );
nand U1251 ( n1194, n1492, n1197 );
nand U1252 ( n1197, n1491, n709 );
nand U1253 ( n1186, n1493, n1198 );
nand U1254 ( n1198, n1199, n1200 );
nand U1255 ( n1200, n1196, n713 );
nand U1256 ( n1199, n1201, n1202 );
not U1257 ( n1202, n1196 );
nand U1258 ( n1201, n1203, n1204 );
nand U1259 ( n1204, n701, n743 );
nor U1260 ( n1203, n1205, n1206 );
nor U1261 ( n1206, n1491, n1509 );
nor U1262 ( n1205, n719, n1207 );
nand U1263 ( n1207, n1492, n706 );
xnor U1264 ( n1184, n744, n1432 );
nor U1265 ( n1182, n1208, n1209 );
nand U1266 ( n1209, n1196, n1432 );
nor U1267 ( n1196, n1492, n1491 );
nand U1268 ( n1208, n1210, n771 );
nor U1269 ( n1210, n1431, n1493 );
nand U1270 ( g6284, n1181, n925 );
xnor U1271 ( n925, n1211, n1212 );
xor U1272 ( n1212, n1213, n1214 );
xnor U1273 ( n1214, n745, new_g6688_ );
xnor U1274 ( n1213, n746, new_g6690_ );
xor U1275 ( n1211, n1215, n1216 );
xnor U1276 ( n1216, n747, new_g6686_ );
xnor U1277 ( n1215, new_g6684_, new_g6685_ );
nor U1278 ( n1181, g6282, n1477 );
nand U1279 ( new_g5630_, n1217, n1218 );
nand U1280 ( n1218, n1517, n701 );
nand U1281 ( n1217, n1219, n707 );
nor U1282 ( n1219, n1220, n1221 );
nor U1283 ( n1220, n765, n1222 );
nand U1284 ( n1222, n1223, n1224 );
nand U1285 ( n1223, n1225, n741 );
nand U1286 ( new_g5629_, n1226, n1227 );
nand U1287 ( n1227, n1516, n701 );
nand U1288 ( n1226, n1228, n708 );
nor U1289 ( n1228, n1229, n1230 );
nor U1290 ( n1229, n766, n1231 );
nand U1291 ( n1231, n1232, n1233 );
nand U1292 ( n1232, n1234, n742 );
nand U1293 ( new_g5628_, n1235, n1236 );
nand U1294 ( n1236, n1517, n709 );
nand U1295 ( n1235, n1237, n707 );
nor U1296 ( n1237, n840, n1238 );
nor U1297 ( n1238, n1239, n1221 );
xor U1298 ( n1239, n1240, n1433 );
nand U1299 ( new_g5627_, n1241, n1242 );
nand U1300 ( n1242, n1243, n1244 );
xnor U1301 ( n1243, n1480, n887 );
nand U1302 ( n1241, n1517, n710 );
nand U1303 ( new_g5626_, n1245, n1246 );
nand U1304 ( n1246, n1516, n709 );
nand U1305 ( n1245, n1247, n708 );
nor U1306 ( n1247, n855, n1248 );
nor U1307 ( n1248, n1249, n1230 );
xor U1308 ( n1249, n1250, n1436 );
nand U1309 ( new_g5625_, n1251, n1252 );
nand U1310 ( n1252, n1244, n1253 );
nand U1311 ( n1253, n1254, n1255 );
nand U1312 ( n1255, n1479, n715 );
not U1313 ( n1254, n886 );
nor U1314 ( n886, n715, n1479 );
nand U1315 ( n1251, n1517, n711 );
nand U1316 ( new_g5624_, n1256, n1257 );
nand U1317 ( n1257, n1258, n1259 );
xnor U1318 ( n1258, n1485, n916 );
nand U1319 ( n1256, n1516, n710 );
nand U1320 ( new_g5622_, n1260, n1261 );
nand U1321 ( n1261, n1259, n1262 );
nand U1322 ( n1262, n1263, n1264 );
nand U1323 ( n1264, n1484, n716 );
not U1324 ( n1263, n915 );
nor U1325 ( n915, n716, n1484 );
nand U1326 ( n1260, n1516, n711 );
nand U1327 ( new_g5535_, n1265, n1266 );
nand U1328 ( n1266, n1517, n713 );
nand U1329 ( n1265, n1267, n707 );
nand U1330 ( n1267, n1268, n1269 );
nor U1331 ( n1268, n840, n1270 );
xnor U1332 ( n1270, n1481, n1225 );
nand U1333 ( new_g5533_, n1271, n1272 );
nand U1334 ( n1272, n1516, n713 );
nand U1335 ( n1271, n1273, n708 );
nand U1336 ( n1273, n1274, n1275 );
nor U1337 ( n1274, n855, n1276 );
xnor U1338 ( n1276, n1486, n1234 );
nand U1339 ( new_g5532_, n1277, n1278 );
nand U1340 ( n1278, n1244, n1478 );
and U1341 ( n1244, n1279, n1269 );
not U1342 ( n1269, n1221 );
nand U1343 ( n1221, n850, n1280 );
nand U1344 ( n1280, n1281, n1282 );
nor U1345 ( n1282, n729, n702 );
nor U1346 ( n1281, n717, n1283 );
nand U1347 ( n850, n1284, n1225 );
nor U1348 ( n1284, n1434, n1481 );
nor U1349 ( n1279, n1517, n840 );
not U1350 ( n840, n1224 );
nand U1351 ( n1224, n1285, n1286 );
nor U1352 ( n1286, n872, n729 );
not U1353 ( n872, n1283 );
nand U1354 ( n1283, n871, n1147 );
nand U1355 ( n1147, n1287, n1481 );
and U1356 ( n1287, n765, n1225 );
nor U1357 ( n1225, n1240, n1433 );
nand U1358 ( n1240, n887, n750 );
nor U1359 ( n887, n1478, n1479 );
xnor U1360 ( n871, n741, n1434 );
nor U1361 ( n1285, n702, n717 );
nand U1362 ( n1277, n1517, n712 );
nand U1363 ( new_g5531_, n1288, n1289 );
nand U1364 ( n1289, n1259, n1483 );
and U1365 ( n1259, n1290, n1275 );
not U1366 ( n1275, n1230 );
nand U1367 ( n1230, n865, n1291 );
nand U1368 ( n1291, n1292, n1293 );
nor U1369 ( n1293, n728, n703 );
nor U1370 ( n1292, n718, n1294 );
nand U1371 ( n865, n1295, n1234 );
nor U1372 ( n1295, n1437, n1486 );
nor U1373 ( n1290, n1516, n855 );
not U1374 ( n855, n1233 );
nand U1375 ( n1233, n1296, n1297 );
nor U1376 ( n1297, n901, n728 );
not U1377 ( n901, n1294 );
nand U1378 ( n1294, n900, n1148 );
nand U1379 ( n1148, n1298, n1486 );
and U1380 ( n1298, n766, n1234 );
nor U1381 ( n1234, n1250, n1436 );
nand U1382 ( n1250, n916, n751 );
nor U1383 ( n916, n1483, n1484 );
xnor U1384 ( n900, n742, n1437 );
nor U1385 ( n1296, n703, n718 );
nand U1386 ( n1288, n1516, n712 );
nand U1387 ( new_g5386_, n1503, n1299 );
nand U1388 ( n1299, n1440, n1300 );
nand U1389 ( g6282, n1301, n1440 );
nor U1390 ( n1301, n1439, n1068 );
nand U1391 ( n1068, g676, n1302 );
nand U1392 ( n1302, n1477, n1303 );
nand U1393 ( new_g5231_, n1504, n1304 );
nand U1394 ( n1304, n1305, n1440 );
and U1395 ( n1305, n1303, n1477 );
xnor U1396 ( n1303, n1306, n1445 );
nor U1397 ( new_g5167_, n1500, n1307 );
xnor U1398 ( n1307, n1497, n1157 );
or U1399 ( n1157, n1308, n1457 );
nor U1400 ( new_g5149_, n1499, n1309 );
xor U1401 ( n1309, n1441, n1310 );
nor U1402 ( n1310, n1456, n1311 );
not U1403 ( new_g5019_, n1300 );
xnor U1404 ( n1300, n1312, n1313 );
xor U1405 ( n1313, n1314, n1315 );
xor U1406 ( n1315, n1444, n1445 );
xor U1407 ( n1314, n1442, n1443 );
xor U1408 ( n1312, n1316, n1317 );
xor U1409 ( n1317, n1446, n1454 );
xor U1410 ( n1316, n1306, n1455 );
xor U1411 ( n1306, n1318, n1319 );
xor U1412 ( n1319, n1320, n1321 );
xor U1413 ( n1321, n1449, n1450 );
xor U1414 ( n1320, n1447, n1448 );
xor U1415 ( n1318, n1322, n1323 );
xor U1416 ( n1323, n1451, n1452 );
xor U1417 ( n1322, g10, n1453 );
nor U1418 ( new_g5017_, n1499, n1324 );
xnor U1419 ( n1324, n1456, n1311 );
nand U1420 ( n1311, n1325, g650 );
nor U1421 ( new_g4872_, n1500, n1326 );
xnor U1422 ( n1326, n1457, n1308 );
or U1423 ( n1308, n1327, n1458 );
nor U1424 ( new_g4761_, n1499, n1328 );
xnor U1425 ( n1328, g650, n1325 );
nor U1426 ( n1325, n1329, n1459 );
nor U1427 ( new_g4687_, n1500, n1330 );
xnor U1428 ( n1330, n1458, n1327 );
or U1429 ( n1327, n1331, n1460 );
nor U1430 ( new_g4501_, n1499, n1332 );
xnor U1431 ( n1332, n1459, n1329 );
or U1432 ( n1329, n1333, n1490 );
nor U1433 ( new_g4460_, n1500, n1334 );
xnor U1434 ( n1334, n1460, n1331 );
or U1435 ( n1331, n1335, n1496 );
nand U1436 ( new_g4458_, n1336, n1337 );
nand U1437 ( n1337, n1338, n730 );
nand U1438 ( n1336, n1339, n736 );
nand U1439 ( new_g4455_, n1340, n1341 );
nand U1440 ( n1341, n1338, n731 );
nand U1441 ( n1340, n1339, n730 );
nand U1442 ( new_g4454_, n1342, n1343 );
nand U1443 ( n1343, n1338, n752 );
nand U1444 ( n1342, n1339, n739 );
nand U1445 ( new_g4451_, n1344, n1345 );
nand U1446 ( n1345, n1338, n732 );
nand U1447 ( n1344, n1339, n731 );
nand U1448 ( new_g4450_, n1346, n1347 );
nand U1449 ( n1347, n1338, n753 );
nand U1450 ( n1346, n1339, n752 );
nand U1451 ( new_g4447_, n1348, n1349 );
nand U1452 ( n1349, n1338, n733 );
nand U1453 ( n1348, n1339, n732 );
nand U1454 ( new_g4446_, n1350, n1351 );
nand U1455 ( n1351, n1338, n734 );
nand U1456 ( n1350, n1339, n753 );
nand U1457 ( new_g4444_, n1352, n1353 );
nand U1458 ( n1353, n1338, n754 );
nand U1459 ( n1352, n1339, n733 );
nand U1460 ( new_g4443_, n1354, n1355 );
nand U1461 ( n1355, n1338, n735 );
nand U1462 ( n1354, n1339, n734 );
nand U1463 ( new_g4441_, n1356, n1357 );
nand U1464 ( n1357, n1338, n755 );
nand U1465 ( n1356, n1339, n754 );
nand U1466 ( new_g4440_, n1358, n1359 );
nand U1467 ( n1359, n1338, n737 );
nand U1468 ( n1358, n1339, n735 );
nand U1469 ( new_g4438_, n1360, n1361 );
nand U1470 ( n1361, n1339, n755 );
nand U1471 ( n1360, n1362, n1338 );
nand U1472 ( n1362, n1363, n1364 );
nand U1473 ( n1364, n1518, n728 );
nand U1474 ( n1363, n700, n729 );
nand U1475 ( new_g4436_, n1365, n1366 );
nand U1476 ( n1366, n1338, n738 );
nand U1477 ( n1365, n1339, n761 );
nand U1478 ( new_g4434_, n1367, n1368 );
nand U1479 ( n1368, n1338, n736 );
nand U1480 ( n1367, n1339, n737 );
nand U1481 ( new_g4433_, n1369, n1370 );
nand U1482 ( n1370, n1338, n740 );
nand U1483 ( n1369, n1339, n738 );
nand U1484 ( new_g4430_, n1371, n1372 );
nand U1485 ( n1372, n1338, n739 );
not U1486 ( n1338, n1339 );
nand U1487 ( n1371, n1339, n740 );
nand U1488 ( n1339, n1165, n1520 );
nor U1489 ( n1165, n834, n756 );
nand U1490 ( n834, n1373, n1374 );
nor U1491 ( n1374, n1375, n1376 );
nand U1492 ( n1376, n1377, n1378 );
xnor U1493 ( n1378, g236, n720 );
xnor U1494 ( n1377, g230, n721 );
nand U1495 ( n1375, n1379, n1380 );
xnor U1496 ( n1380, g242, n722 );
nor U1497 ( n1379, n1381, n1382 );
xnor U1498 ( n1382, n1468, n723 );
xor U1499 ( n1381, n1469, n1470 );
nor U1500 ( n1373, n1383, n1384 );
nand U1501 ( n1384, n1385, n1386 );
xor U1502 ( n1386, g212, n1467 );
xnor U1503 ( n1385, g224, n724 );
nand U1504 ( n1383, n1387, n1388 );
xnor U1505 ( n1388, g254, n725 );
xnor U1506 ( n1387, g248, n726 );
nor U1507 ( new_g4219_, n1499, n1389 );
xnor U1508 ( n1389, n1490, n1333 );
nand U1509 ( n1333, n1390, g642 );
nor U1510 ( new_g4157_, n1500, n1391 );
xnor U1511 ( n1391, n1496, n1335 );
nand U1512 ( n1335, n1392, n1393 );
nor U1513 ( n1392, n1475, n1495 );
nor U1514 ( new_g3910_, n1476, n774 );
nand U1515 ( new_g3844_, n1394, n1395 );
nand U1516 ( n1395, n1396, g642 );
nor U1517 ( n1396, n1499, n1390 );
and U1518 ( n1390, n1397, g634 );
nand U1519 ( n1394, n1398, n1489 );
nor U1520 ( n1398, new_g3599_, n1399 );
nand U1521 ( n1399, g634, g598 );
nand U1522 ( new_g3828_, n1400, n714 );
xor U1523 ( n1400, n1471, n1401 );
nor U1524 ( n1401, n1475, n1474 );
nor U1525 ( new_g3814_, n1476, n764 );
nand U1526 ( new_g3768_, n1402, n1403 );
nand U1527 ( n1403, n1404, n772 );
nand U1528 ( n1404, n1405, n1406 );
nand U1529 ( n1406, n1407, n714 );
nand U1530 ( n1402, n1408, n1495 );
nor U1531 ( n1408, n1407, n1409 );
or U1532 ( n1409, n1500, n1475 );
not U1533 ( n1407, n1393 );
nor U1534 ( n1393, n1471, n1474 );
nand U1535 ( new_g3454_, n1410, n1411 );
nand U1536 ( n1411, n1412, g634 );
nor U1537 ( n1412, n1499, n1397 );
nor U1538 ( n1397, n1472, n1473 );
nand U1539 ( n1410, n1413, n1488 );
nor U1540 ( n1413, n1472, new_g3599_ );
not U1541 ( new_g3599_, n1414 );
not U1542 ( new_g2861_, n1405 );
nand U1543 ( new_g2859_, n1415, n1416 );
nand U1544 ( n1416, n1417, g598 );
nor U1545 ( n1417, n1499, g567 );
nand U1546 ( n1415, n1472, n1414 );
nor U1547 ( n1414, n1473, n1499 );
nand U1548 ( new_g2670_, n1418, n1419 );
or U1549 ( n1419, n1405, n1474 );
nand U1550 ( n1405, n1475, n714 );
nand U1551 ( n1418, n1420, n1474 );
nor U1552 ( n1420, n1475, n1500 );
nor U1553 ( g4809, n1421, n1422 );
nor U1554 ( n1422, n1521, n762 );
nor U1555 ( n1421, n1522, n763 );
nor U1556 ( g2584, g102, n1423 );
not U1557 ( n1423, g89 );
endmodule

