module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule

module fir_ori ( clk, reset, inData_0, inData_1, inData_2, inData_3, inData_4, inData_5, inData_6, inData_7, inData_8, inData_9, inData_10, inData_11, inData_12, inData_13, inData_14, inData_15, inData_16, inData_17, inData_18, inData_19, inData_20, inData_21, inData_22, inData_23, inData_24, inData_25, inData_26, inData_27, inData_28, inData_29, inData_30, inData_31, outData_0, outData_1, outData_2, outData_3, outData_4, outData_5, outData_6, outData_7, outData_8, outData_9, outData_10, outData_11, outData_12, outData_13, outData_14, outData_15, outData_16, outData_17, outData_18, outData_19, outData_20, outData_21, outData_22, outData_23, outData_24, outData_25, outData_26, outData_27, outData_28, outData_29, outData_30, outData_31 );
input clk, reset, inData_0, inData_1, inData_2, inData_3, inData_4, inData_5, inData_6, inData_7, inData_8, inData_9, inData_10, inData_11, inData_12, inData_13, inData_14, inData_15, inData_16, inData_17, inData_18, inData_19, inData_20, inData_21, inData_22, inData_23, inData_24, inData_25, inData_26, inData_27, inData_28, inData_29, inData_30, inData_31;
output outData_0, outData_1, outData_2, outData_3, outData_4, outData_5, outData_6, outData_7, outData_8, outData_9, outData_10, outData_11, outData_12, outData_13, outData_14, outData_15, outData_16, outData_17, outData_18, outData_19, outData_20, outData_21, outData_22, outData_23, outData_24, outData_25, outData_26, outData_27, outData_28, outData_29, outData_30, outData_31;
wire my_FIR_filter_firBlock_left_N288, ex_wire0, my_FIR_filter_firBlock_left_N287,
my_FIR_filter_firBlock_left_N286, my_FIR_filter_firBlock_left_N285,
my_FIR_filter_firBlock_left_N284, my_FIR_filter_firBlock_left_N283,
my_FIR_filter_firBlock_left_N282, my_FIR_filter_firBlock_left_N281,
my_FIR_filter_firBlock_left_N280, my_FIR_filter_firBlock_left_N279,
my_FIR_filter_firBlock_left_N278, my_FIR_filter_firBlock_left_N277,
my_FIR_filter_firBlock_left_N276, my_FIR_filter_firBlock_left_N275,
my_FIR_filter_firBlock_left_N274, my_FIR_filter_firBlock_left_N273,
my_FIR_filter_firBlock_left_N272, my_FIR_filter_firBlock_left_N271,
my_FIR_filter_firBlock_left_N270, my_FIR_filter_firBlock_left_N269,
my_FIR_filter_firBlock_left_N268, my_FIR_filter_firBlock_left_N267,
my_FIR_filter_firBlock_left_N266, my_FIR_filter_firBlock_left_N265,
my_FIR_filter_firBlock_left_N264, my_FIR_filter_firBlock_left_N263,
my_FIR_filter_firBlock_left_N262, my_FIR_filter_firBlock_left_N261,
my_FIR_filter_firBlock_left_N260, my_FIR_filter_firBlock_left_N259,
my_FIR_filter_firBlock_left_N258, my_FIR_filter_firBlock_left_N257,
my_FIR_filter_firBlock_left_N256, my_FIR_filter_firBlock_left_N255,
my_FIR_filter_firBlock_left_N254, my_FIR_filter_firBlock_left_N253,
my_FIR_filter_firBlock_left_N252, my_FIR_filter_firBlock_left_N251,
my_FIR_filter_firBlock_left_N250, my_FIR_filter_firBlock_left_N249,
my_FIR_filter_firBlock_left_N248, my_FIR_filter_firBlock_left_N247,
my_FIR_filter_firBlock_left_N246, my_FIR_filter_firBlock_left_N245,
my_FIR_filter_firBlock_left_N244, my_FIR_filter_firBlock_left_N243,
my_FIR_filter_firBlock_left_N242, my_FIR_filter_firBlock_left_N241,
my_FIR_filter_firBlock_left_N240, my_FIR_filter_firBlock_left_N239,
my_FIR_filter_firBlock_left_N238, my_FIR_filter_firBlock_left_N237,
my_FIR_filter_firBlock_left_N236, my_FIR_filter_firBlock_left_N235,
my_FIR_filter_firBlock_left_N234, my_FIR_filter_firBlock_left_N233,
my_FIR_filter_firBlock_left_N232, my_FIR_filter_firBlock_left_N231,
my_FIR_filter_firBlock_left_N230, my_FIR_filter_firBlock_left_N229,
my_FIR_filter_firBlock_left_N228, my_FIR_filter_firBlock_left_N227,
my_FIR_filter_firBlock_left_N226, my_FIR_filter_firBlock_left_N225,
my_FIR_filter_firBlock_left_N224, my_FIR_filter_firBlock_left_N223,
my_FIR_filter_firBlock_left_N222, my_FIR_filter_firBlock_left_N221,
my_FIR_filter_firBlock_left_N220, my_FIR_filter_firBlock_left_N219,
my_FIR_filter_firBlock_left_N218, my_FIR_filter_firBlock_left_N217,
my_FIR_filter_firBlock_left_N216, my_FIR_filter_firBlock_left_N215,
my_FIR_filter_firBlock_left_N214, my_FIR_filter_firBlock_left_N213,
my_FIR_filter_firBlock_left_N212, my_FIR_filter_firBlock_left_N211,
my_FIR_filter_firBlock_left_N210, my_FIR_filter_firBlock_left_N209,
my_FIR_filter_firBlock_left_N208, my_FIR_filter_firBlock_left_N207,
my_FIR_filter_firBlock_left_N206, my_FIR_filter_firBlock_left_N205,
my_FIR_filter_firBlock_left_N204, my_FIR_filter_firBlock_left_N203,
my_FIR_filter_firBlock_left_N202, my_FIR_filter_firBlock_left_N201,
my_FIR_filter_firBlock_left_N200, my_FIR_filter_firBlock_left_N199,
my_FIR_filter_firBlock_left_N198, my_FIR_filter_firBlock_left_N197,
my_FIR_filter_firBlock_left_N196, my_FIR_filter_firBlock_left_N195,
my_FIR_filter_firBlock_left_N194, my_FIR_filter_firBlock_left_N193,
my_FIR_filter_firBlock_left_N192, my_FIR_filter_firBlock_left_N191,
my_FIR_filter_firBlock_left_N190, my_FIR_filter_firBlock_left_N189,
my_FIR_filter_firBlock_left_N188, my_FIR_filter_firBlock_left_N187,
my_FIR_filter_firBlock_left_N186, my_FIR_filter_firBlock_left_N185,
my_FIR_filter_firBlock_left_N184, my_FIR_filter_firBlock_left_N183,
my_FIR_filter_firBlock_left_N182, my_FIR_filter_firBlock_left_N181,
my_FIR_filter_firBlock_left_N180, my_FIR_filter_firBlock_left_N179,
my_FIR_filter_firBlock_left_N178, my_FIR_filter_firBlock_left_N177,
my_FIR_filter_firBlock_left_N176, my_FIR_filter_firBlock_left_N175,
my_FIR_filter_firBlock_left_N174, my_FIR_filter_firBlock_left_N173,
my_FIR_filter_firBlock_left_N172, my_FIR_filter_firBlock_left_N171,
my_FIR_filter_firBlock_left_N170, my_FIR_filter_firBlock_left_N169,
my_FIR_filter_firBlock_left_N168, my_FIR_filter_firBlock_left_N167,
my_FIR_filter_firBlock_left_N166, my_FIR_filter_firBlock_left_N165,
my_FIR_filter_firBlock_left_N164, my_FIR_filter_firBlock_left_N163,
my_FIR_filter_firBlock_left_N162, my_FIR_filter_firBlock_left_N161,
my_FIR_filter_firBlock_left_N160, my_FIR_filter_firBlock_left_N159,
my_FIR_filter_firBlock_left_N158, my_FIR_filter_firBlock_left_N157,
my_FIR_filter_firBlock_left_N156, my_FIR_filter_firBlock_left_N155,
my_FIR_filter_firBlock_left_N154, my_FIR_filter_firBlock_left_N153,
my_FIR_filter_firBlock_left_N152, my_FIR_filter_firBlock_left_N151,
my_FIR_filter_firBlock_left_N150, my_FIR_filter_firBlock_left_N149,
my_FIR_filter_firBlock_left_N148, my_FIR_filter_firBlock_left_N147,
my_FIR_filter_firBlock_left_N146, my_FIR_filter_firBlock_left_N145,
my_FIR_filter_firBlock_left_N144, my_FIR_filter_firBlock_left_N143,
my_FIR_filter_firBlock_left_N142, my_FIR_filter_firBlock_left_N141,
my_FIR_filter_firBlock_left_N140, my_FIR_filter_firBlock_left_N139,
my_FIR_filter_firBlock_left_N138, my_FIR_filter_firBlock_left_N137,
my_FIR_filter_firBlock_left_N136, my_FIR_filter_firBlock_left_N135,
my_FIR_filter_firBlock_left_N134, my_FIR_filter_firBlock_left_N133,
my_FIR_filter_firBlock_left_N132, my_FIR_filter_firBlock_left_N131,
my_FIR_filter_firBlock_left_N130, my_FIR_filter_firBlock_left_N129,
my_FIR_filter_firBlock_left_N128, my_FIR_filter_firBlock_left_N127,
my_FIR_filter_firBlock_left_N126, my_FIR_filter_firBlock_left_N125,
my_FIR_filter_firBlock_left_N124, my_FIR_filter_firBlock_left_N123,
my_FIR_filter_firBlock_left_N122, my_FIR_filter_firBlock_left_N121,
my_FIR_filter_firBlock_left_N120, my_FIR_filter_firBlock_left_N119,
my_FIR_filter_firBlock_left_N118, my_FIR_filter_firBlock_left_N117,
my_FIR_filter_firBlock_left_N116, my_FIR_filter_firBlock_left_N115,
my_FIR_filter_firBlock_left_N114, my_FIR_filter_firBlock_left_N113,
my_FIR_filter_firBlock_left_N112, my_FIR_filter_firBlock_left_N111,
my_FIR_filter_firBlock_left_N110, my_FIR_filter_firBlock_left_N109,
my_FIR_filter_firBlock_left_N108, my_FIR_filter_firBlock_left_N107,
my_FIR_filter_firBlock_left_N106, my_FIR_filter_firBlock_left_N105,
my_FIR_filter_firBlock_left_N104, my_FIR_filter_firBlock_left_N103,
my_FIR_filter_firBlock_left_N102, my_FIR_filter_firBlock_left_N101,
my_FIR_filter_firBlock_left_N100, my_FIR_filter_firBlock_left_N99,
my_FIR_filter_firBlock_left_N98, my_FIR_filter_firBlock_left_N97,
my_FIR_filter_firBlock_left_N96, my_FIR_filter_firBlock_left_N95,
my_FIR_filter_firBlock_left_N94, my_FIR_filter_firBlock_left_N93,
my_FIR_filter_firBlock_left_N92, my_FIR_filter_firBlock_left_N91,
my_FIR_filter_firBlock_left_N90, my_FIR_filter_firBlock_left_N89,
my_FIR_filter_firBlock_left_N88, my_FIR_filter_firBlock_left_N87,
my_FIR_filter_firBlock_left_N86, my_FIR_filter_firBlock_left_N85,
my_FIR_filter_firBlock_left_N84, my_FIR_filter_firBlock_left_N83,
my_FIR_filter_firBlock_left_N82, my_FIR_filter_firBlock_left_N81,
my_FIR_filter_firBlock_left_N80, my_FIR_filter_firBlock_left_N79,
my_FIR_filter_firBlock_left_N78, my_FIR_filter_firBlock_left_N77,
my_FIR_filter_firBlock_left_N76, my_FIR_filter_firBlock_left_N75,
my_FIR_filter_firBlock_left_N74, my_FIR_filter_firBlock_left_N73,
my_FIR_filter_firBlock_left_N72, my_FIR_filter_firBlock_left_N71,
my_FIR_filter_firBlock_left_N70, my_FIR_filter_firBlock_left_N69,
my_FIR_filter_firBlock_left_N68, my_FIR_filter_firBlock_left_N67,
my_FIR_filter_firBlock_left_N66, my_FIR_filter_firBlock_left_N65,
my_FIR_filter_firBlock_left_N64, my_FIR_filter_firBlock_left_N63,
my_FIR_filter_firBlock_left_N62, my_FIR_filter_firBlock_left_N61,
my_FIR_filter_firBlock_left_N60, my_FIR_filter_firBlock_left_N59,
my_FIR_filter_firBlock_left_N58, my_FIR_filter_firBlock_left_N57,
my_FIR_filter_firBlock_left_N56, my_FIR_filter_firBlock_left_N55,
my_FIR_filter_firBlock_left_N54, my_FIR_filter_firBlock_left_N53,
my_FIR_filter_firBlock_left_N52, my_FIR_filter_firBlock_left_N51,
my_FIR_filter_firBlock_left_N50, my_FIR_filter_firBlock_left_N49,
my_FIR_filter_firBlock_left_N48, my_FIR_filter_firBlock_left_N47,
my_FIR_filter_firBlock_left_N46, my_FIR_filter_firBlock_left_N45,
my_FIR_filter_firBlock_left_N44, my_FIR_filter_firBlock_left_N43,
my_FIR_filter_firBlock_left_N42, my_FIR_filter_firBlock_left_N41,
my_FIR_filter_firBlock_left_N40, my_FIR_filter_firBlock_left_N39,
my_FIR_filter_firBlock_left_N38, my_FIR_filter_firBlock_left_N37,
my_FIR_filter_firBlock_left_N36, my_FIR_filter_firBlock_left_N35,
my_FIR_filter_firBlock_left_N34, my_FIR_filter_firBlock_left_N33,
my_FIR_filter_firBlock_left_N32, my_FIR_filter_firBlock_left_N31,
my_FIR_filter_firBlock_left_N30, my_FIR_filter_firBlock_left_N29,
my_FIR_filter_firBlock_left_N28, my_FIR_filter_firBlock_left_N27,
my_FIR_filter_firBlock_left_N26, my_FIR_filter_firBlock_left_N25,
my_FIR_filter_firBlock_left_N24, my_FIR_filter_firBlock_left_N23,
my_FIR_filter_firBlock_left_N22, my_FIR_filter_firBlock_left_N21,
my_FIR_filter_firBlock_left_N20, my_FIR_filter_firBlock_left_N19,
my_FIR_filter_firBlock_left_N18, my_FIR_filter_firBlock_left_N17,
my_FIR_filter_firBlock_left_N16, my_FIR_filter_firBlock_left_N15,
my_FIR_filter_firBlock_left_N14, my_FIR_filter_firBlock_left_N13,
my_FIR_filter_firBlock_left_N12, my_FIR_filter_firBlock_left_N11,
my_FIR_filter_firBlock_left_N10, my_FIR_filter_firBlock_left_N9,
my_FIR_filter_firBlock_left_N8, my_FIR_filter_firBlock_left_N7,
my_FIR_filter_firBlock_left_N6, my_FIR_filter_firBlock_left_N5,
my_FIR_filter_firBlock_left_N4, my_FIR_filter_firBlock_left_N3,
my_FIR_filter_firBlock_left_N2, my_FIR_filter_firBlock_left_N1,
my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_,
n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
n2303;
wire [5:1] inData_in;
wire [31:1] outData_in;
wire [31:0] leftOut;
wire [31:0] rightOut;
wire [287:0] my_FIR_filter_firBlock_left_firStep;
wire [114:0] my_FIR_filter_firBlock_left_multProducts;
wire [31:0] my_FIR_filter_firBlock_left_Y_in;
wire [38:6] my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192;
wire [31:0] my_FIR_filter_firBlock_right_multProducts;

dff inData_in_reg_31_ ( clk, n98_r, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, inData_31 );
not U_inv0 ( n17, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv1 ( n98_r, n98 );
dff inData_in_reg_16_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[100], inData_16 );
not U_inv2 ( n34, my_FIR_filter_firBlock_left_multProducts[100] );
not U_inv3 ( n97_r, n97 );
dff inData_in_reg_2_ ( clk, n95_r, inData_in[2], inData_2 );
not U_inv4 ( n20, inData_in[2] );
not U_inv5 ( n95_r, n95 );
dff inData_in_reg_0_ ( clk, n95_r, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[6], inData_0 );
not U_inv6 ( n19, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[6] );
not U_inv7 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__0_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[256], my_FIR_filter_firBlock_left_multProducts[90] );
not U_inv8 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__1_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[257], my_FIR_filter_firBlock_left_multProducts[91] );
not U_inv9 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__2_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[258], my_FIR_filter_firBlock_left_multProducts[92] );
not U_inv10 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__3_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[259], my_FIR_filter_firBlock_left_multProducts[93] );
not U_inv11 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__4_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[260], my_FIR_filter_firBlock_left_multProducts[94] );
not U_inv12 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__5_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[261], my_FIR_filter_firBlock_left_multProducts[95] );
not U_inv13 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__6_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[262], my_FIR_filter_firBlock_left_multProducts[96] );
not U_inv14 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__7_ ( clk, n95_r, my_FIR_filter_firBlock_left_firStep[263], my_FIR_filter_firBlock_left_multProducts[97] );
not U_inv15 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__8_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[264], my_FIR_filter_firBlock_left_multProducts[98] );
not U_inv16 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__9_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[265], my_FIR_filter_firBlock_left_multProducts[99] );
not U_inv17 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__10_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[266], my_FIR_filter_firBlock_left_multProducts[100] );
not U_inv18 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__11_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[267], my_FIR_filter_firBlock_left_multProducts[101] );
not U_inv19 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__12_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[268], my_FIR_filter_firBlock_left_multProducts[102] );
not U_inv20 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__13_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[269], my_FIR_filter_firBlock_left_multProducts[103] );
not U_inv21 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__14_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[270], my_FIR_filter_firBlock_left_multProducts[104] );
not U_inv22 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__15_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[271], my_FIR_filter_firBlock_left_multProducts[105] );
not U_inv23 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__16_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[272], my_FIR_filter_firBlock_left_multProducts[106] );
not U_inv24 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__17_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[273], my_FIR_filter_firBlock_left_multProducts[107] );
not U_inv25 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__18_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[274], my_FIR_filter_firBlock_left_multProducts[108] );
not U_inv26 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__19_ ( clk, n94_r, my_FIR_filter_firBlock_left_firStep[275], my_FIR_filter_firBlock_left_multProducts[109] );
not U_inv27 ( n94_r, n94 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__20_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[276], my_FIR_filter_firBlock_left_multProducts[110] );
not U_inv28 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__21_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[277], my_FIR_filter_firBlock_left_multProducts[111] );
not U_inv29 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__22_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[278], my_FIR_filter_firBlock_left_multProducts[112] );
not U_inv30 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__23_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[279], my_FIR_filter_firBlock_left_multProducts[113] );
not U_inv31 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__24_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[280], my_FIR_filter_firBlock_left_multProducts[114] );
not U_inv32 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__25_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[281], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv33 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__26_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[282], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv34 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__27_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[283], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv35 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__28_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[284], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv36 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__29_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[285], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv37 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__30_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[286], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv38 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_0__31_ ( clk, n93_r, my_FIR_filter_firBlock_left_firStep[287], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv39 ( n93_r, n93 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__0_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[224], my_FIR_filter_firBlock_left_N1 );
not U_inv40 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__1_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[225], my_FIR_filter_firBlock_left_N2 );
not U_inv41 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__2_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[226], my_FIR_filter_firBlock_left_N3 );
not U_inv42 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__3_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[227], my_FIR_filter_firBlock_left_N4 );
not U_inv43 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__4_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[228], my_FIR_filter_firBlock_left_N5 );
not U_inv44 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__5_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[229], my_FIR_filter_firBlock_left_N6 );
not U_inv45 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__6_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[230], my_FIR_filter_firBlock_left_N7 );
not U_inv46 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__7_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[231], my_FIR_filter_firBlock_left_N8 );
not U_inv47 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__8_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[232], my_FIR_filter_firBlock_left_N9 );
not U_inv48 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__9_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[233], my_FIR_filter_firBlock_left_N10 );
not U_inv49 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__10_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[234], my_FIR_filter_firBlock_left_N11 );
not U_inv50 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__11_ ( clk, n92_r, my_FIR_filter_firBlock_left_firStep[235], my_FIR_filter_firBlock_left_N12 );
not U_inv51 ( n92_r, n92 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__12_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[236], my_FIR_filter_firBlock_left_N13 );
not U_inv52 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__13_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[237], my_FIR_filter_firBlock_left_N14 );
not U_inv53 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__14_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[238], my_FIR_filter_firBlock_left_N15 );
not U_inv54 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__15_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[239], my_FIR_filter_firBlock_left_N16 );
not U_inv55 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__16_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[240], my_FIR_filter_firBlock_left_N17 );
not U_inv56 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__17_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[241], my_FIR_filter_firBlock_left_N18 );
not U_inv57 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__18_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[242], my_FIR_filter_firBlock_left_N19 );
not U_inv58 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__19_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[243], my_FIR_filter_firBlock_left_N20 );
not U_inv59 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__20_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[244], my_FIR_filter_firBlock_left_N21 );
not U_inv60 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__21_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[245], my_FIR_filter_firBlock_left_N22 );
not U_inv61 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__22_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[246], my_FIR_filter_firBlock_left_N23 );
not U_inv62 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__23_ ( clk, n91_r, my_FIR_filter_firBlock_left_firStep[247], my_FIR_filter_firBlock_left_N24 );
not U_inv63 ( n91_r, n91 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__24_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[248], my_FIR_filter_firBlock_left_N25 );
not U_inv64 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__25_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[249], my_FIR_filter_firBlock_left_N26 );
not U_inv65 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__26_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[250], my_FIR_filter_firBlock_left_N27 );
not U_inv66 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__27_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[251], my_FIR_filter_firBlock_left_N28 );
not U_inv67 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__28_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[252], my_FIR_filter_firBlock_left_N29 );
not U_inv68 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__29_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[253], my_FIR_filter_firBlock_left_N30 );
not U_inv69 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__30_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[254], my_FIR_filter_firBlock_left_N31 );
not U_inv70 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__0_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[192], my_FIR_filter_firBlock_left_N33 );
not U_inv71 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__1_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[193], my_FIR_filter_firBlock_left_N34 );
not U_inv72 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__2_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[194], my_FIR_filter_firBlock_left_N35 );
not U_inv73 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__3_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[195], my_FIR_filter_firBlock_left_N36 );
not U_inv74 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__4_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[196], my_FIR_filter_firBlock_left_N37 );
not U_inv75 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__5_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[197], my_FIR_filter_firBlock_left_N38 );
not U_inv76 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__6_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[198], my_FIR_filter_firBlock_left_N39 );
not U_inv77 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__7_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[199], my_FIR_filter_firBlock_left_N40 );
not U_inv78 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__8_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[200], my_FIR_filter_firBlock_left_N41 );
not U_inv79 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__9_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[201], my_FIR_filter_firBlock_left_N42 );
not U_inv80 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__10_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[202], my_FIR_filter_firBlock_left_N43 );
not U_inv81 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__11_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[203], my_FIR_filter_firBlock_left_N44 );
not U_inv82 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__12_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[204], my_FIR_filter_firBlock_left_N45 );
not U_inv83 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__13_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[205], my_FIR_filter_firBlock_left_N46 );
not U_inv84 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__14_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[206], my_FIR_filter_firBlock_left_N47 );
not U_inv85 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__15_ ( clk, n89_r, my_FIR_filter_firBlock_left_firStep[207], my_FIR_filter_firBlock_left_N48 );
not U_inv86 ( n89_r, n89 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__16_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[208], my_FIR_filter_firBlock_left_N49 );
not U_inv87 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__17_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[209], my_FIR_filter_firBlock_left_N50 );
not U_inv88 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__18_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[210], my_FIR_filter_firBlock_left_N51 );
not U_inv89 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__19_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[211], my_FIR_filter_firBlock_left_N52 );
not U_inv90 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__20_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[212], my_FIR_filter_firBlock_left_N53 );
not U_inv91 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__21_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[213], my_FIR_filter_firBlock_left_N54 );
not U_inv92 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__22_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[214], my_FIR_filter_firBlock_left_N55 );
not U_inv93 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__23_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[215], my_FIR_filter_firBlock_left_N56 );
not U_inv94 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__24_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[216], my_FIR_filter_firBlock_left_N57 );
not U_inv95 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__25_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[217], my_FIR_filter_firBlock_left_N58 );
not U_inv96 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__26_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[218], my_FIR_filter_firBlock_left_N59 );
not U_inv97 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__27_ ( clk, n88_r, my_FIR_filter_firBlock_left_firStep[219], my_FIR_filter_firBlock_left_N60 );
not U_inv98 ( n88_r, n88 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__28_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[220], my_FIR_filter_firBlock_left_N61 );
not U_inv99 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__29_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[221], my_FIR_filter_firBlock_left_N62 );
not U_inv100 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__30_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[222], my_FIR_filter_firBlock_left_N63 );
not U_inv101 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_2__31_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[223], my_FIR_filter_firBlock_left_N64 );
not U_inv102 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__0_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[160], my_FIR_filter_firBlock_left_N65 );
not U_inv103 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__1_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[161], my_FIR_filter_firBlock_left_N66 );
not U_inv104 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__2_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[162], my_FIR_filter_firBlock_left_N67 );
not U_inv105 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__3_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[163], my_FIR_filter_firBlock_left_N68 );
not U_inv106 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__4_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[164], my_FIR_filter_firBlock_left_N69 );
not U_inv107 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__5_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[165], my_FIR_filter_firBlock_left_N70 );
not U_inv108 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__6_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[166], my_FIR_filter_firBlock_left_N71 );
not U_inv109 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__7_ ( clk, n87_r, my_FIR_filter_firBlock_left_firStep[167], my_FIR_filter_firBlock_left_N72 );
not U_inv110 ( n87_r, n87 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__8_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[168], my_FIR_filter_firBlock_left_N73 );
not U_inv111 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__9_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[169], my_FIR_filter_firBlock_left_N74 );
not U_inv112 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__10_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[170], my_FIR_filter_firBlock_left_N75 );
not U_inv113 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__11_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[171], my_FIR_filter_firBlock_left_N76 );
not U_inv114 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__12_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[172], my_FIR_filter_firBlock_left_N77 );
not U_inv115 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__13_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[173], my_FIR_filter_firBlock_left_N78 );
not U_inv116 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__14_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[174], my_FIR_filter_firBlock_left_N79 );
not U_inv117 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__15_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[175], my_FIR_filter_firBlock_left_N80 );
not U_inv118 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__16_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[176], my_FIR_filter_firBlock_left_N81 );
not U_inv119 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__17_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[177], my_FIR_filter_firBlock_left_N82 );
not U_inv120 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__18_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[178], my_FIR_filter_firBlock_left_N83 );
not U_inv121 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__19_ ( clk, n86_r, my_FIR_filter_firBlock_left_firStep[179], my_FIR_filter_firBlock_left_N84 );
not U_inv122 ( n86_r, n86 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__20_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[180], my_FIR_filter_firBlock_left_N85 );
not U_inv123 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__21_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[181], my_FIR_filter_firBlock_left_N86 );
not U_inv124 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__22_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[182], my_FIR_filter_firBlock_left_N87 );
not U_inv125 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__23_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[183], my_FIR_filter_firBlock_left_N88 );
not U_inv126 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__24_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[184], my_FIR_filter_firBlock_left_N89 );
not U_inv127 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__25_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[185], my_FIR_filter_firBlock_left_N90 );
not U_inv128 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__26_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[186], my_FIR_filter_firBlock_left_N91 );
not U_inv129 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__27_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[187], my_FIR_filter_firBlock_left_N92 );
not U_inv130 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__28_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[188], my_FIR_filter_firBlock_left_N93 );
not U_inv131 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__29_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[189], my_FIR_filter_firBlock_left_N94 );
not U_inv132 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__30_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[190], my_FIR_filter_firBlock_left_N95 );
not U_inv133 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_3__31_ ( clk, n85_r, my_FIR_filter_firBlock_left_firStep[191], my_FIR_filter_firBlock_left_N96 );
not U_inv134 ( n85_r, n85 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__0_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[128], my_FIR_filter_firBlock_left_N97 );
not U_inv135 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__1_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[129], my_FIR_filter_firBlock_left_N98 );
not U_inv136 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__2_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[130], my_FIR_filter_firBlock_left_N99 );
not U_inv137 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__3_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[131], my_FIR_filter_firBlock_left_N100 );
not U_inv138 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__4_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[132], my_FIR_filter_firBlock_left_N101 );
not U_inv139 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__5_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[133], my_FIR_filter_firBlock_left_N102 );
not U_inv140 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__6_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[134], my_FIR_filter_firBlock_left_N103 );
not U_inv141 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__7_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[135], my_FIR_filter_firBlock_left_N104 );
not U_inv142 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__8_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[136], my_FIR_filter_firBlock_left_N105 );
not U_inv143 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__9_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[137], my_FIR_filter_firBlock_left_N106 );
not U_inv144 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__10_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[138], my_FIR_filter_firBlock_left_N107 );
not U_inv145 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__11_ ( clk, n84_r, my_FIR_filter_firBlock_left_firStep[139], my_FIR_filter_firBlock_left_N108 );
not U_inv146 ( n84_r, n84 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__12_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[140], my_FIR_filter_firBlock_left_N109 );
not U_inv147 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__13_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[141], my_FIR_filter_firBlock_left_N110 );
not U_inv148 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__14_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[142], my_FIR_filter_firBlock_left_N111 );
not U_inv149 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__15_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[143], my_FIR_filter_firBlock_left_N112 );
not U_inv150 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__16_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[144], my_FIR_filter_firBlock_left_N113 );
not U_inv151 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__17_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[145], my_FIR_filter_firBlock_left_N114 );
not U_inv152 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__18_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[146], my_FIR_filter_firBlock_left_N115 );
not U_inv153 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__19_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[147], my_FIR_filter_firBlock_left_N116 );
not U_inv154 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__20_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[148], my_FIR_filter_firBlock_left_N117 );
not U_inv155 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__21_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[149], my_FIR_filter_firBlock_left_N118 );
not U_inv156 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__22_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[150], my_FIR_filter_firBlock_left_N119 );
not U_inv157 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__23_ ( clk, n83_r, my_FIR_filter_firBlock_left_firStep[151], my_FIR_filter_firBlock_left_N120 );
not U_inv158 ( n83_r, n83 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__24_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[152], my_FIR_filter_firBlock_left_N121 );
not U_inv159 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__25_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[153], my_FIR_filter_firBlock_left_N122 );
not U_inv160 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__26_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[154], my_FIR_filter_firBlock_left_N123 );
not U_inv161 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__27_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[155], my_FIR_filter_firBlock_left_N124 );
not U_inv162 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__28_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[156], my_FIR_filter_firBlock_left_N125 );
not U_inv163 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__29_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[157], my_FIR_filter_firBlock_left_N126 );
not U_inv164 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__30_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[158], my_FIR_filter_firBlock_left_N127 );
not U_inv165 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_4__31_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[159], my_FIR_filter_firBlock_left_N128 );
not U_inv166 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__0_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[96], my_FIR_filter_firBlock_left_N129 );
not U_inv167 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__1_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[97], my_FIR_filter_firBlock_left_N130 );
not U_inv168 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__2_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[98], my_FIR_filter_firBlock_left_N131 );
not U_inv169 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__3_ ( clk, n82_r, my_FIR_filter_firBlock_left_firStep[99], my_FIR_filter_firBlock_left_N132 );
not U_inv170 ( n82_r, n82 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__4_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[100], my_FIR_filter_firBlock_left_N133 );
not U_inv171 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__5_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[101], my_FIR_filter_firBlock_left_N134 );
not U_inv172 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__6_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[102], my_FIR_filter_firBlock_left_N135 );
not U_inv173 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__7_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[103], my_FIR_filter_firBlock_left_N136 );
not U_inv174 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__8_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[104], my_FIR_filter_firBlock_left_N137 );
not U_inv175 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__9_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[105], my_FIR_filter_firBlock_left_N138 );
not U_inv176 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__10_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[106], my_FIR_filter_firBlock_left_N139 );
not U_inv177 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__11_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[107], my_FIR_filter_firBlock_left_N140 );
not U_inv178 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__12_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[108], my_FIR_filter_firBlock_left_N141 );
not U_inv179 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__13_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[109], my_FIR_filter_firBlock_left_N142 );
not U_inv180 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__14_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[110], my_FIR_filter_firBlock_left_N143 );
not U_inv181 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__15_ ( clk, n81_r, my_FIR_filter_firBlock_left_firStep[111], my_FIR_filter_firBlock_left_N144 );
not U_inv182 ( n81_r, n81 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__16_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[112], my_FIR_filter_firBlock_left_N145 );
not U_inv183 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__17_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[113], my_FIR_filter_firBlock_left_N146 );
not U_inv184 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__18_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[114], my_FIR_filter_firBlock_left_N147 );
not U_inv185 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__19_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[115], my_FIR_filter_firBlock_left_N148 );
not U_inv186 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__20_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[116], my_FIR_filter_firBlock_left_N149 );
not U_inv187 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__21_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[117], my_FIR_filter_firBlock_left_N150 );
not U_inv188 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__22_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[118], my_FIR_filter_firBlock_left_N151 );
not U_inv189 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__23_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[119], my_FIR_filter_firBlock_left_N152 );
not U_inv190 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__24_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[120], my_FIR_filter_firBlock_left_N153 );
not U_inv191 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__25_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[121], my_FIR_filter_firBlock_left_N154 );
not U_inv192 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__26_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[122], my_FIR_filter_firBlock_left_N155 );
not U_inv193 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__27_ ( clk, n80_r, my_FIR_filter_firBlock_left_firStep[123], my_FIR_filter_firBlock_left_N156 );
not U_inv194 ( n80_r, n80 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__28_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[124], my_FIR_filter_firBlock_left_N157 );
not U_inv195 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__29_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[125], my_FIR_filter_firBlock_left_N158 );
not U_inv196 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__30_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[126], my_FIR_filter_firBlock_left_N159 );
not U_inv197 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_5__31_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[127], my_FIR_filter_firBlock_left_N160 );
not U_inv198 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__0_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[64], my_FIR_filter_firBlock_left_N161 );
not U_inv199 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__1_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[65], my_FIR_filter_firBlock_left_N162 );
not U_inv200 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__2_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[66], my_FIR_filter_firBlock_left_N163 );
not U_inv201 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__3_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[67], my_FIR_filter_firBlock_left_N164 );
not U_inv202 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__4_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[68], my_FIR_filter_firBlock_left_N165 );
not U_inv203 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__5_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[69], my_FIR_filter_firBlock_left_N166 );
not U_inv204 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__6_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[70], my_FIR_filter_firBlock_left_N167 );
not U_inv205 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__7_ ( clk, n79_r, my_FIR_filter_firBlock_left_firStep[71], my_FIR_filter_firBlock_left_N168 );
not U_inv206 ( n79_r, n79 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__8_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[72], my_FIR_filter_firBlock_left_N169 );
not U_inv207 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__9_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[73], my_FIR_filter_firBlock_left_N170 );
not U_inv208 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__10_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[74], my_FIR_filter_firBlock_left_N171 );
not U_inv209 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__11_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[75], my_FIR_filter_firBlock_left_N172 );
not U_inv210 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__12_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[76], my_FIR_filter_firBlock_left_N173 );
not U_inv211 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__13_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[77], my_FIR_filter_firBlock_left_N174 );
not U_inv212 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__14_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[78], my_FIR_filter_firBlock_left_N175 );
not U_inv213 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__15_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[79], my_FIR_filter_firBlock_left_N176 );
not U_inv214 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__16_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[80], my_FIR_filter_firBlock_left_N177 );
not U_inv215 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__17_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[81], my_FIR_filter_firBlock_left_N178 );
not U_inv216 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__18_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[82], my_FIR_filter_firBlock_left_N179 );
not U_inv217 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__19_ ( clk, n78_r, my_FIR_filter_firBlock_left_firStep[83], my_FIR_filter_firBlock_left_N180 );
not U_inv218 ( n78_r, n78 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__20_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[84], my_FIR_filter_firBlock_left_N181 );
not U_inv219 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__21_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[85], my_FIR_filter_firBlock_left_N182 );
not U_inv220 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__22_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[86], my_FIR_filter_firBlock_left_N183 );
not U_inv221 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__23_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[87], my_FIR_filter_firBlock_left_N184 );
not U_inv222 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__24_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[88], my_FIR_filter_firBlock_left_N185 );
not U_inv223 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__25_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[89], my_FIR_filter_firBlock_left_N186 );
not U_inv224 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__26_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[90], my_FIR_filter_firBlock_left_N187 );
not U_inv225 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__27_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[91], my_FIR_filter_firBlock_left_N188 );
not U_inv226 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__28_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[92], my_FIR_filter_firBlock_left_N189 );
not U_inv227 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__29_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[93], my_FIR_filter_firBlock_left_N190 );
not U_inv228 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__30_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[94], my_FIR_filter_firBlock_left_N191 );
not U_inv229 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_6__31_ ( clk, n77_r, my_FIR_filter_firBlock_left_firStep[95], my_FIR_filter_firBlock_left_N192 );
not U_inv230 ( n77_r, n77 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__0_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[32], my_FIR_filter_firBlock_left_N193 );
not U_inv231 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__1_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[33], my_FIR_filter_firBlock_left_N194 );
not U_inv232 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__2_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[34], my_FIR_filter_firBlock_left_N195 );
not U_inv233 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__3_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[35], my_FIR_filter_firBlock_left_N196 );
not U_inv234 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__4_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[36], my_FIR_filter_firBlock_left_N197 );
not U_inv235 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__5_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[37], my_FIR_filter_firBlock_left_N198 );
not U_inv236 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__6_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[38], my_FIR_filter_firBlock_left_N199 );
not U_inv237 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__7_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[39], my_FIR_filter_firBlock_left_N200 );
not U_inv238 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__8_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[40], my_FIR_filter_firBlock_left_N201 );
not U_inv239 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__9_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[41], my_FIR_filter_firBlock_left_N202 );
not U_inv240 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__10_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[42], my_FIR_filter_firBlock_left_N203 );
not U_inv241 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__11_ ( clk, n76_r, my_FIR_filter_firBlock_left_firStep[43], my_FIR_filter_firBlock_left_N204 );
not U_inv242 ( n76_r, n76 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__12_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[44], my_FIR_filter_firBlock_left_N205 );
not U_inv243 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__13_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[45], my_FIR_filter_firBlock_left_N206 );
not U_inv244 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__14_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[46], my_FIR_filter_firBlock_left_N207 );
not U_inv245 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__15_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[47], my_FIR_filter_firBlock_left_N208 );
not U_inv246 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__16_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[48], my_FIR_filter_firBlock_left_N209 );
not U_inv247 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__17_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[49], my_FIR_filter_firBlock_left_N210 );
not U_inv248 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__18_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[50], my_FIR_filter_firBlock_left_N211 );
not U_inv249 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__19_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[51], my_FIR_filter_firBlock_left_N212 );
not U_inv250 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__20_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[52], my_FIR_filter_firBlock_left_N213 );
not U_inv251 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__21_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[53], my_FIR_filter_firBlock_left_N214 );
not U_inv252 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__22_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[54], my_FIR_filter_firBlock_left_N215 );
not U_inv253 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__23_ ( clk, n75_r, my_FIR_filter_firBlock_left_firStep[55], my_FIR_filter_firBlock_left_N216 );
not U_inv254 ( n75_r, n75 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__24_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[56], my_FIR_filter_firBlock_left_N217 );
not U_inv255 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__25_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[57], my_FIR_filter_firBlock_left_N218 );
not U_inv256 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__26_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[58], my_FIR_filter_firBlock_left_N219 );
not U_inv257 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__27_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[59], my_FIR_filter_firBlock_left_N220 );
not U_inv258 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__28_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[60], my_FIR_filter_firBlock_left_N221 );
not U_inv259 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__29_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[61], my_FIR_filter_firBlock_left_N222 );
not U_inv260 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__30_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[62], my_FIR_filter_firBlock_left_N223 );
not U_inv261 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_7__31_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[63], my_FIR_filter_firBlock_left_N224 );
not U_inv262 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__0_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[0], my_FIR_filter_firBlock_left_N225 );
not U_inv263 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__1_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[1], my_FIR_filter_firBlock_left_N226 );
not U_inv264 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__2_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[2], my_FIR_filter_firBlock_left_N227 );
not U_inv265 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__3_ ( clk, n74_r, my_FIR_filter_firBlock_left_firStep[3], my_FIR_filter_firBlock_left_N228 );
not U_inv266 ( n74_r, n74 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__4_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[4], my_FIR_filter_firBlock_left_N229 );
not U_inv267 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__5_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[5], my_FIR_filter_firBlock_left_N230 );
not U_inv268 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__6_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[6], my_FIR_filter_firBlock_left_N231 );
not U_inv269 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__7_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[7], my_FIR_filter_firBlock_left_N232 );
not U_inv270 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__8_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[8], my_FIR_filter_firBlock_left_N233 );
not U_inv271 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__9_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[9], my_FIR_filter_firBlock_left_N234 );
not U_inv272 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__10_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[10], my_FIR_filter_firBlock_left_N235 );
not U_inv273 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__11_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[11], my_FIR_filter_firBlock_left_N236 );
not U_inv274 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__12_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[12], my_FIR_filter_firBlock_left_N237 );
not U_inv275 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__13_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[13], my_FIR_filter_firBlock_left_N238 );
not U_inv276 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__14_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[14], my_FIR_filter_firBlock_left_N239 );
not U_inv277 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__15_ ( clk, n73_r, my_FIR_filter_firBlock_left_firStep[15], my_FIR_filter_firBlock_left_N240 );
not U_inv278 ( n73_r, n73 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__16_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[16], my_FIR_filter_firBlock_left_N241 );
not U_inv279 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__17_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[17], my_FIR_filter_firBlock_left_N242 );
not U_inv280 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__18_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[18], my_FIR_filter_firBlock_left_N243 );
not U_inv281 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__19_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[19], my_FIR_filter_firBlock_left_N244 );
not U_inv282 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__20_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[20], my_FIR_filter_firBlock_left_N245 );
not U_inv283 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__21_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[21], my_FIR_filter_firBlock_left_N246 );
not U_inv284 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__22_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[22], my_FIR_filter_firBlock_left_N247 );
not U_inv285 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__23_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[23], my_FIR_filter_firBlock_left_N248 );
not U_inv286 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__24_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[24], my_FIR_filter_firBlock_left_N249 );
not U_inv287 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__25_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[25], my_FIR_filter_firBlock_left_N250 );
not U_inv288 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__26_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[26], my_FIR_filter_firBlock_left_N251 );
not U_inv289 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__27_ ( clk, n72_r, my_FIR_filter_firBlock_left_firStep[27], my_FIR_filter_firBlock_left_N252 );
not U_inv290 ( n72_r, n72 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__28_ ( clk, n71_r, my_FIR_filter_firBlock_left_firStep[28], my_FIR_filter_firBlock_left_N253 );
not U_inv291 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__29_ ( clk, n71_r, my_FIR_filter_firBlock_left_firStep[29], my_FIR_filter_firBlock_left_N254 );
not U_inv292 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__30_ ( clk, n71_r, my_FIR_filter_firBlock_left_firStep[30], my_FIR_filter_firBlock_left_N255 );
not U_inv293 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__0_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[0], my_FIR_filter_firBlock_left_N257 );
not U_inv294 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__1_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[1], my_FIR_filter_firBlock_left_N258 );
not U_inv295 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__2_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[2], my_FIR_filter_firBlock_left_N259 );
not U_inv296 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__3_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[3], my_FIR_filter_firBlock_left_N260 );
not U_inv297 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__4_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[4], my_FIR_filter_firBlock_left_N261 );
not U_inv298 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__5_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[5], my_FIR_filter_firBlock_left_N262 );
not U_inv299 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__6_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[6], my_FIR_filter_firBlock_left_N263 );
not U_inv300 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__7_ ( clk, n71_r, my_FIR_filter_firBlock_left_Y_in[7], my_FIR_filter_firBlock_left_N264 );
not U_inv301 ( n71_r, n71 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__8_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[8], my_FIR_filter_firBlock_left_N265 );
not U_inv302 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__9_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[9], my_FIR_filter_firBlock_left_N266 );
not U_inv303 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__10_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[10], my_FIR_filter_firBlock_left_N267 );
not U_inv304 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__11_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[11], my_FIR_filter_firBlock_left_N268 );
not U_inv305 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__12_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[12], my_FIR_filter_firBlock_left_N269 );
not U_inv306 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__13_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[13], my_FIR_filter_firBlock_left_N270 );
not U_inv307 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__14_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[14], my_FIR_filter_firBlock_left_N271 );
not U_inv308 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__15_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[15], my_FIR_filter_firBlock_left_N272 );
not U_inv309 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__16_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[16], my_FIR_filter_firBlock_left_N273 );
not U_inv310 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__17_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[17], my_FIR_filter_firBlock_left_N274 );
not U_inv311 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__18_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[18], my_FIR_filter_firBlock_left_N275 );
not U_inv312 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__19_ ( clk, n70_r, my_FIR_filter_firBlock_left_Y_in[19], my_FIR_filter_firBlock_left_N276 );
not U_inv313 ( n70_r, n70 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__20_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[20], my_FIR_filter_firBlock_left_N277 );
not U_inv314 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__21_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[21], my_FIR_filter_firBlock_left_N278 );
not U_inv315 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__22_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[22], my_FIR_filter_firBlock_left_N279 );
not U_inv316 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__23_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[23], my_FIR_filter_firBlock_left_N280 );
not U_inv317 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__24_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[24], my_FIR_filter_firBlock_left_N281 );
not U_inv318 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__25_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[25], my_FIR_filter_firBlock_left_N282 );
not U_inv319 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__26_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[26], my_FIR_filter_firBlock_left_N283 );
not U_inv320 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__27_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[27], my_FIR_filter_firBlock_left_N284 );
not U_inv321 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__28_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[28], my_FIR_filter_firBlock_left_N285 );
not U_inv322 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__29_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[29], my_FIR_filter_firBlock_left_N286 );
not U_inv323 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__30_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[30], my_FIR_filter_firBlock_left_N287 );
not U_inv324 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_firStep_reg_9__31_ ( clk, n69_r, my_FIR_filter_firBlock_left_Y_in[31], my_FIR_filter_firBlock_left_N288 );
not U_inv325 ( n69_r, n69 );
dff my_FIR_filter_firBlock_left_Y_reg_0_ ( clk, n68_r, leftOut[0], my_FIR_filter_firBlock_left_Y_in[0] );
not U_inv326 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_1_ ( clk, n68_r, leftOut[1], my_FIR_filter_firBlock_left_Y_in[1] );
not U_inv327 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_2_ ( clk, n68_r, leftOut[2], my_FIR_filter_firBlock_left_Y_in[2] );
not U_inv328 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_3_ ( clk, n68_r, leftOut[3], my_FIR_filter_firBlock_left_Y_in[3] );
not U_inv329 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_4_ ( clk, n68_r, leftOut[4], my_FIR_filter_firBlock_left_Y_in[4] );
not U_inv330 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_5_ ( clk, n68_r, leftOut[5], my_FIR_filter_firBlock_left_Y_in[5] );
not U_inv331 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_6_ ( clk, n68_r, leftOut[6], my_FIR_filter_firBlock_left_Y_in[6] );
not U_inv332 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_7_ ( clk, n68_r, leftOut[7], my_FIR_filter_firBlock_left_Y_in[7] );
not U_inv333 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_8_ ( clk, n68_r, leftOut[8], my_FIR_filter_firBlock_left_Y_in[8] );
not U_inv334 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_9_ ( clk, n68_r, leftOut[9], my_FIR_filter_firBlock_left_Y_in[9] );
not U_inv335 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_10_ ( clk, n68_r, leftOut[10], my_FIR_filter_firBlock_left_Y_in[10] );
not U_inv336 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_11_ ( clk, n68_r, leftOut[11], my_FIR_filter_firBlock_left_Y_in[11] );
not U_inv337 ( n68_r, n68 );
dff my_FIR_filter_firBlock_left_Y_reg_12_ ( clk, n67_r, leftOut[12], my_FIR_filter_firBlock_left_Y_in[12] );
not U_inv338 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_13_ ( clk, n67_r, leftOut[13], my_FIR_filter_firBlock_left_Y_in[13] );
not U_inv339 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_14_ ( clk, n67_r, leftOut[14], my_FIR_filter_firBlock_left_Y_in[14] );
not U_inv340 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_15_ ( clk, n67_r, leftOut[15], my_FIR_filter_firBlock_left_Y_in[15] );
not U_inv341 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_16_ ( clk, n67_r, leftOut[16], my_FIR_filter_firBlock_left_Y_in[16] );
not U_inv342 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_17_ ( clk, n67_r, leftOut[17], my_FIR_filter_firBlock_left_Y_in[17] );
not U_inv343 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_18_ ( clk, n67_r, leftOut[18], my_FIR_filter_firBlock_left_Y_in[18] );
not U_inv344 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_19_ ( clk, n67_r, leftOut[19], my_FIR_filter_firBlock_left_Y_in[19] );
not U_inv345 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_20_ ( clk, n67_r, leftOut[20], my_FIR_filter_firBlock_left_Y_in[20] );
not U_inv346 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_21_ ( clk, n67_r, leftOut[21], my_FIR_filter_firBlock_left_Y_in[21] );
not U_inv347 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_22_ ( clk, n67_r, leftOut[22], my_FIR_filter_firBlock_left_Y_in[22] );
not U_inv348 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_23_ ( clk, n67_r, leftOut[23], my_FIR_filter_firBlock_left_Y_in[23] );
not U_inv349 ( n67_r, n67 );
dff my_FIR_filter_firBlock_left_Y_reg_24_ ( clk, n66_r, leftOut[24], my_FIR_filter_firBlock_left_Y_in[24] );
not U_inv350 ( n66_r, n66 );
dff my_FIR_filter_firBlock_left_Y_reg_25_ ( clk, n66_r, leftOut[25], my_FIR_filter_firBlock_left_Y_in[25] );
not U_inv351 ( n66_r, n66 );
dff my_FIR_filter_firBlock_left_Y_reg_26_ ( clk, n66_r, leftOut[26], my_FIR_filter_firBlock_left_Y_in[26] );
not U_inv352 ( n66_r, n66 );
dff my_FIR_filter_firBlock_left_Y_reg_27_ ( clk, n66_r, leftOut[27], my_FIR_filter_firBlock_left_Y_in[27] );
not U_inv353 ( n66_r, n66 );
dff my_FIR_filter_firBlock_left_Y_reg_28_ ( clk, n66_r, leftOut[28], my_FIR_filter_firBlock_left_Y_in[28] );
not U_inv354 ( n66_r, n66 );
dff my_FIR_filter_firBlock_left_Y_reg_29_ ( clk, n66_r, leftOut[29], my_FIR_filter_firBlock_left_Y_in[29] );
not U_inv355 ( n66_r, n66 );
dff my_FIR_filter_firBlock_left_Y_reg_30_ ( clk, n66_r, leftOut[30], my_FIR_filter_firBlock_left_Y_in[30] );
not U_inv356 ( n66_r, n66 );
dff my_FIR_filter_firBlock_left_Y_reg_31_ ( clk, n66_r, leftOut[31], my_FIR_filter_firBlock_left_Y_in[31] );
not U_inv357 ( n66_r, n66 );
dff my_FIR_filter_firBlock_right_Y_reg_31_ ( clk, n66_r, rightOut[31], my_FIR_filter_firBlock_right_multProducts[31] );
not U_inv358 ( n66_r, n66 );
dff outData_reg_0_ ( clk, n66_r, outData_0, my_FIR_filter_firBlock_right_multProducts[0] );
not U_inv359 ( n66_r, n66 );
dff outData_reg_1_ ( clk, n66_r, outData_1, outData_in[1] );
not U_inv360 ( n66_r, n66 );
dff outData_reg_2_ ( clk, n66_r, outData_2, outData_in[2] );
not U_inv361 ( n66_r, n66 );
dff outData_reg_3_ ( clk, n65_r, outData_3, outData_in[3] );
not U_inv362 ( n65_r, n65 );
dff outData_reg_4_ ( clk, n65_r, outData_4, outData_in[4] );
not U_inv363 ( n65_r, n65 );
dff outData_reg_5_ ( clk, n65_r, outData_5, outData_in[5] );
not U_inv364 ( n65_r, n65 );
dff outData_reg_6_ ( clk, n65_r, outData_6, outData_in[6] );
not U_inv365 ( n65_r, n65 );
dff outData_reg_7_ ( clk, n65_r, outData_7, outData_in[7] );
not U_inv366 ( n65_r, n65 );
dff outData_reg_8_ ( clk, n65_r, outData_8, outData_in[8] );
not U_inv367 ( n65_r, n65 );
dff outData_reg_9_ ( clk, n65_r, outData_9, outData_in[9] );
not U_inv368 ( n65_r, n65 );
dff outData_reg_10_ ( clk, n65_r, outData_10, outData_in[10] );
not U_inv369 ( n65_r, n65 );
dff outData_reg_11_ ( clk, n65_r, outData_11, outData_in[11] );
not U_inv370 ( n65_r, n65 );
dff outData_reg_12_ ( clk, n65_r, outData_12, outData_in[12] );
not U_inv371 ( n65_r, n65 );
dff outData_reg_13_ ( clk, n65_r, outData_13, outData_in[13] );
not U_inv372 ( n65_r, n65 );
dff outData_reg_14_ ( clk, n65_r, outData_14, outData_in[14] );
not U_inv373 ( n65_r, n65 );
dff outData_reg_15_ ( clk, n64_r, outData_15, outData_in[15] );
not U_inv374 ( n64_r, n64 );
dff outData_reg_16_ ( clk, n64_r, outData_16, outData_in[16] );
not U_inv375 ( n64_r, n64 );
dff outData_reg_17_ ( clk, n64_r, outData_17, outData_in[17] );
not U_inv376 ( n64_r, n64 );
dff outData_reg_18_ ( clk, n64_r, outData_18, outData_in[18] );
not U_inv377 ( n64_r, n64 );
dff outData_reg_19_ ( clk, n64_r, outData_19, outData_in[19] );
not U_inv378 ( n64_r, n64 );
dff outData_reg_20_ ( clk, n64_r, outData_20, outData_in[20] );
not U_inv379 ( n64_r, n64 );
dff outData_reg_21_ ( clk, n64_r, outData_21, outData_in[21] );
not U_inv380 ( n64_r, n64 );
dff outData_reg_22_ ( clk, n64_r, outData_22, outData_in[22] );
not U_inv381 ( n64_r, n64 );
dff outData_reg_23_ ( clk, n64_r, outData_23, outData_in[23] );
not U_inv382 ( n64_r, n64 );
dff outData_reg_24_ ( clk, n64_r, outData_24, outData_in[24] );
not U_inv383 ( n64_r, n64 );
dff outData_reg_25_ ( clk, n64_r, outData_25, outData_in[25] );
not U_inv384 ( n64_r, n64 );
dff outData_reg_26_ ( clk, n64_r, outData_26, outData_in[26] );
not U_inv385 ( n64_r, n64 );
dff outData_reg_27_ ( clk, n63_r, outData_27, outData_in[27] );
not U_inv386 ( n63_r, n63 );
dff outData_reg_28_ ( clk, n63_r, outData_28, outData_in[28] );
not U_inv387 ( n63_r, n63 );
dff outData_reg_29_ ( clk, n63_r, outData_29, outData_in[29] );
not U_inv388 ( n63_r, n63 );
dff outData_reg_30_ ( clk, n63_r, outData_30, outData_in[30] );
not U_inv389 ( n63_r, n63 );
dff outData_reg_31_ ( clk, n63_r, outData_31, outData_in[31] );
not U_inv390 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_0_ ( clk, n63_r, rightOut[0], my_FIR_filter_firBlock_right_multProducts[0] );
not U_inv391 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_1_ ( clk, n63_r, rightOut[1], my_FIR_filter_firBlock_right_multProducts[1] );
not U_inv392 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_2_ ( clk, n63_r, rightOut[2], my_FIR_filter_firBlock_right_multProducts[2] );
not U_inv393 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_3_ ( clk, n63_r, rightOut[3], my_FIR_filter_firBlock_right_multProducts[3] );
not U_inv394 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_4_ ( clk, n63_r, rightOut[4], my_FIR_filter_firBlock_right_multProducts[4] );
not U_inv395 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_5_ ( clk, n63_r, rightOut[5], my_FIR_filter_firBlock_right_multProducts[5] );
not U_inv396 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_6_ ( clk, n63_r, rightOut[6], my_FIR_filter_firBlock_right_multProducts[6] );
not U_inv397 ( n63_r, n63 );
dff my_FIR_filter_firBlock_right_Y_reg_7_ ( clk, n62_r, rightOut[7], my_FIR_filter_firBlock_right_multProducts[7] );
not U_inv398 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_8_ ( clk, n62_r, rightOut[8], my_FIR_filter_firBlock_right_multProducts[8] );
not U_inv399 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_9_ ( clk, n62_r, rightOut[9], my_FIR_filter_firBlock_right_multProducts[9] );
not U_inv400 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_10_ ( clk, n62_r, rightOut[10], my_FIR_filter_firBlock_right_multProducts[10] );
not U_inv401 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_11_ ( clk, n62_r, rightOut[11], my_FIR_filter_firBlock_right_multProducts[11] );
not U_inv402 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_12_ ( clk, n62_r, rightOut[12], my_FIR_filter_firBlock_right_multProducts[12] );
not U_inv403 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_13_ ( clk, n62_r, rightOut[13], my_FIR_filter_firBlock_right_multProducts[13] );
not U_inv404 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_14_ ( clk, n62_r, rightOut[14], my_FIR_filter_firBlock_right_multProducts[14] );
not U_inv405 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_15_ ( clk, n62_r, rightOut[15], my_FIR_filter_firBlock_right_multProducts[15] );
not U_inv406 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_16_ ( clk, n62_r, rightOut[16], my_FIR_filter_firBlock_right_multProducts[16] );
not U_inv407 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_17_ ( clk, n62_r, rightOut[17], my_FIR_filter_firBlock_right_multProducts[17] );
not U_inv408 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_18_ ( clk, n62_r, rightOut[18], my_FIR_filter_firBlock_right_multProducts[18] );
not U_inv409 ( n62_r, n62 );
dff my_FIR_filter_firBlock_right_Y_reg_19_ ( clk, n61_r, rightOut[19], my_FIR_filter_firBlock_right_multProducts[19] );
not U_inv410 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_20_ ( clk, n61_r, rightOut[20], my_FIR_filter_firBlock_right_multProducts[20] );
not U_inv411 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_21_ ( clk, n61_r, rightOut[21], my_FIR_filter_firBlock_right_multProducts[21] );
not U_inv412 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_22_ ( clk, n61_r, rightOut[22], my_FIR_filter_firBlock_right_multProducts[22] );
not U_inv413 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_23_ ( clk, n61_r, rightOut[23], my_FIR_filter_firBlock_right_multProducts[23] );
not U_inv414 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_24_ ( clk, n61_r, rightOut[24], my_FIR_filter_firBlock_right_multProducts[24] );
not U_inv415 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_25_ ( clk, n61_r, rightOut[25], my_FIR_filter_firBlock_right_multProducts[25] );
not U_inv416 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_26_ ( clk, n61_r, rightOut[26], my_FIR_filter_firBlock_right_multProducts[26] );
not U_inv417 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_27_ ( clk, n61_r, rightOut[27], my_FIR_filter_firBlock_right_multProducts[27] );
not U_inv418 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_28_ ( clk, n61_r, rightOut[28], my_FIR_filter_firBlock_right_multProducts[28] );
not U_inv419 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_29_ ( clk, n61_r, rightOut[29], my_FIR_filter_firBlock_right_multProducts[29] );
not U_inv420 ( n61_r, n61 );
dff my_FIR_filter_firBlock_right_Y_reg_30_ ( clk, n61_r, ex_wire0, my_FIR_filter_firBlock_right_multProducts[30] );
not U_inv421 ( n49, ex_wire0 );
not U_inv422 ( n61_r, n61 );
dff inData_in_reg_1_ ( clk, n95_r, inData_in[1], inData_1 );
not U_inv423 ( n18, inData_in[1] );
not U_inv424 ( n95_r, n95 );
dff my_FIR_filter_firBlock_left_firStep_reg_1__31_ ( clk, n90_r, my_FIR_filter_firBlock_left_firStep[255], my_FIR_filter_firBlock_left_N32 );
not U_inv425 ( n90_r, n90 );
dff my_FIR_filter_firBlock_left_firStep_reg_8__31_ ( clk, n71_r, my_FIR_filter_firBlock_left_firStep[31], my_FIR_filter_firBlock_left_N256 );
not U_inv426 ( n71_r, n71 );
dff inData_in_reg_30_ ( clk, n98_r, my_FIR_filter_firBlock_left_multProducts[114], inData_30 );
not U_inv427 ( n48, my_FIR_filter_firBlock_left_multProducts[114] );
not U_inv428 ( n98_r, n98 );
dff inData_in_reg_29_ ( clk, n98_r, my_FIR_filter_firBlock_left_multProducts[113], inData_29 );
not U_inv429 ( n47, my_FIR_filter_firBlock_left_multProducts[113] );
not U_inv430 ( n98_r, n98 );
dff inData_in_reg_28_ ( clk, n98_r, my_FIR_filter_firBlock_left_multProducts[112], inData_28 );
not U_inv431 ( n46, my_FIR_filter_firBlock_left_multProducts[112] );
not U_inv432 ( n98_r, n98 );
dff inData_in_reg_27_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[111], inData_27 );
not U_inv433 ( n45, my_FIR_filter_firBlock_left_multProducts[111] );
not U_inv434 ( n97_r, n97 );
dff inData_in_reg_26_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[110], inData_26 );
not U_inv435 ( n44, my_FIR_filter_firBlock_left_multProducts[110] );
not U_inv436 ( n97_r, n97 );
dff inData_in_reg_25_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[109], inData_25 );
not U_inv437 ( n43, my_FIR_filter_firBlock_left_multProducts[109] );
not U_inv438 ( n97_r, n97 );
dff inData_in_reg_24_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[108], inData_24 );
not U_inv439 ( n42, my_FIR_filter_firBlock_left_multProducts[108] );
not U_inv440 ( n97_r, n97 );
dff inData_in_reg_23_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[107], inData_23 );
not U_inv441 ( n41, my_FIR_filter_firBlock_left_multProducts[107] );
not U_inv442 ( n97_r, n97 );
dff inData_in_reg_22_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[106], inData_22 );
not U_inv443 ( n40, my_FIR_filter_firBlock_left_multProducts[106] );
not U_inv444 ( n97_r, n97 );
dff inData_in_reg_21_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[105], inData_21 );
not U_inv445 ( n39, my_FIR_filter_firBlock_left_multProducts[105] );
not U_inv446 ( n97_r, n97 );
dff inData_in_reg_20_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[104], inData_20 );
not U_inv447 ( n38, my_FIR_filter_firBlock_left_multProducts[104] );
not U_inv448 ( n97_r, n97 );
dff inData_in_reg_19_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[103], inData_19 );
not U_inv449 ( n37, my_FIR_filter_firBlock_left_multProducts[103] );
not U_inv450 ( n97_r, n97 );
dff inData_in_reg_18_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[102], inData_18 );
not U_inv451 ( n36, my_FIR_filter_firBlock_left_multProducts[102] );
not U_inv452 ( n97_r, n97 );
dff inData_in_reg_17_ ( clk, n97_r, my_FIR_filter_firBlock_left_multProducts[101], inData_17 );
not U_inv453 ( n35, my_FIR_filter_firBlock_left_multProducts[101] );
not U_inv454 ( n97_r, n97 );
dff inData_in_reg_15_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[99], inData_15 );
not U_inv455 ( n33, my_FIR_filter_firBlock_left_multProducts[99] );
not U_inv456 ( n96_r, n96 );
dff inData_in_reg_14_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[98], inData_14 );
not U_inv457 ( n32, my_FIR_filter_firBlock_left_multProducts[98] );
not U_inv458 ( n96_r, n96 );
dff inData_in_reg_13_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[97], inData_13 );
not U_inv459 ( n31, my_FIR_filter_firBlock_left_multProducts[97] );
not U_inv460 ( n96_r, n96 );
dff inData_in_reg_12_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[96], inData_12 );
not U_inv461 ( n30, my_FIR_filter_firBlock_left_multProducts[96] );
not U_inv462 ( n96_r, n96 );
dff inData_in_reg_11_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[95], inData_11 );
not U_inv463 ( n29, my_FIR_filter_firBlock_left_multProducts[95] );
not U_inv464 ( n96_r, n96 );
dff inData_in_reg_10_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[94], inData_10 );
not U_inv465 ( n28, my_FIR_filter_firBlock_left_multProducts[94] );
not U_inv466 ( n96_r, n96 );
dff inData_in_reg_9_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[93], inData_9 );
not U_inv467 ( n27, my_FIR_filter_firBlock_left_multProducts[93] );
not U_inv468 ( n96_r, n96 );
dff inData_in_reg_8_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[92], inData_8 );
not U_inv469 ( n26, my_FIR_filter_firBlock_left_multProducts[92] );
not U_inv470 ( n96_r, n96 );
dff inData_in_reg_7_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[91], inData_7 );
not U_inv471 ( n25, my_FIR_filter_firBlock_left_multProducts[91] );
not U_inv472 ( n96_r, n96 );
dff inData_in_reg_6_ ( clk, n96_r, my_FIR_filter_firBlock_left_multProducts[90], inData_6 );
not U_inv473 ( n24, my_FIR_filter_firBlock_left_multProducts[90] );
not U_inv474 ( n96_r, n96 );
dff inData_in_reg_5_ ( clk, n96_r, inData_in[5], inData_5 );
not U_inv475 ( n23, inData_in[5] );
not U_inv476 ( n96_r, n96 );
dff inData_in_reg_4_ ( clk, n96_r, inData_in[4], inData_4 );
not U_inv477 ( n22, inData_in[4] );
not U_inv478 ( n96_r, n96 );
dff inData_in_reg_3_ ( clk, n95_r, inData_in[3], inData_3 );
not U_inv479 ( n21, inData_in[3] );
not U_inv480 ( n95_r, n95 );
buf U19 ( n108, n113 );
buf U20 ( n107, n113 );
buf U21 ( n106, n113 );
buf U22 ( n105, n114 );
buf U23 ( n104, n114 );
buf U24 ( n103, n114 );
buf U25 ( n102, n115 );
buf U26 ( n101, n115 );
buf U27 ( n100, n115 );
buf U28 ( n110, n112 );
buf U29 ( n109, n112 );
and U30 ( n52, n50, n51 );
nand U31 ( n50, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[38], n1344 );
nand U32 ( n51, n1345, n58 );
buf U33 ( n113, n118 );
buf U34 ( n114, n117 );
buf U35 ( n115, n117 );
buf U36 ( n112, n118 );
buf U37 ( n99, n116 );
buf U38 ( n117, reset );
buf U39 ( n71, n108 );
buf U40 ( n90, n101 );
buf U41 ( n95, n100 );
buf U42 ( n63, n110 );
buf U43 ( n64, n110 );
buf U44 ( n65, n110 );
buf U45 ( n66, n109 );
buf U46 ( n67, n109 );
buf U47 ( n68, n109 );
buf U48 ( n69, n108 );
buf U49 ( n70, n108 );
buf U50 ( n72, n107 );
buf U51 ( n73, n107 );
buf U52 ( n74, n107 );
buf U53 ( n75, n106 );
buf U54 ( n76, n106 );
buf U55 ( n77, n106 );
buf U56 ( n78, n105 );
buf U57 ( n79, n105 );
buf U58 ( n80, n105 );
buf U59 ( n81, n104 );
buf U60 ( n82, n104 );
buf U61 ( n83, n104 );
buf U62 ( n84, n103 );
buf U63 ( n85, n103 );
buf U64 ( n86, n103 );
buf U65 ( n87, n102 );
buf U66 ( n88, n102 );
buf U67 ( n89, n102 );
buf U68 ( n91, n101 );
buf U69 ( n92, n101 );
buf U70 ( n93, n100 );
buf U71 ( n94, n100 );
buf U72 ( n61, n111 );
buf U73 ( n62, n111 );
nand U74 ( n1344, n1343, n1342 );
nand U75 ( n1342, n1341, n57 );
xor U76 ( my_FIR_filter_firBlock_left_multProducts[29], n1340, n1339 );
nand U77 ( n2303, n2302, n125 );
xor U78 ( my_FIR_filter_firBlock_right_multProducts[29], n125, n2302 );
xor U79 ( my_FIR_filter_firBlock_right_multProducts[25], n124, n2297 );
xor U80 ( my_FIR_filter_firBlock_right_multProducts[21], n123, n2291 );
xor U81 ( my_FIR_filter_firBlock_right_multProducts[17], n122, n2285 );
not U82 ( n59, n17 );
buf U83 ( n57, n60 );
xor U84 ( my_FIR_filter_firBlock_right_multProducts[13], n121, n2279 );
buf U85 ( n58, n60 );
nand U86 ( n2264, n2262, n128 );
xor U87 ( my_FIR_filter_firBlock_right_multProducts[9], n126, n2273 );
xor U88 ( my_FIR_filter_firBlock_right_multProducts[5], n127, n2267 );
xor U89 ( my_FIR_filter_firBlock_right_multProducts[2], n128, n2262 );
buf U90 ( n111, n112 );
buf U91 ( n96, n99 );
buf U92 ( n97, n99 );
buf U93 ( n98, n99 );
nand U94 ( n418, n281, n20 );
xor U95 ( n410, n47, n59 );
xor U96 ( n1348, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[9], n27 );
nand U97 ( n1199, n1198, n26 );
xor U98 ( my_FIR_filter_firBlock_left_multProducts[2], n1205, n1204 );
nand U99 ( n1205, n1203, n1202 );
xor U100 ( n1209, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[11], n29 );
nand U101 ( my_FIR_filter_firBlock_left_multProducts[89], n574, n573 );
xor U102 ( n1214, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[12], n30 );
nand U103 ( n1215, n1213, n1212 );
nand U104 ( n1212, n1211, n29 );
xor U105 ( n1219, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[13], n31 );
nand U106 ( n1220, n1218, n1217 );
nand U107 ( n1217, n1216, n30 );
nand U108 ( n1235, n1233, n1232 );
nand U109 ( n1232, n1231, n33 );
nand U110 ( n1240, n1238, n1237 );
nand U111 ( n1237, n1236, n34 );
nand U112 ( n1225, n1223, n1222 );
nand U113 ( n1222, n1221, n31 );
nand U114 ( n1230, n1228, n1227 );
nand U115 ( n1227, n1226, n32 );
xor U116 ( n1229, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[15], n33 );
nand U117 ( n1250, n1248, n1247 );
nand U118 ( n1247, n1246, n36 );
nand U119 ( n1245, n1243, n1242 );
nand U120 ( n1242, n1241, n35 );
xor U121 ( my_FIR_filter_firBlock_left_multProducts[12], n1255, n1254 );
nand U122 ( n1255, n1253, n1252 );
nand U123 ( n1252, n1251, n37 );
nand U124 ( n1302, n1301, n47 );
nand U125 ( n1335, n1333, n1332 );
nand U126 ( n1332, n1331, n58 );
nand U127 ( n1330, n1328, n1327 );
nand U128 ( n1327, n1326, n57 );
nand U129 ( n1340, n1338, n1337 );
nand U130 ( n1337, n1336, n57 );
nand U131 ( n1320, n1318, n1317 );
nand U132 ( n1317, n1316, n58 );
nand U133 ( n1325, n1323, n1322 );
nand U134 ( n1322, n1321, n58 );
nand U135 ( n1315, n1313, n1312 );
nand U136 ( n1312, n1311, n58 );
nand U137 ( n1295, n1293, n1292 );
nand U138 ( n1292, n1291, n45 );
nand U139 ( n1290, n1288, n1287 );
nand U140 ( n1287, n1286, n44 );
nand U141 ( n1280, n1278, n1277 );
nand U142 ( n1277, n1276, n42 );
nand U143 ( n1285, n1283, n1282 );
nand U144 ( n1282, n1281, n43 );
nand U145 ( n1265, n1263, n1262 );
nand U146 ( n1262, n1261, n39 );
nand U147 ( n1260, n1258, n1257 );
nand U148 ( n1257, n1256, n38 );
nand U149 ( n1310, n1308, n1307 );
nand U150 ( n1307, n1306, n48 );
nand U151 ( n1275, n1273, n1272 );
nand U152 ( n1272, n1271, n41 );
nand U153 ( n1270, n1268, n1267 );
nand U154 ( n1267, n1266, n40 );
nand U155 ( n1300, n1298, n1297 );
nand U156 ( n1297, n1296, n46 );
xor U157 ( n1264, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[22], n40 );
xor U158 ( n53, n1344, n54 );
xnor U159 ( n54, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[38], n58 );
xor U160 ( n1269, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[23], n41 );
xor U161 ( n1299, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[29], n47 );
xnor U162 ( my_FIR_filter_firBlock_right_multProducts[31], n55, outData_in[31] );
nor U163 ( n55, n2303, outData_in[30] );
xor U164 ( n1279, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[25], n43 );
xor U165 ( n1284, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[26], n44 );
xor U166 ( n1289, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[27], n45 );
xor U167 ( n1294, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[28], n46 );
xor U168 ( n1274, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[24], n42 );
xor U169 ( n1304, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[30], n48 );
xor U170 ( n1314, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[32], n57 );
xor U171 ( my_FIR_filter_firBlock_left_multProducts[28], n1335, n1334 );
xor U172 ( my_FIR_filter_firBlock_left_multProducts[25], n1320, n1319 );
xor U173 ( n1319, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[33], n57 );
xor U174 ( n1309, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[31], n57 );
xor U175 ( n1324, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[34], n57 );
xor U176 ( my_FIR_filter_firBlock_left_multProducts[27], n1330, n1329 );
xor U177 ( n1329, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[35], n57 );
not U178 ( n119, my_FIR_filter_firBlock_left_multProducts[60] );
xor U179 ( my_FIR_filter_firBlock_right_multProducts[30], n2303, outData_in[30] );
not U180 ( n125, outData_in[29] );
nor U181 ( n2302, n2301, n2300 );
or U182 ( n2301, outData_in[28], outData_in[27] );
nand U183 ( n2300, n2298, n2297 );
nor U184 ( n2298, outData_in[26], outData_in[25] );
xnor U185 ( my_FIR_filter_firBlock_right_multProducts[28], outData_in[28], n2299 );
nor U186 ( n2299, outData_in[27], n2300 );
xor U187 ( my_FIR_filter_firBlock_right_multProducts[27], n2300, outData_in[27] );
nor U188 ( n2297, n2295, n2294 );
or U189 ( n2295, outData_in[24], outData_in[23] );
xor U190 ( my_FIR_filter_firBlock_right_multProducts[26], n2296, outData_in[26] );
nand U191 ( n2296, n2297, n124 );
not U192 ( n124, outData_in[25] );
nand U193 ( n2294, n2292, n2291 );
nor U194 ( n2292, outData_in[22], outData_in[21] );
xnor U195 ( my_FIR_filter_firBlock_right_multProducts[24], outData_in[24], n2293 );
nor U196 ( n2293, outData_in[23], n2294 );
nor U197 ( n2291, n2289, n2288 );
or U198 ( n2289, outData_in[20], outData_in[19] );
xor U199 ( my_FIR_filter_firBlock_right_multProducts[23], n2294, outData_in[23] );
nand U200 ( n2288, n2286, n2285 );
nor U201 ( n2286, outData_in[18], outData_in[17] );
xor U202 ( my_FIR_filter_firBlock_right_multProducts[22], n2290, outData_in[22] );
nand U203 ( n2290, n2291, n123 );
not U204 ( n123, outData_in[21] );
nor U205 ( n2285, n2283, n2282 );
or U206 ( n2283, outData_in[16], outData_in[15] );
xnor U207 ( my_FIR_filter_firBlock_right_multProducts[20], outData_in[20], n2287 );
nor U208 ( n2287, outData_in[19], n2288 );
nand U209 ( n2282, n2280, n2279 );
nor U210 ( n2280, outData_in[14], outData_in[13] );
xor U211 ( my_FIR_filter_firBlock_right_multProducts[19], n2288, outData_in[19] );
xor U212 ( my_FIR_filter_firBlock_right_multProducts[18], n2284, outData_in[18] );
nand U213 ( n2284, n2285, n122 );
nor U214 ( n2279, n2277, n2276 );
or U215 ( n2277, outData_in[12], outData_in[11] );
not U216 ( n122, outData_in[17] );
nand U217 ( n2276, n2274, n2273 );
nor U218 ( n2274, outData_in[10], outData_in[9] );
xnor U219 ( my_FIR_filter_firBlock_right_multProducts[16], outData_in[16], n2281 );
nor U220 ( n2281, outData_in[15], n2282 );
xor U221 ( my_FIR_filter_firBlock_right_multProducts[15], n2282, outData_in[15] );
nor U222 ( n2273, n2271, n2270 );
or U223 ( n2271, outData_in[8], outData_in[7] );
xor U224 ( my_FIR_filter_firBlock_right_multProducts[14], n2278, outData_in[14] );
nand U225 ( n2278, n2279, n121 );
buf U226 ( n60, n17 );
not U227 ( n121, outData_in[13] );
nand U228 ( n2270, n2268, n2267 );
nor U229 ( n2268, outData_in[6], outData_in[5] );
xnor U230 ( my_FIR_filter_firBlock_right_multProducts[12], outData_in[12], n2275 );
nor U231 ( n2275, outData_in[11], n2276 );
nor U232 ( n2267, n2265, n2264 );
or U233 ( n2265, outData_in[4], outData_in[3] );
xor U234 ( my_FIR_filter_firBlock_right_multProducts[11], n2276, outData_in[11] );
xor U235 ( my_FIR_filter_firBlock_right_multProducts[10], n2272, outData_in[10] );
nand U236 ( n2272, n2273, n126 );
not U237 ( n128, outData_in[2] );
nor U238 ( n2262, my_FIR_filter_firBlock_right_multProducts[0], outData_in[1] );
not U239 ( n126, outData_in[9] );
xnor U240 ( my_FIR_filter_firBlock_right_multProducts[8], outData_in[8], n2269 );
nor U241 ( n2269, outData_in[7], n2270 );
xor U242 ( my_FIR_filter_firBlock_right_multProducts[7], n2270, outData_in[7] );
xor U243 ( my_FIR_filter_firBlock_right_multProducts[6], n2266, outData_in[6] );
nand U244 ( n2266, n2267, n127 );
not U245 ( n127, outData_in[5] );
xnor U246 ( my_FIR_filter_firBlock_right_multProducts[4], outData_in[4], n2263 );
nor U247 ( n2263, outData_in[3], n2264 );
xor U248 ( my_FIR_filter_firBlock_right_multProducts[3], n2264, outData_in[3] );
xor U249 ( my_FIR_filter_firBlock_right_multProducts[1], outData_in[1], my_FIR_filter_firBlock_right_multProducts[0] );
buf U250 ( n116, n117 );
nand U251 ( n2013, my_FIR_filter_firBlock_left_multProducts[76], n2012 );
nand U252 ( n2019, my_FIR_filter_firBlock_left_firStep[48], n2016 );
nand U253 ( n2001, n1999, n1998 );
nand U254 ( n1998, my_FIR_filter_firBlock_left_multProducts[73], n1997 );
nand U255 ( n1963, my_FIR_filter_firBlock_left_firStep[34], n2084 );
nand U256 ( n1962, my_FIR_filter_firBlock_left_multProducts[63], n1961 );
or U257 ( n1961, n2084, my_FIR_filter_firBlock_left_firStep[34] );
nand U258 ( n2084, n1960, n1959 );
nand U259 ( n1969, my_FIR_filter_firBlock_left_firStep[36], n2099 );
nand U260 ( n1989, my_FIR_filter_firBlock_left_firStep[42], n1986 );
nand U261 ( n1983, my_FIR_filter_firBlock_left_multProducts[70], n1982 );
nand U262 ( n445, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[13], n576 );
or U263 ( n443, n576, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[13] );
nand U264 ( n576, n442, n441 );
nand U265 ( n442, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[12], n439 );
nand U266 ( n441, inData_in[3], n440 );
or U267 ( n440, n439, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[12] );
nand U268 ( n439, n438, n437 );
nand U269 ( n438, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[11], n435 );
nand U270 ( n437, inData_in[2], n436 );
or U271 ( n436, n435, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[11] );
nand U272 ( n435, n434, n433 );
and U273 ( n432, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[9], n431 );
nand U274 ( n1996, n1994, n1993 );
nand U275 ( n1993, my_FIR_filter_firBlock_left_multProducts[72], n1992 );
nand U276 ( n2103, n1972, n1971 );
nand U277 ( n2104, n1975, n1974 );
nand U278 ( n2048, n2046, n2045 );
nand U279 ( n2045, my_FIR_filter_firBlock_left_multProducts[82], n2044 );
nand U280 ( n2063, n2061, n2060 );
nand U281 ( n2085, n2081, n2080 );
nand U282 ( n2091, n2088, n2087 );
nand U283 ( n708, n704, n703 );
nand U284 ( n701, n699, n698 );
xor U285 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[23], n339, n338 );
xor U286 ( n338, n33, my_FIR_filter_firBlock_left_multProducts[101] );
xor U287 ( my_FIR_filter_firBlock_left_multProducts[71], n488, n487 );
xor U288 ( n487, my_FIR_filter_firBlock_left_multProducts[98], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[23] );
nand U289 ( n631, my_FIR_filter_firBlock_left_multProducts[75], n630 );
nand U290 ( n622, my_FIR_filter_firBlock_left_firStep[268], n619 );
or U291 ( n620, n619, my_FIR_filter_firBlock_left_firStep[268] );
nand U292 ( n637, my_FIR_filter_firBlock_left_firStep[271], n634 );
nand U293 ( n619, n617, n616 );
nand U294 ( n641, my_FIR_filter_firBlock_left_multProducts[77], n640 );
nand U295 ( n649, n647, n646 );
nand U296 ( n646, my_FIR_filter_firBlock_left_multProducts[78], n645 );
nand U297 ( n319, n317, n316 );
nand U298 ( n316, n315, n30 );
nand U299 ( n426, n293, n292 );
nand U300 ( n292, n291, n24 );
nand U301 ( n614, n612, n611 );
nand U302 ( n611, my_FIR_filter_firBlock_left_multProducts[71], n610 );
nand U303 ( n324, n322, n321 );
nand U304 ( n651, my_FIR_filter_firBlock_left_multProducts[79], n650 );
nand U305 ( n659, my_FIR_filter_firBlock_left_firStep[275], n656 );
nand U306 ( n361, n360, n39 );
nand U307 ( n346, n345, n36 );
nand U308 ( n341, n340, n35 );
nand U309 ( n379, n377, n376 );
nand U310 ( n374, n372, n371 );
nand U311 ( n371, n370, n41 );
nand U312 ( n359, n357, n356 );
nand U313 ( n356, n355, n38 );
nand U314 ( n381, n380, n43 );
nand U315 ( n394, n392, n391 );
nand U316 ( n391, n390, n45 );
nand U317 ( n401, n397, n396 );
nand U318 ( n396, n395, n46 );
nand U319 ( n406, n404, n403 );
nand U320 ( n403, n402, n47 );
xor U321 ( n542, my_FIR_filter_firBlock_left_multProducts[109], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[34] );
nand U322 ( n408, n407, n48 );
xor U323 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[38], n416, n415 );
xor U324 ( n415, n48, n59 );
nand U325 ( n416, n414, n413 );
nand U326 ( n414, my_FIR_filter_firBlock_left_multProducts[113], n411 );
nand U327 ( n413, n412, n57 );
or U328 ( n412, n411, my_FIR_filter_firBlock_left_multProducts[113] );
xor U329 ( n393, n44, my_FIR_filter_firBlock_left_multProducts[112] );
xor U330 ( n482, my_FIR_filter_firBlock_left_multProducts[97], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[22] );
xor U331 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[22], n334, n333 );
xor U332 ( n333, n32, my_FIR_filter_firBlock_left_multProducts[100] );
nand U333 ( n607, my_FIR_filter_firBlock_left_firStep[265], n731 );
xor U334 ( n398, n45, my_FIR_filter_firBlock_left_multProducts[113] );
xor U335 ( n547, my_FIR_filter_firBlock_left_multProducts[110], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[35] );
nand U336 ( n468, n466, n465 );
nand U337 ( n465, my_FIR_filter_firBlock_left_multProducts[93], n464 );
nand U338 ( n453, n451, n450 );
xor U339 ( n343, n34, my_FIR_filter_firBlock_left_multProducts[102] );
xor U340 ( n492, my_FIR_filter_firBlock_left_multProducts[99], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[24] );
nand U341 ( n491, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[23], n488 );
nand U342 ( n498, n496, n495 );
nand U343 ( n495, my_FIR_filter_firBlock_left_multProducts[99], n494 );
nand U344 ( n501, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[25], n498 );
xor U345 ( n507, my_FIR_filter_firBlock_left_multProducts[102], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[27] );
nand U346 ( n505, my_FIR_filter_firBlock_left_multProducts[101], n504 );
nand U347 ( n586, my_FIR_filter_firBlock_left_firStep[258], n707 );
or U348 ( n584, n707, my_FIR_filter_firBlock_left_firStep[258] );
nand U349 ( n707, n583, n582 );
nand U350 ( n583, my_FIR_filter_firBlock_left_firStep[257], n655 );
or U351 ( n581, my_FIR_filter_firBlock_left_firStep[257], n655 );
nand U352 ( n595, my_FIR_filter_firBlock_left_firStep[261], n723 );
nand U353 ( n723, n592, n591 );
xor U354 ( my_FIR_filter_firBlock_left_multProducts[67], n468, n467 );
xor U355 ( n358, n37, my_FIR_filter_firBlock_left_multProducts[105] );
xor U356 ( n427, n24, my_FIR_filter_firBlock_left_multProducts[92] );
xor U357 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[30], n374, n373 );
xor U358 ( n373, n40, my_FIR_filter_firBlock_left_multProducts[108] );
xor U359 ( my_FIR_filter_firBlock_left_multProducts[78], n523, n522 );
xor U360 ( n522, my_FIR_filter_firBlock_left_multProducts[105], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[30] );
xor U361 ( n388, n43, my_FIR_filter_firBlock_left_multProducts[111] );
xor U362 ( n537, my_FIR_filter_firBlock_left_multProducts[108], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[33] );
xor U363 ( my_FIR_filter_firBlock_left_multProducts[84], n553, n552 );
nand U364 ( n526, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[30], n523 );
nand U365 ( n523, n521, n520 );
nand U366 ( n520, my_FIR_filter_firBlock_left_multProducts[104], n519 );
nand U367 ( n553, n551, n550 );
nand U368 ( n550, my_FIR_filter_firBlock_left_multProducts[110], n549 );
nand U369 ( n538, n536, n535 );
nand U370 ( n535, my_FIR_filter_firBlock_left_multProducts[107], n534 );
xor U371 ( n512, my_FIR_filter_firBlock_left_multProducts[103], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[28] );
xor U372 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[28], n364, n363 );
xor U373 ( n363, n38, my_FIR_filter_firBlock_left_multProducts[106] );
xor U374 ( n405, n48, my_FIR_filter_firBlock_left_multProducts[112] );
xor U375 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[13], n426, n425 );
xor U376 ( n425, n23, my_FIR_filter_firBlock_left_multProducts[91] );
and U377 ( n655, my_FIR_filter_firBlock_left_multProducts[61], my_FIR_filter_firBlock_left_firStep[256] );
xor U378 ( n502, my_FIR_filter_firBlock_left_multProducts[101], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[26] );
xor U379 ( n532, my_FIR_filter_firBlock_left_multProducts[107], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[32] );
xor U380 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[32], n384, n383 );
xor U381 ( n383, n42, my_FIR_filter_firBlock_left_multProducts[110] );
nand U382 ( n563, n561, n560 );
xor U383 ( n567, my_FIR_filter_firBlock_left_multProducts[114], n59 );
xor U384 ( n353, n36, my_FIR_filter_firBlock_left_multProducts[104] );
xor U385 ( n378, n41, my_FIR_filter_firBlock_left_multProducts[109] );
xor U386 ( n527, my_FIR_filter_firBlock_left_multProducts[106], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[31] );
xor U387 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[19], n319, n318 );
xor U388 ( n318, n31, my_FIR_filter_firBlock_left_multProducts[95] );
xor U389 ( n429, n25, my_FIR_filter_firBlock_left_multProducts[93] );
xor U390 ( n368, n39, my_FIR_filter_firBlock_left_multProducts[107] );
xor U391 ( n517, my_FIR_filter_firBlock_left_multProducts[104], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[29] );
nand U392 ( n1455, n1453, n1452 );
nand U393 ( n1440, n1438, n1437 );
nand U394 ( n1403, n1401, n1400 );
nand U395 ( n1400, my_FIR_filter_firBlock_left_multProducts[14], n1399 );
xnor U396 ( n1487, n52, my_FIR_filter_firBlock_left_firStep[191] );
nor U397 ( n1486, n1485, n1484 );
nand U398 ( n1460, n1458, n1457 );
nand U399 ( n1458, my_FIR_filter_firBlock_left_firStep[185], n1455 );
nand U400 ( n1457, my_FIR_filter_firBlock_left_multProducts[25], n1456 );
or U401 ( n1456, n1455, my_FIR_filter_firBlock_left_firStep[185] );
nand U402 ( n1425, n1421, n1420 );
nand U403 ( n1430, n1428, n1427 );
nand U404 ( n1428, my_FIR_filter_firBlock_left_firStep[179], n1425 );
nand U405 ( n1408, n1406, n1405 );
nand U406 ( n1406, my_FIR_filter_firBlock_left_firStep[175], n1403 );
nand U407 ( n1405, my_FIR_filter_firBlock_left_multProducts[15], n1404 );
or U408 ( n1404, n1403, my_FIR_filter_firBlock_left_firStep[175] );
nand U409 ( n1398, n1396, n1395 );
nand U410 ( n1435, n1433, n1432 );
nand U411 ( n1433, my_FIR_filter_firBlock_left_firStep[180], n1430 );
nand U412 ( n1413, n1411, n1410 );
nand U413 ( n1411, my_FIR_filter_firBlock_left_firStep[176], n1408 );
nand U414 ( n1450, n1448, n1447 );
nand U415 ( n1445, n1443, n1442 );
nand U416 ( n1443, my_FIR_filter_firBlock_left_firStep[182], n1440 );
nand U417 ( n1442, my_FIR_filter_firBlock_left_multProducts[22], n1441 );
or U418 ( n1441, n1440, my_FIR_filter_firBlock_left_firStep[182] );
nand U419 ( n1465, n1463, n1462 );
nand U420 ( n1463, my_FIR_filter_firBlock_left_firStep[186], n1460 );
nand U421 ( n1462, my_FIR_filter_firBlock_left_multProducts[26], n1461 );
or U422 ( n1461, n1460, my_FIR_filter_firBlock_left_firStep[186] );
nand U423 ( n1418, n1416, n1415 );
nand U424 ( n1415, my_FIR_filter_firBlock_left_multProducts[17], n1414 );
nand U425 ( n1470, n1468, n1467 );
nand U426 ( n1467, my_FIR_filter_firBlock_left_multProducts[27], n1466 );
nand U427 ( n1483, n1480, n1479 );
nand U428 ( n1480, my_FIR_filter_firBlock_left_firStep[189], n1477 );
nand U429 ( n1479, my_FIR_filter_firBlock_left_multProducts[29], n1478 );
or U430 ( n1478, n1477, my_FIR_filter_firBlock_left_firStep[189] );
nand U431 ( n1388, n1386, n1385 );
nand U432 ( n1492, n1361, n1360 );
nand U433 ( n1361, my_FIR_filter_firBlock_left_firStep[164], n1491 );
nand U434 ( n1360, my_FIR_filter_firBlock_left_multProducts[4], n1359 );
or U435 ( n1359, n1491, my_FIR_filter_firBlock_left_firStep[164] );
nand U436 ( n1495, n1364, n1363 );
nand U437 ( n1364, my_FIR_filter_firBlock_left_firStep[165], n1492 );
nand U438 ( n1378, n1376, n1375 );
nand U439 ( n1375, my_FIR_filter_firBlock_left_multProducts[9], n1374 );
nand U440 ( n1491, n1358, n1357 );
nand U441 ( n1357, my_FIR_filter_firBlock_left_multProducts[3], n1356 );
nand U442 ( n1476, n1352, n1351 );
nand U443 ( n1352, my_FIR_filter_firBlock_left_firStep[161], n1424 );
or U444 ( n1350, my_FIR_filter_firBlock_left_firStep[161], n1424 );
nand U445 ( n1500, n1373, n1372 );
nand U446 ( n1499, n1370, n1369 );
nand U447 ( n1347, n1197, n1196 );
nand U448 ( n1197, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[7], n1194 );
or U449 ( n1196, my_FIR_filter_firBlock_left_multProducts[91], n1195 );
nor U450 ( n1195, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[7], n1194 );
nand U451 ( n1383, n1381, n1380 );
nand U452 ( n1381, my_FIR_filter_firBlock_left_firStep[170], n1378 );
nand U453 ( n1380, my_FIR_filter_firBlock_left_multProducts[10], n1379 );
or U454 ( n1379, n1378, my_FIR_filter_firBlock_left_firStep[170] );
nand U455 ( n1191, n1187, n1186 );
nor U456 ( n1187, inData_in[3], inData_in[2] );
nand U457 ( n1393, n1391, n1390 );
nand U458 ( n1391, my_FIR_filter_firBlock_left_firStep[172], n1388 );
nand U459 ( n1390, my_FIR_filter_firBlock_left_multProducts[12], n1389 );
or U460 ( n1389, n1388, my_FIR_filter_firBlock_left_firStep[172] );
nand U461 ( n1488, n1355, n1354 );
nand U462 ( n1355, my_FIR_filter_firBlock_left_firStep[162], n1476 );
or U463 ( n1353, n1476, my_FIR_filter_firBlock_left_firStep[162] );
or U464 ( n1194, n1193, n1192 );
nor U465 ( n1193, n1191, n1190 );
nand U466 ( n1496, n1367, n1366 );
nand U467 ( n1367, my_FIR_filter_firBlock_left_firStep[166], n1495 );
nand U468 ( n1366, my_FIR_filter_firBlock_left_multProducts[6], n1365 );
or U469 ( n1365, n1495, my_FIR_filter_firBlock_left_firStep[166] );
xor U470 ( n323, n30, my_FIR_filter_firBlock_left_multProducts[98] );
xnor U471 ( my_FIR_filter_firBlock_left_multProducts[0], n1347, n1346 );
xor U472 ( n1346, my_FIR_filter_firBlock_left_multProducts[92], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[8] );
and U473 ( n1424, my_FIR_filter_firBlock_left_multProducts[0], my_FIR_filter_firBlock_left_firStep[160] );
xor U474 ( n348, n35, my_FIR_filter_firBlock_left_multProducts[103] );
xor U475 ( n328, n31, my_FIR_filter_firBlock_left_multProducts[99] );
nand U476 ( n746, inData_in[5], n745 );
nand U477 ( n876, n738, n737 );
nand U478 ( n737, inData_in[2], n736 );
nand U479 ( n779, n777, n776 );
nand U480 ( n777, my_FIR_filter_firBlock_left_multProducts[95], n774 );
nand U481 ( n776, my_FIR_filter_firBlock_left_multProducts[99], n775 );
nand U482 ( n879, n741, n740 );
nand U483 ( n741, my_FIR_filter_firBlock_left_multProducts[91], n876 );
nand U484 ( n740, inData_in[3], n739 );
or U485 ( n739, n876, my_FIR_filter_firBlock_left_multProducts[91] );
nand U486 ( n774, n772, n771 );
nand U487 ( n772, my_FIR_filter_firBlock_left_multProducts[94], n769 );
nand U488 ( n771, my_FIR_filter_firBlock_left_multProducts[98], n770 );
nand U489 ( n759, n757, n756 );
nand U490 ( n756, my_FIR_filter_firBlock_left_multProducts[95], n755 );
nand U491 ( n769, n767, n766 );
nand U492 ( n766, my_FIR_filter_firBlock_left_multProducts[97], n765 );
nand U493 ( n754, n752, n751 );
nand U494 ( n751, my_FIR_filter_firBlock_left_multProducts[94], n750 );
nand U495 ( n764, n762, n761 );
nand U496 ( n762, my_FIR_filter_firBlock_left_multProducts[92], n759 );
nand U497 ( n761, my_FIR_filter_firBlock_left_multProducts[96], n760 );
nand U498 ( n880, n744, n743 );
nand U499 ( n744, my_FIR_filter_firBlock_left_multProducts[92], n879 );
or U500 ( n742, n879, my_FIR_filter_firBlock_left_multProducts[92] );
nand U501 ( n875, n735, n734 );
nand U502 ( n734, inData_in[5], n733 );
nand U503 ( n789, n787, n786 );
nand U504 ( n786, my_FIR_filter_firBlock_left_multProducts[101], n785 );
nand U505 ( n782, my_FIR_filter_firBlock_left_multProducts[96], n779 );
nand U506 ( n781, my_FIR_filter_firBlock_left_multProducts[100], n780 );
or U507 ( n780, n779, my_FIR_filter_firBlock_left_multProducts[96] );
nand U508 ( n794, n792, n791 );
nand U509 ( n792, my_FIR_filter_firBlock_left_multProducts[98], n789 );
nand U510 ( n791, my_FIR_filter_firBlock_left_multProducts[102], n790 );
or U511 ( n790, n789, my_FIR_filter_firBlock_left_multProducts[98] );
nand U512 ( n801, my_FIR_filter_firBlock_left_multProducts[104], n800 );
nand U513 ( n829, n827, n826 );
nand U514 ( n827, my_FIR_filter_firBlock_left_multProducts[105], n824 );
nand U515 ( n826, my_FIR_filter_firBlock_left_multProducts[109], n825 );
nand U516 ( n859, n857, n856 );
nand U517 ( n857, my_FIR_filter_firBlock_left_multProducts[111], n854 );
nand U518 ( n856, n59, n855 );
nand U519 ( n819, n817, n816 );
nand U520 ( n816, my_FIR_filter_firBlock_left_multProducts[107], n815 );
nand U521 ( n824, n822, n821 );
nand U522 ( n822, my_FIR_filter_firBlock_left_multProducts[104], n819 );
nand U523 ( n821, my_FIR_filter_firBlock_left_multProducts[108], n820 );
or U524 ( n820, n819, my_FIR_filter_firBlock_left_multProducts[104] );
nand U525 ( n854, n852, n851 );
nand U526 ( n851, my_FIR_filter_firBlock_left_multProducts[114], n850 );
nand U527 ( n809, n807, n806 );
nand U528 ( n806, my_FIR_filter_firBlock_left_multProducts[105], n805 );
nand U529 ( n844, n842, n841 );
nand U530 ( n842, my_FIR_filter_firBlock_left_multProducts[108], n839 );
nand U531 ( n841, my_FIR_filter_firBlock_left_multProducts[112], n840 );
nand U532 ( n814, n812, n811 );
nand U533 ( n812, my_FIR_filter_firBlock_left_multProducts[102], n809 );
nand U534 ( n811, my_FIR_filter_firBlock_left_multProducts[106], n810 );
nand U535 ( n834, n832, n831 );
nand U536 ( n832, my_FIR_filter_firBlock_left_multProducts[106], n829 );
nand U537 ( n831, my_FIR_filter_firBlock_left_multProducts[110], n830 );
or U538 ( n830, n829, my_FIR_filter_firBlock_left_multProducts[106] );
nand U539 ( n849, n847, n846 );
nand U540 ( n846, my_FIR_filter_firBlock_left_multProducts[113], n845 );
nand U541 ( n799, n797, n796 );
nand U542 ( n796, my_FIR_filter_firBlock_left_multProducts[103], n795 );
nand U543 ( n863, n862, n861 );
nand U544 ( n862, my_FIR_filter_firBlock_left_multProducts[112], n859 );
nand U545 ( n861, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n860 );
or U546 ( n860, n859, my_FIR_filter_firBlock_left_multProducts[112] );
xor U547 ( my_FIR_filter_firBlock_left_multProducts[59], n868, n867 );
xor U548 ( n867, n59, my_FIR_filter_firBlock_left_multProducts[114] );
nand U549 ( n1933, n1929, n1928 );
nand U550 ( n1929, my_FIR_filter_firBlock_left_firStep[92], n1926 );
nand U551 ( n1928, my_FIR_filter_firBlock_left_multProducts[59], n1927 );
or U552 ( n1927, n1926, my_FIR_filter_firBlock_left_firStep[92] );
nand U553 ( n868, n866, n865 );
nand U554 ( n866, my_FIR_filter_firBlock_left_multProducts[113], n863 );
nand U555 ( n865, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n864 );
or U556 ( n864, n863, my_FIR_filter_firBlock_left_multProducts[113] );
nand U557 ( n1936, my_FIR_filter_firBlock_left_firStep[93], n1933 );
nand U558 ( n1935, my_FIR_filter_firBlock_left_multProducts[60], n1934 );
or U559 ( n1934, n1933, my_FIR_filter_firBlock_left_firStep[93] );
xor U560 ( my_FIR_filter_firBlock_left_N224, n1943, n1942 );
xnor U561 ( n1943, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, my_FIR_filter_firBlock_left_firStep[95] );
nor U562 ( n1942, n1941, n1940 );
nor U563 ( n1941, n1938, n57 );
nand U564 ( n1009, n1005, n1004 );
nand U565 ( n1005, my_FIR_filter_firBlock_left_firStep[252], n1002 );
nand U566 ( n1012, my_FIR_filter_firBlock_left_firStep[253], n1009 );
or U567 ( n1010, n1009, my_FIR_filter_firBlock_left_firStep[253] );
xor U568 ( my_FIR_filter_firBlock_left_N64, n1019, n1018 );
xnor U569 ( n1019, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, my_FIR_filter_firBlock_left_firStep[255] );
nor U570 ( n1018, n1017, n1016 );
and U571 ( n1016, n1015, my_FIR_filter_firBlock_left_firStep[254] );
nor U572 ( n1017, n1014, n57 );
xor U573 ( n421, n21, inData_in[5] );
xor U574 ( my_FIR_filter_firBlock_left_multProducts[57], n859, n858 );
xor U575 ( n858, n59, my_FIR_filter_firBlock_left_multProducts[112] );
nand U576 ( n1924, my_FIR_filter_firBlock_left_firStep[91], n1921 );
or U577 ( n1922, n1921, my_FIR_filter_firBlock_left_firStep[91] );
nand U578 ( n1921, n1919, n1918 );
nand U579 ( n1919, my_FIR_filter_firBlock_left_firStep[90], n1916 );
xnor U580 ( my_FIR_filter_firBlock_left_multProducts[52], n833, n834 );
xnor U581 ( n833, my_FIR_filter_firBlock_left_multProducts[107], my_FIR_filter_firBlock_left_multProducts[111] );
nand U582 ( n1901, n1899, n1898 );
nand U583 ( n1899, my_FIR_filter_firBlock_left_firStep[86], n1896 );
nand U584 ( n1911, n1909, n1908 );
nand U585 ( n1909, my_FIR_filter_firBlock_left_firStep[88], n1906 );
nand U586 ( n1896, n1894, n1893 );
nand U587 ( n1894, my_FIR_filter_firBlock_left_firStep[85], n1891 );
nand U588 ( n1906, n1904, n1903 );
nand U589 ( n1904, my_FIR_filter_firBlock_left_firStep[87], n1901 );
nand U590 ( n1903, my_FIR_filter_firBlock_left_multProducts[54], n1902 );
or U591 ( n1902, n1901, my_FIR_filter_firBlock_left_firStep[87] );
nand U592 ( n1916, n1914, n1913 );
nand U593 ( n1914, my_FIR_filter_firBlock_left_firStep[89], n1911 );
nand U594 ( n1913, my_FIR_filter_firBlock_left_multProducts[56], n1912 );
or U595 ( n1912, n1911, my_FIR_filter_firBlock_left_firStep[89] );
xor U596 ( my_FIR_filter_firBlock_left_multProducts[53], n839, n838 );
xor U597 ( n838, my_FIR_filter_firBlock_left_multProducts[112], my_FIR_filter_firBlock_left_multProducts[108] );
xor U598 ( n308, n27, my_FIR_filter_firBlock_left_multProducts[95] );
xor U599 ( n313, n30, my_FIR_filter_firBlock_left_multProducts[94] );
xnor U600 ( my_FIR_filter_firBlock_left_multProducts[54], n843, n844 );
xnor U601 ( n843, my_FIR_filter_firBlock_left_multProducts[109], my_FIR_filter_firBlock_left_multProducts[113] );
xor U602 ( my_FIR_filter_firBlock_left_multProducts[55], n849, n848 );
xor U603 ( n848, my_FIR_filter_firBlock_left_multProducts[114], my_FIR_filter_firBlock_left_multProducts[110] );
xor U604 ( n303, n26, my_FIR_filter_firBlock_left_multProducts[94] );
xnor U605 ( my_FIR_filter_firBlock_left_multProducts[56], n853, n854 );
xnor U606 ( n853, my_FIR_filter_firBlock_left_multProducts[111], n59 );
xor U607 ( my_FIR_filter_firBlock_left_multProducts[51], n829, n828 );
xor U608 ( n828, my_FIR_filter_firBlock_left_multProducts[110], my_FIR_filter_firBlock_left_multProducts[106] );
nand U609 ( n1891, n1889, n1888 );
nand U610 ( n1889, my_FIR_filter_firBlock_left_firStep[84], n1886 );
nand U611 ( my_FIR_filter_firBlock_left_multProducts[88], n571, n570 );
xor U612 ( my_FIR_filter_firBlock_left_multProducts[45], n799, n798 );
xor U613 ( n798, my_FIR_filter_firBlock_left_multProducts[104], my_FIR_filter_firBlock_left_multProducts[100] );
nand U614 ( n1881, n1877, n1876 );
nand U615 ( n1877, my_FIR_filter_firBlock_left_firStep[82], n1874 );
nand U616 ( n1869, n1867, n1866 );
nand U617 ( n1867, my_FIR_filter_firBlock_left_firStep[80], n1864 );
nand U618 ( n1859, n1857, n1856 );
nand U619 ( n1857, my_FIR_filter_firBlock_left_firStep[78], n1854 );
nand U620 ( n1886, n1884, n1883 );
nand U621 ( n1884, my_FIR_filter_firBlock_left_firStep[83], n1881 );
nand U622 ( n1883, my_FIR_filter_firBlock_left_multProducts[50], n1882 );
or U623 ( n1882, n1881, my_FIR_filter_firBlock_left_firStep[83] );
nand U624 ( n1874, n1872, n1871 );
nand U625 ( n1872, my_FIR_filter_firBlock_left_firStep[81], n1869 );
nand U626 ( n1871, my_FIR_filter_firBlock_left_multProducts[48], n1870 );
or U627 ( n1870, n1869, my_FIR_filter_firBlock_left_firStep[81] );
nand U628 ( n1864, n1862, n1861 );
nand U629 ( n1862, my_FIR_filter_firBlock_left_firStep[79], n1859 );
nand U630 ( n1861, my_FIR_filter_firBlock_left_multProducts[46], n1860 );
or U631 ( n1860, n1859, my_FIR_filter_firBlock_left_firStep[79] );
nand U632 ( n997, n995, n994 );
nand U633 ( n995, my_FIR_filter_firBlock_left_firStep[250], n992 );
nand U634 ( n1002, n1000, n999 );
nand U635 ( n1000, my_FIR_filter_firBlock_left_firStep[251], n997 );
or U636 ( n998, n997, my_FIR_filter_firBlock_left_firStep[251] );
xor U637 ( my_FIR_filter_firBlock_left_multProducts[49], n819, n818 );
xor U638 ( n818, my_FIR_filter_firBlock_left_multProducts[108], my_FIR_filter_firBlock_left_multProducts[104] );
xnor U639 ( my_FIR_filter_firBlock_left_multProducts[44], n793, n794 );
xnor U640 ( n793, my_FIR_filter_firBlock_left_multProducts[99], my_FIR_filter_firBlock_left_multProducts[103] );
nand U641 ( n1854, n1852, n1851 );
nand U642 ( n1852, my_FIR_filter_firBlock_left_firStep[77], n1849 );
nand U643 ( n1851, my_FIR_filter_firBlock_left_multProducts[44], n1850 );
or U644 ( n1850, n1849, my_FIR_filter_firBlock_left_firStep[77] );
xor U645 ( my_FIR_filter_firBlock_left_multProducts[43], n789, n788 );
xor U646 ( n788, my_FIR_filter_firBlock_left_multProducts[102], my_FIR_filter_firBlock_left_multProducts[98] );
nand U647 ( n1849, n1847, n1846 );
nand U648 ( n1847, my_FIR_filter_firBlock_left_firStep[76], n1844 );
xor U649 ( my_FIR_filter_firBlock_left_multProducts[47], n809, n808 );
xor U650 ( n808, my_FIR_filter_firBlock_left_multProducts[106], my_FIR_filter_firBlock_left_multProducts[102] );
xnor U651 ( my_FIR_filter_firBlock_left_multProducts[50], n823, n824 );
xnor U652 ( n823, my_FIR_filter_firBlock_left_multProducts[105], my_FIR_filter_firBlock_left_multProducts[109] );
xor U653 ( my_FIR_filter_firBlock_left_multProducts[58], n56, n863 );
xor U654 ( n56, my_FIR_filter_firBlock_left_multProducts[113], n59 );
xnor U655 ( my_FIR_filter_firBlock_left_multProducts[48], n813, n814 );
xnor U656 ( n813, my_FIR_filter_firBlock_left_multProducts[103], my_FIR_filter_firBlock_left_multProducts[107] );
xnor U657 ( my_FIR_filter_firBlock_left_multProducts[46], n803, n804 );
xnor U658 ( n803, my_FIR_filter_firBlock_left_multProducts[101], my_FIR_filter_firBlock_left_multProducts[105] );
xnor U659 ( my_FIR_filter_firBlock_left_multProducts[32], n877, n876 );
xnor U660 ( n877, inData_in[3], my_FIR_filter_firBlock_left_multProducts[91] );
nand U661 ( n1956, n1829, n1828 );
nand U662 ( n1829, my_FIR_filter_firBlock_left_firStep[72], n1955 );
nand U663 ( n1948, n1817, n1816 );
nand U664 ( n1817, my_FIR_filter_firBlock_left_firStep[68], n1947 );
nand U665 ( n1952, n1823, n1822 );
nand U666 ( n1823, my_FIR_filter_firBlock_left_firStep[70], n1951 );
nand U667 ( n1944, n1811, n1810 );
nand U668 ( n1811, my_FIR_filter_firBlock_left_firStep[66], n1932 );
nand U669 ( n1810, my_FIR_filter_firBlock_left_multProducts[33], n1809 );
or U670 ( n1809, n1932, my_FIR_filter_firBlock_left_firStep[66] );
nand U671 ( n1932, n1808, n1807 );
nand U672 ( n1808, my_FIR_filter_firBlock_left_firStep[65], n1880 );
nand U673 ( n1807, my_FIR_filter_firBlock_left_multProducts[32], n1806 );
or U674 ( n1806, my_FIR_filter_firBlock_left_firStep[65], n1880 );
nand U675 ( n1839, n1837, n1836 );
nand U676 ( n1837, my_FIR_filter_firBlock_left_firStep[74], n1834 );
nand U677 ( n1844, n1842, n1841 );
nand U678 ( n1842, my_FIR_filter_firBlock_left_firStep[75], n1839 );
nand U679 ( n1947, n1814, n1813 );
nand U680 ( n1814, my_FIR_filter_firBlock_left_firStep[67], n1944 );
nand U681 ( n1813, my_FIR_filter_firBlock_left_multProducts[34], n1812 );
or U682 ( n1812, n1944, my_FIR_filter_firBlock_left_firStep[67] );
nand U683 ( n1834, n1832, n1831 );
nand U684 ( n1832, my_FIR_filter_firBlock_left_firStep[73], n1956 );
nand U685 ( n1831, my_FIR_filter_firBlock_left_multProducts[40], n1830 );
or U686 ( n1830, n1956, my_FIR_filter_firBlock_left_firStep[73] );
nand U687 ( n1951, n1820, n1819 );
nand U688 ( n1820, my_FIR_filter_firBlock_left_firStep[69], n1948 );
nand U689 ( n1819, my_FIR_filter_firBlock_left_multProducts[36], n1818 );
or U690 ( n1818, n1948, my_FIR_filter_firBlock_left_firStep[69] );
nand U691 ( n1955, n1826, n1825 );
nand U692 ( n1826, my_FIR_filter_firBlock_left_firStep[71], n1952 );
nand U693 ( n1825, my_FIR_filter_firBlock_left_multProducts[38], n1824 );
or U694 ( n1824, n1952, my_FIR_filter_firBlock_left_firStep[71] );
nand U695 ( n977, n975, n974 );
nand U696 ( n975, my_FIR_filter_firBlock_left_firStep[246], n972 );
nand U697 ( n987, n985, n984 );
nand U698 ( n985, my_FIR_filter_firBlock_left_firStep[248], n982 );
nand U699 ( n992, n990, n989 );
nand U700 ( n990, my_FIR_filter_firBlock_left_firStep[249], n987 );
nand U701 ( n982, n980, n979 );
nand U702 ( n980, my_FIR_filter_firBlock_left_firStep[247], n977 );
nand U703 ( n979, my_FIR_filter_firBlock_left_multProducts[54], n978 );
or U704 ( n978, n977, my_FIR_filter_firBlock_left_firStep[247] );
nand U705 ( n972, n970, n969 );
nand U706 ( n970, my_FIR_filter_firBlock_left_firStep[245], n967 );
nand U707 ( n969, my_FIR_filter_firBlock_left_multProducts[52], n968 );
or U708 ( n968, n967, my_FIR_filter_firBlock_left_firStep[245] );
xor U709 ( my_FIR_filter_firBlock_left_multProducts[33], n879, n878 );
nand U710 ( n967, n965, n964 );
nand U711 ( n965, my_FIR_filter_firBlock_left_firStep[244], n962 );
nand U712 ( n957, n953, n952 );
nand U713 ( n953, my_FIR_filter_firBlock_left_firStep[242], n950 );
nand U714 ( n962, n960, n959 );
nand U715 ( n960, my_FIR_filter_firBlock_left_firStep[243], n957 );
nand U716 ( n959, my_FIR_filter_firBlock_left_multProducts[50], n958 );
or U717 ( n958, n957, my_FIR_filter_firBlock_left_firStep[243] );
xnor U718 ( my_FIR_filter_firBlock_left_multProducts[42], n783, n784 );
xnor U719 ( n783, my_FIR_filter_firBlock_left_multProducts[97], my_FIR_filter_firBlock_left_multProducts[101] );
nand U720 ( n945, n943, n942 );
nand U721 ( n943, my_FIR_filter_firBlock_left_firStep[240], n940 );
nand U722 ( n950, n948, n947 );
nand U723 ( n948, my_FIR_filter_firBlock_left_firStep[241], n945 );
nand U724 ( n947, my_FIR_filter_firBlock_left_multProducts[48], n946 );
or U725 ( n946, n945, my_FIR_filter_firBlock_left_firStep[241] );
nand U726 ( n1032, n905, n904 );
nand U727 ( n905, my_FIR_filter_firBlock_left_firStep[232], n1031 );
nand U728 ( n925, n923, n922 );
nand U729 ( n923, my_FIR_filter_firBlock_left_firStep[236], n920 );
nand U730 ( n1028, n899, n898 );
nand U731 ( n899, my_FIR_filter_firBlock_left_firStep[230], n1027 );
nand U732 ( n915, n913, n912 );
nand U733 ( n913, my_FIR_filter_firBlock_left_firStep[234], n910 );
nand U734 ( n1020, n887, n886 );
nand U735 ( n887, my_FIR_filter_firBlock_left_firStep[226], n1008 );
nand U736 ( n886, my_FIR_filter_firBlock_left_multProducts[33], n885 );
or U737 ( n885, n1008, my_FIR_filter_firBlock_left_firStep[226] );
nand U738 ( n1008, n884, n883 );
nand U739 ( n884, my_FIR_filter_firBlock_left_firStep[225], n956 );
nand U740 ( n883, my_FIR_filter_firBlock_left_multProducts[32], n882 );
or U741 ( n882, my_FIR_filter_firBlock_left_firStep[225], n956 );
nand U742 ( n1023, n890, n889 );
nand U743 ( n890, my_FIR_filter_firBlock_left_firStep[227], n1020 );
nand U744 ( n889, my_FIR_filter_firBlock_left_multProducts[34], n888 );
or U745 ( n888, n1020, my_FIR_filter_firBlock_left_firStep[227] );
nand U746 ( n935, n933, n932 );
nand U747 ( n933, my_FIR_filter_firBlock_left_firStep[238], n930 );
nand U748 ( n940, n938, n937 );
nand U749 ( n938, my_FIR_filter_firBlock_left_firStep[239], n935 );
nand U750 ( n1027, n896, n895 );
nand U751 ( n896, my_FIR_filter_firBlock_left_firStep[229], n1024 );
nand U752 ( n1024, n893, n892 );
nand U753 ( n893, my_FIR_filter_firBlock_left_firStep[228], n1023 );
nand U754 ( n892, my_FIR_filter_firBlock_left_multProducts[35], n891 );
or U755 ( n891, n1023, my_FIR_filter_firBlock_left_firStep[228] );
nand U756 ( n930, n928, n927 );
nand U757 ( n928, my_FIR_filter_firBlock_left_firStep[237], n925 );
nand U758 ( n927, my_FIR_filter_firBlock_left_multProducts[44], n926 );
or U759 ( n926, n925, my_FIR_filter_firBlock_left_firStep[237] );
nand U760 ( n910, n908, n907 );
nand U761 ( n908, my_FIR_filter_firBlock_left_firStep[233], n1032 );
nand U762 ( n907, my_FIR_filter_firBlock_left_multProducts[40], n906 );
or U763 ( n906, n1032, my_FIR_filter_firBlock_left_firStep[233] );
nand U764 ( n920, n918, n917 );
nand U765 ( n918, my_FIR_filter_firBlock_left_firStep[235], n915 );
nand U766 ( n917, my_FIR_filter_firBlock_left_multProducts[42], n916 );
or U767 ( n916, n915, my_FIR_filter_firBlock_left_firStep[235] );
nand U768 ( n1031, n902, n901 );
nand U769 ( n902, my_FIR_filter_firBlock_left_firStep[231], n1028 );
nand U770 ( n901, my_FIR_filter_firBlock_left_multProducts[38], n900 );
or U771 ( n900, n1028, my_FIR_filter_firBlock_left_firStep[231] );
xor U772 ( my_FIR_filter_firBlock_left_multProducts[41], n779, n778 );
xor U773 ( n778, my_FIR_filter_firBlock_left_multProducts[100], my_FIR_filter_firBlock_left_multProducts[96] );
xor U774 ( my_FIR_filter_firBlock_left_multProducts[31], n875, n874 );
and U775 ( n1880, my_FIR_filter_firBlock_left_multProducts[31], my_FIR_filter_firBlock_left_firStep[64] );
xnor U776 ( my_FIR_filter_firBlock_left_multProducts[34], n881, n880 );
xnor U777 ( n881, inData_in[5], my_FIR_filter_firBlock_left_multProducts[93] );
xor U778 ( my_FIR_filter_firBlock_left_multProducts[39], n769, n768 );
xor U779 ( n768, my_FIR_filter_firBlock_left_multProducts[98], my_FIR_filter_firBlock_left_multProducts[94] );
xnor U780 ( my_FIR_filter_firBlock_left_multProducts[40], n773, n774 );
xnor U781 ( n773, my_FIR_filter_firBlock_left_multProducts[95], my_FIR_filter_firBlock_left_multProducts[99] );
xor U782 ( my_FIR_filter_firBlock_left_multProducts[37], n759, n758 );
xor U783 ( n758, my_FIR_filter_firBlock_left_multProducts[96], my_FIR_filter_firBlock_left_multProducts[92] );
xor U784 ( my_FIR_filter_firBlock_left_multProducts[35], n749, n748 );
xnor U785 ( my_FIR_filter_firBlock_left_multProducts[38], n763, n764 );
xnor U786 ( n763, my_FIR_filter_firBlock_left_multProducts[97], my_FIR_filter_firBlock_left_multProducts[93] );
xnor U787 ( my_FIR_filter_firBlock_left_multProducts[36], n753, n754 );
xnor U788 ( n753, my_FIR_filter_firBlock_left_multProducts[95], my_FIR_filter_firBlock_left_multProducts[91] );
and U789 ( n956, my_FIR_filter_firBlock_left_multProducts[31], my_FIR_filter_firBlock_left_firStep[224] );
xnor U790 ( n1639, n52, my_FIR_filter_firBlock_left_firStep[159] );
xnor U791 ( n2089, n120, my_FIR_filter_firBlock_left_firStep[62] );
xnor U792 ( n712, n120, my_FIR_filter_firBlock_left_firStep[286] );
xor U793 ( outData_in[31], n266, n265 );
xnor U794 ( n266, rightOut[31], leftOut[31] );
nor U795 ( n265, n264, n263 );
and U796 ( n263, n262, leftOut[30] );
nand U797 ( n262, n259, n258 );
nand U798 ( n259, leftOut[29], n256 );
nand U799 ( n258, rightOut[29], n257 );
or U800 ( n257, n256, leftOut[29] );
nand U801 ( n267, n134, n133 );
nand U802 ( n134, leftOut[2], n255 );
nand U803 ( n133, rightOut[2], n132 );
or U804 ( n132, n255, leftOut[2] );
nand U805 ( n275, n146, n145 );
nand U806 ( n146, leftOut[6], n274 );
nand U807 ( n145, rightOut[6], n144 );
or U808 ( n144, n274, leftOut[6] );
nand U809 ( n279, n152, n151 );
nand U810 ( n152, leftOut[8], n278 );
nand U811 ( n151, rightOut[8], n150 );
or U812 ( n150, n278, leftOut[8] );
nand U813 ( n162, n160, n159 );
nand U814 ( n160, leftOut[10], n157 );
nand U815 ( n159, rightOut[10], n158 );
or U816 ( n158, n157, leftOut[10] );
nand U817 ( n172, n170, n169 );
nand U818 ( n170, leftOut[12], n167 );
nand U819 ( n169, rightOut[12], n168 );
or U820 ( n168, n167, leftOut[12] );
nand U821 ( n182, n180, n179 );
nand U822 ( n180, leftOut[14], n177 );
nand U823 ( n179, rightOut[14], n178 );
or U824 ( n178, n177, leftOut[14] );
nand U825 ( n192, n190, n189 );
nand U826 ( n190, leftOut[16], n187 );
nand U827 ( n189, rightOut[16], n188 );
or U828 ( n188, n187, leftOut[16] );
nand U829 ( n204, n200, n199 );
nand U830 ( n200, leftOut[18], n197 );
nand U831 ( n199, rightOut[18], n198 );
or U832 ( n198, n197, leftOut[18] );
nand U833 ( n214, n212, n211 );
nand U834 ( n212, leftOut[20], n209 );
nand U835 ( n211, rightOut[20], n210 );
or U836 ( n210, n209, leftOut[20] );
nand U837 ( n224, n222, n221 );
nand U838 ( n222, leftOut[22], n219 );
nand U839 ( n221, rightOut[22], n220 );
or U840 ( n220, n219, leftOut[22] );
nand U841 ( n234, n232, n231 );
nand U842 ( n232, leftOut[24], n229 );
nand U843 ( n231, rightOut[24], n230 );
or U844 ( n230, n229, leftOut[24] );
nand U845 ( n244, n242, n241 );
nand U846 ( n242, leftOut[26], n239 );
nand U847 ( n241, rightOut[26], n240 );
or U848 ( n240, n239, leftOut[26] );
nand U849 ( n256, n252, n251 );
nand U850 ( n252, leftOut[28], n249 );
nand U851 ( n251, rightOut[28], n250 );
or U852 ( n250, n249, leftOut[28] );
nand U853 ( n255, n131, n130 );
nand U854 ( n131, leftOut[1], n203 );
nand U855 ( n130, rightOut[1], n129 );
or U856 ( n129, leftOut[1], n203 );
nand U857 ( n270, n137, n136 );
nand U858 ( n137, leftOut[3], n267 );
nand U859 ( n136, rightOut[3], n135 );
or U860 ( n135, n267, leftOut[3] );
nand U861 ( n274, n143, n142 );
nand U862 ( n143, leftOut[5], n271 );
nand U863 ( n142, rightOut[5], n141 );
or U864 ( n141, n271, leftOut[5] );
nand U865 ( n278, n149, n148 );
nand U866 ( n149, leftOut[7], n275 );
nand U867 ( n148, rightOut[7], n147 );
or U868 ( n147, n275, leftOut[7] );
nand U869 ( n157, n155, n154 );
nand U870 ( n155, leftOut[9], n279 );
nand U871 ( n154, rightOut[9], n153 );
or U872 ( n153, n279, leftOut[9] );
nand U873 ( n167, n165, n164 );
nand U874 ( n165, leftOut[11], n162 );
nand U875 ( n164, rightOut[11], n163 );
or U876 ( n163, n162, leftOut[11] );
nand U877 ( n177, n175, n174 );
nand U878 ( n175, leftOut[13], n172 );
nand U879 ( n174, rightOut[13], n173 );
or U880 ( n173, n172, leftOut[13] );
nand U881 ( n187, n185, n184 );
nand U882 ( n185, leftOut[15], n182 );
nand U883 ( n184, rightOut[15], n183 );
or U884 ( n183, n182, leftOut[15] );
nand U885 ( n197, n195, n194 );
nand U886 ( n195, leftOut[17], n192 );
nand U887 ( n194, rightOut[17], n193 );
or U888 ( n193, n192, leftOut[17] );
nand U889 ( n209, n207, n206 );
nand U890 ( n207, leftOut[19], n204 );
nand U891 ( n206, rightOut[19], n205 );
or U892 ( n205, n204, leftOut[19] );
nand U893 ( n219, n217, n216 );
nand U894 ( n217, leftOut[21], n214 );
nand U895 ( n216, rightOut[21], n215 );
or U896 ( n215, n214, leftOut[21] );
nand U897 ( n229, n227, n226 );
nand U898 ( n227, leftOut[23], n224 );
nand U899 ( n226, rightOut[23], n225 );
or U900 ( n225, n224, leftOut[23] );
nand U901 ( n239, n237, n236 );
nand U902 ( n237, leftOut[25], n234 );
nand U903 ( n236, rightOut[25], n235 );
or U904 ( n235, n234, leftOut[25] );
nand U905 ( n249, n247, n246 );
nand U906 ( n247, leftOut[27], n244 );
nand U907 ( n246, rightOut[27], n245 );
or U908 ( n245, n244, leftOut[27] );
nor U909 ( n264, n261, n49 );
nor U910 ( n261, leftOut[30], n262 );
and U911 ( n203, rightOut[0], leftOut[0] );
nand U912 ( n271, n140, n139 );
nand U913 ( n140, leftOut[4], n270 );
nand U914 ( n139, rightOut[4], n138 );
or U915 ( n138, n270, leftOut[4] );
nand U916 ( n1602, n1600, n1599 );
nand U917 ( n1582, n1580, n1579 );
nand U918 ( n1560, n1558, n1557 );
nand U919 ( n1557, my_FIR_filter_firBlock_left_multProducts[15], n1556 );
nand U920 ( n1550, n1548, n1547 );
nand U921 ( n1547, my_FIR_filter_firBlock_left_multProducts[13], n1546 );
nand U922 ( n1612, n1610, n1609 );
nand U923 ( n1609, my_FIR_filter_firBlock_left_multProducts[25], n1608 );
nand U924 ( n1617, n1615, n1614 );
nand U925 ( n1615, my_FIR_filter_firBlock_left_firStep[154], n1612 );
nand U926 ( n1555, n1553, n1552 );
nand U927 ( n1553, my_FIR_filter_firBlock_left_firStep[142], n1550 );
nand U928 ( n1607, n1605, n1604 );
nand U929 ( n1605, my_FIR_filter_firBlock_left_firStep[152], n1602 );
nand U930 ( n1587, n1585, n1584 );
nand U931 ( n1585, my_FIR_filter_firBlock_left_firStep[148], n1582 );
nand U932 ( n1565, n1563, n1562 );
nand U933 ( n1563, my_FIR_filter_firBlock_left_firStep[144], n1560 );
nand U934 ( n1597, n1595, n1594 );
nand U935 ( n1594, my_FIR_filter_firBlock_left_multProducts[22], n1593 );
nand U936 ( n1577, n1573, n1572 );
nand U937 ( n1573, my_FIR_filter_firBlock_left_firStep[146], n1570 );
nand U938 ( n1572, my_FIR_filter_firBlock_left_multProducts[18], n1571 );
or U939 ( n1571, n1570, my_FIR_filter_firBlock_left_firStep[146] );
nand U940 ( n1592, n1590, n1589 );
nand U941 ( n1589, my_FIR_filter_firBlock_left_multProducts[21], n1588 );
nand U942 ( n1629, n1625, n1624 );
nand U943 ( n1625, my_FIR_filter_firBlock_left_firStep[156], n1622 );
nand U944 ( n1624, my_FIR_filter_firBlock_left_multProducts[28], n1623 );
or U945 ( n1623, n1622, my_FIR_filter_firBlock_left_firStep[156] );
nand U946 ( n1635, n1632, n1631 );
nand U947 ( n1631, my_FIR_filter_firBlock_left_multProducts[29], n1630 );
nand U948 ( n1644, n1513, n1512 );
nand U949 ( n1647, n1516, n1515 );
nand U950 ( n1651, n1522, n1521 );
nand U951 ( n1533, my_FIR_filter_firBlock_left_firStep[138], n1530 );
nand U952 ( n1628, n1504, n1503 );
nand U953 ( n1504, my_FIR_filter_firBlock_left_firStep[129], n1576 );
or U954 ( n1502, my_FIR_filter_firBlock_left_firStep[129], n1576 );
nand U955 ( n1530, n1528, n1527 );
nand U956 ( n1527, my_FIR_filter_firBlock_left_multProducts[9], n1526 );
nand U957 ( n1643, n1510, n1509 );
nand U958 ( n1648, n1519, n1518 );
nand U959 ( n1519, my_FIR_filter_firBlock_left_firStep[134], n1647 );
nand U960 ( n1518, my_FIR_filter_firBlock_left_multProducts[6], n1517 );
or U961 ( n1517, n1647, my_FIR_filter_firBlock_left_firStep[134] );
nand U962 ( n1652, n1525, n1524 );
nand U963 ( n1525, my_FIR_filter_firBlock_left_firStep[136], n1651 );
nand U964 ( n1524, my_FIR_filter_firBlock_left_multProducts[8], n1523 );
or U965 ( n1523, n1651, my_FIR_filter_firBlock_left_firStep[136] );
nand U966 ( n1540, n1538, n1537 );
nand U967 ( n1537, my_FIR_filter_firBlock_left_multProducts[11], n1536 );
nand U968 ( n1545, n1543, n1542 );
nand U969 ( n1542, my_FIR_filter_firBlock_left_multProducts[12], n1541 );
nand U970 ( n1640, n1507, n1506 );
nand U971 ( n1507, my_FIR_filter_firBlock_left_firStep[130], n1628 );
or U972 ( n1505, n1628, my_FIR_filter_firBlock_left_firStep[130] );
and U973 ( n1576, my_FIR_filter_firBlock_left_multProducts[0], my_FIR_filter_firBlock_left_firStep[128] );
nand U974 ( n1164, my_FIR_filter_firBlock_left_firStep[221], n1161 );
xor U975 ( my_FIR_filter_firBlock_left_N96, n1171, n1170 );
xnor U976 ( n1171, n59, my_FIR_filter_firBlock_left_firStep[223] );
nor U977 ( n1170, n1169, n1168 );
and U978 ( n1168, n1167, my_FIR_filter_firBlock_left_firStep[222] );
nor U979 ( n1169, n1166, n119 );
nor U980 ( n1166, my_FIR_filter_firBlock_left_firStep[222], n1167 );
nand U981 ( n2243, n2240, n2239 );
nand U982 ( n2240, my_FIR_filter_firBlock_left_firStep[29], n2237 );
nand U983 ( n2239, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2238 );
or U984 ( n2238, n2237, my_FIR_filter_firBlock_left_firStep[29] );
nand U985 ( n2143, n2141, n2140 );
nand U986 ( n2141, my_FIR_filter_firBlock_left_firStep[10], n2138 );
nand U987 ( n2140, my_FIR_filter_firBlock_left_multProducts[100], n2139 );
or U988 ( n2139, n2138, my_FIR_filter_firBlock_left_firStep[10] );
nand U989 ( n2205, n2203, n2202 );
nand U990 ( n2203, my_FIR_filter_firBlock_left_firStep[22], n2200 );
nand U991 ( n2202, my_FIR_filter_firBlock_left_multProducts[112], n2201 );
or U992 ( n2201, n2200, my_FIR_filter_firBlock_left_firStep[22] );
nand U993 ( n2256, n2127, n2126 );
nand U994 ( n2127, my_FIR_filter_firBlock_left_firStep[6], n2255 );
nand U995 ( n2126, my_FIR_filter_firBlock_left_multProducts[96], n2125 );
or U996 ( n2125, n2255, my_FIR_filter_firBlock_left_firStep[6] );
nand U997 ( n2260, n2133, n2132 );
nand U998 ( n2133, my_FIR_filter_firBlock_left_firStep[8], n2259 );
nand U999 ( n2132, my_FIR_filter_firBlock_left_multProducts[98], n2131 );
or U1000 ( n2131, n2259, my_FIR_filter_firBlock_left_firStep[8] );
nand U1001 ( n2153, n2151, n2150 );
nand U1002 ( n2151, my_FIR_filter_firBlock_left_firStep[12], n2148 );
nand U1003 ( n2150, my_FIR_filter_firBlock_left_multProducts[102], n2149 );
or U1004 ( n2149, n2148, my_FIR_filter_firBlock_left_firStep[12] );
nand U1005 ( n2163, n2161, n2160 );
nand U1006 ( n2161, my_FIR_filter_firBlock_left_firStep[14], n2158 );
nand U1007 ( n2160, my_FIR_filter_firBlock_left_multProducts[104], n2159 );
or U1008 ( n2159, n2158, my_FIR_filter_firBlock_left_firStep[14] );
nand U1009 ( n2173, n2171, n2170 );
nand U1010 ( n2171, my_FIR_filter_firBlock_left_firStep[16], n2168 );
nand U1011 ( n2170, my_FIR_filter_firBlock_left_multProducts[106], n2169 );
or U1012 ( n2169, n2168, my_FIR_filter_firBlock_left_firStep[16] );
nand U1013 ( n2185, n2181, n2180 );
nand U1014 ( n2181, my_FIR_filter_firBlock_left_firStep[18], n2178 );
nand U1015 ( n2180, my_FIR_filter_firBlock_left_multProducts[108], n2179 );
or U1016 ( n2179, n2178, my_FIR_filter_firBlock_left_firStep[18] );
nand U1017 ( n2195, n2193, n2192 );
nand U1018 ( n2193, my_FIR_filter_firBlock_left_firStep[20], n2190 );
nand U1019 ( n2192, my_FIR_filter_firBlock_left_multProducts[110], n2191 );
or U1020 ( n2191, n2190, my_FIR_filter_firBlock_left_firStep[20] );
nand U1021 ( n2215, n2213, n2212 );
nand U1022 ( n2213, my_FIR_filter_firBlock_left_firStep[24], n2210 );
nand U1023 ( n2212, my_FIR_filter_firBlock_left_multProducts[114], n2211 );
or U1024 ( n2211, n2210, my_FIR_filter_firBlock_left_firStep[24] );
nand U1025 ( n2225, n2223, n2222 );
nand U1026 ( n2223, my_FIR_filter_firBlock_left_firStep[26], n2220 );
nand U1027 ( n2222, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2221 );
or U1028 ( n2221, n2220, my_FIR_filter_firBlock_left_firStep[26] );
nand U1029 ( n2237, n2233, n2232 );
nand U1030 ( n2233, my_FIR_filter_firBlock_left_firStep[28], n2230 );
nand U1031 ( n2232, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2231 );
or U1032 ( n2231, n2230, my_FIR_filter_firBlock_left_firStep[28] );
nand U1033 ( n2236, n2112, n2111 );
nand U1034 ( n2112, my_FIR_filter_firBlock_left_firStep[1], n2184 );
nand U1035 ( n2111, my_FIR_filter_firBlock_left_multProducts[91], n2110 );
or U1036 ( n2110, my_FIR_filter_firBlock_left_firStep[1], n2184 );
nand U1037 ( n2251, n2118, n2117 );
nand U1038 ( n2118, my_FIR_filter_firBlock_left_firStep[3], n2248 );
nand U1039 ( n2117, my_FIR_filter_firBlock_left_multProducts[93], n2116 );
or U1040 ( n2116, n2248, my_FIR_filter_firBlock_left_firStep[3] );
nand U1041 ( n2255, n2124, n2123 );
nand U1042 ( n2124, my_FIR_filter_firBlock_left_firStep[5], n2252 );
nand U1043 ( n2123, my_FIR_filter_firBlock_left_multProducts[95], n2122 );
or U1044 ( n2122, n2252, my_FIR_filter_firBlock_left_firStep[5] );
nand U1045 ( n2138, n2136, n2135 );
nand U1046 ( n2136, my_FIR_filter_firBlock_left_firStep[9], n2260 );
nand U1047 ( n2135, my_FIR_filter_firBlock_left_multProducts[99], n2134 );
or U1048 ( n2134, n2260, my_FIR_filter_firBlock_left_firStep[9] );
nand U1049 ( n2148, n2146, n2145 );
nand U1050 ( n2146, my_FIR_filter_firBlock_left_firStep[11], n2143 );
nand U1051 ( n2145, my_FIR_filter_firBlock_left_multProducts[101], n2144 );
or U1052 ( n2144, n2143, my_FIR_filter_firBlock_left_firStep[11] );
nand U1053 ( n2158, n2156, n2155 );
nand U1054 ( n2156, my_FIR_filter_firBlock_left_firStep[13], n2153 );
nand U1055 ( n2155, my_FIR_filter_firBlock_left_multProducts[103], n2154 );
or U1056 ( n2154, n2153, my_FIR_filter_firBlock_left_firStep[13] );
nand U1057 ( n2168, n2166, n2165 );
nand U1058 ( n2166, my_FIR_filter_firBlock_left_firStep[15], n2163 );
nand U1059 ( n2165, my_FIR_filter_firBlock_left_multProducts[105], n2164 );
or U1060 ( n2164, n2163, my_FIR_filter_firBlock_left_firStep[15] );
nand U1061 ( n2178, n2176, n2175 );
nand U1062 ( n2176, my_FIR_filter_firBlock_left_firStep[17], n2173 );
nand U1063 ( n2175, my_FIR_filter_firBlock_left_multProducts[107], n2174 );
or U1064 ( n2174, n2173, my_FIR_filter_firBlock_left_firStep[17] );
nand U1065 ( n2190, n2188, n2187 );
nand U1066 ( n2188, my_FIR_filter_firBlock_left_firStep[19], n2185 );
nand U1067 ( n2187, my_FIR_filter_firBlock_left_multProducts[109], n2186 );
or U1068 ( n2186, n2185, my_FIR_filter_firBlock_left_firStep[19] );
nand U1069 ( n2200, n2198, n2197 );
nand U1070 ( n2198, my_FIR_filter_firBlock_left_firStep[21], n2195 );
nand U1071 ( n2197, my_FIR_filter_firBlock_left_multProducts[111], n2196 );
or U1072 ( n2196, n2195, my_FIR_filter_firBlock_left_firStep[21] );
nand U1073 ( n2210, n2208, n2207 );
nand U1074 ( n2208, my_FIR_filter_firBlock_left_firStep[23], n2205 );
nand U1075 ( n2207, my_FIR_filter_firBlock_left_multProducts[113], n2206 );
or U1076 ( n2206, n2205, my_FIR_filter_firBlock_left_firStep[23] );
nand U1077 ( n2259, n2130, n2129 );
nand U1078 ( n2130, my_FIR_filter_firBlock_left_firStep[7], n2256 );
nand U1079 ( n2129, my_FIR_filter_firBlock_left_multProducts[97], n2128 );
or U1080 ( n2128, n2256, my_FIR_filter_firBlock_left_firStep[7] );
nand U1081 ( n2220, n2218, n2217 );
nand U1082 ( n2218, my_FIR_filter_firBlock_left_firStep[25], n2215 );
nand U1083 ( n2217, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2216 );
or U1084 ( n2216, n2215, my_FIR_filter_firBlock_left_firStep[25] );
nand U1085 ( n2230, n2228, n2227 );
nand U1086 ( n2228, my_FIR_filter_firBlock_left_firStep[27], n2225 );
nand U1087 ( n2227, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2226 );
or U1088 ( n2226, n2225, my_FIR_filter_firBlock_left_firStep[27] );
nor U1089 ( n2245, n2242, n57 );
nor U1090 ( n2242, my_FIR_filter_firBlock_left_firStep[30], n2243 );
xor U1091 ( my_FIR_filter_firBlock_left_N288, n2247, n2246 );
xnor U1092 ( n2247, n59, my_FIR_filter_firBlock_left_firStep[31] );
nor U1093 ( n2246, n2245, n2244 );
and U1094 ( n2244, n2243, my_FIR_filter_firBlock_left_firStep[30] );
nand U1095 ( n2248, n2115, n2114 );
nand U1096 ( n2115, my_FIR_filter_firBlock_left_firStep[2], n2236 );
nand U1097 ( n2114, my_FIR_filter_firBlock_left_multProducts[92], n2113 );
or U1098 ( n2113, n2236, my_FIR_filter_firBlock_left_firStep[2] );
nand U1099 ( n2252, n2121, n2120 );
nand U1100 ( n2121, my_FIR_filter_firBlock_left_firStep[4], n2251 );
nand U1101 ( n2120, my_FIR_filter_firBlock_left_multProducts[94], n2119 );
or U1102 ( n2119, n2251, my_FIR_filter_firBlock_left_firStep[4] );
nand U1103 ( my_FIR_filter_firBlock_left_multProducts[60], n871, n870 );
nand U1104 ( n871, my_FIR_filter_firBlock_left_multProducts[114], n868 );
nand U1105 ( n870, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n869 );
or U1106 ( n869, n868, my_FIR_filter_firBlock_left_multProducts[114] );
nand U1107 ( n1149, n1147, n1146 );
nand U1108 ( n1147, my_FIR_filter_firBlock_left_firStep[218], n1144 );
nand U1109 ( n1154, n1152, n1151 );
nand U1110 ( n1152, my_FIR_filter_firBlock_left_firStep[219], n1149 );
nand U1111 ( n1151, my_FIR_filter_firBlock_left_multProducts[57], n1150 );
or U1112 ( n1150, n1149, my_FIR_filter_firBlock_left_firStep[219] );
nand U1113 ( n1161, n1157, n1156 );
nand U1114 ( n1157, my_FIR_filter_firBlock_left_firStep[220], n1154 );
or U1115 ( n1155, n1154, my_FIR_filter_firBlock_left_firStep[220] );
nand U1116 ( n1737, my_FIR_filter_firBlock_left_firStep[116], n1734 );
nand U1117 ( n1720, my_FIR_filter_firBlock_left_firStep[113], n1717 );
nand U1118 ( n1787, n1784, n1783 );
nand U1119 ( n1784, my_FIR_filter_firBlock_left_firStep[125], n1781 );
or U1120 ( n1782, n1781, my_FIR_filter_firBlock_left_firStep[125] );
nand U1121 ( n1707, n1705, n1704 );
nand U1122 ( n1705, my_FIR_filter_firBlock_left_firStep[110], n1702 );
nand U1123 ( n1744, n1742, n1741 );
nand U1124 ( n1742, my_FIR_filter_firBlock_left_firStep[117], n1739 );
nand U1125 ( n1741, my_FIR_filter_firBlock_left_multProducts[51], n1740 );
or U1126 ( n1740, n1739, my_FIR_filter_firBlock_left_firStep[117] );
nand U1127 ( n1702, n1700, n1699 );
nand U1128 ( n1700, my_FIR_filter_firBlock_left_firStep[109], n1697 );
nand U1129 ( n1699, my_FIR_filter_firBlock_left_multProducts[43], n1698 );
or U1130 ( n1698, n1697, my_FIR_filter_firBlock_left_firStep[109] );
nand U1131 ( n1749, n1747, n1746 );
nand U1132 ( n1747, my_FIR_filter_firBlock_left_firStep[118], n1744 );
nand U1133 ( n1746, my_FIR_filter_firBlock_left_multProducts[52], n1745 );
or U1134 ( n1745, n1744, my_FIR_filter_firBlock_left_firStep[118] );
nand U1135 ( n1729, n1725, n1724 );
nand U1136 ( n1725, my_FIR_filter_firBlock_left_firStep[114], n1722 );
nand U1137 ( n1724, my_FIR_filter_firBlock_left_multProducts[48], n1723 );
or U1138 ( n1723, n1722, my_FIR_filter_firBlock_left_firStep[114] );
nand U1139 ( n1697, n1695, n1694 );
nand U1140 ( n1695, my_FIR_filter_firBlock_left_firStep[108], n1692 );
nand U1141 ( n1694, my_FIR_filter_firBlock_left_multProducts[42], n1693 );
or U1142 ( n1693, n1692, my_FIR_filter_firBlock_left_firStep[108] );
nand U1143 ( n1774, n1772, n1771 );
nand U1144 ( n1772, my_FIR_filter_firBlock_left_firStep[123], n1769 );
nand U1145 ( n1764, n1762, n1761 );
nand U1146 ( n1762, my_FIR_filter_firBlock_left_firStep[121], n1759 );
nand U1147 ( n1781, n1777, n1776 );
nand U1148 ( n1777, my_FIR_filter_firBlock_left_firStep[124], n1774 );
or U1149 ( n1775, n1774, my_FIR_filter_firBlock_left_firStep[124] );
xnor U1150 ( n1791, n59, my_FIR_filter_firBlock_left_firStep[127] );
and U1151 ( n1788, n1787, my_FIR_filter_firBlock_left_firStep[126] );
nand U1152 ( n1712, n1710, n1709 );
nand U1153 ( n1710, my_FIR_filter_firBlock_left_firStep[111], n1707 );
nand U1154 ( n1709, my_FIR_filter_firBlock_left_multProducts[45], n1708 );
or U1155 ( n1708, n1707, my_FIR_filter_firBlock_left_firStep[111] );
nand U1156 ( n1692, n1690, n1689 );
nand U1157 ( n1690, my_FIR_filter_firBlock_left_firStep[107], n1687 );
nand U1158 ( n1689, my_FIR_filter_firBlock_left_multProducts[41], n1688 );
or U1159 ( n1688, n1687, my_FIR_filter_firBlock_left_firStep[107] );
nand U1160 ( n1759, n1757, n1756 );
nand U1161 ( n1757, my_FIR_filter_firBlock_left_firStep[120], n1754 );
nand U1162 ( n1769, n1767, n1766 );
nand U1163 ( n1767, my_FIR_filter_firBlock_left_firStep[122], n1764 );
nand U1164 ( n1766, my_FIR_filter_firBlock_left_multProducts[56], n1765 );
or U1165 ( n1765, n1764, my_FIR_filter_firBlock_left_firStep[122] );
nand U1166 ( n1717, n1715, n1714 );
nand U1167 ( n1715, my_FIR_filter_firBlock_left_firStep[112], n1712 );
nand U1168 ( n1714, my_FIR_filter_firBlock_left_multProducts[46], n1713 );
or U1169 ( n1713, n1712, my_FIR_filter_firBlock_left_firStep[112] );
nand U1170 ( n1754, n1752, n1751 );
nand U1171 ( n1752, my_FIR_filter_firBlock_left_firStep[119], n1749 );
nand U1172 ( n1751, my_FIR_filter_firBlock_left_multProducts[53], n1750 );
or U1173 ( n1750, n1749, my_FIR_filter_firBlock_left_firStep[119] );
nand U1174 ( n1734, n1732, n1731 );
nand U1175 ( n1732, my_FIR_filter_firBlock_left_firStep[115], n1729 );
nand U1176 ( n1731, my_FIR_filter_firBlock_left_multProducts[49], n1730 );
or U1177 ( n1730, n1729, my_FIR_filter_firBlock_left_firStep[115] );
nor U1178 ( n1789, n1786, n119 );
nor U1179 ( n1786, my_FIR_filter_firBlock_left_firStep[126], n1787 );
nand U1180 ( n1687, n1685, n1684 );
nand U1181 ( n1685, my_FIR_filter_firBlock_left_firStep[106], n1682 );
nand U1182 ( n1682, n1680, n1679 );
nand U1183 ( n1680, my_FIR_filter_firBlock_left_firStep[105], n1804 );
nand U1184 ( n1679, my_FIR_filter_firBlock_left_multProducts[39], n1678 );
or U1185 ( n1678, n1804, my_FIR_filter_firBlock_left_firStep[105] );
nand U1186 ( n1134, n1132, n1131 );
nand U1187 ( n1132, my_FIR_filter_firBlock_left_firStep[215], n1129 );
nand U1188 ( n1139, n1137, n1136 );
nand U1189 ( n1137, my_FIR_filter_firBlock_left_firStep[216], n1134 );
nand U1190 ( n1136, my_FIR_filter_firBlock_left_multProducts[54], n1135 );
or U1191 ( n1135, n1134, my_FIR_filter_firBlock_left_firStep[216] );
nand U1192 ( n1129, n1127, n1126 );
nand U1193 ( n1127, my_FIR_filter_firBlock_left_firStep[214], n1124 );
nand U1194 ( n1126, my_FIR_filter_firBlock_left_multProducts[52], n1125 );
or U1195 ( n1125, n1124, my_FIR_filter_firBlock_left_firStep[214] );
nand U1196 ( n1144, n1142, n1141 );
nand U1197 ( n1142, my_FIR_filter_firBlock_left_firStep[217], n1139 );
nand U1198 ( n1124, n1122, n1121 );
nand U1199 ( n1122, my_FIR_filter_firBlock_left_firStep[213], n1119 );
nand U1200 ( n1804, n1677, n1676 );
nand U1201 ( n1677, my_FIR_filter_firBlock_left_firStep[104], n1803 );
nand U1202 ( n1799, n1668, n1667 );
nand U1203 ( n1668, my_FIR_filter_firBlock_left_firStep[101], n1796 );
nand U1204 ( n1780, n1656, n1655 );
nand U1205 ( n1656, my_FIR_filter_firBlock_left_firStep[97], n1728 );
nand U1206 ( n1655, my_FIR_filter_firBlock_left_multProducts[31], n1654 );
or U1207 ( n1654, my_FIR_filter_firBlock_left_firStep[97], n1728 );
nand U1208 ( n1796, n1665, n1664 );
nand U1209 ( n1665, my_FIR_filter_firBlock_left_firStep[100], n1795 );
nand U1210 ( n1795, n1662, n1661 );
nand U1211 ( n1662, my_FIR_filter_firBlock_left_firStep[99], n1792 );
nand U1212 ( n1803, n1674, n1673 );
nand U1213 ( n1674, my_FIR_filter_firBlock_left_firStep[103], n1800 );
nand U1214 ( n1800, n1671, n1670 );
nand U1215 ( n1671, my_FIR_filter_firBlock_left_firStep[102], n1799 );
nand U1216 ( n1670, my_FIR_filter_firBlock_left_multProducts[36], n1669 );
or U1217 ( n1669, n1799, my_FIR_filter_firBlock_left_firStep[102] );
and U1218 ( n1728, my_FIR_filter_firBlock_left_multProducts[30], my_FIR_filter_firBlock_left_firStep[96] );
nand U1219 ( n1792, n1659, n1658 );
nand U1220 ( n1659, my_FIR_filter_firBlock_left_firStep[98], n1780 );
nand U1221 ( n1658, my_FIR_filter_firBlock_left_multProducts[32], n1657 );
or U1222 ( n1657, n1780, my_FIR_filter_firBlock_left_firStep[98] );
nand U1223 ( n1114, n1112, n1111 );
nand U1224 ( n1112, my_FIR_filter_firBlock_left_firStep[211], n1109 );
nand U1225 ( n1119, n1117, n1116 );
nand U1226 ( n1117, my_FIR_filter_firBlock_left_firStep[212], n1114 );
nand U1227 ( n1116, my_FIR_filter_firBlock_left_multProducts[50], n1115 );
or U1228 ( n1115, n1114, my_FIR_filter_firBlock_left_firStep[212] );
nand U1229 ( n1082, n1080, n1079 );
nand U1230 ( n1080, my_FIR_filter_firBlock_left_firStep[205], n1077 );
nand U1231 ( n1062, n1060, n1059 );
nand U1232 ( n1060, my_FIR_filter_firBlock_left_firStep[201], n1184 );
nand U1233 ( n1097, n1095, n1094 );
nand U1234 ( n1095, my_FIR_filter_firBlock_left_firStep[208], n1092 );
nand U1235 ( n1180, n1051, n1050 );
nand U1236 ( n1051, my_FIR_filter_firBlock_left_firStep[198], n1179 );
nand U1237 ( n1160, n1036, n1035 );
nand U1238 ( n1036, my_FIR_filter_firBlock_left_firStep[193], n1108 );
nand U1239 ( n1035, my_FIR_filter_firBlock_left_multProducts[31], n1034 );
or U1240 ( n1034, my_FIR_filter_firBlock_left_firStep[193], n1108 );
nand U1241 ( n1175, n1042, n1041 );
nand U1242 ( n1042, my_FIR_filter_firBlock_left_firStep[195], n1172 );
nand U1243 ( n1041, my_FIR_filter_firBlock_left_multProducts[33], n1040 );
or U1244 ( n1040, n1172, my_FIR_filter_firBlock_left_firStep[195] );
nand U1245 ( n1109, n1105, n1104 );
nand U1246 ( n1105, my_FIR_filter_firBlock_left_firStep[210], n1102 );
nand U1247 ( n1184, n1057, n1056 );
nand U1248 ( n1057, my_FIR_filter_firBlock_left_firStep[200], n1183 );
nand U1249 ( n1092, n1090, n1089 );
nand U1250 ( n1090, my_FIR_filter_firBlock_left_firStep[207], n1087 );
nand U1251 ( n1179, n1048, n1047 );
nand U1252 ( n1048, my_FIR_filter_firBlock_left_firStep[197], n1176 );
nand U1253 ( n1087, n1085, n1084 );
nand U1254 ( n1085, my_FIR_filter_firBlock_left_firStep[206], n1082 );
nand U1255 ( n1084, my_FIR_filter_firBlock_left_multProducts[44], n1083 );
or U1256 ( n1083, n1082, my_FIR_filter_firBlock_left_firStep[206] );
nand U1257 ( n1077, n1075, n1074 );
nand U1258 ( n1075, my_FIR_filter_firBlock_left_firStep[204], n1072 );
nand U1259 ( n1074, my_FIR_filter_firBlock_left_multProducts[42], n1073 );
or U1260 ( n1073, n1072, my_FIR_filter_firBlock_left_firStep[204] );
nand U1261 ( n1176, n1045, n1044 );
nand U1262 ( n1045, my_FIR_filter_firBlock_left_firStep[196], n1175 );
nand U1263 ( n1044, my_FIR_filter_firBlock_left_multProducts[34], n1043 );
or U1264 ( n1043, n1175, my_FIR_filter_firBlock_left_firStep[196] );
nand U1265 ( n1067, n1065, n1064 );
nand U1266 ( n1065, my_FIR_filter_firBlock_left_firStep[202], n1062 );
nand U1267 ( n1064, my_FIR_filter_firBlock_left_multProducts[40], n1063 );
or U1268 ( n1063, n1062, my_FIR_filter_firBlock_left_firStep[202] );
nand U1269 ( n1102, n1100, n1099 );
nand U1270 ( n1100, my_FIR_filter_firBlock_left_firStep[209], n1097 );
nand U1271 ( n1099, my_FIR_filter_firBlock_left_multProducts[47], n1098 );
or U1272 ( n1098, n1097, my_FIR_filter_firBlock_left_firStep[209] );
and U1273 ( n1108, my_FIR_filter_firBlock_left_multProducts[30], my_FIR_filter_firBlock_left_firStep[192] );
nand U1274 ( n1072, n1070, n1069 );
nand U1275 ( n1070, my_FIR_filter_firBlock_left_firStep[203], n1067 );
nand U1276 ( n1172, n1039, n1038 );
nand U1277 ( n1039, my_FIR_filter_firBlock_left_firStep[194], n1160 );
nand U1278 ( n1038, my_FIR_filter_firBlock_left_multProducts[32], n1037 );
or U1279 ( n1037, n1160, my_FIR_filter_firBlock_left_firStep[194] );
nand U1280 ( n1183, n1054, n1053 );
nand U1281 ( n1054, my_FIR_filter_firBlock_left_firStep[199], n1180 );
nand U1282 ( n1053, my_FIR_filter_firBlock_left_multProducts[37], n1052 );
or U1283 ( n1052, n1180, my_FIR_filter_firBlock_left_firStep[199] );
xor U1284 ( my_FIR_filter_firBlock_left_N63, n1015, n1013 );
xnor U1285 ( n1013, n57, my_FIR_filter_firBlock_left_firStep[254] );
xnor U1286 ( n700, n120, my_FIR_filter_firBlock_left_firStep[284] );
xnor U1287 ( n2077, n120, my_FIR_filter_firBlock_left_firStep[60] );
xnor U1288 ( n1937, n57, my_FIR_filter_firBlock_left_firStep[94] );
xor U1289 ( outData_in[30], n262, n260 );
xnor U1290 ( n260, n49, leftOut[30] );
xor U1291 ( my_FIR_filter_firBlock_left_N95, n1167, n1165 );
xnor U1292 ( n1165, n119, my_FIR_filter_firBlock_left_firStep[222] );
xor U1293 ( my_FIR_filter_firBlock_left_N191, n1787, n1785 );
xnor U1294 ( n1785, n119, my_FIR_filter_firBlock_left_firStep[126] );
xnor U1295 ( my_FIR_filter_firBlock_left_N126, n1474, n1477 );
xnor U1296 ( n1474, my_FIR_filter_firBlock_left_firStep[189], my_FIR_filter_firBlock_left_multProducts[29] );
xnor U1297 ( n1626, my_FIR_filter_firBlock_left_firStep[157], my_FIR_filter_firBlock_left_multProducts[29] );
xnor U1298 ( outData_in[29], n253, n256 );
xnor U1299 ( n253, leftOut[29], rightOut[29] );
xor U1300 ( my_FIR_filter_firBlock_left_N287, n2243, n2241 );
xnor U1301 ( n2241, n57, my_FIR_filter_firBlock_left_firStep[30] );
xnor U1302 ( my_FIR_filter_firBlock_left_N222, n1930, n1933 );
xnor U1303 ( n1930, my_FIR_filter_firBlock_left_firStep[93], my_FIR_filter_firBlock_left_multProducts[60] );
xnor U1304 ( my_FIR_filter_firBlock_left_N62, n1006, n1009 );
xnor U1305 ( n1006, my_FIR_filter_firBlock_left_firStep[253], my_FIR_filter_firBlock_left_multProducts[60] );
xor U1306 ( my_FIR_filter_firBlock_left_N221, n1926, n1925 );
xor U1307 ( n1925, my_FIR_filter_firBlock_left_multProducts[59], my_FIR_filter_firBlock_left_firStep[92] );
xor U1308 ( my_FIR_filter_firBlock_left_N61, n1002, n1001 );
xor U1309 ( n1001, my_FIR_filter_firBlock_left_multProducts[59], my_FIR_filter_firBlock_left_firStep[252] );
xnor U1310 ( my_FIR_filter_firBlock_left_N190, n1778, n1781 );
xnor U1311 ( n1778, my_FIR_filter_firBlock_left_firStep[125], my_FIR_filter_firBlock_left_multProducts[59] );
xnor U1312 ( my_FIR_filter_firBlock_left_N94, n1158, n1161 );
xnor U1313 ( n1158, my_FIR_filter_firBlock_left_firStep[221], my_FIR_filter_firBlock_left_multProducts[59] );
xor U1314 ( outData_in[28], n249, n248 );
xor U1315 ( n248, rightOut[28], leftOut[28] );
xor U1316 ( my_FIR_filter_firBlock_left_N157, n1622, n1621 );
xor U1317 ( n1621, my_FIR_filter_firBlock_left_multProducts[28], my_FIR_filter_firBlock_left_firStep[156] );
xor U1318 ( n1469, my_FIR_filter_firBlock_left_multProducts[28], my_FIR_filter_firBlock_left_firStep[188] );
xnor U1319 ( my_FIR_filter_firBlock_left_N286, n2234, n2237 );
xnor U1320 ( n2234, my_FIR_filter_firBlock_left_firStep[29], n59 );
xnor U1321 ( outData_in[27], n243, n244 );
xnor U1322 ( n243, leftOut[27], rightOut[27] );
xor U1323 ( my_FIR_filter_firBlock_left_N189, n1774, n1773 );
xor U1324 ( my_FIR_filter_firBlock_left_N93, n1154, n1153 );
xnor U1325 ( my_FIR_filter_firBlock_left_N220, n1920, n1921 );
xnor U1326 ( my_FIR_filter_firBlock_left_N60, n996, n997 );
xnor U1327 ( n1616, my_FIR_filter_firBlock_left_firStep[155], my_FIR_filter_firBlock_left_multProducts[27] );
xnor U1328 ( n1464, my_FIR_filter_firBlock_left_firStep[187], my_FIR_filter_firBlock_left_multProducts[27] );
xor U1329 ( outData_in[26], n239, n238 );
xor U1330 ( n238, rightOut[26], leftOut[26] );
xor U1331 ( my_FIR_filter_firBlock_left_N219, n1916, n1915 );
xor U1332 ( n1915, my_FIR_filter_firBlock_left_multProducts[57], my_FIR_filter_firBlock_left_firStep[90] );
xor U1333 ( my_FIR_filter_firBlock_left_N59, n992, n991 );
xor U1334 ( n991, my_FIR_filter_firBlock_left_multProducts[57], my_FIR_filter_firBlock_left_firStep[250] );
xor U1335 ( my_FIR_filter_firBlock_left_N285, n2230, n2229 );
xnor U1336 ( n2229, n57, my_FIR_filter_firBlock_left_firStep[28] );
xnor U1337 ( my_FIR_filter_firBlock_left_N92, n1148, n1149 );
xnor U1338 ( n1148, my_FIR_filter_firBlock_left_firStep[219], my_FIR_filter_firBlock_left_multProducts[57] );
xnor U1339 ( my_FIR_filter_firBlock_left_N188, n1768, n1769 );
xnor U1340 ( n1768, my_FIR_filter_firBlock_left_firStep[123], my_FIR_filter_firBlock_left_multProducts[57] );
xor U1341 ( my_FIR_filter_firBlock_left_N155, n1612, n1611 );
xor U1342 ( n1611, my_FIR_filter_firBlock_left_multProducts[26], my_FIR_filter_firBlock_left_firStep[154] );
xor U1343 ( my_FIR_filter_firBlock_left_N123, n1460, n1459 );
xor U1344 ( n1459, my_FIR_filter_firBlock_left_multProducts[26], my_FIR_filter_firBlock_left_firStep[186] );
xnor U1345 ( outData_in[25], n233, n234 );
xnor U1346 ( n233, leftOut[25], rightOut[25] );
xor U1347 ( my_FIR_filter_firBlock_left_N187, n1764, n1763 );
xor U1348 ( n1763, my_FIR_filter_firBlock_left_multProducts[56], my_FIR_filter_firBlock_left_firStep[122] );
xor U1349 ( my_FIR_filter_firBlock_left_N91, n1144, n1143 );
xor U1350 ( n1143, my_FIR_filter_firBlock_left_multProducts[56], my_FIR_filter_firBlock_left_firStep[218] );
xnor U1351 ( my_FIR_filter_firBlock_left_N58, n986, n987 );
xnor U1352 ( n986, my_FIR_filter_firBlock_left_firStep[249], my_FIR_filter_firBlock_left_multProducts[56] );
xnor U1353 ( my_FIR_filter_firBlock_left_N218, n1910, n1911 );
xnor U1354 ( n1910, my_FIR_filter_firBlock_left_firStep[89], my_FIR_filter_firBlock_left_multProducts[56] );
xnor U1355 ( my_FIR_filter_firBlock_left_N284, n2224, n2225 );
xnor U1356 ( n2224, my_FIR_filter_firBlock_left_firStep[27], n59 );
xor U1357 ( outData_in[24], n229, n228 );
xor U1358 ( n228, rightOut[24], leftOut[24] );
xnor U1359 ( my_FIR_filter_firBlock_left_N122, n1454, n1455 );
xnor U1360 ( n1454, my_FIR_filter_firBlock_left_firStep[185], my_FIR_filter_firBlock_left_multProducts[25] );
xnor U1361 ( n1606, my_FIR_filter_firBlock_left_firStep[153], my_FIR_filter_firBlock_left_multProducts[25] );
xor U1362 ( my_FIR_filter_firBlock_left_N217, n1906, n1905 );
xor U1363 ( n1905, my_FIR_filter_firBlock_left_multProducts[55], my_FIR_filter_firBlock_left_firStep[88] );
xor U1364 ( my_FIR_filter_firBlock_left_N57, n982, n981 );
xor U1365 ( n981, my_FIR_filter_firBlock_left_multProducts[55], my_FIR_filter_firBlock_left_firStep[248] );
xor U1366 ( n670, my_FIR_filter_firBlock_left_multProducts[83], my_FIR_filter_firBlock_left_firStep[278] );
xor U1367 ( n2047, my_FIR_filter_firBlock_left_multProducts[83], my_FIR_filter_firBlock_left_firStep[54] );
xor U1368 ( my_FIR_filter_firBlock_left_N283, n2220, n2219 );
xnor U1369 ( n2219, n57, my_FIR_filter_firBlock_left_firStep[26] );
xor U1370 ( my_FIR_filter_firBlock_left_N153, n1602, n1601 );
xor U1371 ( n1601, my_FIR_filter_firBlock_left_multProducts[24], my_FIR_filter_firBlock_left_firStep[152] );
xnor U1372 ( my_FIR_filter_firBlock_left_N186, n1758, n1759 );
xnor U1373 ( n1758, my_FIR_filter_firBlock_left_firStep[121], my_FIR_filter_firBlock_left_multProducts[55] );
xnor U1374 ( my_FIR_filter_firBlock_left_N90, n1138, n1139 );
xnor U1375 ( n1138, my_FIR_filter_firBlock_left_firStep[217], my_FIR_filter_firBlock_left_multProducts[55] );
xnor U1376 ( outData_in[23], n223, n224 );
xnor U1377 ( n223, leftOut[23], rightOut[23] );
xor U1378 ( n1449, my_FIR_filter_firBlock_left_multProducts[24], my_FIR_filter_firBlock_left_firStep[184] );
xor U1379 ( outData_in[22], n219, n218 );
xor U1380 ( n218, rightOut[22], leftOut[22] );
xor U1381 ( my_FIR_filter_firBlock_left_N185, n1754, n1753 );
xor U1382 ( n1753, my_FIR_filter_firBlock_left_multProducts[54], my_FIR_filter_firBlock_left_firStep[120] );
xor U1383 ( my_FIR_filter_firBlock_left_N89, n1134, n1133 );
xor U1384 ( n1133, my_FIR_filter_firBlock_left_multProducts[54], my_FIR_filter_firBlock_left_firStep[216] );
xnor U1385 ( n665, my_FIR_filter_firBlock_left_firStep[277], my_FIR_filter_firBlock_left_multProducts[82] );
xnor U1386 ( n2042, my_FIR_filter_firBlock_left_firStep[53], my_FIR_filter_firBlock_left_multProducts[82] );
xnor U1387 ( my_FIR_filter_firBlock_left_N216, n1900, n1901 );
xnor U1388 ( n1900, my_FIR_filter_firBlock_left_firStep[87], my_FIR_filter_firBlock_left_multProducts[54] );
xnor U1389 ( my_FIR_filter_firBlock_left_N56, n976, n977 );
xnor U1390 ( n976, my_FIR_filter_firBlock_left_firStep[247], my_FIR_filter_firBlock_left_multProducts[54] );
xnor U1391 ( my_FIR_filter_firBlock_left_N282, n2214, n2215 );
xnor U1392 ( n2214, my_FIR_filter_firBlock_left_firStep[25], n59 );
xnor U1393 ( n1596, my_FIR_filter_firBlock_left_firStep[151], my_FIR_filter_firBlock_left_multProducts[23] );
xnor U1394 ( n1444, my_FIR_filter_firBlock_left_firStep[183], my_FIR_filter_firBlock_left_multProducts[23] );
xnor U1395 ( outData_in[21], n213, n214 );
xnor U1396 ( n213, leftOut[21], rightOut[21] );
xor U1397 ( n2037, my_FIR_filter_firBlock_left_multProducts[81], my_FIR_filter_firBlock_left_firStep[52] );
xor U1398 ( n660, my_FIR_filter_firBlock_left_multProducts[81], my_FIR_filter_firBlock_left_firStep[276] );
xor U1399 ( my_FIR_filter_firBlock_left_N119, n1440, n1439 );
xor U1400 ( n1439, my_FIR_filter_firBlock_left_multProducts[22], my_FIR_filter_firBlock_left_firStep[182] );
xor U1401 ( my_FIR_filter_firBlock_left_N215, n1896, n1895 );
xor U1402 ( n1895, my_FIR_filter_firBlock_left_multProducts[53], my_FIR_filter_firBlock_left_firStep[86] );
xor U1403 ( my_FIR_filter_firBlock_left_N55, n972, n971 );
xor U1404 ( n971, my_FIR_filter_firBlock_left_multProducts[53], my_FIR_filter_firBlock_left_firStep[246] );
xor U1405 ( n1591, my_FIR_filter_firBlock_left_multProducts[22], my_FIR_filter_firBlock_left_firStep[150] );
xnor U1406 ( my_FIR_filter_firBlock_left_N184, n1748, n1749 );
xnor U1407 ( n1748, my_FIR_filter_firBlock_left_firStep[119], my_FIR_filter_firBlock_left_multProducts[53] );
xnor U1408 ( my_FIR_filter_firBlock_left_N88, n1128, n1129 );
xnor U1409 ( n1128, my_FIR_filter_firBlock_left_firStep[215], my_FIR_filter_firBlock_left_multProducts[53] );
xor U1410 ( my_FIR_filter_firBlock_left_N281, n2210, n2209 );
xor U1411 ( n2209, my_FIR_filter_firBlock_left_multProducts[114], my_FIR_filter_firBlock_left_firStep[24] );
xor U1412 ( outData_in[20], n209, n208 );
xor U1413 ( n208, rightOut[20], leftOut[20] );
xor U1414 ( my_FIR_filter_firBlock_left_N183, n1744, n1743 );
xor U1415 ( n1743, my_FIR_filter_firBlock_left_multProducts[52], my_FIR_filter_firBlock_left_firStep[118] );
xor U1416 ( my_FIR_filter_firBlock_left_N87, n1124, n1123 );
xor U1417 ( n1123, my_FIR_filter_firBlock_left_multProducts[52], my_FIR_filter_firBlock_left_firStep[214] );
xnor U1418 ( my_FIR_filter_firBlock_left_N54, n966, n967 );
xnor U1419 ( n966, my_FIR_filter_firBlock_left_firStep[245], my_FIR_filter_firBlock_left_multProducts[52] );
xnor U1420 ( my_FIR_filter_firBlock_left_N214, n1890, n1891 );
xnor U1421 ( n1890, my_FIR_filter_firBlock_left_firStep[85], my_FIR_filter_firBlock_left_multProducts[52] );
xnor U1422 ( n1586, my_FIR_filter_firBlock_left_firStep[149], my_FIR_filter_firBlock_left_multProducts[21] );
xnor U1423 ( n1434, my_FIR_filter_firBlock_left_firStep[181], my_FIR_filter_firBlock_left_multProducts[21] );
xnor U1424 ( my_FIR_filter_firBlock_left_N20, n653, n656 );
xnor U1425 ( my_FIR_filter_firBlock_left_N280, n2204, n2205 );
xnor U1426 ( n2204, my_FIR_filter_firBlock_left_firStep[23], my_FIR_filter_firBlock_left_multProducts[113] );
xnor U1427 ( outData_in[19], n201, n204 );
xnor U1428 ( n201, leftOut[19], rightOut[19] );
xor U1429 ( n648, my_FIR_filter_firBlock_left_multProducts[79], my_FIR_filter_firBlock_left_firStep[274] );
xor U1430 ( n2025, my_FIR_filter_firBlock_left_multProducts[79], my_FIR_filter_firBlock_left_firStep[50] );
xor U1431 ( my_FIR_filter_firBlock_left_N149, n1582, n1581 );
xor U1432 ( n1581, my_FIR_filter_firBlock_left_multProducts[20], my_FIR_filter_firBlock_left_firStep[148] );
xor U1433 ( my_FIR_filter_firBlock_left_N117, n1430, n1429 );
xor U1434 ( n1429, my_FIR_filter_firBlock_left_multProducts[20], my_FIR_filter_firBlock_left_firStep[180] );
xor U1435 ( outData_in[18], n197, n196 );
xor U1436 ( n196, rightOut[18], leftOut[18] );
xor U1437 ( my_FIR_filter_firBlock_left_N213, n1886, n1885 );
xor U1438 ( n1885, my_FIR_filter_firBlock_left_multProducts[51], my_FIR_filter_firBlock_left_firStep[84] );
xor U1439 ( my_FIR_filter_firBlock_left_N53, n962, n961 );
xor U1440 ( n961, my_FIR_filter_firBlock_left_multProducts[51], my_FIR_filter_firBlock_left_firStep[244] );
xnor U1441 ( my_FIR_filter_firBlock_left_N182, n1738, n1739 );
xnor U1442 ( n1738, my_FIR_filter_firBlock_left_firStep[117], my_FIR_filter_firBlock_left_multProducts[51] );
xnor U1443 ( my_FIR_filter_firBlock_left_N86, n1118, n1119 );
xnor U1444 ( n1118, my_FIR_filter_firBlock_left_firStep[213], my_FIR_filter_firBlock_left_multProducts[51] );
xor U1445 ( my_FIR_filter_firBlock_left_N279, n2200, n2199 );
xor U1446 ( n2199, my_FIR_filter_firBlock_left_multProducts[112], my_FIR_filter_firBlock_left_firStep[22] );
xor U1447 ( my_FIR_filter_firBlock_left_N85, n1114, n1113 );
xor U1448 ( n1113, my_FIR_filter_firBlock_left_multProducts[50], my_FIR_filter_firBlock_left_firStep[212] );
xor U1449 ( my_FIR_filter_firBlock_left_N181, n1734, n1733 );
xor U1450 ( n1733, my_FIR_filter_firBlock_left_multProducts[50], my_FIR_filter_firBlock_left_firStep[116] );
xnor U1451 ( my_FIR_filter_firBlock_left_N116, n1422, n1425 );
xnor U1452 ( n1422, my_FIR_filter_firBlock_left_firStep[179], my_FIR_filter_firBlock_left_multProducts[19] );
xnor U1453 ( n2020, my_FIR_filter_firBlock_left_firStep[49], my_FIR_filter_firBlock_left_multProducts[78] );
xnor U1454 ( n643, my_FIR_filter_firBlock_left_firStep[273], my_FIR_filter_firBlock_left_multProducts[78] );
xnor U1455 ( outData_in[17], n191, n192 );
xnor U1456 ( n191, leftOut[17], rightOut[17] );
xnor U1457 ( n1574, my_FIR_filter_firBlock_left_firStep[147], my_FIR_filter_firBlock_left_multProducts[19] );
xnor U1458 ( my_FIR_filter_firBlock_left_N212, n1878, n1881 );
xnor U1459 ( n1878, my_FIR_filter_firBlock_left_firStep[83], my_FIR_filter_firBlock_left_multProducts[50] );
xnor U1460 ( my_FIR_filter_firBlock_left_N52, n954, n957 );
xnor U1461 ( n954, my_FIR_filter_firBlock_left_firStep[243], my_FIR_filter_firBlock_left_multProducts[50] );
xor U1462 ( my_FIR_filter_firBlock_left_N241, n2016, n2015 );
xor U1463 ( n2015, my_FIR_filter_firBlock_left_multProducts[77], my_FIR_filter_firBlock_left_firStep[48] );
xnor U1464 ( my_FIR_filter_firBlock_left_N278, n2194, n2195 );
xnor U1465 ( n2194, my_FIR_filter_firBlock_left_firStep[21], my_FIR_filter_firBlock_left_multProducts[111] );
xor U1466 ( outData_in[16], n187, n186 );
xor U1467 ( n186, rightOut[16], leftOut[16] );
xor U1468 ( n638, my_FIR_filter_firBlock_left_multProducts[77], my_FIR_filter_firBlock_left_firStep[272] );
xor U1469 ( my_FIR_filter_firBlock_left_N147, n1570, n1569 );
xor U1470 ( n1569, my_FIR_filter_firBlock_left_multProducts[18], my_FIR_filter_firBlock_left_firStep[146] );
xor U1471 ( n1417, my_FIR_filter_firBlock_left_multProducts[18], my_FIR_filter_firBlock_left_firStep[178] );
xor U1472 ( my_FIR_filter_firBlock_left_N211, n1874, n1873 );
xor U1473 ( n1873, my_FIR_filter_firBlock_left_multProducts[49], my_FIR_filter_firBlock_left_firStep[82] );
xor U1474 ( my_FIR_filter_firBlock_left_N51, n950, n949 );
xor U1475 ( n949, my_FIR_filter_firBlock_left_multProducts[49], my_FIR_filter_firBlock_left_firStep[242] );
xnor U1476 ( my_FIR_filter_firBlock_left_N180, n1726, n1729 );
xnor U1477 ( n1726, my_FIR_filter_firBlock_left_firStep[115], my_FIR_filter_firBlock_left_multProducts[49] );
xnor U1478 ( my_FIR_filter_firBlock_left_N84, n1106, n1109 );
xnor U1479 ( n1106, my_FIR_filter_firBlock_left_firStep[211], my_FIR_filter_firBlock_left_multProducts[49] );
xor U1480 ( my_FIR_filter_firBlock_left_N277, n2190, n2189 );
xor U1481 ( n2189, my_FIR_filter_firBlock_left_multProducts[110], my_FIR_filter_firBlock_left_firStep[20] );
xnor U1482 ( outData_in[15], n181, n182 );
xnor U1483 ( n181, leftOut[15], rightOut[15] );
xnor U1484 ( my_FIR_filter_firBlock_left_N16, n633, n634 );
xnor U1485 ( n633, my_FIR_filter_firBlock_left_firStep[271], my_FIR_filter_firBlock_left_multProducts[76] );
xnor U1486 ( n2010, my_FIR_filter_firBlock_left_firStep[47], my_FIR_filter_firBlock_left_multProducts[76] );
xnor U1487 ( n1564, my_FIR_filter_firBlock_left_firStep[145], my_FIR_filter_firBlock_left_multProducts[17] );
xnor U1488 ( n1412, my_FIR_filter_firBlock_left_firStep[177], my_FIR_filter_firBlock_left_multProducts[17] );
xor U1489 ( my_FIR_filter_firBlock_left_N179, n1722, n1721 );
xor U1490 ( n1721, my_FIR_filter_firBlock_left_multProducts[48], my_FIR_filter_firBlock_left_firStep[114] );
xor U1491 ( my_FIR_filter_firBlock_left_N83, n1102, n1101 );
xor U1492 ( n1101, my_FIR_filter_firBlock_left_multProducts[48], my_FIR_filter_firBlock_left_firStep[210] );
xnor U1493 ( my_FIR_filter_firBlock_left_N210, n1868, n1869 );
xnor U1494 ( n1868, my_FIR_filter_firBlock_left_firStep[81], my_FIR_filter_firBlock_left_multProducts[48] );
xnor U1495 ( my_FIR_filter_firBlock_left_N50, n944, n945 );
xnor U1496 ( n944, my_FIR_filter_firBlock_left_firStep[241], my_FIR_filter_firBlock_left_multProducts[48] );
xor U1497 ( outData_in[14], n177, n176 );
xor U1498 ( n176, rightOut[14], leftOut[14] );
xor U1499 ( n628, my_FIR_filter_firBlock_left_multProducts[75], my_FIR_filter_firBlock_left_firStep[270] );
xor U1500 ( n2005, my_FIR_filter_firBlock_left_multProducts[75], my_FIR_filter_firBlock_left_firStep[46] );
xnor U1501 ( my_FIR_filter_firBlock_left_N276, n2182, n2185 );
xnor U1502 ( n2182, my_FIR_filter_firBlock_left_firStep[19], my_FIR_filter_firBlock_left_multProducts[109] );
xor U1503 ( my_FIR_filter_firBlock_left_N145, n1560, n1559 );
xor U1504 ( n1559, my_FIR_filter_firBlock_left_multProducts[16], my_FIR_filter_firBlock_left_firStep[144] );
xor U1505 ( my_FIR_filter_firBlock_left_N113, n1408, n1407 );
xor U1506 ( n1407, my_FIR_filter_firBlock_left_multProducts[16], my_FIR_filter_firBlock_left_firStep[176] );
xor U1507 ( my_FIR_filter_firBlock_left_N209, n1864, n1863 );
xor U1508 ( n1863, my_FIR_filter_firBlock_left_multProducts[47], my_FIR_filter_firBlock_left_firStep[80] );
xor U1509 ( my_FIR_filter_firBlock_left_N49, n940, n939 );
xor U1510 ( n939, my_FIR_filter_firBlock_left_multProducts[47], my_FIR_filter_firBlock_left_firStep[240] );
xnor U1511 ( outData_in[13], n171, n172 );
xnor U1512 ( n171, leftOut[13], rightOut[13] );
xnor U1513 ( my_FIR_filter_firBlock_left_N178, n1716, n1717 );
xnor U1514 ( n1716, my_FIR_filter_firBlock_left_firStep[113], my_FIR_filter_firBlock_left_multProducts[47] );
xnor U1515 ( my_FIR_filter_firBlock_left_N82, n1096, n1097 );
xnor U1516 ( n1096, my_FIR_filter_firBlock_left_firStep[209], my_FIR_filter_firBlock_left_multProducts[47] );
xnor U1517 ( n2000, my_FIR_filter_firBlock_left_firStep[45], my_FIR_filter_firBlock_left_multProducts[74] );
xnor U1518 ( n623, my_FIR_filter_firBlock_left_firStep[269], my_FIR_filter_firBlock_left_multProducts[74] );
xor U1519 ( my_FIR_filter_firBlock_left_N275, n2178, n2177 );
xor U1520 ( n2177, my_FIR_filter_firBlock_left_multProducts[108], my_FIR_filter_firBlock_left_firStep[18] );
xnor U1521 ( my_FIR_filter_firBlock_left_N112, n1402, n1403 );
xnor U1522 ( n1402, my_FIR_filter_firBlock_left_firStep[175], my_FIR_filter_firBlock_left_multProducts[15] );
xor U1523 ( outData_in[12], n167, n166 );
xor U1524 ( n166, rightOut[12], leftOut[12] );
xnor U1525 ( n1554, my_FIR_filter_firBlock_left_firStep[143], my_FIR_filter_firBlock_left_multProducts[15] );
xor U1526 ( my_FIR_filter_firBlock_left_N177, n1712, n1711 );
xor U1527 ( n1711, my_FIR_filter_firBlock_left_multProducts[46], my_FIR_filter_firBlock_left_firStep[112] );
xor U1528 ( my_FIR_filter_firBlock_left_N81, n1092, n1091 );
xor U1529 ( n1091, my_FIR_filter_firBlock_left_multProducts[46], my_FIR_filter_firBlock_left_firStep[208] );
xnor U1530 ( my_FIR_filter_firBlock_left_N208, n1858, n1859 );
xnor U1531 ( n1858, my_FIR_filter_firBlock_left_firStep[79], my_FIR_filter_firBlock_left_multProducts[46] );
xnor U1532 ( my_FIR_filter_firBlock_left_N48, n934, n935 );
xnor U1533 ( n934, my_FIR_filter_firBlock_left_firStep[239], my_FIR_filter_firBlock_left_multProducts[46] );
xor U1534 ( my_FIR_filter_firBlock_left_N13, n619, n618 );
xor U1535 ( n618, my_FIR_filter_firBlock_left_multProducts[73], my_FIR_filter_firBlock_left_firStep[268] );
xor U1536 ( n1995, my_FIR_filter_firBlock_left_multProducts[73], my_FIR_filter_firBlock_left_firStep[44] );
xor U1537 ( my_FIR_filter_firBlock_left_N143, n1550, n1549 );
xor U1538 ( n1549, my_FIR_filter_firBlock_left_multProducts[14], my_FIR_filter_firBlock_left_firStep[142] );
xnor U1539 ( outData_in[11], n161, n162 );
xnor U1540 ( n161, leftOut[11], rightOut[11] );
xor U1541 ( n1397, my_FIR_filter_firBlock_left_multProducts[14], my_FIR_filter_firBlock_left_firStep[174] );
xnor U1542 ( my_FIR_filter_firBlock_left_N274, n2172, n2173 );
xnor U1543 ( n2172, my_FIR_filter_firBlock_left_firStep[17], my_FIR_filter_firBlock_left_multProducts[107] );
xnor U1544 ( n1990, my_FIR_filter_firBlock_left_firStep[43], my_FIR_filter_firBlock_left_multProducts[72] );
xnor U1545 ( n613, my_FIR_filter_firBlock_left_firStep[267], my_FIR_filter_firBlock_left_multProducts[72] );
xor U1546 ( my_FIR_filter_firBlock_left_N207, n1854, n1853 );
xor U1547 ( n1853, my_FIR_filter_firBlock_left_multProducts[45], my_FIR_filter_firBlock_left_firStep[78] );
xor U1548 ( my_FIR_filter_firBlock_left_N47, n930, n929 );
xor U1549 ( n929, my_FIR_filter_firBlock_left_multProducts[45], my_FIR_filter_firBlock_left_firStep[238] );
xnor U1550 ( my_FIR_filter_firBlock_left_N176, n1706, n1707 );
xnor U1551 ( n1706, my_FIR_filter_firBlock_left_firStep[111], my_FIR_filter_firBlock_left_multProducts[45] );
xnor U1552 ( my_FIR_filter_firBlock_left_N80, n1086, n1087 );
xnor U1553 ( n1086, my_FIR_filter_firBlock_left_firStep[207], my_FIR_filter_firBlock_left_multProducts[45] );
xor U1554 ( outData_in[10], n157, n156 );
xor U1555 ( n156, rightOut[10], leftOut[10] );
xnor U1556 ( n1544, my_FIR_filter_firBlock_left_firStep[141], my_FIR_filter_firBlock_left_multProducts[13] );
xnor U1557 ( n1392, my_FIR_filter_firBlock_left_firStep[173], my_FIR_filter_firBlock_left_multProducts[13] );
xor U1558 ( my_FIR_filter_firBlock_left_N273, n2168, n2167 );
xor U1559 ( n2167, my_FIR_filter_firBlock_left_multProducts[106], my_FIR_filter_firBlock_left_firStep[16] );
xor U1560 ( my_FIR_filter_firBlock_left_N79, n1082, n1081 );
xor U1561 ( n1081, my_FIR_filter_firBlock_left_multProducts[44], my_FIR_filter_firBlock_left_firStep[206] );
xor U1562 ( my_FIR_filter_firBlock_left_N175, n1702, n1701 );
xor U1563 ( n1701, my_FIR_filter_firBlock_left_multProducts[44], my_FIR_filter_firBlock_left_firStep[110] );
xor U1564 ( my_FIR_filter_firBlock_left_N235, n1986, n1985 );
xor U1565 ( n1985, my_FIR_filter_firBlock_left_multProducts[71], my_FIR_filter_firBlock_left_firStep[42] );
xnor U1566 ( my_FIR_filter_firBlock_left_N206, n1848, n1849 );
xnor U1567 ( n1848, my_FIR_filter_firBlock_left_firStep[77], my_FIR_filter_firBlock_left_multProducts[44] );
xnor U1568 ( my_FIR_filter_firBlock_left_N46, n924, n925 );
xnor U1569 ( n924, my_FIR_filter_firBlock_left_firStep[237], my_FIR_filter_firBlock_left_multProducts[44] );
xor U1570 ( n608, my_FIR_filter_firBlock_left_multProducts[71], my_FIR_filter_firBlock_left_firStep[266] );
xnor U1571 ( outData_in[9], n280, n279 );
xnor U1572 ( n280, leftOut[9], rightOut[9] );
xor U1573 ( my_FIR_filter_firBlock_left_N109, n1388, n1387 );
xor U1574 ( n1387, my_FIR_filter_firBlock_left_multProducts[12], my_FIR_filter_firBlock_left_firStep[172] );
xor U1575 ( n1539, my_FIR_filter_firBlock_left_multProducts[12], my_FIR_filter_firBlock_left_firStep[140] );
xor U1576 ( outData_in[8], n278, n277 );
xor U1577 ( n277, rightOut[8], leftOut[8] );
xnor U1578 ( my_FIR_filter_firBlock_left_N272, n2162, n2163 );
xnor U1579 ( n2162, my_FIR_filter_firBlock_left_firStep[15], my_FIR_filter_firBlock_left_multProducts[105] );
xnor U1580 ( my_FIR_filter_firBlock_left_N10, n732, n731 );
xnor U1581 ( n732, my_FIR_filter_firBlock_left_firStep[265], my_FIR_filter_firBlock_left_multProducts[70] );
xnor U1582 ( n2109, my_FIR_filter_firBlock_left_firStep[41], my_FIR_filter_firBlock_left_multProducts[70] );
xor U1583 ( my_FIR_filter_firBlock_left_N205, n1844, n1843 );
xor U1584 ( n1843, my_FIR_filter_firBlock_left_multProducts[43], my_FIR_filter_firBlock_left_firStep[76] );
xor U1585 ( my_FIR_filter_firBlock_left_N45, n920, n919 );
xor U1586 ( n919, my_FIR_filter_firBlock_left_multProducts[43], my_FIR_filter_firBlock_left_firStep[236] );
xnor U1587 ( my_FIR_filter_firBlock_left_N174, n1696, n1697 );
xnor U1588 ( n1696, my_FIR_filter_firBlock_left_firStep[109], my_FIR_filter_firBlock_left_multProducts[43] );
xnor U1589 ( my_FIR_filter_firBlock_left_N78, n1076, n1077 );
xnor U1590 ( n1076, my_FIR_filter_firBlock_left_firStep[205], my_FIR_filter_firBlock_left_multProducts[43] );
xnor U1591 ( n1534, my_FIR_filter_firBlock_left_firStep[139], my_FIR_filter_firBlock_left_multProducts[11] );
xnor U1592 ( n1382, my_FIR_filter_firBlock_left_firStep[171], my_FIR_filter_firBlock_left_multProducts[11] );
xnor U1593 ( outData_in[7], n276, n275 );
xnor U1594 ( n276, leftOut[7], rightOut[7] );
xor U1595 ( my_FIR_filter_firBlock_left_N271, n2158, n2157 );
xor U1596 ( n2157, my_FIR_filter_firBlock_left_multProducts[104], my_FIR_filter_firBlock_left_firStep[14] );
xor U1597 ( my_FIR_filter_firBlock_left_N173, n1692, n1691 );
xor U1598 ( n1691, my_FIR_filter_firBlock_left_multProducts[42], my_FIR_filter_firBlock_left_firStep[108] );
xor U1599 ( my_FIR_filter_firBlock_left_N77, n1072, n1071 );
xor U1600 ( n1071, my_FIR_filter_firBlock_left_multProducts[42], my_FIR_filter_firBlock_left_firStep[204] );
xnor U1601 ( my_FIR_filter_firBlock_left_N204, n1838, n1839 );
xnor U1602 ( n1838, my_FIR_filter_firBlock_left_firStep[75], my_FIR_filter_firBlock_left_multProducts[42] );
xnor U1603 ( my_FIR_filter_firBlock_left_N44, n914, n915 );
xnor U1604 ( n914, my_FIR_filter_firBlock_left_firStep[235], my_FIR_filter_firBlock_left_multProducts[42] );
xor U1605 ( outData_in[6], n274, n273 );
xor U1606 ( n273, rightOut[6], leftOut[6] );
xor U1607 ( my_FIR_filter_firBlock_left_N107, n1378, n1377 );
xor U1608 ( n1377, my_FIR_filter_firBlock_left_multProducts[10], my_FIR_filter_firBlock_left_firStep[170] );
xor U1609 ( my_FIR_filter_firBlock_left_N139, n1530, n1529 );
xor U1610 ( n1529, my_FIR_filter_firBlock_left_multProducts[10], my_FIR_filter_firBlock_left_firStep[138] );
xnor U1611 ( my_FIR_filter_firBlock_left_N270, n2152, n2153 );
xnor U1612 ( n2152, my_FIR_filter_firBlock_left_firStep[13], my_FIR_filter_firBlock_left_multProducts[103] );
xor U1613 ( my_FIR_filter_firBlock_left_N203, n1834, n1833 );
xor U1614 ( n1833, my_FIR_filter_firBlock_left_multProducts[41], my_FIR_filter_firBlock_left_firStep[74] );
xor U1615 ( my_FIR_filter_firBlock_left_N43, n910, n909 );
xor U1616 ( n909, my_FIR_filter_firBlock_left_multProducts[41], my_FIR_filter_firBlock_left_firStep[234] );
xnor U1617 ( my_FIR_filter_firBlock_left_N172, n1686, n1687 );
xnor U1618 ( n1686, my_FIR_filter_firBlock_left_firStep[107], my_FIR_filter_firBlock_left_multProducts[41] );
xnor U1619 ( my_FIR_filter_firBlock_left_N76, n1066, n1067 );
xnor U1620 ( n1066, my_FIR_filter_firBlock_left_firStep[203], my_FIR_filter_firBlock_left_multProducts[41] );
xnor U1621 ( outData_in[5], n272, n271 );
xnor U1622 ( n272, leftOut[5], rightOut[5] );
xnor U1623 ( n1653, my_FIR_filter_firBlock_left_firStep[137], my_FIR_filter_firBlock_left_multProducts[9] );
xnor U1624 ( n1501, my_FIR_filter_firBlock_left_firStep[169], my_FIR_filter_firBlock_left_multProducts[9] );
xor U1625 ( outData_in[4], n270, n269 );
xor U1626 ( n269, rightOut[4], leftOut[4] );
xor U1627 ( my_FIR_filter_firBlock_left_N269, n2148, n2147 );
xor U1628 ( n2147, my_FIR_filter_firBlock_left_multProducts[102], my_FIR_filter_firBlock_left_firStep[12] );
xor U1629 ( my_FIR_filter_firBlock_left_N75, n1062, n1061 );
xor U1630 ( n1061, my_FIR_filter_firBlock_left_multProducts[40], my_FIR_filter_firBlock_left_firStep[202] );
xor U1631 ( my_FIR_filter_firBlock_left_N171, n1682, n1681 );
xor U1632 ( n1681, my_FIR_filter_firBlock_left_multProducts[40], my_FIR_filter_firBlock_left_firStep[106] );
xnor U1633 ( my_FIR_filter_firBlock_left_N202, n1957, n1956 );
xnor U1634 ( n1957, my_FIR_filter_firBlock_left_firStep[73], my_FIR_filter_firBlock_left_multProducts[40] );
xnor U1635 ( my_FIR_filter_firBlock_left_N42, n1033, n1032 );
xnor U1636 ( n1033, my_FIR_filter_firBlock_left_firStep[233], my_FIR_filter_firBlock_left_multProducts[40] );
xor U1637 ( my_FIR_filter_firBlock_left_N137, n1651, n1650 );
xor U1638 ( n1650, my_FIR_filter_firBlock_left_multProducts[8], my_FIR_filter_firBlock_left_firStep[136] );
xor U1639 ( n1498, my_FIR_filter_firBlock_left_multProducts[8], my_FIR_filter_firBlock_left_firStep[168] );
xnor U1640 ( my_FIR_filter_firBlock_left_N6, n724, n723 );
xnor U1641 ( outData_in[3], n268, n267 );
xnor U1642 ( n268, leftOut[3], rightOut[3] );
xnor U1643 ( my_FIR_filter_firBlock_left_N268, n2142, n2143 );
xnor U1644 ( n2142, my_FIR_filter_firBlock_left_firStep[11], my_FIR_filter_firBlock_left_multProducts[101] );
xor U1645 ( my_FIR_filter_firBlock_left_N201, n1955, n1954 );
xor U1646 ( n1954, my_FIR_filter_firBlock_left_multProducts[39], my_FIR_filter_firBlock_left_firStep[72] );
xor U1647 ( my_FIR_filter_firBlock_left_N41, n1031, n1030 );
xor U1648 ( n1030, my_FIR_filter_firBlock_left_multProducts[39], my_FIR_filter_firBlock_left_firStep[232] );
xnor U1649 ( my_FIR_filter_firBlock_left_N170, n1805, n1804 );
xnor U1650 ( n1805, my_FIR_filter_firBlock_left_firStep[105], my_FIR_filter_firBlock_left_multProducts[39] );
xnor U1651 ( my_FIR_filter_firBlock_left_N74, n1185, n1184 );
xnor U1652 ( n1185, my_FIR_filter_firBlock_left_firStep[201], my_FIR_filter_firBlock_left_multProducts[39] );
xnor U1653 ( n1649, my_FIR_filter_firBlock_left_firStep[135], my_FIR_filter_firBlock_left_multProducts[7] );
xnor U1654 ( n1497, my_FIR_filter_firBlock_left_firStep[167], my_FIR_filter_firBlock_left_multProducts[7] );
xor U1655 ( my_FIR_filter_firBlock_left_N229, n2099, n2098 );
xor U1656 ( outData_in[2], n255, n254 );
xor U1657 ( n254, rightOut[2], leftOut[2] );
xor U1658 ( my_FIR_filter_firBlock_left_N267, n2138, n2137 );
xor U1659 ( n2137, my_FIR_filter_firBlock_left_multProducts[100], my_FIR_filter_firBlock_left_firStep[10] );
xor U1660 ( outData_in[1], n203, n202 );
xor U1661 ( n202, rightOut[1], leftOut[1] );
xor U1662 ( my_FIR_filter_firBlock_left_N135, n1647, n1646 );
xor U1663 ( n1646, my_FIR_filter_firBlock_left_multProducts[6], my_FIR_filter_firBlock_left_firStep[134] );
xor U1664 ( my_FIR_filter_firBlock_left_N103, n1495, n1494 );
xor U1665 ( n1494, my_FIR_filter_firBlock_left_multProducts[6], my_FIR_filter_firBlock_left_firStep[166] );
xor U1666 ( my_FIR_filter_firBlock_left_N169, n1803, n1802 );
xor U1667 ( n1802, my_FIR_filter_firBlock_left_multProducts[38], my_FIR_filter_firBlock_left_firStep[104] );
xor U1668 ( my_FIR_filter_firBlock_left_N73, n1183, n1182 );
xor U1669 ( n1182, my_FIR_filter_firBlock_left_multProducts[38], my_FIR_filter_firBlock_left_firStep[200] );
xnor U1670 ( my_FIR_filter_firBlock_left_N200, n1953, n1952 );
xnor U1671 ( n1953, my_FIR_filter_firBlock_left_firStep[71], my_FIR_filter_firBlock_left_multProducts[38] );
xnor U1672 ( my_FIR_filter_firBlock_left_N40, n1029, n1028 );
xnor U1673 ( n1029, my_FIR_filter_firBlock_left_firStep[231], my_FIR_filter_firBlock_left_multProducts[38] );
xor U1674 ( my_FIR_filter_firBlock_right_multProducts[0], rightOut[0], leftOut[0] );
xor U1675 ( my_FIR_filter_firBlock_left_N227, n2084, n2083 );
xor U1676 ( n2083, my_FIR_filter_firBlock_left_multProducts[63], my_FIR_filter_firBlock_left_firStep[34] );
xor U1677 ( my_FIR_filter_firBlock_left_N3, n707, n706 );
xor U1678 ( n706, my_FIR_filter_firBlock_left_multProducts[63], my_FIR_filter_firBlock_left_firStep[258] );
xor U1679 ( my_FIR_filter_firBlock_left_N199, n1951, n1950 );
xor U1680 ( n1950, my_FIR_filter_firBlock_left_multProducts[37], my_FIR_filter_firBlock_left_firStep[70] );
xor U1681 ( my_FIR_filter_firBlock_left_N39, n1027, n1026 );
xor U1682 ( n1026, my_FIR_filter_firBlock_left_multProducts[37], my_FIR_filter_firBlock_left_firStep[230] );
xnor U1683 ( my_FIR_filter_firBlock_left_N266, n2261, n2260 );
xnor U1684 ( n2261, my_FIR_filter_firBlock_left_firStep[9], my_FIR_filter_firBlock_left_multProducts[99] );
xnor U1685 ( my_FIR_filter_firBlock_left_N102, n1493, n1492 );
xnor U1686 ( n1493, my_FIR_filter_firBlock_left_firStep[165], my_FIR_filter_firBlock_left_multProducts[5] );
xnor U1687 ( my_FIR_filter_firBlock_left_N168, n1801, n1800 );
xnor U1688 ( n1801, my_FIR_filter_firBlock_left_firStep[103], my_FIR_filter_firBlock_left_multProducts[37] );
xnor U1689 ( my_FIR_filter_firBlock_left_N72, n1181, n1180 );
xnor U1690 ( n1181, my_FIR_filter_firBlock_left_firStep[199], my_FIR_filter_firBlock_left_multProducts[37] );
xnor U1691 ( n1645, my_FIR_filter_firBlock_left_firStep[133], my_FIR_filter_firBlock_left_multProducts[5] );
xor U1692 ( my_FIR_filter_firBlock_left_N101, n1491, n1490 );
xor U1693 ( n1490, my_FIR_filter_firBlock_left_multProducts[4], my_FIR_filter_firBlock_left_firStep[164] );
xor U1694 ( my_FIR_filter_firBlock_left_N167, n1799, n1798 );
xor U1695 ( n1798, my_FIR_filter_firBlock_left_multProducts[36], my_FIR_filter_firBlock_left_firStep[102] );
xor U1696 ( my_FIR_filter_firBlock_left_N71, n1179, n1178 );
xor U1697 ( n1178, my_FIR_filter_firBlock_left_multProducts[36], my_FIR_filter_firBlock_left_firStep[198] );
xor U1698 ( n1642, my_FIR_filter_firBlock_left_multProducts[4], my_FIR_filter_firBlock_left_firStep[132] );
xor U1699 ( my_FIR_filter_firBlock_left_N2, n655, n654 );
xor U1700 ( my_FIR_filter_firBlock_left_N265, n2259, n2258 );
xor U1701 ( n2258, my_FIR_filter_firBlock_left_multProducts[98], my_FIR_filter_firBlock_left_firStep[8] );
xnor U1702 ( my_FIR_filter_firBlock_left_N198, n1949, n1948 );
xnor U1703 ( n1949, my_FIR_filter_firBlock_left_firStep[69], my_FIR_filter_firBlock_left_multProducts[36] );
xnor U1704 ( my_FIR_filter_firBlock_left_N38, n1025, n1024 );
xnor U1705 ( n1025, my_FIR_filter_firBlock_left_firStep[229], my_FIR_filter_firBlock_left_multProducts[36] );
xnor U1706 ( n1641, my_FIR_filter_firBlock_left_firStep[131], my_FIR_filter_firBlock_left_multProducts[3] );
xnor U1707 ( n1489, my_FIR_filter_firBlock_left_firStep[163], my_FIR_filter_firBlock_left_multProducts[3] );
xor U1708 ( my_FIR_filter_firBlock_left_N197, n1947, n1946 );
xor U1709 ( n1946, my_FIR_filter_firBlock_left_multProducts[35], my_FIR_filter_firBlock_left_firStep[68] );
xor U1710 ( my_FIR_filter_firBlock_left_N37, n1023, n1022 );
xor U1711 ( n1022, my_FIR_filter_firBlock_left_multProducts[35], my_FIR_filter_firBlock_left_firStep[228] );
xnor U1712 ( my_FIR_filter_firBlock_left_N264, n2257, n2256 );
xnor U1713 ( n2257, my_FIR_filter_firBlock_left_firStep[7], my_FIR_filter_firBlock_left_multProducts[97] );
xnor U1714 ( my_FIR_filter_firBlock_left_N166, n1797, n1796 );
xnor U1715 ( n1797, my_FIR_filter_firBlock_left_firStep[101], my_FIR_filter_firBlock_left_multProducts[35] );
xnor U1716 ( my_FIR_filter_firBlock_left_N70, n1177, n1176 );
xnor U1717 ( n1177, my_FIR_filter_firBlock_left_firStep[197], my_FIR_filter_firBlock_left_multProducts[35] );
xor U1718 ( my_FIR_filter_firBlock_left_N131, n1628, n1627 );
xor U1719 ( my_FIR_filter_firBlock_left_N99, n1476, n1475 );
xor U1720 ( my_FIR_filter_firBlock_left_N165, n1795, n1794 );
xor U1721 ( n1794, my_FIR_filter_firBlock_left_multProducts[34], my_FIR_filter_firBlock_left_firStep[100] );
xor U1722 ( my_FIR_filter_firBlock_left_N69, n1175, n1174 );
xor U1723 ( n1174, my_FIR_filter_firBlock_left_multProducts[34], my_FIR_filter_firBlock_left_firStep[196] );
xnor U1724 ( my_FIR_filter_firBlock_left_N196, n1945, n1944 );
xnor U1725 ( n1945, my_FIR_filter_firBlock_left_firStep[67], my_FIR_filter_firBlock_left_multProducts[34] );
xnor U1726 ( my_FIR_filter_firBlock_left_N36, n1021, n1020 );
xnor U1727 ( n1021, my_FIR_filter_firBlock_left_firStep[227], my_FIR_filter_firBlock_left_multProducts[34] );
xor U1728 ( my_FIR_filter_firBlock_left_N263, n2255, n2254 );
xor U1729 ( n2254, my_FIR_filter_firBlock_left_multProducts[96], my_FIR_filter_firBlock_left_firStep[6] );
xor U1730 ( my_FIR_filter_firBlock_left_N195, n1932, n1931 );
xor U1731 ( n1931, my_FIR_filter_firBlock_left_multProducts[33], my_FIR_filter_firBlock_left_firStep[66] );
xor U1732 ( my_FIR_filter_firBlock_left_N35, n1008, n1007 );
xor U1733 ( n1007, my_FIR_filter_firBlock_left_multProducts[33], my_FIR_filter_firBlock_left_firStep[226] );
xor U1734 ( my_FIR_filter_firBlock_left_N130, n1576, n1575 );
xor U1735 ( my_FIR_filter_firBlock_left_N98, n1424, n1423 );
xnor U1736 ( my_FIR_filter_firBlock_left_N164, n1793, n1792 );
xnor U1737 ( n1793, my_FIR_filter_firBlock_left_firStep[99], my_FIR_filter_firBlock_left_multProducts[33] );
xnor U1738 ( my_FIR_filter_firBlock_left_N68, n1173, n1172 );
xnor U1739 ( n1173, my_FIR_filter_firBlock_left_firStep[195], my_FIR_filter_firBlock_left_multProducts[33] );
xnor U1740 ( my_FIR_filter_firBlock_left_N262, n2253, n2252 );
xnor U1741 ( n2253, my_FIR_filter_firBlock_left_firStep[5], my_FIR_filter_firBlock_left_multProducts[95] );
xor U1742 ( my_FIR_filter_firBlock_left_N194, n1880, n1879 );
xor U1743 ( n1879, my_FIR_filter_firBlock_left_multProducts[32], my_FIR_filter_firBlock_left_firStep[65] );
xor U1744 ( my_FIR_filter_firBlock_left_N163, n1780, n1779 );
xor U1745 ( n1779, my_FIR_filter_firBlock_left_multProducts[32], my_FIR_filter_firBlock_left_firStep[98] );
xor U1746 ( my_FIR_filter_firBlock_left_N67, n1160, n1159 );
xor U1747 ( n1159, my_FIR_filter_firBlock_left_multProducts[32], my_FIR_filter_firBlock_left_firStep[194] );
xor U1748 ( my_FIR_filter_firBlock_left_N34, n956, n955 );
xor U1749 ( n955, my_FIR_filter_firBlock_left_multProducts[32], my_FIR_filter_firBlock_left_firStep[225] );
xor U1750 ( my_FIR_filter_firBlock_left_N261, n2251, n2250 );
xor U1751 ( n2250, my_FIR_filter_firBlock_left_multProducts[94], my_FIR_filter_firBlock_left_firStep[4] );
xor U1752 ( my_FIR_filter_firBlock_left_N129, my_FIR_filter_firBlock_left_multProducts[0], my_FIR_filter_firBlock_left_firStep[128] );
xor U1753 ( my_FIR_filter_firBlock_left_N97, my_FIR_filter_firBlock_left_multProducts[0], my_FIR_filter_firBlock_left_firStep[160] );
xor U1754 ( my_FIR_filter_firBlock_left_N162, n1728, n1727 );
xor U1755 ( n1727, my_FIR_filter_firBlock_left_multProducts[31], my_FIR_filter_firBlock_left_firStep[97] );
xor U1756 ( my_FIR_filter_firBlock_left_N66, n1108, n1107 );
xor U1757 ( n1107, my_FIR_filter_firBlock_left_multProducts[31], my_FIR_filter_firBlock_left_firStep[193] );
xnor U1758 ( my_FIR_filter_firBlock_left_N260, n2249, n2248 );
xnor U1759 ( n2249, my_FIR_filter_firBlock_left_firStep[3], my_FIR_filter_firBlock_left_multProducts[93] );
xor U1760 ( my_FIR_filter_firBlock_left_N193, my_FIR_filter_firBlock_left_multProducts[31], my_FIR_filter_firBlock_left_firStep[64] );
xor U1761 ( my_FIR_filter_firBlock_left_N33, my_FIR_filter_firBlock_left_multProducts[31], my_FIR_filter_firBlock_left_firStep[224] );
xor U1762 ( my_FIR_filter_firBlock_left_N259, n2236, n2235 );
xor U1763 ( n2235, my_FIR_filter_firBlock_left_multProducts[92], my_FIR_filter_firBlock_left_firStep[2] );
xor U1764 ( my_FIR_filter_firBlock_left_N161, my_FIR_filter_firBlock_left_multProducts[30], my_FIR_filter_firBlock_left_firStep[96] );
xor U1765 ( my_FIR_filter_firBlock_left_N65, my_FIR_filter_firBlock_left_multProducts[30], my_FIR_filter_firBlock_left_firStep[192] );
xor U1766 ( my_FIR_filter_firBlock_left_N258, n2184, n2183 );
xor U1767 ( n2183, my_FIR_filter_firBlock_left_multProducts[91], my_FIR_filter_firBlock_left_firStep[1] );
buf U1768 ( n118, reset );
xor U1769 ( n729, my_FIR_filter_firBlock_left_multProducts[69], my_FIR_filter_firBlock_left_firStep[264] );
xor U1770 ( n2106, my_FIR_filter_firBlock_left_multProducts[69], my_FIR_filter_firBlock_left_firStep[40] );
xor U1771 ( n1259, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[21], n39 );
nand U1772 ( n603, my_FIR_filter_firBlock_left_multProducts[69], n602 );
xor U1773 ( n477, my_FIR_filter_firBlock_left_multProducts[96], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[21] );
xor U1774 ( my_FIR_filter_firBlock_left_N128, n1487, n1486 );
nand U1775 ( n1323, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[33], n1320 );
or U1776 ( n1321, n1320, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[33] );
nand U1777 ( n1308, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[30], n1305 );
xor U1778 ( my_FIR_filter_firBlock_left_multProducts[22], n1305, n1304 );
or U1779 ( n1306, n1305, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[30] );
nand U1780 ( n1305, n1303, n1302 );
xor U1781 ( my_FIR_filter_firBlock_left_multProducts[21], n1300, n1299 );
nand U1782 ( n1303, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[29], n1300 );
or U1783 ( n1301, n1300, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[29] );
xor U1784 ( my_FIR_filter_firBlock_left_multProducts[17], n1280, n1279 );
nand U1785 ( n1283, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[25], n1280 );
or U1786 ( n1281, n1280, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[25] );
xor U1787 ( my_FIR_filter_firBlock_left_multProducts[15], n1270, n1269 );
nand U1788 ( n1273, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[23], n1270 );
or U1789 ( n1271, n1270, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[23] );
xor U1790 ( my_FIR_filter_firBlock_left_multProducts[9], n1240, n1239 );
xor U1791 ( my_FIR_filter_firBlock_left_multProducts[6], n1225, n1224 );
nand U1792 ( n1213, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[11], n1210 );
or U1793 ( n1211, n1210, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[11] );
nand U1794 ( n1200, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[8], n1347 );
or U1795 ( n1198, n1347, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[8] );
nand U1796 ( n488, n486, n485 );
nand U1797 ( n485, my_FIR_filter_firBlock_left_multProducts[97], n484 );
nand U1798 ( n490, my_FIR_filter_firBlock_left_multProducts[98], n489 );
nand U1799 ( n560, my_FIR_filter_firBlock_left_multProducts[112], n559 );
nand U1800 ( n540, my_FIR_filter_firBlock_left_multProducts[108], n539 );
xnor U1801 ( my_FIR_filter_firBlock_left_N26, n685, n686 );
nand U1802 ( n689, my_FIR_filter_firBlock_left_firStep[281], n686 );
nand U1803 ( n727, n598, n597 );
nand U1804 ( n722, n589, n588 );
xor U1805 ( my_FIR_filter_firBlock_left_N245, n2038, n2037 );
xnor U1806 ( n2030, my_FIR_filter_firBlock_left_firStep[51], my_FIR_filter_firBlock_left_multProducts[80] );
xnor U1807 ( n653, my_FIR_filter_firBlock_left_firStep[275], my_FIR_filter_firBlock_left_multProducts[80] );
nand U1808 ( n2041, my_FIR_filter_firBlock_left_firStep[52], n2038 );
nand U1809 ( n2035, my_FIR_filter_firBlock_left_multProducts[80], n2034 );
nand U1810 ( n376, n375, n42 );
xor U1811 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[29], n369, n368 );
nand U1812 ( n351, n350, n37 );
nand U1813 ( n321, n320, n31 );
nand U1814 ( n422, n287, n286 );
nand U1815 ( n455, my_FIR_filter_firBlock_left_multProducts[91], n454 );
nand U1816 ( n636, my_FIR_filter_firBlock_left_multProducts[76], n635 );
nand U1817 ( n508, n506, n505 );
xor U1818 ( n2102, my_FIR_filter_firBlock_left_multProducts[67], my_FIR_filter_firBlock_left_firStep[38] );
xor U1819 ( n725, my_FIR_filter_firBlock_left_multProducts[67], my_FIR_filter_firBlock_left_firStep[262] );
nand U1820 ( n686, n684, n683 );
xor U1821 ( n1249, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[19], n37 );
nand U1822 ( n1974, my_FIR_filter_firBlock_left_multProducts[67], n1973 );
nand U1823 ( n597, my_FIR_filter_firBlock_left_multProducts[67], n596 );
nand U1824 ( n471, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[19], n468 );
xor U1825 ( n467, my_FIR_filter_firBlock_left_multProducts[94], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[19] );
nand U1826 ( n1141, my_FIR_filter_firBlock_left_multProducts[55], n1140 );
or U1827 ( n1140, n1139, my_FIR_filter_firBlock_left_firStep[217] );
nand U1828 ( n1146, my_FIR_filter_firBlock_left_multProducts[56], n1145 );
or U1829 ( n1145, n1144, my_FIR_filter_firBlock_left_firStep[218] );
nand U1830 ( n1094, my_FIR_filter_firBlock_left_multProducts[46], n1093 );
or U1831 ( n1093, n1092, my_FIR_filter_firBlock_left_firStep[208] );
nand U1832 ( n1056, my_FIR_filter_firBlock_left_multProducts[38], n1055 );
or U1833 ( n1055, n1183, my_FIR_filter_firBlock_left_firStep[200] );
nand U1834 ( n1050, my_FIR_filter_firBlock_left_multProducts[36], n1049 );
or U1835 ( n1049, n1179, my_FIR_filter_firBlock_left_firStep[198] );
nand U1836 ( n1163, my_FIR_filter_firBlock_left_multProducts[59], n1162 );
or U1837 ( n1162, n1161, my_FIR_filter_firBlock_left_firStep[221] );
nand U1838 ( n1121, my_FIR_filter_firBlock_left_multProducts[51], n1120 );
or U1839 ( n1120, n1119, my_FIR_filter_firBlock_left_firStep[213] );
nand U1840 ( n1131, my_FIR_filter_firBlock_left_multProducts[53], n1130 );
or U1841 ( n1130, n1129, my_FIR_filter_firBlock_left_firStep[215] );
nand U1842 ( n1069, my_FIR_filter_firBlock_left_multProducts[41], n1068 );
or U1843 ( n1068, n1067, my_FIR_filter_firBlock_left_firStep[203] );
nand U1844 ( n1111, my_FIR_filter_firBlock_left_multProducts[49], n1110 );
or U1845 ( n1110, n1109, my_FIR_filter_firBlock_left_firStep[211] );
nand U1846 ( n1089, my_FIR_filter_firBlock_left_multProducts[45], n1088 );
or U1847 ( n1088, n1087, my_FIR_filter_firBlock_left_firStep[207] );
nand U1848 ( n1079, my_FIR_filter_firBlock_left_multProducts[43], n1078 );
or U1849 ( n1078, n1077, my_FIR_filter_firBlock_left_firStep[205] );
nand U1850 ( n1059, my_FIR_filter_firBlock_left_multProducts[39], n1058 );
or U1851 ( n1058, n1184, my_FIR_filter_firBlock_left_firStep[201] );
nand U1852 ( n1047, my_FIR_filter_firBlock_left_multProducts[35], n1046 );
or U1853 ( n1046, n1176, my_FIR_filter_firBlock_left_firStep[197] );
nand U1854 ( n1104, my_FIR_filter_firBlock_left_multProducts[48], n1103 );
or U1855 ( n1103, n1102, my_FIR_filter_firBlock_left_firStep[210] );
nand U1856 ( n1167, n1164, n1163 );
xor U1857 ( my_FIR_filter_firBlock_left_multProducts[30], n873, n872 );
xor U1858 ( my_FIR_filter_firBlock_left_N192, n1791, n1790 );
nor U1859 ( n1790, n1789, n1788 );
nand U1860 ( n1722, n1720, n1719 );
nand U1861 ( n1719, my_FIR_filter_firBlock_left_multProducts[47], n1718 );
nand U1862 ( n1739, n1737, n1736 );
nand U1863 ( n1736, my_FIR_filter_firBlock_left_multProducts[50], n1735 );
nand U1864 ( n1761, my_FIR_filter_firBlock_left_multProducts[55], n1760 );
or U1865 ( n1760, n1759, my_FIR_filter_firBlock_left_firStep[121] );
nand U1866 ( n1771, my_FIR_filter_firBlock_left_multProducts[57], n1770 );
or U1867 ( n1770, n1769, my_FIR_filter_firBlock_left_firStep[123] );
or U1868 ( n1718, n1717, my_FIR_filter_firBlock_left_firStep[113] );
nand U1869 ( n1673, my_FIR_filter_firBlock_left_multProducts[37], n1672 );
or U1870 ( n1672, n1800, my_FIR_filter_firBlock_left_firStep[103] );
nand U1871 ( n1756, my_FIR_filter_firBlock_left_multProducts[54], n1755 );
or U1872 ( n1755, n1754, my_FIR_filter_firBlock_left_firStep[120] );
or U1873 ( n1735, n1734, my_FIR_filter_firBlock_left_firStep[116] );
nand U1874 ( n1704, my_FIR_filter_firBlock_left_multProducts[44], n1703 );
or U1875 ( n1703, n1702, my_FIR_filter_firBlock_left_firStep[110] );
nand U1876 ( n1676, my_FIR_filter_firBlock_left_multProducts[38], n1675 );
or U1877 ( n1675, n1803, my_FIR_filter_firBlock_left_firStep[104] );
nand U1878 ( n1684, my_FIR_filter_firBlock_left_multProducts[40], n1683 );
or U1879 ( n1683, n1682, my_FIR_filter_firBlock_left_firStep[106] );
nand U1880 ( n1664, my_FIR_filter_firBlock_left_multProducts[34], n1663 );
or U1881 ( n1663, n1795, my_FIR_filter_firBlock_left_firStep[100] );
nand U1882 ( n1667, my_FIR_filter_firBlock_left_multProducts[35], n1666 );
or U1883 ( n1666, n1796, my_FIR_filter_firBlock_left_firStep[101] );
nand U1884 ( n1661, my_FIR_filter_firBlock_left_multProducts[33], n1660 );
or U1885 ( n1660, n1792, my_FIR_filter_firBlock_left_firStep[99] );
nand U1886 ( n1783, my_FIR_filter_firBlock_left_multProducts[59], n1782 );
nand U1887 ( n804, n802, n801 );
nand U1888 ( n839, n837, n836 );
or U1889 ( n770, n769, my_FIR_filter_firBlock_left_multProducts[94] );
or U1890 ( n810, n809, my_FIR_filter_firBlock_left_multProducts[102] );
or U1891 ( n760, n759, my_FIR_filter_firBlock_left_multProducts[92] );
or U1892 ( n840, n839, my_FIR_filter_firBlock_left_multProducts[108] );
or U1893 ( n855, n854, my_FIR_filter_firBlock_left_multProducts[111] );
or U1894 ( n825, n824, my_FIR_filter_firBlock_left_multProducts[105] );
or U1895 ( n775, n774, my_FIR_filter_firBlock_left_multProducts[95] );
nor U1896 ( n1014, my_FIR_filter_firBlock_left_firStep[254], n1015 );
nand U1897 ( n354, n352, n351 );
nand U1898 ( n369, n367, n366 );
nand U1899 ( n344, n342, n341 );
nand U1900 ( n295, n294, n25 );
xor U1901 ( my_FIR_filter_firBlock_left_multProducts[85], n558, n557 );
xor U1902 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[37], n411, n410 );
xnor U1903 ( n728, my_FIR_filter_firBlock_left_firStep[263], my_FIR_filter_firBlock_left_multProducts[68] );
xnor U1904 ( n2105, my_FIR_filter_firBlock_left_firStep[39], my_FIR_filter_firBlock_left_multProducts[68] );
nand U1905 ( n681, n679, n678 );
nand U1906 ( n639, n637, n636 );
nand U1907 ( n1258, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[20], n1255 );
or U1908 ( n1256, n1255, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[20] );
xor U1909 ( n1254, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[20], n38 );
xor U1910 ( n472, my_FIR_filter_firBlock_left_multProducts[95], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[20] );
xor U1911 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[16], n304, n303 );
nand U1912 ( n1535, n1533, n1532 );
nand U1913 ( n1532, my_FIR_filter_firBlock_left_multProducts[10], n1531 );
xor U1914 ( my_FIR_filter_firBlock_left_N160, n1639, n1638 );
nor U1915 ( n1638, n1637, n1636 );
nand U1916 ( n1622, n1620, n1619 );
nand U1917 ( n1619, my_FIR_filter_firBlock_left_multProducts[27], n1618 );
nand U1918 ( n1570, n1568, n1567 );
nand U1919 ( n1567, my_FIR_filter_firBlock_left_multProducts[17], n1566 );
nand U1920 ( n1604, my_FIR_filter_firBlock_left_multProducts[24], n1603 );
or U1921 ( n1603, n1602, my_FIR_filter_firBlock_left_firStep[152] );
nand U1922 ( n1584, my_FIR_filter_firBlock_left_multProducts[20], n1583 );
or U1923 ( n1583, n1582, my_FIR_filter_firBlock_left_firStep[148] );
nand U1924 ( n1562, my_FIR_filter_firBlock_left_multProducts[16], n1561 );
or U1925 ( n1561, n1560, my_FIR_filter_firBlock_left_firStep[144] );
nand U1926 ( n1599, my_FIR_filter_firBlock_left_multProducts[23], n1598 );
nand U1927 ( n1579, my_FIR_filter_firBlock_left_multProducts[19], n1578 );
nand U1928 ( n1515, my_FIR_filter_firBlock_left_multProducts[5], n1514 );
nand U1929 ( n1521, my_FIR_filter_firBlock_left_multProducts[7], n1520 );
nand U1930 ( n1614, my_FIR_filter_firBlock_left_multProducts[26], n1613 );
or U1931 ( n1613, n1612, my_FIR_filter_firBlock_left_firStep[154] );
nand U1932 ( n1552, my_FIR_filter_firBlock_left_multProducts[14], n1551 );
or U1933 ( n1551, n1550, my_FIR_filter_firBlock_left_firStep[142] );
or U1934 ( n1531, n1530, my_FIR_filter_firBlock_left_firStep[138] );
nand U1935 ( n1512, my_FIR_filter_firBlock_left_multProducts[4], n1511 );
nand U1936 ( n1509, my_FIR_filter_firBlock_left_multProducts[3], n1508 );
nor U1937 ( n1634, my_FIR_filter_firBlock_left_firStep[158], n1635 );
nand U1938 ( n1349, n1200, n1199 );
xnor U1939 ( n695, my_FIR_filter_firBlock_left_firStep[283], my_FIR_filter_firBlock_left_multProducts[88] );
xnor U1940 ( n2072, my_FIR_filter_firBlock_left_firStep[59], my_FIR_filter_firBlock_left_multProducts[88] );
xnor U1941 ( n705, my_FIR_filter_firBlock_left_firStep[285], my_FIR_filter_firBlock_left_multProducts[89] );
xnor U1942 ( n2082, my_FIR_filter_firBlock_left_firStep[61], my_FIR_filter_firBlock_left_multProducts[89] );
xnor U1943 ( n718, my_FIR_filter_firBlock_left_multProducts[89], my_FIR_filter_firBlock_left_firStep[287] );
xnor U1944 ( n2095, my_FIR_filter_firBlock_left_multProducts[89], my_FIR_filter_firBlock_left_firStep[63] );
not U1945 ( n120, my_FIR_filter_firBlock_left_multProducts[89] );
nand U1946 ( n2087, my_FIR_filter_firBlock_left_multProducts[89], n2086 );
nand U1947 ( n703, my_FIR_filter_firBlock_left_multProducts[89], n702 );
nand U1948 ( n2080, my_FIR_filter_firBlock_left_multProducts[89], n2079 );
nand U1949 ( n698, my_FIR_filter_firBlock_left_multProducts[88], n697 );
nand U1950 ( n574, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, my_FIR_filter_firBlock_left_multProducts[88] );
or U1951 ( n572, my_FIR_filter_firBlock_left_multProducts[88], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
nand U1952 ( n571, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n568 );
or U1953 ( n569, n568, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
nand U1954 ( n543, n541, n540 );
nand U1955 ( n528, n526, n525 );
nand U1956 ( n496, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[24], n493 );
xor U1957 ( my_FIR_filter_firBlock_left_multProducts[72], n493, n492 );
xor U1958 ( my_FIR_filter_firBlock_left_multProducts[62], n578, n577 );
xnor U1959 ( my_FIR_filter_firBlock_left_N232, n2105, n2104 );
xor U1960 ( my_FIR_filter_firBlock_left_N231, n2103, n2102 );
xor U1961 ( my_FIR_filter_firBlock_left_N233, n2107, n2106 );
nand U1962 ( n2073, n2071, n2070 );
nand U1963 ( n2053, n2051, n2050 );
nand U1964 ( n2043, n2041, n2040 );
nand U1965 ( n2038, n2036, n2035 );
nand U1966 ( n2016, n2014, n2013 );
nand U1967 ( n2011, n2009, n2008 );
nand U1968 ( n1986, n1984, n1983 );
nand U1969 ( n1981, my_FIR_filter_firBlock_left_firStep[40], n2107 );
nand U1970 ( n1978, my_FIR_filter_firBlock_left_firStep[39], n2104 );
nand U1971 ( n1975, my_FIR_filter_firBlock_left_firStep[38], n2103 );
or U1972 ( n1973, n2103, my_FIR_filter_firBlock_left_firStep[38] );
nand U1973 ( n2099, n1966, n1965 );
nand U1974 ( n1210, n1208, n1207 );
nand U1975 ( n1207, n1206, n28 );
nand U1976 ( n1477, n1473, n1472 );
nand U1977 ( n1472, my_FIR_filter_firBlock_left_multProducts[28], n1471 );
nand U1978 ( n1452, my_FIR_filter_firBlock_left_multProducts[24], n1451 );
nand U1979 ( n1432, my_FIR_filter_firBlock_left_multProducts[20], n1431 );
or U1980 ( n1431, n1430, my_FIR_filter_firBlock_left_firStep[180] );
nand U1981 ( n1410, my_FIR_filter_firBlock_left_multProducts[16], n1409 );
or U1982 ( n1409, n1408, my_FIR_filter_firBlock_left_firStep[176] );
nand U1983 ( n1420, my_FIR_filter_firBlock_left_multProducts[18], n1419 );
nand U1984 ( n1372, my_FIR_filter_firBlock_left_multProducts[8], n1371 );
nand U1985 ( n1447, my_FIR_filter_firBlock_left_multProducts[23], n1446 );
nand U1986 ( n1427, my_FIR_filter_firBlock_left_multProducts[19], n1426 );
or U1987 ( n1426, n1425, my_FIR_filter_firBlock_left_firStep[179] );
nand U1988 ( n1385, my_FIR_filter_firBlock_left_multProducts[11], n1384 );
nand U1989 ( n1395, my_FIR_filter_firBlock_left_multProducts[13], n1394 );
nand U1990 ( n1369, my_FIR_filter_firBlock_left_multProducts[7], n1368 );
nand U1991 ( n1363, my_FIR_filter_firBlock_left_multProducts[5], n1362 );
or U1992 ( n1362, n1492, my_FIR_filter_firBlock_left_firStep[165] );
nor U1993 ( n1482, my_FIR_filter_firBlock_left_firStep[190], n1483 );
xor U1994 ( my_FIR_filter_firBlock_left_multProducts[3], n1210, n1209 );
nor U1995 ( n713, my_FIR_filter_firBlock_left_firStep[286], n714 );
or U1996 ( n1345, n1344, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[38] );
xor U1997 ( n562, my_FIR_filter_firBlock_left_multProducts[113], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[38] );
nand U1998 ( n386, n385, n44 );
nand U1999 ( n377, my_FIR_filter_firBlock_left_multProducts[106], n374 );
or U2000 ( n375, n374, my_FIR_filter_firBlock_left_multProducts[106] );
nand U2001 ( n366, n365, n40 );
xor U2002 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[24], n344, n343 );
nand U2003 ( n304, n302, n301 );
nand U2004 ( n1893, my_FIR_filter_firBlock_left_multProducts[52], n1892 );
or U2005 ( n1892, n1891, my_FIR_filter_firBlock_left_firStep[85] );
nand U2006 ( n1841, my_FIR_filter_firBlock_left_multProducts[42], n1840 );
or U2007 ( n1840, n1839, my_FIR_filter_firBlock_left_firStep[75] );
nand U2008 ( n1908, my_FIR_filter_firBlock_left_multProducts[55], n1907 );
or U2009 ( n1907, n1906, my_FIR_filter_firBlock_left_firStep[88] );
nand U2010 ( n1918, my_FIR_filter_firBlock_left_multProducts[57], n1917 );
or U2011 ( n1917, n1916, my_FIR_filter_firBlock_left_firStep[90] );
nand U2012 ( n1898, my_FIR_filter_firBlock_left_multProducts[53], n1897 );
or U2013 ( n1897, n1896, my_FIR_filter_firBlock_left_firStep[86] );
nand U2014 ( n1876, my_FIR_filter_firBlock_left_multProducts[49], n1875 );
or U2015 ( n1875, n1874, my_FIR_filter_firBlock_left_firStep[82] );
nand U2016 ( n1888, my_FIR_filter_firBlock_left_multProducts[51], n1887 );
or U2017 ( n1887, n1886, my_FIR_filter_firBlock_left_firStep[84] );
nand U2018 ( n1856, my_FIR_filter_firBlock_left_multProducts[45], n1855 );
or U2019 ( n1855, n1854, my_FIR_filter_firBlock_left_firStep[78] );
nand U2020 ( n1866, my_FIR_filter_firBlock_left_multProducts[47], n1865 );
or U2021 ( n1865, n1864, my_FIR_filter_firBlock_left_firStep[80] );
nand U2022 ( n1846, my_FIR_filter_firBlock_left_multProducts[43], n1845 );
or U2023 ( n1845, n1844, my_FIR_filter_firBlock_left_firStep[76] );
nand U2024 ( n1828, my_FIR_filter_firBlock_left_multProducts[39], n1827 );
or U2025 ( n1827, n1955, my_FIR_filter_firBlock_left_firStep[72] );
nand U2026 ( n1836, my_FIR_filter_firBlock_left_multProducts[41], n1835 );
or U2027 ( n1835, n1834, my_FIR_filter_firBlock_left_firStep[74] );
nand U2028 ( n1822, my_FIR_filter_firBlock_left_multProducts[37], n1821 );
or U2029 ( n1821, n1951, my_FIR_filter_firBlock_left_firStep[70] );
nand U2030 ( n1816, my_FIR_filter_firBlock_left_multProducts[35], n1815 );
or U2031 ( n1815, n1947, my_FIR_filter_firBlock_left_firStep[68] );
nor U2032 ( n1938, my_FIR_filter_firBlock_left_firStep[94], n1939 );
nand U2033 ( n1939, n1936, n1935 );
xor U2034 ( my_FIR_filter_firBlock_left_N21, n661, n660 );
xor U2035 ( my_FIR_filter_firBlock_left_N7, n726, n725 );
xor U2036 ( my_FIR_filter_firBlock_left_N1, my_FIR_filter_firBlock_left_multProducts[61], my_FIR_filter_firBlock_left_firStep[256] );
xor U2037 ( my_FIR_filter_firBlock_left_N225, my_FIR_filter_firBlock_left_multProducts[61], my_FIR_filter_firBlock_left_firStep[32] );
nand U2038 ( n714, n711, n710 );
nand U2039 ( n664, my_FIR_filter_firBlock_left_firStep[276], n661 );
or U2040 ( n662, n661, my_FIR_filter_firBlock_left_firStep[276] );
nand U2041 ( n661, n659, n658 );
nand U2042 ( n609, n607, n606 );
nand U2043 ( n598, my_FIR_filter_firBlock_left_firStep[262], n726 );
or U2044 ( n596, n726, my_FIR_filter_firBlock_left_firStep[262] );
and U2045 ( n2032, my_FIR_filter_firBlock_left_multProducts[61], my_FIR_filter_firBlock_left_firStep[32] );
nand U2046 ( n286, n285, n22 );
nand U2047 ( n989, my_FIR_filter_firBlock_left_multProducts[56], n988 );
or U2048 ( n988, n987, my_FIR_filter_firBlock_left_firStep[249] );
nand U2049 ( n937, my_FIR_filter_firBlock_left_multProducts[46], n936 );
or U2050 ( n936, n935, my_FIR_filter_firBlock_left_firStep[239] );
nand U2051 ( n895, my_FIR_filter_firBlock_left_multProducts[36], n894 );
or U2052 ( n894, n1024, my_FIR_filter_firBlock_left_firStep[229] );
nand U2053 ( n1004, my_FIR_filter_firBlock_left_multProducts[59], n1003 );
or U2054 ( n1003, n1002, my_FIR_filter_firBlock_left_firStep[252] );
nand U2055 ( n994, my_FIR_filter_firBlock_left_multProducts[57], n993 );
or U2056 ( n993, n992, my_FIR_filter_firBlock_left_firStep[250] );
nand U2057 ( n974, my_FIR_filter_firBlock_left_multProducts[53], n973 );
or U2058 ( n973, n972, my_FIR_filter_firBlock_left_firStep[246] );
nand U2059 ( n984, my_FIR_filter_firBlock_left_multProducts[55], n983 );
or U2060 ( n983, n982, my_FIR_filter_firBlock_left_firStep[248] );
nand U2061 ( n952, my_FIR_filter_firBlock_left_multProducts[49], n951 );
or U2062 ( n951, n950, my_FIR_filter_firBlock_left_firStep[242] );
nand U2063 ( n964, my_FIR_filter_firBlock_left_multProducts[51], n963 );
or U2064 ( n963, n962, my_FIR_filter_firBlock_left_firStep[244] );
nand U2065 ( n942, my_FIR_filter_firBlock_left_multProducts[47], n941 );
or U2066 ( n941, n940, my_FIR_filter_firBlock_left_firStep[240] );
nand U2067 ( n922, my_FIR_filter_firBlock_left_multProducts[43], n921 );
or U2068 ( n921, n920, my_FIR_filter_firBlock_left_firStep[236] );
nand U2069 ( n932, my_FIR_filter_firBlock_left_multProducts[45], n931 );
or U2070 ( n931, n930, my_FIR_filter_firBlock_left_firStep[238] );
nand U2071 ( n904, my_FIR_filter_firBlock_left_multProducts[39], n903 );
or U2072 ( n903, n1031, my_FIR_filter_firBlock_left_firStep[232] );
nand U2073 ( n912, my_FIR_filter_firBlock_left_multProducts[41], n911 );
or U2074 ( n911, n910, my_FIR_filter_firBlock_left_firStep[234] );
nand U2075 ( n898, my_FIR_filter_firBlock_left_multProducts[37], n897 );
or U2076 ( n897, n1027, my_FIR_filter_firBlock_left_firStep[230] );
nand U2077 ( n1015, n1012, n1011 );
nand U2078 ( n1011, my_FIR_filter_firBlock_left_multProducts[60], n1010 );
xor U2079 ( my_FIR_filter_firBlock_left_N223, n1939, n1937 );
xnor U2080 ( n996, my_FIR_filter_firBlock_left_firStep[251], my_FIR_filter_firBlock_left_multProducts[58] );
xnor U2081 ( n1920, my_FIR_filter_firBlock_left_firStep[91], my_FIR_filter_firBlock_left_multProducts[58] );
xor U2082 ( n1153, my_FIR_filter_firBlock_left_multProducts[58], my_FIR_filter_firBlock_left_firStep[220] );
xor U2083 ( n1773, my_FIR_filter_firBlock_left_multProducts[58], my_FIR_filter_firBlock_left_firStep[124] );
and U2084 ( n1940, n1939, my_FIR_filter_firBlock_left_firStep[94] );
nand U2085 ( n1156, my_FIR_filter_firBlock_left_multProducts[58], n1155 );
nand U2086 ( n1776, my_FIR_filter_firBlock_left_multProducts[58], n1775 );
nand U2087 ( n1926, n1924, n1923 );
nand U2088 ( n999, my_FIR_filter_firBlock_left_multProducts[58], n998 );
nand U2089 ( n1923, my_FIR_filter_firBlock_left_multProducts[58], n1922 );
nand U2090 ( n852, my_FIR_filter_firBlock_left_multProducts[110], n849 );
or U2091 ( n850, n849, my_FIR_filter_firBlock_left_multProducts[110] );
nand U2092 ( n847, my_FIR_filter_firBlock_left_multProducts[109], n844 );
or U2093 ( n845, n844, my_FIR_filter_firBlock_left_multProducts[109] );
nand U2094 ( n836, my_FIR_filter_firBlock_left_multProducts[111], n835 );
nand U2095 ( n837, my_FIR_filter_firBlock_left_multProducts[107], n834 );
or U2096 ( n835, n834, my_FIR_filter_firBlock_left_multProducts[107] );
nand U2097 ( n817, my_FIR_filter_firBlock_left_multProducts[103], n814 );
or U2098 ( n815, n814, my_FIR_filter_firBlock_left_multProducts[103] );
nand U2099 ( n807, my_FIR_filter_firBlock_left_multProducts[101], n804 );
or U2100 ( n805, n804, my_FIR_filter_firBlock_left_multProducts[101] );
nand U2101 ( n802, my_FIR_filter_firBlock_left_multProducts[100], n799 );
or U2102 ( n800, n799, my_FIR_filter_firBlock_left_multProducts[100] );
nand U2103 ( n797, my_FIR_filter_firBlock_left_multProducts[99], n794 );
or U2104 ( n795, n794, my_FIR_filter_firBlock_left_multProducts[99] );
nand U2105 ( n787, my_FIR_filter_firBlock_left_multProducts[97], n784 );
or U2106 ( n785, n784, my_FIR_filter_firBlock_left_multProducts[97] );
nand U2107 ( n784, n782, n781 );
nand U2108 ( n767, my_FIR_filter_firBlock_left_multProducts[93], n764 );
or U2109 ( n765, n764, my_FIR_filter_firBlock_left_multProducts[93] );
nand U2110 ( n757, my_FIR_filter_firBlock_left_multProducts[91], n754 );
or U2111 ( n755, n754, my_FIR_filter_firBlock_left_multProducts[91] );
nand U2112 ( n749, n747, n746 );
nand U2113 ( n747, my_FIR_filter_firBlock_left_multProducts[93], n880 );
or U2114 ( n745, n880, my_FIR_filter_firBlock_left_multProducts[93] );
xor U2115 ( my_FIR_filter_firBlock_left_N253, n2078, n2077 );
nand U2116 ( n2081, my_FIR_filter_firBlock_left_firStep[60], n2078 );
nand U2117 ( n568, n566, n565 );
nand U2118 ( n558, n556, n555 );
nand U2119 ( n548, n546, n545 );
nand U2120 ( n536, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[32], n533 );
xor U2121 ( my_FIR_filter_firBlock_left_multProducts[80], n533, n532 );
nand U2122 ( n518, n516, n515 );
nand U2123 ( n516, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[28], n513 );
xor U2124 ( my_FIR_filter_firBlock_left_multProducts[76], n513, n512 );
nand U2125 ( n493, n491, n490 );
xor U2126 ( my_FIR_filter_firBlock_left_multProducts[70], n483, n482 );
nand U2127 ( n486, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[22], n483 );
or U2128 ( n484, n483, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[22] );
nand U2129 ( n478, n476, n475 );
nand U2130 ( n473, n471, n470 );
nand U2131 ( n451, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[15], n580 );
nand U2132 ( n710, my_FIR_filter_firBlock_left_multProducts[89], n709 );
nand U2133 ( n626, my_FIR_filter_firBlock_left_multProducts[74], n625 );
nand U2134 ( n600, my_FIR_filter_firBlock_left_multProducts[68], n599 );
nand U2135 ( n726, n595, n594 );
nand U2136 ( n621, my_FIR_filter_firBlock_left_multProducts[73], n620 );
nand U2137 ( n585, my_FIR_filter_firBlock_left_multProducts[63], n584 );
nand U2138 ( n428, n296, n295 );
xor U2139 ( my_FIR_filter_firBlock_left_N257, my_FIR_filter_firBlock_left_multProducts[90], my_FIR_filter_firBlock_left_firStep[0] );
xnor U2140 ( n1481, n53, my_FIR_filter_firBlock_left_firStep[190] );
xnor U2141 ( n1633, n53, my_FIR_filter_firBlock_left_firStep[158] );
nor U2142 ( n1485, n1482, n53 );
nor U2143 ( n1637, n1634, n53 );
nand U2144 ( n1333, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[35], n1330 );
or U2145 ( n1331, n1330, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[35] );
xor U2146 ( my_FIR_filter_firBlock_left_multProducts[26], n1325, n1324 );
nand U2147 ( n1328, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[34], n1325 );
or U2148 ( n1326, n1325, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[34] );
xor U2149 ( my_FIR_filter_firBlock_left_multProducts[24], n1315, n1314 );
nand U2150 ( n1318, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[32], n1315 );
or U2151 ( n1316, n1315, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[32] );
xor U2152 ( my_FIR_filter_firBlock_left_multProducts[23], n1310, n1309 );
nand U2153 ( n1313, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[31], n1310 );
or U2154 ( n1311, n1310, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[31] );
xor U2155 ( my_FIR_filter_firBlock_left_multProducts[20], n1295, n1294 );
nand U2156 ( n1298, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[28], n1295 );
or U2157 ( n1296, n1295, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[28] );
xor U2158 ( my_FIR_filter_firBlock_left_multProducts[19], n1290, n1289 );
nand U2159 ( n1293, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[27], n1290 );
or U2160 ( n1291, n1290, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[27] );
xor U2161 ( my_FIR_filter_firBlock_left_multProducts[18], n1285, n1284 );
nand U2162 ( n1288, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[26], n1285 );
or U2163 ( n1286, n1285, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[26] );
xor U2164 ( my_FIR_filter_firBlock_left_multProducts[16], n1275, n1274 );
nand U2165 ( n1278, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[24], n1275 );
or U2166 ( n1276, n1275, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[24] );
xor U2167 ( my_FIR_filter_firBlock_left_multProducts[14], n1265, n1264 );
nand U2168 ( n1268, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[22], n1265 );
or U2169 ( n1266, n1265, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[22] );
xor U2170 ( my_FIR_filter_firBlock_left_multProducts[13], n1260, n1259 );
nand U2171 ( n1263, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[21], n1260 );
or U2172 ( n1261, n1260, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[21] );
xor U2173 ( my_FIR_filter_firBlock_left_multProducts[11], n1250, n1249 );
nand U2174 ( n1253, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[19], n1250 );
or U2175 ( n1251, n1250, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[19] );
xor U2176 ( my_FIR_filter_firBlock_left_multProducts[10], n1245, n1244 );
xor U2177 ( my_FIR_filter_firBlock_left_multProducts[8], n1235, n1234 );
xor U2178 ( my_FIR_filter_firBlock_left_multProducts[7], n1230, n1229 );
nand U2179 ( n1233, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[15], n1230 );
or U2180 ( n1231, n1230, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[15] );
xor U2181 ( my_FIR_filter_firBlock_left_multProducts[5], n1220, n1219 );
nand U2182 ( n1223, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[13], n1220 );
or U2183 ( n1221, n1220, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[13] );
nand U2184 ( n450, my_FIR_filter_firBlock_left_multProducts[90], n449 );
xor U2185 ( my_FIR_filter_firBlock_left_multProducts[4], n1215, n1214 );
nand U2186 ( n1218, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[12], n1215 );
or U2187 ( n1216, n1215, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[12] );
nand U2188 ( n752, my_FIR_filter_firBlock_left_multProducts[90], n749 );
or U2189 ( n750, n749, my_FIR_filter_firBlock_left_multProducts[90] );
xor U2190 ( n748, my_FIR_filter_firBlock_left_multProducts[94], my_FIR_filter_firBlock_left_multProducts[90] );
xor U2191 ( n423, n22, my_FIR_filter_firBlock_left_multProducts[90] );
and U2192 ( n2184, my_FIR_filter_firBlock_left_multProducts[90], my_FIR_filter_firBlock_left_firStep[0] );
nand U2193 ( n738, my_FIR_filter_firBlock_left_multProducts[90], n875 );
or U2194 ( n736, n875, my_FIR_filter_firBlock_left_multProducts[90] );
xor U2195 ( n874, inData_in[2], my_FIR_filter_firBlock_left_multProducts[90] );
nand U2196 ( n1190, n1189, n1188 );
xnor U2197 ( n2062, my_FIR_filter_firBlock_left_firStep[57], my_FIR_filter_firBlock_left_multProducts[86] );
xnor U2198 ( n685, my_FIR_filter_firBlock_left_firStep[281], my_FIR_filter_firBlock_left_multProducts[86] );
nand U2199 ( n688, my_FIR_filter_firBlock_left_multProducts[86], n687 );
nand U2200 ( n404, my_FIR_filter_firBlock_left_multProducts[111], n401 );
xor U2201 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[35], n401, n398 );
or U2202 ( n402, n401, my_FIR_filter_firBlock_left_multProducts[111] );
nand U2203 ( n372, my_FIR_filter_firBlock_left_multProducts[105], n369 );
or U2204 ( n370, n369, my_FIR_filter_firBlock_left_multProducts[105] );
nand U2205 ( n337, my_FIR_filter_firBlock_left_multProducts[98], n334 );
or U2206 ( n335, n334, my_FIR_filter_firBlock_left_multProducts[98] );
xor U2207 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[14], n428, n427 );
xor U2208 ( my_FIR_filter_firBlock_left_N11, n609, n608 );
xor U2209 ( my_FIR_filter_firBlock_left_N17, n639, n638 );
xnor U2210 ( n720, my_FIR_filter_firBlock_left_firStep[259], my_FIR_filter_firBlock_left_multProducts[64] );
xnor U2211 ( n2097, my_FIR_filter_firBlock_left_firStep[35], my_FIR_filter_firBlock_left_multProducts[64] );
nand U2212 ( n696, n694, n693 );
nand U2213 ( n642, my_FIR_filter_firBlock_left_firStep[272], n639 );
or U2214 ( n640, n639, my_FIR_filter_firBlock_left_firStep[272] );
nand U2215 ( n612, my_FIR_filter_firBlock_left_firStep[266], n609 );
or U2216 ( n610, n609, my_FIR_filter_firBlock_left_firStep[266] );
nand U2217 ( n1238, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[16], n1235 );
xor U2218 ( n1234, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[16], n34 );
or U2219 ( n1236, n1235, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[16] );
nand U2220 ( n1965, my_FIR_filter_firBlock_left_multProducts[64], n1964 );
nand U2221 ( n588, my_FIR_filter_firBlock_left_multProducts[64], n587 );
nand U2222 ( n456, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[16], n453 );
xor U2223 ( my_FIR_filter_firBlock_left_multProducts[64], n453, n452 );
or U2224 ( n454, n453, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[16] );
xor U2225 ( n452, my_FIR_filter_firBlock_left_multProducts[91], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[16] );
xnor U2226 ( my_FIR_filter_firBlock_left_N228, n2097, n2096 );
xnor U2227 ( my_FIR_filter_firBlock_left_N230, n2101, n2100 );
xor U2228 ( my_FIR_filter_firBlock_left_N226, n2032, n2031 );
xor U2229 ( my_FIR_filter_firBlock_left_N239, n2006, n2005 );
xor U2230 ( my_FIR_filter_firBlock_left_N256, n2095, n2094 );
xor U2231 ( my_FIR_filter_firBlock_left_N243, n2026, n2025 );
xor U2232 ( my_FIR_filter_firBlock_left_N249, n2058, n2057 );
nand U2233 ( n2061, my_FIR_filter_firBlock_left_firStep[56], n2058 );
or U2234 ( n2059, n2058, my_FIR_filter_firBlock_left_firStep[56] );
nand U2235 ( n2033, n2029, n2028 );
nand U2236 ( n2029, my_FIR_filter_firBlock_left_firStep[50], n2026 );
nand U2237 ( n2021, n2019, n2018 );
nand U2238 ( n2009, my_FIR_filter_firBlock_left_firStep[46], n2006 );
nand U2239 ( n2006, n2004, n2003 );
nand U2240 ( n1991, n1989, n1988 );
nand U2241 ( n2108, n1981, n1980 );
nand U2242 ( n2107, n1978, n1977 );
nand U2243 ( n1972, my_FIR_filter_firBlock_left_firStep[37], n2100 );
or U2244 ( n1970, n2100, my_FIR_filter_firBlock_left_firStep[37] );
nand U2245 ( n1966, my_FIR_filter_firBlock_left_firStep[35], n2096 );
or U2246 ( n1964, n2096, my_FIR_filter_firBlock_left_firStep[35] );
nand U2247 ( n2096, n1963, n1962 );
nand U2248 ( n1960, my_FIR_filter_firBlock_left_firStep[33], n2032 );
or U2249 ( n1958, my_FIR_filter_firBlock_left_firStep[33], n2032 );
xor U2250 ( my_FIR_filter_firBlock_left_multProducts[61], n576, n575 );
nand U2251 ( n329, n327, n326 );
nand U2252 ( n326, n325, n32 );
nand U2253 ( n339, n337, n336 );
nand U2254 ( n336, n335, n34 );
nand U2255 ( n306, my_FIR_filter_firBlock_left_multProducts[92], n305 );
nand U2256 ( n298, n297, n26 );
nand U2257 ( n283, n282, n21 );
nand U2258 ( n311, my_FIR_filter_firBlock_left_multProducts[93], n310 );
nand U2259 ( n334, n332, n331 );
nand U2260 ( n331, n330, n33 );
nand U2261 ( n658, my_FIR_filter_firBlock_left_multProducts[80], n657 );
nand U2262 ( n673, my_FIR_filter_firBlock_left_multProducts[83], n672 );
nand U2263 ( n663, my_FIR_filter_firBlock_left_multProducts[81], n662 );
xor U2264 ( my_FIR_filter_firBlock_left_multProducts[73], n498, n497 );
xor U2265 ( n497, my_FIR_filter_firBlock_left_multProducts[100], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[25] );
xor U2266 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[25], n349, n348 );
nand U2267 ( n349, n347, n346 );
xnor U2268 ( my_FIR_filter_firBlock_left_N100, n1489, n1488 );
xnor U2269 ( my_FIR_filter_firBlock_left_N104, n1497, n1496 );
xnor U2270 ( my_FIR_filter_firBlock_left_N108, n1382, n1383 );
xnor U2271 ( my_FIR_filter_firBlock_left_N106, n1501, n1500 );
xnor U2272 ( my_FIR_filter_firBlock_left_N110, n1392, n1393 );
xnor U2273 ( my_FIR_filter_firBlock_left_N114, n1412, n1413 );
xnor U2274 ( my_FIR_filter_firBlock_left_N118, n1434, n1435 );
xnor U2275 ( my_FIR_filter_firBlock_left_N120, n1444, n1445 );
xnor U2276 ( my_FIR_filter_firBlock_left_N124, n1464, n1465 );
xor U2277 ( my_FIR_filter_firBlock_left_N105, n1499, n1498 );
xor U2278 ( my_FIR_filter_firBlock_left_N111, n1398, n1397 );
xor U2279 ( my_FIR_filter_firBlock_left_N115, n1418, n1417 );
xor U2280 ( my_FIR_filter_firBlock_left_N121, n1450, n1449 );
xor U2281 ( my_FIR_filter_firBlock_left_N125, n1470, n1469 );
xor U2282 ( my_FIR_filter_firBlock_left_N127, n1483, n1481 );
xor U2283 ( n1475, my_FIR_filter_firBlock_left_multProducts[2], my_FIR_filter_firBlock_left_firStep[162] );
xor U2284 ( n1627, my_FIR_filter_firBlock_left_multProducts[2], my_FIR_filter_firBlock_left_firStep[130] );
and U2285 ( n1484, n1483, my_FIR_filter_firBlock_left_firStep[190] );
nand U2286 ( n1473, my_FIR_filter_firBlock_left_firStep[188], n1470 );
or U2287 ( n1471, n1470, my_FIR_filter_firBlock_left_firStep[188] );
nand U2288 ( n1468, my_FIR_filter_firBlock_left_firStep[187], n1465 );
or U2289 ( n1466, n1465, my_FIR_filter_firBlock_left_firStep[187] );
nand U2290 ( n1453, my_FIR_filter_firBlock_left_firStep[184], n1450 );
or U2291 ( n1451, n1450, my_FIR_filter_firBlock_left_firStep[184] );
nand U2292 ( n1448, my_FIR_filter_firBlock_left_firStep[183], n1445 );
or U2293 ( n1446, n1445, my_FIR_filter_firBlock_left_firStep[183] );
nand U2294 ( n1438, my_FIR_filter_firBlock_left_firStep[181], n1435 );
nand U2295 ( n1437, my_FIR_filter_firBlock_left_multProducts[21], n1436 );
or U2296 ( n1436, n1435, my_FIR_filter_firBlock_left_firStep[181] );
nand U2297 ( n1421, my_FIR_filter_firBlock_left_firStep[178], n1418 );
or U2298 ( n1419, n1418, my_FIR_filter_firBlock_left_firStep[178] );
nand U2299 ( n1416, my_FIR_filter_firBlock_left_firStep[177], n1413 );
or U2300 ( n1414, n1413, my_FIR_filter_firBlock_left_firStep[177] );
nand U2301 ( n1401, my_FIR_filter_firBlock_left_firStep[174], n1398 );
or U2302 ( n1399, n1398, my_FIR_filter_firBlock_left_firStep[174] );
nand U2303 ( n1396, my_FIR_filter_firBlock_left_firStep[173], n1393 );
or U2304 ( n1394, n1393, my_FIR_filter_firBlock_left_firStep[173] );
nand U2305 ( n1386, my_FIR_filter_firBlock_left_firStep[171], n1383 );
or U2306 ( n1384, n1383, my_FIR_filter_firBlock_left_firStep[171] );
nand U2307 ( n1376, my_FIR_filter_firBlock_left_firStep[169], n1500 );
or U2308 ( n1374, n1500, my_FIR_filter_firBlock_left_firStep[169] );
nand U2309 ( n1373, my_FIR_filter_firBlock_left_firStep[168], n1499 );
or U2310 ( n1371, n1499, my_FIR_filter_firBlock_left_firStep[168] );
nand U2311 ( n1370, my_FIR_filter_firBlock_left_firStep[167], n1496 );
or U2312 ( n1368, n1496, my_FIR_filter_firBlock_left_firStep[167] );
nand U2313 ( n1506, my_FIR_filter_firBlock_left_multProducts[2], n1505 );
nand U2314 ( n1358, my_FIR_filter_firBlock_left_firStep[163], n1488 );
or U2315 ( n1356, n1488, my_FIR_filter_firBlock_left_firStep[163] );
nand U2316 ( n1354, my_FIR_filter_firBlock_left_multProducts[2], n1353 );
nand U2317 ( n1202, n1201, n27 );
nand U2318 ( n1203, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[9], n1349 );
xor U2319 ( my_FIR_filter_firBlock_left_multProducts[1], n1349, n1348 );
or U2320 ( n1201, n1349, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[9] );
xnor U2321 ( my_FIR_filter_firBlock_left_N132, n1641, n1640 );
xnor U2322 ( my_FIR_filter_firBlock_left_N136, n1649, n1648 );
xnor U2323 ( my_FIR_filter_firBlock_left_N134, n1645, n1644 );
xnor U2324 ( my_FIR_filter_firBlock_left_N140, n1534, n1535 );
xnor U2325 ( my_FIR_filter_firBlock_left_N138, n1653, n1652 );
xnor U2326 ( my_FIR_filter_firBlock_left_N142, n1544, n1545 );
xnor U2327 ( my_FIR_filter_firBlock_left_N146, n1564, n1565 );
xnor U2328 ( my_FIR_filter_firBlock_left_N144, n1554, n1555 );
xnor U2329 ( my_FIR_filter_firBlock_left_N150, n1586, n1587 );
xnor U2330 ( my_FIR_filter_firBlock_left_N148, n1574, n1577 );
xnor U2331 ( my_FIR_filter_firBlock_left_N152, n1596, n1597 );
xnor U2332 ( my_FIR_filter_firBlock_left_N156, n1616, n1617 );
xnor U2333 ( my_FIR_filter_firBlock_left_N154, n1606, n1607 );
xnor U2334 ( my_FIR_filter_firBlock_left_N158, n1626, n1629 );
xor U2335 ( my_FIR_filter_firBlock_left_N133, n1643, n1642 );
xor U2336 ( my_FIR_filter_firBlock_left_N141, n1540, n1539 );
xor U2337 ( my_FIR_filter_firBlock_left_N151, n1592, n1591 );
xor U2338 ( my_FIR_filter_firBlock_left_N159, n1635, n1633 );
xor U2339 ( n1423, my_FIR_filter_firBlock_left_multProducts[1], my_FIR_filter_firBlock_left_firStep[161] );
xor U2340 ( n1575, my_FIR_filter_firBlock_left_multProducts[1], my_FIR_filter_firBlock_left_firStep[129] );
and U2341 ( n1636, n1635, my_FIR_filter_firBlock_left_firStep[158] );
nand U2342 ( n1632, my_FIR_filter_firBlock_left_firStep[157], n1629 );
or U2343 ( n1630, n1629, my_FIR_filter_firBlock_left_firStep[157] );
nand U2344 ( n1620, my_FIR_filter_firBlock_left_firStep[155], n1617 );
or U2345 ( n1618, n1617, my_FIR_filter_firBlock_left_firStep[155] );
nand U2346 ( n1610, my_FIR_filter_firBlock_left_firStep[153], n1607 );
or U2347 ( n1608, n1607, my_FIR_filter_firBlock_left_firStep[153] );
nand U2348 ( n1600, my_FIR_filter_firBlock_left_firStep[151], n1597 );
or U2349 ( n1598, n1597, my_FIR_filter_firBlock_left_firStep[151] );
nand U2350 ( n1595, my_FIR_filter_firBlock_left_firStep[150], n1592 );
or U2351 ( n1593, n1592, my_FIR_filter_firBlock_left_firStep[150] );
nand U2352 ( n1590, my_FIR_filter_firBlock_left_firStep[149], n1587 );
or U2353 ( n1588, n1587, my_FIR_filter_firBlock_left_firStep[149] );
nand U2354 ( n1580, my_FIR_filter_firBlock_left_firStep[147], n1577 );
or U2355 ( n1578, n1577, my_FIR_filter_firBlock_left_firStep[147] );
nand U2356 ( n1568, my_FIR_filter_firBlock_left_firStep[145], n1565 );
or U2357 ( n1566, n1565, my_FIR_filter_firBlock_left_firStep[145] );
nand U2358 ( n1558, my_FIR_filter_firBlock_left_firStep[143], n1555 );
or U2359 ( n1556, n1555, my_FIR_filter_firBlock_left_firStep[143] );
nand U2360 ( n1548, my_FIR_filter_firBlock_left_firStep[141], n1545 );
or U2361 ( n1546, n1545, my_FIR_filter_firBlock_left_firStep[141] );
nand U2362 ( n1543, my_FIR_filter_firBlock_left_firStep[140], n1540 );
or U2363 ( n1541, n1540, my_FIR_filter_firBlock_left_firStep[140] );
nand U2364 ( n1538, my_FIR_filter_firBlock_left_firStep[139], n1535 );
or U2365 ( n1536, n1535, my_FIR_filter_firBlock_left_firStep[139] );
nand U2366 ( n1528, my_FIR_filter_firBlock_left_firStep[137], n1652 );
or U2367 ( n1526, n1652, my_FIR_filter_firBlock_left_firStep[137] );
nand U2368 ( n1522, my_FIR_filter_firBlock_left_firStep[135], n1648 );
or U2369 ( n1520, n1648, my_FIR_filter_firBlock_left_firStep[135] );
nand U2370 ( n1516, my_FIR_filter_firBlock_left_firStep[133], n1644 );
or U2371 ( n1514, n1644, my_FIR_filter_firBlock_left_firStep[133] );
nand U2372 ( n1513, my_FIR_filter_firBlock_left_firStep[132], n1643 );
or U2373 ( n1511, n1643, my_FIR_filter_firBlock_left_firStep[132] );
nand U2374 ( n1510, my_FIR_filter_firBlock_left_firStep[131], n1640 );
or U2375 ( n1508, n1640, my_FIR_filter_firBlock_left_firStep[131] );
nand U2376 ( n743, inData_in[4], n742 );
nand U2377 ( n1351, my_FIR_filter_firBlock_left_multProducts[1], n1350 );
nand U2378 ( n1503, my_FIR_filter_firBlock_left_multProducts[1], n1502 );
xor U2379 ( n878, inData_in[4], my_FIR_filter_firBlock_left_multProducts[92] );
xor U2380 ( n419, n20, inData_in[4] );
nor U2381 ( n1186, inData_in[5], inData_in[4] );
nand U2382 ( n606, my_FIR_filter_firBlock_left_multProducts[70], n605 );
nand U2383 ( n624, n622, n621 );
or U2384 ( n687, n686, my_FIR_filter_firBlock_left_firStep[281] );
or U2385 ( n593, n723, my_FIR_filter_firBlock_left_firStep[261] );
nand U2386 ( n676, n674, n673 );
nand U2387 ( n666, n664, n663 );
nand U2388 ( n719, n586, n585 );
or U2389 ( n657, n656, my_FIR_filter_firBlock_left_firStep[275] );
or U2390 ( n635, n634, my_FIR_filter_firBlock_left_firStep[271] );
or U2391 ( n605, n731, my_FIR_filter_firBlock_left_firStep[265] );
xor U2392 ( n575, inData_in[4], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[13] );
nand U2393 ( n545, my_FIR_filter_firBlock_left_multProducts[109], n544 );
nand U2394 ( n515, my_FIR_filter_firBlock_left_multProducts[103], n514 );
nand U2395 ( n565, my_FIR_filter_firBlock_left_multProducts[113], n564 );
nand U2396 ( n525, my_FIR_filter_firBlock_left_multProducts[105], n524 );
nand U2397 ( n513, n511, n510 );
nand U2398 ( n510, my_FIR_filter_firBlock_left_multProducts[102], n509 );
nand U2399 ( n475, my_FIR_filter_firBlock_left_multProducts[95], n474 );
nand U2400 ( n470, my_FIR_filter_firBlock_left_multProducts[94], n469 );
nand U2401 ( n460, my_FIR_filter_firBlock_left_multProducts[92], n459 );
nand U2402 ( n500, my_FIR_filter_firBlock_left_multProducts[100], n499 );
nand U2403 ( n483, n481, n480 );
nand U2404 ( n480, my_FIR_filter_firBlock_left_multProducts[96], n479 );
nand U2405 ( n447, inData_in[5], n446 );
nand U2406 ( n555, my_FIR_filter_firBlock_left_multProducts[111], n554 );
nand U2407 ( n444, inData_in[4], n443 );
or U2408 ( n499, n498, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[25] );
nand U2409 ( n573, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w3_38_, n572 );
nand U2410 ( n530, my_FIR_filter_firBlock_left_multProducts[106], n529 );
nand U2411 ( n570, my_FIR_filter_firBlock_left_multProducts[114], n569 );
nand U2412 ( n420, n284, n283 );
xor U2413 ( n680, my_FIR_filter_firBlock_left_multProducts[85], my_FIR_filter_firBlock_left_firStep[280] );
xor U2414 ( n2057, my_FIR_filter_firBlock_left_multProducts[85], my_FIR_filter_firBlock_left_firStep[56] );
nand U2415 ( n1343, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[37], n1340 );
or U2416 ( n1341, n1340, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[37] );
xor U2417 ( n1339, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[37], n58 );
nand U2418 ( n2060, my_FIR_filter_firBlock_left_multProducts[85], n2059 );
nand U2419 ( n683, my_FIR_filter_firBlock_left_multProducts[85], n682 );
nand U2420 ( n561, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[37], n558 );
xor U2421 ( n557, my_FIR_filter_firBlock_left_multProducts[112], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[37] );
nand U2422 ( n411, n409, n408 );
xor U2423 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[36], n406, n405 );
nand U2424 ( n409, my_FIR_filter_firBlock_left_multProducts[112], n406 );
or U2425 ( n407, n406, my_FIR_filter_firBlock_left_multProducts[112] );
nand U2426 ( n389, n387, n386 );
nand U2427 ( n387, my_FIR_filter_firBlock_left_multProducts[108], n384 );
or U2428 ( n385, n384, my_FIR_filter_firBlock_left_multProducts[108] );
nand U2429 ( n364, n362, n361 );
nand U2430 ( n357, my_FIR_filter_firBlock_left_multProducts[102], n354 );
xor U2431 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[26], n354, n353 );
or U2432 ( n355, n354, my_FIR_filter_firBlock_left_multProducts[102] );
nand U2433 ( n347, my_FIR_filter_firBlock_left_multProducts[100], n344 );
or U2434 ( n345, n344, my_FIR_filter_firBlock_left_multProducts[100] );
nand U2435 ( n342, my_FIR_filter_firBlock_left_multProducts[99], n339 );
or U2436 ( n340, n339, my_FIR_filter_firBlock_left_multProducts[99] );
xor U2437 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[21], n329, n328 );
nand U2438 ( n332, my_FIR_filter_firBlock_left_multProducts[97], n329 );
or U2439 ( n330, n329, my_FIR_filter_firBlock_left_multProducts[97] );
nand U2440 ( n301, n300, n27 );
nand U2441 ( n533, n531, n530 );
nand U2442 ( n463, n461, n460 );
or U2443 ( n489, n488, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[23] );
or U2444 ( n524, n523, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[30] );
or U2445 ( n559, n558, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[37] );
or U2446 ( n469, n468, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[19] );
or U2447 ( n494, n493, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[24] );
xor U2448 ( my_FIR_filter_firBlock_left_multProducts[87], n568, n567 );
or U2449 ( n534, n533, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[32] );
or U2450 ( n514, n513, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[28] );
or U2451 ( n449, n580, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[15] );
or U2452 ( n2079, n2078, my_FIR_filter_firBlock_left_firStep[60] );
nor U2453 ( n2094, n2093, n2092 );
xor U2454 ( my_FIR_filter_firBlock_left_N27, n691, n690 );
xor U2455 ( my_FIR_filter_firBlock_left_N23, n671, n670 );
xor U2456 ( my_FIR_filter_firBlock_left_N32, n718, n717 );
nor U2457 ( n717, n716, n715 );
xor U2458 ( n721, my_FIR_filter_firBlock_left_multProducts[65], my_FIR_filter_firBlock_left_firStep[260] );
xor U2459 ( n2098, my_FIR_filter_firBlock_left_multProducts[65], my_FIR_filter_firBlock_left_firStep[36] );
nand U2460 ( n694, my_FIR_filter_firBlock_left_firStep[282], n691 );
or U2461 ( n692, n691, my_FIR_filter_firBlock_left_firStep[282] );
nand U2462 ( n691, n689, n688 );
nand U2463 ( n674, my_FIR_filter_firBlock_left_firStep[278], n671 );
or U2464 ( n672, n671, my_FIR_filter_firBlock_left_firStep[278] );
nand U2465 ( n671, n669, n668 );
nand U2466 ( n656, n652, n651 );
nand U2467 ( n644, n642, n641 );
nand U2468 ( n634, n632, n631 );
nand U2469 ( n629, n627, n626 );
nand U2470 ( n731, n604, n603 );
nand U2471 ( n730, n601, n600 );
nand U2472 ( n1243, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[17], n1240 );
or U2473 ( n1241, n1240, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[17] );
xor U2474 ( n1239, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[17], n35 );
nand U2475 ( n591, my_FIR_filter_firBlock_left_multProducts[65], n590 );
xor U2476 ( n457, my_FIR_filter_firBlock_left_multProducts[92], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[17] );
nand U2477 ( n309, n307, n306 );
nand U2478 ( n307, n304, n28 );
or U2479 ( n305, n28, n304 );
nand U2480 ( n293, inData_in[4], n424 );
xor U2481 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[12], n424, n423 );
or U2482 ( n291, n424, inData_in[4] );
nand U2483 ( n1988, my_FIR_filter_firBlock_left_multProducts[71], n1987 );
or U2484 ( n1987, n1986, my_FIR_filter_firBlock_left_firStep[42] );
nand U2485 ( n424, n290, n289 );
nand U2486 ( n289, n288, n23 );
nand U2487 ( n2078, n2076, n2075 );
nand U2488 ( n2075, my_FIR_filter_firBlock_left_multProducts[88], n2074 );
nand U2489 ( n2058, n2056, n2055 );
nand U2490 ( n2026, n2024, n2023 );
nand U2491 ( n2023, my_FIR_filter_firBlock_left_multProducts[78], n2022 );
nand U2492 ( n2065, my_FIR_filter_firBlock_left_multProducts[86], n2064 );
nand U2493 ( n2100, n1969, n1968 );
nand U2494 ( n1968, my_FIR_filter_firBlock_left_multProducts[65], n1967 );
nand U2495 ( n2040, my_FIR_filter_firBlock_left_multProducts[81], n2039 );
or U2496 ( n2039, n2038, my_FIR_filter_firBlock_left_firStep[52] );
nand U2497 ( n2050, my_FIR_filter_firBlock_left_multProducts[83], n2049 );
nand U2498 ( n2028, my_FIR_filter_firBlock_left_multProducts[79], n2027 );
or U2499 ( n2027, n2026, my_FIR_filter_firBlock_left_firStep[50] );
nand U2500 ( n2008, my_FIR_filter_firBlock_left_multProducts[75], n2007 );
or U2501 ( n2007, n2006, my_FIR_filter_firBlock_left_firStep[46] );
nand U2502 ( n2018, my_FIR_filter_firBlock_left_multProducts[77], n2017 );
or U2503 ( n2017, n2016, my_FIR_filter_firBlock_left_firStep[48] );
nand U2504 ( n1980, my_FIR_filter_firBlock_left_multProducts[69], n1979 );
or U2505 ( n1979, n2107, my_FIR_filter_firBlock_left_firStep[40] );
or U2506 ( n1967, n2099, my_FIR_filter_firBlock_left_firStep[36] );
nand U2507 ( n2003, my_FIR_filter_firBlock_left_multProducts[74], n2002 );
nand U2508 ( n1977, my_FIR_filter_firBlock_left_multProducts[68], n1976 );
or U2509 ( n1976, n2104, my_FIR_filter_firBlock_left_firStep[39] );
nor U2510 ( n2090, my_FIR_filter_firBlock_left_firStep[62], n2091 );
xor U2511 ( my_FIR_filter_firBlock_left_multProducts[63], n580, n579 );
xor U2512 ( n579, my_FIR_filter_firBlock_left_multProducts[90], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[15] );
xor U2513 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[15], n430, n429 );
nand U2514 ( n430, n299, n298 );
xor U2515 ( my_FIR_filter_firBlock_left_N251, n2068, n2067 );
xnor U2516 ( n675, my_FIR_filter_firBlock_left_firStep[279], my_FIR_filter_firBlock_left_multProducts[84] );
xnor U2517 ( n2052, my_FIR_filter_firBlock_left_firStep[55], my_FIR_filter_firBlock_left_multProducts[84] );
nor U2518 ( n2093, n2090, n120 );
nand U2519 ( n1338, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[36], n1335 );
or U2520 ( n1336, n1335, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[36] );
xor U2521 ( n1334, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[36], n58 );
nand U2522 ( n2071, my_FIR_filter_firBlock_left_firStep[58], n2068 );
or U2523 ( n2069, n2068, my_FIR_filter_firBlock_left_firStep[58] );
nand U2524 ( n2068, n2066, n2065 );
nand U2525 ( n678, my_FIR_filter_firBlock_left_multProducts[84], n677 );
nand U2526 ( n2055, my_FIR_filter_firBlock_left_multProducts[84], n2054 );
nand U2527 ( n556, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[36], n553 );
or U2528 ( n554, n553, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[36] );
xor U2529 ( n552, my_FIR_filter_firBlock_left_multProducts[111], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[36] );
nand U2530 ( n397, my_FIR_filter_firBlock_left_multProducts[110], n394 );
xor U2531 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[34], n394, n393 );
or U2532 ( n395, n394, my_FIR_filter_firBlock_left_multProducts[110] );
nand U2533 ( n392, my_FIR_filter_firBlock_left_multProducts[109], n389 );
xor U2534 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[33], n389, n388 );
or U2535 ( n390, n389, my_FIR_filter_firBlock_left_multProducts[109] );
nand U2536 ( n384, n382, n381 );
xor U2537 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[31], n379, n378 );
nand U2538 ( n382, my_FIR_filter_firBlock_left_multProducts[107], n379 );
or U2539 ( n380, n379, my_FIR_filter_firBlock_left_multProducts[107] );
nand U2540 ( n367, my_FIR_filter_firBlock_left_multProducts[104], n364 );
or U2541 ( n365, n364, my_FIR_filter_firBlock_left_multProducts[104] );
nand U2542 ( n362, my_FIR_filter_firBlock_left_multProducts[103], n359 );
xor U2543 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[27], n359, n358 );
or U2544 ( n360, n359, my_FIR_filter_firBlock_left_multProducts[103] );
nand U2545 ( n352, my_FIR_filter_firBlock_left_multProducts[101], n349 );
or U2546 ( n350, n349, my_FIR_filter_firBlock_left_multProducts[101] );
xor U2547 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[20], n324, n323 );
nand U2548 ( n327, my_FIR_filter_firBlock_left_multProducts[96], n324 );
or U2549 ( n325, n324, my_FIR_filter_firBlock_left_multProducts[96] );
nand U2550 ( n322, my_FIR_filter_firBlock_left_multProducts[95], n319 );
or U2551 ( n320, n319, my_FIR_filter_firBlock_left_multProducts[95] );
nand U2552 ( n314, n312, n311 );
xor U2553 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[17], n309, n308 );
nand U2554 ( n312, n309, n29 );
or U2555 ( n310, n29, n309 );
nand U2556 ( n302, my_FIR_filter_firBlock_left_multProducts[91], n430 );
or U2557 ( n300, n430, my_FIR_filter_firBlock_left_multProducts[91] );
xor U2558 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[8], n400, n399 );
xor U2559 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[10], n420, n419 );
nand U2560 ( n287, inData_in[2], n420 );
or U2561 ( n285, n420, inData_in[2] );
xnor U2562 ( my_FIR_filter_firBlock_left_N30, n705, n708 );
xor U2563 ( n690, my_FIR_filter_firBlock_left_multProducts[87], my_FIR_filter_firBlock_left_firStep[282] );
xor U2564 ( n2067, my_FIR_filter_firBlock_left_multProducts[87], my_FIR_filter_firBlock_left_firStep[58] );
nor U2565 ( n716, n713, n120 );
nand U2566 ( n711, my_FIR_filter_firBlock_left_firStep[285], n708 );
or U2567 ( n709, n708, my_FIR_filter_firBlock_left_firStep[285] );
nand U2568 ( n2070, my_FIR_filter_firBlock_left_multProducts[87], n2069 );
nand U2569 ( n693, my_FIR_filter_firBlock_left_multProducts[87], n692 );
nand U2570 ( n566, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[38], n563 );
xor U2571 ( my_FIR_filter_firBlock_left_multProducts[86], n563, n562 );
or U2572 ( n564, n563, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[38] );
nand U2573 ( n551, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[35], n548 );
xor U2574 ( my_FIR_filter_firBlock_left_multProducts[83], n548, n547 );
or U2575 ( n549, n548, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[35] );
nand U2576 ( n546, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[34], n543 );
xor U2577 ( my_FIR_filter_firBlock_left_multProducts[82], n543, n542 );
or U2578 ( n544, n543, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[34] );
xor U2579 ( my_FIR_filter_firBlock_left_multProducts[81], n538, n537 );
nand U2580 ( n541, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[33], n538 );
or U2581 ( n539, n538, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[33] );
xor U2582 ( my_FIR_filter_firBlock_left_multProducts[79], n528, n527 );
nand U2583 ( n531, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[31], n528 );
or U2584 ( n529, n528, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[31] );
xor U2585 ( my_FIR_filter_firBlock_left_multProducts[77], n518, n517 );
nand U2586 ( n521, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[29], n518 );
or U2587 ( n519, n518, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[29] );
xor U2588 ( my_FIR_filter_firBlock_left_multProducts[75], n508, n507 );
nand U2589 ( n511, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[27], n508 );
or U2590 ( n509, n508, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[27] );
xor U2591 ( my_FIR_filter_firBlock_left_multProducts[74], n503, n502 );
nand U2592 ( n506, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[26], n503 );
or U2593 ( n504, n503, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[26] );
nand U2594 ( n503, n501, n500 );
xor U2595 ( my_FIR_filter_firBlock_left_multProducts[69], n478, n477 );
nand U2596 ( n481, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[21], n478 );
or U2597 ( n479, n478, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[21] );
xor U2598 ( my_FIR_filter_firBlock_left_multProducts[68], n473, n472 );
nand U2599 ( n476, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[20], n473 );
or U2600 ( n474, n473, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[20] );
xor U2601 ( my_FIR_filter_firBlock_left_multProducts[65], n458, n457 );
nand U2602 ( n461, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[17], n458 );
or U2603 ( n459, n458, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[17] );
nand U2604 ( n458, n456, n455 );
nand U2605 ( n1208, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[10], n1205 );
or U2606 ( n1206, n1205, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[10] );
nand U2607 ( n580, n448, n447 );
xor U2608 ( n1204, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[10], n28 );
nand U2609 ( n578, n445, n444 );
xor U2610 ( n872, inData_in[5], inData_in[1] );
nand U2611 ( n735, inData_in[1], n873 );
or U2612 ( n733, inData_in[1], n873 );
nand U2613 ( n434, inData_in[1], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[10] );
or U2614 ( n431, inData_in[1], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[10] );
xor U2615 ( n417, inData_in[3], inData_in[1] );
xnor U2616 ( my_FIR_filter_firBlock_left_N4, n720, n719 );
xnor U2617 ( my_FIR_filter_firBlock_left_N8, n728, n727 );
xnor U2618 ( my_FIR_filter_firBlock_left_N12, n613, n614 );
xnor U2619 ( my_FIR_filter_firBlock_left_N14, n623, n624 );
xnor U2620 ( my_FIR_filter_firBlock_left_N18, n643, n644 );
xnor U2621 ( my_FIR_filter_firBlock_left_N22, n665, n666 );
xnor U2622 ( my_FIR_filter_firBlock_left_N24, n675, n676 );
xnor U2623 ( my_FIR_filter_firBlock_left_N28, n695, n696 );
xor U2624 ( my_FIR_filter_firBlock_left_N5, n722, n721 );
xor U2625 ( my_FIR_filter_firBlock_left_N9, n730, n729 );
xor U2626 ( my_FIR_filter_firBlock_left_N15, n629, n628 );
xor U2627 ( my_FIR_filter_firBlock_left_N19, n649, n648 );
xor U2628 ( my_FIR_filter_firBlock_left_N25, n681, n680 );
xor U2629 ( my_FIR_filter_firBlock_left_N29, n701, n700 );
xor U2630 ( my_FIR_filter_firBlock_left_N31, n714, n712 );
xor U2631 ( n654, my_FIR_filter_firBlock_left_multProducts[62], my_FIR_filter_firBlock_left_firStep[257] );
xor U2632 ( n2031, my_FIR_filter_firBlock_left_multProducts[62], my_FIR_filter_firBlock_left_firStep[33] );
and U2633 ( n715, n714, my_FIR_filter_firBlock_left_firStep[286] );
nand U2634 ( n704, my_FIR_filter_firBlock_left_firStep[284], n701 );
or U2635 ( n702, n701, my_FIR_filter_firBlock_left_firStep[284] );
nand U2636 ( n699, my_FIR_filter_firBlock_left_firStep[283], n696 );
or U2637 ( n697, n696, my_FIR_filter_firBlock_left_firStep[283] );
nand U2638 ( n684, my_FIR_filter_firBlock_left_firStep[280], n681 );
or U2639 ( n682, n681, my_FIR_filter_firBlock_left_firStep[280] );
nand U2640 ( n679, my_FIR_filter_firBlock_left_firStep[279], n676 );
or U2641 ( n677, n676, my_FIR_filter_firBlock_left_firStep[279] );
nand U2642 ( n669, my_FIR_filter_firBlock_left_firStep[277], n666 );
nand U2643 ( n668, my_FIR_filter_firBlock_left_multProducts[82], n667 );
or U2644 ( n667, n666, my_FIR_filter_firBlock_left_firStep[277] );
nand U2645 ( n652, my_FIR_filter_firBlock_left_firStep[274], n649 );
or U2646 ( n650, n649, my_FIR_filter_firBlock_left_firStep[274] );
nand U2647 ( n647, my_FIR_filter_firBlock_left_firStep[273], n644 );
or U2648 ( n645, n644, my_FIR_filter_firBlock_left_firStep[273] );
nand U2649 ( n632, my_FIR_filter_firBlock_left_firStep[270], n629 );
or U2650 ( n630, n629, my_FIR_filter_firBlock_left_firStep[270] );
nand U2651 ( n627, my_FIR_filter_firBlock_left_firStep[269], n624 );
or U2652 ( n625, n624, my_FIR_filter_firBlock_left_firStep[269] );
nand U2653 ( n617, my_FIR_filter_firBlock_left_firStep[267], n614 );
nand U2654 ( n616, my_FIR_filter_firBlock_left_multProducts[72], n615 );
or U2655 ( n615, n614, my_FIR_filter_firBlock_left_firStep[267] );
nand U2656 ( n604, my_FIR_filter_firBlock_left_firStep[264], n730 );
or U2657 ( n602, n730, my_FIR_filter_firBlock_left_firStep[264] );
nand U2658 ( n601, my_FIR_filter_firBlock_left_firStep[263], n727 );
or U2659 ( n599, n727, my_FIR_filter_firBlock_left_firStep[263] );
nand U2660 ( n1228, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[14], n1225 );
or U2661 ( n1226, n1225, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[14] );
xor U2662 ( n1224, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[14], n32 );
nand U2663 ( n592, my_FIR_filter_firBlock_left_firStep[260], n722 );
or U2664 ( n590, n722, my_FIR_filter_firBlock_left_firStep[260] );
nand U2665 ( n589, my_FIR_filter_firBlock_left_firStep[259], n719 );
or U2666 ( n587, n719, my_FIR_filter_firBlock_left_firStep[259] );
nand U2667 ( n1959, my_FIR_filter_firBlock_left_multProducts[62], n1958 );
nand U2668 ( n582, my_FIR_filter_firBlock_left_multProducts[62], n581 );
nand U2669 ( n448, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[14], n578 );
or U2670 ( n446, n578, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[14] );
xor U2671 ( n577, inData_in[5], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[14] );
xor U2672 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[11], n422, n421 );
nand U2673 ( n290, inData_in[3], n422 );
or U2674 ( n288, n422, inData_in[3] );
xor U2675 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[9], n418, n417 );
or U2676 ( n284, n18, n418 );
nand U2677 ( n282, n418, n18 );
xnor U2678 ( my_FIR_filter_firBlock_left_N254, n2082, n2085 );
xnor U2679 ( my_FIR_filter_firBlock_left_N236, n1990, n1991 );
xnor U2680 ( my_FIR_filter_firBlock_left_N234, n2109, n2108 );
xnor U2681 ( my_FIR_filter_firBlock_left_N238, n2000, n2001 );
xnor U2682 ( my_FIR_filter_firBlock_left_N242, n2020, n2021 );
xnor U2683 ( my_FIR_filter_firBlock_left_N240, n2010, n2011 );
xnor U2684 ( my_FIR_filter_firBlock_left_N246, n2042, n2043 );
xnor U2685 ( my_FIR_filter_firBlock_left_N244, n2030, n2033 );
xnor U2686 ( my_FIR_filter_firBlock_left_N248, n2052, n2053 );
xnor U2687 ( my_FIR_filter_firBlock_left_N252, n2072, n2073 );
xnor U2688 ( my_FIR_filter_firBlock_left_N250, n2062, n2063 );
xor U2689 ( my_FIR_filter_firBlock_left_N237, n1996, n1995 );
xor U2690 ( my_FIR_filter_firBlock_left_N247, n2048, n2047 );
xor U2691 ( my_FIR_filter_firBlock_left_N255, n2091, n2089 );
xnor U2692 ( n724, my_FIR_filter_firBlock_left_firStep[261], my_FIR_filter_firBlock_left_multProducts[66] );
xnor U2693 ( n2101, my_FIR_filter_firBlock_left_firStep[37], my_FIR_filter_firBlock_left_multProducts[66] );
and U2694 ( n2092, n2091, my_FIR_filter_firBlock_left_firStep[62] );
nand U2695 ( n2088, my_FIR_filter_firBlock_left_firStep[61], n2085 );
or U2696 ( n2086, n2085, my_FIR_filter_firBlock_left_firStep[61] );
nand U2697 ( n2076, my_FIR_filter_firBlock_left_firStep[59], n2073 );
or U2698 ( n2074, n2073, my_FIR_filter_firBlock_left_firStep[59] );
nand U2699 ( n2066, my_FIR_filter_firBlock_left_firStep[57], n2063 );
or U2700 ( n2064, n2063, my_FIR_filter_firBlock_left_firStep[57] );
nand U2701 ( n2056, my_FIR_filter_firBlock_left_firStep[55], n2053 );
or U2702 ( n2054, n2053, my_FIR_filter_firBlock_left_firStep[55] );
nand U2703 ( n2051, my_FIR_filter_firBlock_left_firStep[54], n2048 );
or U2704 ( n2049, n2048, my_FIR_filter_firBlock_left_firStep[54] );
nand U2705 ( n2046, my_FIR_filter_firBlock_left_firStep[53], n2043 );
or U2706 ( n2044, n2043, my_FIR_filter_firBlock_left_firStep[53] );
nand U2707 ( n2036, my_FIR_filter_firBlock_left_firStep[51], n2033 );
or U2708 ( n2034, n2033, my_FIR_filter_firBlock_left_firStep[51] );
nand U2709 ( n2024, my_FIR_filter_firBlock_left_firStep[49], n2021 );
or U2710 ( n2022, n2021, my_FIR_filter_firBlock_left_firStep[49] );
nand U2711 ( n2014, my_FIR_filter_firBlock_left_firStep[47], n2011 );
or U2712 ( n2012, n2011, my_FIR_filter_firBlock_left_firStep[47] );
nand U2713 ( n2004, my_FIR_filter_firBlock_left_firStep[45], n2001 );
or U2714 ( n2002, n2001, my_FIR_filter_firBlock_left_firStep[45] );
nand U2715 ( n1999, my_FIR_filter_firBlock_left_firStep[44], n1996 );
or U2716 ( n1997, n1996, my_FIR_filter_firBlock_left_firStep[44] );
nand U2717 ( n1994, my_FIR_filter_firBlock_left_firStep[43], n1991 );
or U2718 ( n1992, n1991, my_FIR_filter_firBlock_left_firStep[43] );
nand U2719 ( n1248, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[18], n1245 );
or U2720 ( n1246, n1245, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[18] );
nand U2721 ( n1984, my_FIR_filter_firBlock_left_firStep[41], n2108 );
xor U2722 ( n1244, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[18], n36 );
or U2723 ( n1982, n2108, my_FIR_filter_firBlock_left_firStep[41] );
nand U2724 ( n594, my_FIR_filter_firBlock_left_multProducts[66], n593 );
nand U2725 ( n1971, my_FIR_filter_firBlock_left_multProducts[66], n1970 );
nand U2726 ( n466, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[18], n463 );
xor U2727 ( my_FIR_filter_firBlock_left_multProducts[66], n463, n462 );
or U2728 ( n464, n463, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[18] );
xor U2729 ( n462, my_FIR_filter_firBlock_left_multProducts[93], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[18] );
nand U2730 ( n317, my_FIR_filter_firBlock_left_multProducts[94], n314 );
xor U2731 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[18], n314, n313 );
or U2732 ( n315, n314, my_FIR_filter_firBlock_left_multProducts[94] );
nand U2733 ( n299, my_FIR_filter_firBlock_left_multProducts[90], n428 );
or U2734 ( n297, n428, my_FIR_filter_firBlock_left_multProducts[90] );
nand U2735 ( n296, inData_in[5], n426 );
or U2736 ( n294, n426, inData_in[5] );
xor U2737 ( n399, inData_in[2], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[6] );
xor U2738 ( my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[7], inData_in[1], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nor U2739 ( n1192, my_FIR_filter_firBlock_left_multProducts[90], n19 );
and U2740 ( n873, inData_in[4], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nor U2741 ( n1189, inData_in[1], my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nand U2742 ( n1188, my_FIR_filter_firBlock_left_multProducts[90], n19 );
nand U2743 ( n433, n432, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nand U2744 ( n281, n19, n400 );
nand U2745 ( n400, n19, n18 );
endmodule

