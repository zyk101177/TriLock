
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule


module s15850_ori ( clk, reset, g18, g27, g109, g741, g742, g743, g744, g872, g873,
g877, g881, g1960, g1961, g2355, g2601, g2602, g2603, g2604,
g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648, g2986,
g3007, g3069, g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179,
g4180, g4181, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920,
g6926, g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313,
g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352,
g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977, g8978, g8979,
g8980, g8981, g8982, g8983, g8984, g8985, g8986, g9451, g9961, g10377,
g10379, g10455, g10457, g10459, g10461, g10463, g10465, g10628, g10801,
g11163, g11206, g11489 );
input clk, reset, g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, g881, g1960, g1961;
output g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609,
g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172, g4173, g4174,
g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4887, g4888, g5101,
g5105, g5658, g5659, g5816, g6920, g6926, g6932, g6942, g6949, g6955,
g7744, g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331,
g8335, g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565,
g8566, g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984,
g8985, g8986, g9451, g9961, g10377, g10379, g10455, g10457, g10459,
g10461, g10463, g10465, g10628, g10801, g11163, g11206, g11489;
wire g4178, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, ex_wire30, ex_wire31, ex_wire32, ex_wire33, ex_wire34, ex_wire35, ex_wire36, ex_wire37, ex_wire38, ex_wire39, ex_wire40, ex_wire41, ex_wire42, ex_wire43, ex_wire44, ex_wire45, ex_wire46, ex_wire47, ex_wire48, ex_wire49, ex_wire50, ex_wire51, ex_wire52, ex_wire53, ex_wire54, ex_wire55, ex_wire56, ex_wire57, ex_wire58, ex_wire59, ex_wire60, ex_wire61, ex_wire62, ex_wire63, ex_wire64, ex_wire65, ex_wire66, ex_wire67, ex_wire68, ex_wire69, ex_wire70, ex_wire71, ex_wire72, ex_wire73, ex_wire74, ex_wire75, ex_wire76, ex_wire77, ex_wire78, ex_wire79, ex_wire80, ex_wire81, ex_wire82, ex_wire83, ex_wire84, ex_wire85, ex_wire86, ex_wire87, ex_wire88, ex_wire89, ex_wire90, ex_wire91, ex_wire92, ex_wire93, ex_wire94, ex_wire95, ex_wire96, ex_wire97, ex_wire98, ex_wire99, ex_wire100, ex_wire101, ex_wire102, ex_wire103, ex_wire104, ex_wire105, ex_wire106, ex_wire107, ex_wire108, ex_wire109, ex_wire110, ex_wire111, ex_wire112, ex_wire113, ex_wire114, ex_wire115, ex_wire116, ex_wire117, ex_wire118, ex_wire119, ex_wire120, ex_wire121, ex_wire122, ex_wire123, ex_wire124, ex_wire125, ex_wire126, ex_wire127, ex_wire128, ex_wire129, ex_wire130, ex_wire131, ex_wire132, ex_wire133, ex_wire134, ex_wire135, ex_wire136, ex_wire137, ex_wire138, ex_wire139, ex_wire140, ex_wire141, ex_wire142, ex_wire143, ex_wire144, ex_wire145, ex_wire146, ex_wire147, ex_wire148, ex_wire149, ex_wire150, ex_wire151, ex_wire152, ex_wire153, ex_wire154, ex_wire155, ex_wire156, ex_wire157, ex_wire158, ex_wire159, ex_wire160, ex_wire161, ex_wire162, ex_wire163, ex_wire164, ex_wire165, ex_wire166, ex_wire167, ex_wire168, ex_wire169, g18, g27, g872, g873, g1960, g1961, g794, g798, g802, g806, g810,
g814, g818, g822, g1958, g108, g253, g256, g257, g258, g259, g260,
g261, g262, g254, g1170, g1173, g1176, g1854, g1179, g1182, g1185,
g1188, g1191, g1194, g38, g42, g30, g40, g43, g31, g44, g82, g45, g46,
g746, g47, g83, g101, g48, g102, g103, g41, g104, g28, g925, g1713,
g757, g756, g29, g886, g889, g892, g895, g636, g898, g901, g904, g907,
g910, g913, g916, g919, g922, g255, g826, g1197, g1200, g1203,
new_g2478_, new_g2791_, new_g3524_, g6920, g6926, g6932, g6942, g6949,
g6955, new_g4076_, new_g4089_, new_g3462_, new_g4114_, new_g4117_,
new_g3506_, new_g3381_, new_g4231_, new_g4238_, new_g4239_,
new_g4255_, new_g4264_, new_g4274_, new_g4283_, new_g4293_,
new_g4309_, new_g4325_, new_g4330_, new_g4334_, new_g4338_,
new_g4340_, new_g4342_, new_g4465_, new_g4471_, new_g4473_,
new_g4477_, new_g4480_, new_g4484_, new_g4556_, new_g4490_,
new_g4498_, new_g4500_, new_g4506_, new_g4890_, new_g4891_,
new_g4893_, new_g4902_, new_g4903_, new_g4904_, new_g4905_,
new_g5392_, new_g4940_, new_g5445_, new_g5421_, new_g5556_,
new_g5083_, new_g5126_, new_g5148_, new_g5173_, new_g5194_,
new_g5287_, new_g5396_, new_g5404_, new_g5390_, new_g5529_,
new_g5536_, new_g5543_, new_g6126_, new_g6163_, new_g6243_,
new_g6179_, new_g6180_, new_g6193_, new_g6198_, new_g6205_,
new_g6216_, new_g6224_, new_g6244_, new_g5755_, new_g5770_,
new_g5849_, new_g6049_, new_g6155_, new_g5910_, new_g5914_,
new_g5763_, new_g5996_, new_g6000_, new_g6002_, new_g6015_,
new_g6026_, new_g6035_, new_g6038_, new_g6042_, new_g6045_,
new_g6054_, new_g6059_, new_g6068_, new_g6071_, new_g6080_,
new_g6088_, new_g6093_, new_g6096_, new_g6099_, new_g6123_,
new_g6331_, new_g6332_, new_g6333_, new_g6334_, new_g6728_,
new_g6733_, new_g6755_, new_g6747_, new_g6757_, new_g6759_,
new_g6786_, new_g6795_, new_g6656_, new_g6679_, new_g6439_,
new_g6468_, new_g6469_, new_g6470_, new_g6478_, new_g6479_,
new_g6480_, new_g6481_, new_g6500_, new_g6501_, new_g6506_,
new_g6507_, new_g6513_, new_g6514_, new_g6515_, new_g6522_,
new_g6523_, new_g6524_, new_g6528_, new_g6529_, new_g6533_,
new_g6534_, new_g6471_, new_g6537_, new_g6538_, new_g6541_,
new_g6542_, new_g6545_, new_g6546_, new_g6502_, new_g6551_,
new_g6508_, new_g6516_, new_g6525_, new_g6526_, new_g6531_,
new_g6672_, new_g6621_, new_g6627_, new_g6638_, new_g6653_,
new_g6819_, new_g6820_, new_g6821_, new_g6822_, new_g6823_,
new_g6824_, new_g6826_, new_g6827_, new_g6828_, new_g6829_,
new_g6830_, new_g6831_, new_g6832_, new_g6833_, new_g6834_,
new_g6838_, new_g6839_, new_g6840_, new_g6841_, new_g7032_,
new_g7191_, new_g7244_, new_g7202_, new_g7257_, new_g6894_,
new_g6895_, new_g6898_, new_g6897_, new_g6902_, new_g6900_,
new_g6901_, new_g6908_, new_g6909_, new_g6906_, new_g6907_,
new_g6912_, new_g6910_, new_g6911_, new_g6918_, new_g6915_,
new_g6916_, new_g6924_, new_g6922_, new_g6923_, new_g6930_,
new_g6928_, new_g6929_, new_g6934_, new_g6983_, new_g7133_,
new_g7143_, new_g7183_, new_g7134_, new_g7189_, new_g7137_,
new_g7204_, new_g7219_, new_g7705_, new_g7709_, new_g7441_,
new_g7626_, new_g7541_, new_g7581_, new_g7586_, new_g7590_,
new_g7660_, new_g7632_, new_g8019_, new_g8024_, new_g8039_,
new_g8040_, new_g8041_, new_g8042_, new_g8043_, new_g8044_,
new_g8045_, new_g8046_, new_g8047_, new_g8048_, new_g8049_,
new_g8050_, new_g8051_, new_g8052_, new_g8053_, new_g8054_,
new_g8055_, new_g8059_, new_g8060_, new_g7843_, new_g7930_,
new_g8244_, new_g8245_, new_g8250_, new_g8254_, new_g8260_,
new_g8147_, new_g8173_, new_g8193_, new_g8194_, new_g8384_,
new_g8559_, new_g8505_, new_g8631_, new_g8649_, new_g8770_,
new_g8771_, new_g8773_, new_g8774_, new_g8776_, new_g8765_,
new_g8777_, new_g8766_, new_g8779_, new_g8767_, new_g8768_,
new_g8769_, new_g8772_, new_g8775_, new_g8820_, new_g8937_,
new_g8938_, new_g8939_, new_g8940_, new_g8941_, new_g8944_,
new_g8945_, new_g8973_, new_g8922_, new_g8921_, new_g8943_,
new_g8883_, new_g8885_, new_g8887_, new_g8889_, new_g8920_,
new_g8923_, new_g8926_, new_g9272_, new_g9110_, new_g9124_,
new_g9150_, new_g9266_, new_g9269_, new_g9555_, new_g9721_, g9961,
new_g10663_, new_g10664_, new_g10765_, new_g10767_, new_g10770_,
new_g10771_, new_g10773_, new_g10707_, new_g10711_, new_g10717_,
new_g10718_, new_g10719_, new_g10720_, new_g10721_, new_g10722_,
new_g10726_, new_g10858_, new_g10859_, new_g10860_, new_g10861_,
new_g10862_, new_g10863_, new_g10864_, new_g10865_, new_g10866_,
new_g10776_, new_g10791_, new_g10793_, new_g10795_, new_g10780_,
new_g10797_, new_g10782_, new_g10798_, new_g10784_, new_g10799_,
new_g10785_, new_g10800_, new_g10788_, new_g10855_, new_g10898_,
new_g10936_, new_g11305_, new_g11306_, new_g11308_, new_g11310_,
new_g11312_, new_g11314_, new_g11320_, new_g11294_, new_g11293_,
new_g11290_, new_g11291_, new_g11292_, new_g11298_, new_g11300_,
new_g11303_, new_g11391_, new_g11392_, new_g11393_, new_g11340_,
new_g11349_, new_g11372_, new_g11376_, new_g11380_, new_g11478_,
new_g11481_, new_g11482_, new_g11483_, new_g11484_, new_g11485_,
new_g11486_, new_g11487_, new_g11488_, new_g11514_, new_g11561_,
new_g11579_, new_g11602_, new_g11603_, new_g11604_, new_g11605_,
new_g11606_, new_g11607_, new_g11608_, new_g11609_, new_g11610_,
new_g11625_, new_g11639_, new_g11640_, new_g11641_, new_g11636_,
new_g11647_, g1765, g1710, g632, g1850, g8, g17, g1317, n2181, n2186,
n2191, n2196, n2201, n2206, n2141, n2146, n2151, n2156, n2161, n2166,
n2171, n2176, n1810, n1815, n1820, n1825, n1830, n1835, n1840, n1845,
n1184, n1189, n1194, n1199, n1204, n1209, n1214, n1219, n1379, n1424,
n1429, n1434, n1439, n1444, n1449, n1384, n1389, n1394, n1399, n1404,
n1409, n1414, n1419, n1234, n1279, n1284, n1289, n1294, n1299, n1304,
n1239, n1244, n1249, n1254, n1259, n1264, n1269, n1274, n2136, g1737,
n596, n765, n774, n1588, n1597, n1601, n1605, n1864, n2102, n2111,
n2235, N41, n3, n7, n44, n68, n122, g8271, n186, n192, n2187, n2188,
n2189, n2190, n2192, n2194, n2195, n2197, n2198, n2199, n2200, n2202,
n2203, n2204, n2205, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
n2234, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773;
assign g2355 = g18;
assign g7744 = g27;
assign g8061 = g872;
assign g5101 = g872;
assign g8062 = g873;
assign g5105 = g873;
assign g4888 = g1960;
assign g4887 = g1961;
assign g8561 = g6920;
assign g8562 = g6926;
assign g8563 = g6932;
assign g8564 = g6942;
assign g8565 = g6949;
assign g8566 = g6955;
assign g9451 = g9961;
assign g5816 = g8271;
assign g11489 = 1'b0;

dff g30_reg ( clk, reset, g30, g30 );
dff g31_reg ( clk, reset, g31, g31 );
not U_inv0 ( n4639, g31 );
dff g41_reg ( clk, reset, g41, g41 );
not U_inv1 ( n4638, g41 );
dff g42_reg ( clk, reset, g42, g42 );
not U_inv2 ( n4658, g42 );
dff g43_reg ( clk, reset, g43, g43 );
not U_inv3 ( n4659, g43 );
dff g44_reg ( clk, reset, g44, g44 );
not U_inv4 ( n4660, g44 );
dff g45_reg ( clk, reset, g45, g45 );
not U_inv5 ( n4661, g45 );
dff g46_reg ( clk, reset, g46, g46 );
not U_inv6 ( n4640, g46 );
dff g47_reg ( clk, reset, g47, g47 );
not U_inv7 ( n4662, g47 );
dff g48_reg ( clk, reset, g48, g48 );
not U_inv8 ( n4663, g48 );
dff g82_reg ( clk, reset, g82, g82 );
not U_inv9 ( n4664, g82 );
dff g83_reg ( clk, reset, g83, g83 );
dff g101_reg ( clk, reset, g101, g101 );
dff g102_reg ( clk, reset, g102, g102 );
dff g103_reg ( clk, reset, g103, g103 );
dff g104_reg ( clk, reset, g104, g104 );
dff g28_reg ( clk, reset, g28, g28 );
dff g29_reg ( clk, reset, g29, g29 );
dff g898_reg ( clk, reset, g898, g898 );
not U_inv10 ( n4582, g898 );
dff g901_reg ( clk, reset, g901, g901 );
dff g904_reg ( clk, reset, g904, g904 );
dff g907_reg ( clk, reset, g907, g907 );
dff g910_reg ( clk, reset, g910, g910 );
not U_inv11 ( n4586, g910 );
dff g913_reg ( clk, reset, g913, g913 );
not U_inv12 ( n4572, g913 );
dff g916_reg ( clk, reset, g916, g916 );
not U_inv13 ( n4629, g916 );
dff g919_reg ( clk, reset, g919, g919 );
not U_inv14 ( n4575, g919 );
dff g922_reg ( clk, reset, g922, g922 );
not U_inv15 ( n4581, g922 );
dff g925_reg ( clk, reset, g925, g925 );
dff g886_reg ( clk, reset, g886, g886 );
dff g889_reg ( clk, reset, g889, g889 );
dff g892_reg ( clk, reset, g892, g892 );
not U_inv16 ( n4610, g892 );
dff g895_reg ( clk, reset, g895, g895 );
not U_inv17 ( n4600, g895 );
dff g755_reg ( clk, reset, n596, g83 );
dff g756_reg ( clk, reset, g756, n596 );
dff g746_reg ( clk, reset, g746, g756 );
not U_inv18 ( n4670, g746 );
dff g745_reg ( clk, reset, ex_wire0, g746 );
not U_inv19 ( n4477, ex_wire0 );
dff g750_reg ( clk, reset, ex_wire1, new_g2791_ );
not U_inv20 ( n4671, ex_wire1 );
dff g754_reg ( clk, reset, g4172, new_g3462_ );
dff g794_reg ( clk, reset, g794, new_g5849_ );
not U_inv21 ( n4476, g794 );
dff g798_reg ( clk, reset, g798, new_g6243_ );
not U_inv22 ( n4475, g798 );
dff g802_reg ( clk, reset, g802, new_g5543_ );
not U_inv23 ( n4676, g802 );
dff g806_reg ( clk, reset, g806, new_g6126_ );
not U_inv24 ( n4677, g806 );
dff g810_reg ( clk, reset, g810, new_g6733_ );
not U_inv25 ( n4678, g810 );
dff g814_reg ( clk, reset, g814, new_g7202_ );
not U_inv26 ( n4443, g814 );
dff g818_reg ( clk, reset, g818, new_g7709_ );
not U_inv27 ( n4442, g818 );
dff g822_reg ( clk, reset, g822, new_g8024_ );
not U_inv28 ( n4679, g822 );
dff g826_reg ( clk, reset, g826, new_g8245_ );
not U_inv29 ( n4440, g826 );
dff g829_reg ( clk, reset, n2430, g794 );
dff g833_reg ( clk, reset, n2240, g798 );
dff g837_reg ( clk, reset, ex_wire2, g802 );
not U_inv30 ( n4641, ex_wire2 );
dff g841_reg ( clk, reset, n2239, g806 );
dff g845_reg ( clk, reset, ex_wire3, g810 );
not U_inv31 ( n4561, ex_wire3 );
dff g849_reg ( clk, reset, ex_wire4, g814 );
not U_inv32 ( n4562, ex_wire4 );
dff g853_reg ( clk, reset, ex_wire5, g818 );
not U_inv33 ( n4680, ex_wire5 );
dff g857_reg ( clk, reset, ex_wire6, g822 );
not U_inv34 ( n4563, ex_wire6 );
dff g861_reg ( clk, reset, n2431, g826 );
dff g874_reg ( clk, reset, n765, n2190 );
dff g868_reg ( clk, reset, ex_wire7, n765 );
not U_inv35 ( n4499, ex_wire7 );
dff g875_reg ( clk, reset, n774, n2189 );
dff g869_reg ( clk, reset, ex_wire8, n774 );
not U_inv36 ( n4502, ex_wire8 );
dff g584_reg ( clk, reset, g2610, g101 );
dff g585_reg ( clk, reset, g2611, g102 );
dff g586_reg ( clk, reset, g2612, g103 );
dff g587_reg ( clk, reset, g2602, g104 );
dff g588_reg ( clk, reset, g2603, g28 );
dff g589_reg ( clk, reset, g2604, g29 );
dff g578_reg ( clk, reset, g2601, g101 );
dff g579_reg ( clk, reset, g2605, g102 );
dff g580_reg ( clk, reset, g2606, g103 );
dff g581_reg ( clk, reset, g2607, g104 );
dff g582_reg ( clk, reset, g2608, g28 );
dff g583_reg ( clk, reset, g2609, g29 );
dff g736_reg ( clk, reset, n2456, n1219 );
not U_inv37 ( n4695, n2456 );
dff g731_reg ( clk, reset, n2454, new_g8926_ );
not U_inv38 ( n4435, n2454 );
dff g622_reg ( clk, reset, n2450, new_g8820_ );
not U_inv39 ( n4439, n2450 );
dff g605_reg ( clk, reset, n2265, new_g9150_ );
not U_inv40 ( n4685, n2265 );
dff g599_reg ( clk, reset, n2199, new_g9124_ );
not U_inv41 ( n4684, n2199 );
dff g591_reg ( clk, reset, n2208, new_g9110_ );
not U_inv42 ( n4683, n2208 );
dff g643_reg ( clk, reset, ex_wire9, new_g7441_ );
not U_inv43 ( n4653, ex_wire9 );
dff g650_reg ( clk, reset, ex_wire10, new_g7137_ );
not U_inv44 ( n4654, ex_wire10 );
dff g646_reg ( clk, reset, ex_wire11, new_g7134_ );
not U_inv45 ( n4688, ex_wire11 );
dff g654_reg ( clk, reset, ex_wire12, new_g7660_ );
not U_inv46 ( n4655, ex_wire12 );
dff g664_reg ( clk, reset, n2331, new_g8649_ );
not U_inv47 ( n4652, n2331 );
dff g617_reg ( clk, reset, n2449, new_g8505_ );
not U_inv48 ( n4682, n2449 );
dff g611_reg ( clk, reset, n2245, new_g9721_ );
not U_inv49 ( n4681, n2245 );
dff g631_reg ( clk, reset, ex_wire13, new_g4890_ );
not U_inv50 ( n4483, ex_wire13 );
dff g632_reg ( clk, reset, g632, new_g4891_ );
dff g635_reg ( clk, reset, ex_wire14, n68 );
not U_inv51 ( n4482, ex_wire14 );
dff g627_reg ( clk, reset, n2446, new_g4893_ );
not U_inv52 ( n4686, n2446 );
dff g630_reg ( clk, reset, ex_wire15, new_g6672_ );
not U_inv53 ( n4484, ex_wire15 );
dff g673_reg ( clk, reset, n2249, n1184 );
dff g682_reg ( clk, reset, n2289, n1189 );
dff g691_reg ( clk, reset, n2340, n1194 );
not U_inv54 ( n4651, n2340 );
dff g700_reg ( clk, reset, n2339, n1199 );
not U_inv55 ( n4650, n2339 );
dff g709_reg ( clk, reset, n2288, n1204 );
dff g718_reg ( clk, reset, n2338, n1209 );
not U_inv56 ( n4649, n2338 );
dff g727_reg ( clk, reset, n2330, n1214 );
not U_inv57 ( n4648, n2330 );
dff g639_reg ( clk, reset, n2281, new_g7626_ );
not U_inv58 ( n4687, n2281 );
dff g658_reg ( clk, reset, ex_wire16, new_g8973_ );
not U_inv59 ( n4689, ex_wire16 );
dff g668_reg ( clk, reset, n2305, new_g8922_ );
not U_inv60 ( n4690, n2305 );
dff g677_reg ( clk, reset, n2195, new_g8883_ );
not U_inv61 ( n4691, n2195 );
dff g686_reg ( clk, reset, n2230, new_g8885_ );
not U_inv62 ( n4692, n2230 );
dff g695_reg ( clk, reset, n2312, new_g8887_ );
not U_inv63 ( n4693, n2312 );
dff g704_reg ( clk, reset, n2294, new_g8889_ );
not U_inv64 ( n4437, n2294 );
dff g713_reg ( clk, reset, ex_wire17, new_g8920_ );
not U_inv65 ( n4694, ex_wire17 );
dff g722_reg ( clk, reset, ex_wire18, new_g8923_ );
not U_inv66 ( n4436, ex_wire18 );
dff g17_reg ( clk, reset, g17, new_g4117_ );
dff g49_reg ( clk, reset, g8976, new_g7143_ );
not U_inv67 ( n2444, g8976 );
dff g52_reg ( clk, reset, g8977, new_g6621_ );
not U_inv68 ( n2437, g8977 );
dff g55_reg ( clk, reset, g8978, new_g7183_ );
not U_inv69 ( n2443, g8978 );
dff g58_reg ( clk, reset, g8979, new_g6627_ );
not U_inv70 ( n2436, g8979 );
dff g61_reg ( clk, reset, g8980, new_g7189_ );
not U_inv71 ( n2442, g8980 );
dff g64_reg ( clk, reset, g8981, new_g6638_ );
not U_inv72 ( n2435, g8981 );
dff g67_reg ( clk, reset, g8982, new_g7204_ );
not U_inv73 ( n2441, g8982 );
dff g70_reg ( clk, reset, g8983, new_g6653_ );
not U_inv74 ( n2434, g8983 );
dff g73_reg ( clk, reset, g8984, new_g7219_ );
not U_inv75 ( n2440, g8984 );
dff g76_reg ( clk, reset, g8985, new_g6526_ );
not U_inv76 ( n2439, g8985 );
dff g79_reg ( clk, reset, g8986, new_g6531_ );
not U_inv77 ( n2438, g8986 );
dff g114_reg ( clk, reset, ex_wire19, n1588 );
not U_inv78 ( n4441, ex_wire19 );
dff g940_reg ( clk, reset, ex_wire20, new_g8260_ );
not U_inv79 ( n4669, ex_wire20 );
dff g936_reg ( clk, reset, ex_wire21, new_g8254_ );
not U_inv80 ( n4668, ex_wire21 );
dff g932_reg ( clk, reset, ex_wire22, new_g8250_ );
not U_inv81 ( n4667, ex_wire22 );
dff g928_reg ( clk, reset, ex_wire23, new_g8147_ );
not U_inv82 ( n4666, ex_wire23 );
dff g883_reg ( clk, reset, g2986, new_g3381_ );
dff g882_reg ( clk, reset, ex_wire24, g2986 );
not U_inv83 ( n4531, ex_wire24 );
dff g113_reg ( clk, reset, n1588, n44 );
dff g1955_reg ( clk, reset, n1597, g83 );
dff g1956_reg ( clk, reset, n1601, n1597 );
dff g1957_reg ( clk, reset, n1605, n1601 );
dff g1700_reg ( clk, reset, n2451, n1605 );
not U_inv84 ( n122, n2451 );
dff g1959_reg ( clk, reset, ex_wire25, n122 );
not U_inv85 ( n4485, ex_wire25 );
dff g1710_reg ( clk, reset, g1710, new_g4089_ );
dff g1696_reg ( clk, reset, n2250, new_g5287_ );
not U_inv86 ( n4708, n2250 );
dff g1703_reg ( clk, reset, ex_wire26, new_g5083_ );
not U_inv87 ( n4546, ex_wire26 );
dff g1610_reg ( clk, reset, n2259, new_g5194_ );
not U_inv88 ( n4529, n2259 );
dff g1736_reg ( clk, reset, n1864, new_g5392_ );
dff g1737_reg ( clk, reset, g1737, n1864 );
dff g1765_reg ( clk, reset, g1765, new_g2478_ );
dff g1645_reg ( clk, reset, ex_wire27, new_g10785_ );
not U_inv89 ( n4522, ex_wire27 );
dff g1642_reg ( clk, reset, ex_wire28, new_g10784_ );
not U_inv90 ( n4523, ex_wire28 );
dff g1651_reg ( clk, reset, ex_wire29, new_g10782_ );
not U_inv91 ( n4524, ex_wire29 );
dff g1648_reg ( clk, reset, ex_wire30, new_g10780_ );
not U_inv92 ( n4525, ex_wire30 );
dff g1713_reg ( clk, reset, g1713, new_g5396_ );
not U_inv93 ( n4709, g1713 );
dff g590_reg ( clk, reset, ex_wire31, g1713 );
not U_inv94 ( n4532, ex_wire31 );
dff g758_reg ( clk, reset, g4173, new_g4940_ );
not U_inv95 ( n4672, g4173 );
dff g762_reg ( clk, reset, g4174, new_g5529_ );
not U_inv96 ( n4673, g4174 );
dff g766_reg ( clk, reset, g4175, new_g5536_ );
not U_inv97 ( n4536, g4175 );
dff g770_reg ( clk, reset, g4176, new_g6123_ );
not U_inv98 ( n4674, g4176 );
dff g774_reg ( clk, reset, g4177, new_g6728_ );
not U_inv99 ( n4535, g4177 );
dff g778_reg ( clk, reset, g4178, new_g7191_ );
not U_inv100 ( n4534, g4178 );
dff g782_reg ( clk, reset, g4179, new_g7705_ );
not U_inv101 ( n4675, g4179 );
dff g786_reg ( clk, reset, g4180, new_g8019_ );
not U_inv102 ( n4533, g4180 );
dff g790_reg ( clk, reset, g4181, new_g8244_ );
dff g865_reg ( clk, reset, g2648, n2192 );
dff g1766_reg ( clk, reset, n2218, new_g7133_ );
not U_inv103 ( n4500, n2218 );
dff g1738_reg ( clk, reset, ex_wire32, new_g4231_ );
not U_inv104 ( n4623, ex_wire32 );
dff g1771_reg ( clk, reset, n2241, new_g6502_ );
not U_inv105 ( n4711, n2241 );
dff g1776_reg ( clk, reset, n2270, new_g6508_ );
not U_inv106 ( n4712, n2270 );
dff g1781_reg ( clk, reset, n2198, new_g6516_ );
dff g1747_reg ( clk, reset, n2417, new_g4255_ );
dff g1744_reg ( clk, reset, ex_wire33, new_g4239_ );
not U_inv107 ( n4577, ex_wire33 );
dff g1786_reg ( clk, reset, n2285, new_g6525_ );
not U_inv108 ( n4713, n2285 );
dff g1791_reg ( clk, reset, n2217, new_g6983_ );
dff g1796_reg ( clk, reset, n2200, new_g7541_ );
dff g1756_reg ( clk, reset, ex_wire34, new_g4283_ );
not U_inv109 ( n4594, ex_wire34 );
dff g1753_reg ( clk, reset, n2410, new_g4274_ );
dff g1801_reg ( clk, reset, n2276, new_g7930_ );
not U_inv110 ( n4714, n2276 );
dff g1806_reg ( clk, reset, n2263, new_g8173_ );
not U_inv111 ( n4501, n2263 );
dff g1762_reg ( clk, reset, ex_wire35, new_g4309_ );
not U_inv112 ( n4624, ex_wire35 );
dff g1759_reg ( clk, reset, ex_wire36, new_g4293_ );
not U_inv113 ( n4570, ex_wire36 );
dff g1750_reg ( clk, reset, n2423, new_g4264_ );
dff g1741_reg ( clk, reset, n2398, new_g4238_ );
dff g1718_reg ( clk, reset, n2267, new_g5404_ );
not U_inv114 ( n4710, n2267 );
dff g1707_reg ( clk, reset, n2318, new_g4076_ );
not U_inv115 ( n4486, n2318 );
dff g1690_reg ( clk, reset, n2197, new_g6155_ );
not U_inv116 ( n4730, n2197 );
dff g1958_reg ( clk, reset, g1958, new_g5556_ );
dff g1810_reg ( clk, reset, ex_wire37, g1958 );
not U_inv117 ( g8271, ex_wire37 );
dff g1170_reg ( clk, reset, g1170, g1170 );
not U_inv118 ( n4578, g1170 );
dff g1173_reg ( clk, reset, g1173, g1173 );
not U_inv119 ( n4633, g1173 );
dff g1176_reg ( clk, reset, g1176, g1176 );
not U_inv120 ( n4614, g1176 );
dff g1179_reg ( clk, reset, g1179, g1179 );
not U_inv121 ( n4603, g1179 );
dff g1182_reg ( clk, reset, g1182, g1182 );
not U_inv122 ( n4592, g1182 );
dff g1185_reg ( clk, reset, g1185, g1185 );
not U_inv123 ( n4567, g1185 );
dff g1188_reg ( clk, reset, g1188, g1188 );
dff g1191_reg ( clk, reset, g1191, g1191 );
dff g1194_reg ( clk, reset, g1194, g1194 );
dff g1197_reg ( clk, reset, g1197, g1197 );
not U_inv124 ( n4632, g1197 );
dff g1200_reg ( clk, reset, g1200, g1200 );
not U_inv125 ( n4613, g1200 );
dff g1203_reg ( clk, reset, g1203, g1203 );
not U_inv126 ( n4602, g1203 );
dff g1360_reg ( clk, reset, n2102, n2188 );
dff g1216_reg ( clk, reset, ex_wire38, n2102 );
not U_inv127 ( n4478, ex_wire38 );
dff g1217_reg ( clk, reset, n2111, n2187 );
dff g1212_reg ( clk, reset, ex_wire39, n2111 );
not U_inv128 ( n4487, ex_wire39 );
dff g1357_reg ( clk, reset, ex_wire40, new_g4500_ );
not U_inv129 ( n4526, ex_wire40 );
dff g1289_reg ( clk, reset, ex_wire41, new_g4556_ );
not U_inv130 ( n4545, ex_wire41 );
dff g1231_reg ( clk, reset, n2467, new_g7590_ );
not U_inv131 ( n4542, n2467 );
dff g1218_reg ( clk, reset, n2301, new_g7632_ );
not U_inv132 ( n4541, n2301 );
dff g1223_reg ( clk, reset, ex_wire42, new_g7581_ );
not U_inv133 ( n4735, ex_wire42 );
dff g1227_reg ( clk, reset, ex_wire43, new_g7586_ );
not U_inv134 ( n4543, ex_wire43 );
dff g1117_reg ( clk, reset, ex_wire44, new_g4465_ );
not U_inv135 ( n4494, ex_wire44 );
dff g1121_reg ( clk, reset, n2295, new_g4471_ );
not U_inv136 ( n4736, n2295 );
dff g1125_reg ( clk, reset, ex_wire45, new_g4473_ );
not U_inv137 ( n4737, ex_wire45 );
dff g1129_reg ( clk, reset, ex_wire46, new_g4477_ );
not U_inv138 ( n4495, ex_wire46 );
dff g1133_reg ( clk, reset, ex_wire47, new_g4480_ );
not U_inv139 ( n4738, ex_wire47 );
dff g1137_reg ( clk, reset, ex_wire48, new_g4484_ );
not U_inv140 ( n4739, ex_wire48 );
dff g1141_reg ( clk, reset, ex_wire49, new_g4490_ );
not U_inv141 ( n4488, ex_wire49 );
dff g1145_reg ( clk, reset, ex_wire50, new_g4498_ );
not U_inv142 ( n4489, ex_wire50 );
dff g1113_reg ( clk, reset, ex_wire51, new_g4506_ );
not U_inv143 ( n4740, ex_wire51 );
dff g1166_reg ( clk, reset, ex_wire52, new_g4325_ );
not U_inv144 ( n4491, ex_wire52 );
dff g1163_reg ( clk, reset, n2466, new_g4330_ );
not U_inv145 ( n4490, n2466 );
dff g1160_reg ( clk, reset, n2465, new_g4334_ );
not U_inv146 ( n4493, n2465 );
dff g1157_reg ( clk, reset, ex_wire53, new_g4338_ );
not U_inv147 ( n4492, ex_wire53 );
dff g1153_reg ( clk, reset, n2296, new_g4340_ );
not U_inv148 ( n4741, n2296 );
dff g1149_reg ( clk, reset, n2457, new_g4342_ );
not U_inv149 ( n4742, n2457 );
dff g1101_reg ( clk, reset, n2448, new_g5390_ );
not U_inv150 ( n4743, n2448 );
dff g1104_reg ( clk, reset, n2251, new_g5126_ );
not U_inv151 ( n4744, n2251 );
dff g1107_reg ( clk, reset, n2268, new_g5148_ );
not U_inv152 ( n4745, n2268 );
dff g1110_reg ( clk, reset, ex_wire54, new_g5173_ );
not U_inv153 ( n4746, ex_wire54 );
dff g1639_reg ( clk, reset, n2386, new_g8193_ );
dff g1512_reg ( clk, reset, n2375, new_g8194_ );
dff g1386_reg ( clk, reset, n2468, new_g6833_ );
not U_inv154 ( n4772, n2468 );
dff g201_reg ( clk, reset, n2247, new_g5755_ );
not U_inv155 ( n4497, n2247 );
dff g1374_reg ( clk, reset, n2463, new_g6331_ );
not U_inv156 ( n4752, n2463 );
dff g197_reg ( clk, reset, ex_wire55, new_g6332_ );
not U_inv157 ( n4753, ex_wire55 );
dff g1389_reg ( clk, reset, ex_wire56, new_g6333_ );
not U_inv158 ( n4754, ex_wire56 );
dff g192_reg ( clk, reset, n2319, new_g6334_ );
not U_inv159 ( n4755, n2319 );
dff g1397_reg ( clk, reset, ex_wire57, new_g6838_ );
not U_inv160 ( n4474, ex_wire57 );
dff g248_reg ( clk, reset, n2459, new_g6839_ );
not U_inv161 ( n4512, n2459 );
dff g1400_reg ( clk, reset, ex_wire58, new_g6840_ );
not U_inv162 ( n4756, ex_wire58 );
dff g243_reg ( clk, reset, n2458, new_g6841_ );
not U_inv163 ( n4757, n2458 );
dff g1362_reg ( clk, reset, n2464, new_g6819_ );
not U_inv164 ( n4758, n2464 );
dff g237_reg ( clk, reset, ex_wire59, new_g6820_ );
not U_inv165 ( n4759, ex_wire59 );
dff g1365_reg ( clk, reset, ex_wire60, new_g6821_ );
not U_inv166 ( n4760, ex_wire60 );
dff g231_reg ( clk, reset, n2321, new_g6834_ );
not U_inv167 ( n4761, n2321 );
dff g1368_reg ( clk, reset, ex_wire61, new_g6822_ );
not U_inv168 ( n4762, ex_wire61 );
dff g225_reg ( clk, reset, ex_wire62, new_g6823_ );
not U_inv169 ( n4763, ex_wire62 );
dff g1371_reg ( clk, reset, n2461, new_g6826_ );
not U_inv170 ( n4764, n2461 );
dff g219_reg ( clk, reset, ex_wire63, new_g6824_ );
not U_inv171 ( n4765, ex_wire63 );
dff g1377_reg ( clk, reset, ex_wire64, new_g6827_ );
not U_inv172 ( n4766, ex_wire64 );
dff g213_reg ( clk, reset, n2320, new_g6828_ );
not U_inv173 ( n4767, n2320 );
dff g1380_reg ( clk, reset, ex_wire65, new_g6829_ );
not U_inv174 ( n4768, ex_wire65 );
dff g207_reg ( clk, reset, ex_wire66, new_g6830_ );
not U_inv175 ( n4769, ex_wire66 );
dff g1383_reg ( clk, reset, n2462, new_g6831_ );
not U_inv176 ( n4770, n2462 );
dff g186_reg ( clk, reset, ex_wire67, new_g6832_ );
not U_inv177 ( n4771, ex_wire67 );
dff g1615_reg ( clk, reset, n2384, new_g8770_ );
dff g1621_reg ( clk, reset, n2382, new_g8771_ );
dff g1624_reg ( clk, reset, n2380, new_g8773_ );
dff g1627_reg ( clk, reset, n2390, new_g8774_ );
dff g1630_reg ( clk, reset, n2396, new_g8776_ );
dff g1633_reg ( clk, reset, n2394, new_g8777_ );
dff g1636_reg ( clk, reset, n2377, new_g8779_ );
dff g1393_reg ( clk, reset, ex_wire68, new_g6163_ );
not U_inv178 ( n4449, ex_wire68 );
dff g115_reg ( clk, reset, n2460, new_g6179_ );
not U_inv179 ( n4657, n2460 );
dff g1394_reg ( clk, reset, ex_wire69, new_g6747_ );
not U_inv180 ( n4470, ex_wire69 );
dff g119_reg ( clk, reset, n2317, N41 );
not U_inv181 ( n4656, n2317 );
dff g12_reg ( clk, reset, n2328, new_g5445_ );
not U_inv182 ( n4773, n2328 );
dff g9_reg ( clk, reset, n2426, new_g5421_ );
dff g549_reg ( clk, reset, n2374, new_g10855_ );
dff g255_reg ( clk, reset, g255, new_g6049_ );
not U_inv183 ( n4438, g255 );
dff g312_reg ( clk, reset, ex_wire70, g255 );
not U_inv184 ( n4521, ex_wire70 );
dff g636_reg ( clk, reset, g636, new_g8631_ );
dff g8_reg ( clk, reset, g8, g636 );
dff g139_reg ( clk, reset, n2222, new_g8049_ );
dff g296_reg ( clk, reset, n2414, new_g6916_ );
dff g36_reg ( clk, reset, ex_wire71, new_g10722_ );
not U_inv185 ( n4608, ex_wire71 );
dff g1681_reg ( clk, reset, n2367, new_g10864_ );
dff g560_reg ( clk, reset, n2381, new_g10797_ );
dff g258_reg ( clk, reset, g258, new_g6015_ );
dff g321_reg ( clk, reset, ex_wire72, g258 );
not U_inv186 ( n4515, ex_wire72 );
dff g1811_reg ( clk, reset, n2447, new_g10936_ );
dff g1618_reg ( clk, reset, n2388, new_g11579_ );
dff g1499_reg ( clk, reset, n2316, new_g8041_ );
not U_inv187 ( n4472, n2316 );
dff g1531_reg ( clk, reset, ex_wire73, new_g6528_ );
not U_inv188 ( n4618, ex_wire73 );
dff g1504_reg ( clk, reset, ex_wire74, new_g6198_ );
not U_inv189 ( n4469, ex_wire74 );
dff g1528_reg ( clk, reset, n2422, new_g6522_ );
dff g1508_reg ( clk, reset, ex_wire75, n192 );
not U_inv190 ( n4473, ex_wire75 );
dff g1524_reg ( clk, reset, n2407, new_g6513_ );
dff g1453_reg ( clk, reset, n2452, new_g5770_ );
not U_inv191 ( n4749, n2452 );
dff g1458_reg ( clk, reset, n2323, new_g6180_ );
not U_inv192 ( n4451, n2323 );
dff g1462_reg ( clk, reset, ex_wire76, new_g8042_ );
not U_inv193 ( n4452, ex_wire76 );
dff g1466_reg ( clk, reset, n2324, new_g8045_ );
not U_inv194 ( n4453, n2324 );
dff g1470_reg ( clk, reset, ex_wire77, new_g8051_ );
not U_inv195 ( n4750, ex_wire77 );
dff g1474_reg ( clk, reset, ex_wire78, new_g8039_ );
not U_inv196 ( n4455, ex_wire78 );
dff g1478_reg ( clk, reset, ex_wire79, new_g8040_ );
not U_inv197 ( n4450, ex_wire79 );
dff g1482_reg ( clk, reset, n2224, new_g8043_ );
dff g1486_reg ( clk, reset, n2225, new_g8046_ );
dff g1490_reg ( clk, reset, ex_wire80, new_g8052_ );
not U_inv198 ( n4751, ex_wire80 );
dff g1494_reg ( clk, reset, n2252, new_g8055_ );
not U_inv199 ( n4471, n2252 );
dff g1534_reg ( clk, reset, ex_wire81, new_g6533_ );
not U_inv200 ( n4607, ex_wire81 );
dff g1537_reg ( clk, reset, ex_wire82, new_g6537_ );
not U_inv201 ( n4591, ex_wire82 );
dff g1540_reg ( clk, reset, n2416, new_g6541_ );
dff g1543_reg ( clk, reset, ex_wire83, new_g6545_ );
not U_inv202 ( n4627, ex_wire83 );
dff g1546_reg ( clk, reset, n2400, new_g6551_ );
dff g1549_reg ( clk, reset, ex_wire84, new_g6523_ );
not U_inv203 ( n4579, ex_wire84 );
dff g1552_reg ( clk, reset, ex_wire85, new_g6529_ );
not U_inv204 ( n4637, ex_wire85 );
dff g1555_reg ( clk, reset, ex_wire86, new_g6534_ );
not U_inv205 ( n4617, ex_wire86 );
dff g1558_reg ( clk, reset, ex_wire87, new_g6538_ );
not U_inv206 ( n4606, ex_wire87 );
dff g4_reg ( clk, reset, n2418, new_g6656_ );
dff g1561_reg ( clk, reset, ex_wire88, new_g6542_ );
not U_inv207 ( n4587, ex_wire88 );
dff g1564_reg ( clk, reset, ex_wire89, new_g6546_ );
not U_inv208 ( n4565, ex_wire89 );
dff g1448_reg ( clk, reset, n2254, new_g11514_ );
not U_inv209 ( n4498, n2254 );
dff g1444_reg ( clk, reset, ex_wire90, new_g8766_ );
not U_inv210 ( n4456, ex_wire90 );
dff g1440_reg ( clk, reset, ex_wire91, new_g8768_ );
not U_inv211 ( n4457, ex_wire91 );
dff g1436_reg ( clk, reset, ex_wire92, new_g8772_ );
not U_inv212 ( n4458, ex_wire92 );
dff g1432_reg ( clk, reset, ex_wire93, new_g8775_ );
not U_inv213 ( n4459, ex_wire93 );
dff g1403_reg ( clk, reset, ex_wire94, new_g8765_ );
not U_inv214 ( n4460, ex_wire94 );
dff g1428_reg ( clk, reset, ex_wire95, new_g8767_ );
not U_inv215 ( n4454, ex_wire95 );
dff g1407_reg ( clk, reset, n2341, new_g8769_ );
not U_inv216 ( n4468, n2341 );
dff g1586_reg ( clk, reset, n2409, new_g6514_ );
dff g1424_reg ( clk, reset, ex_wire96, new_g6216_ );
not U_inv217 ( n4466, ex_wire96 );
dff g1583_reg ( clk, reset, ex_wire97, new_g6506_ );
not U_inv218 ( n4571, ex_wire97 );
dff g1411_reg ( clk, reset, ex_wire98, n186 );
not U_inv219 ( n4465, ex_wire98 );
dff g1580_reg ( clk, reset, ex_wire99, new_g6500_ );
not U_inv220 ( n4590, ex_wire99 );
dff g1419_reg ( clk, reset, n2226, new_g6244_ );
not U_inv221 ( n4747, n2226 );
dff g1515_reg ( clk, reset, n2277, new_g6193_ );
not U_inv222 ( n4748, n2277 );
dff g1520_reg ( clk, reset, ex_wire100, new_g6205_ );
not U_inv223 ( n4467, ex_wire100 );
dff g1571_reg ( clk, reset, n2421, new_g6469_ );
dff g1415_reg ( clk, reset, n2238, new_g6224_ );
not U_inv224 ( n4496, n2238 );
dff g1567_reg ( clk, reset, n2406, new_g6468_ );
dff g1574_reg ( clk, reset, ex_wire101, new_g6478_ );
not U_inv225 ( n4620, ex_wire101 );
dff g1577_reg ( clk, reset, ex_wire102, new_g6480_ );
not U_inv226 ( n4609, ex_wire102 );
dff g1589_reg ( clk, reset, n2399, new_g6524_ );
dff g1592_reg ( clk, reset, ex_wire103, new_g6470_ );
not U_inv227 ( n4580, ex_wire103 );
dff g1595_reg ( clk, reset, ex_wire104, new_g6479_ );
not U_inv228 ( n4636, ex_wire104 );
dff g1598_reg ( clk, reset, ex_wire105, new_g6481_ );
not U_inv229 ( n4616, ex_wire105 );
dff g1601_reg ( clk, reset, ex_wire106, new_g6501_ );
not U_inv230 ( n4605, ex_wire106 );
dff g1604_reg ( clk, reset, ex_wire107, new_g6507_ );
not U_inv231 ( n4597, ex_wire107 );
dff g1_reg ( clk, reset, n2427, new_g6679_ );
dff g1607_reg ( clk, reset, ex_wire108, new_g6515_ );
not U_inv232 ( n4568, ex_wire108 );
dff g38_reg ( clk, reset, g38, new_g10726_ );
dff g566_reg ( clk, reset, n2378, new_g10799_ );
dff g260_reg ( clk, reset, g260, new_g6035_ );
dff g327_reg ( clk, reset, ex_wire109, g260 );
not U_inv233 ( n4513, ex_wire109 );
dff g1687_reg ( clk, reset, n2389, new_g10776_ );
dff g369_reg ( clk, reset, ex_wire110, new_g11320_ );
not U_inv234 ( n4559, ex_wire110 );
dff g374_reg ( clk, reset, n2302, new_g11290_ );
not U_inv235 ( n4558, n2302 );
dff g378_reg ( clk, reset, ex_wire111, new_g11291_ );
not U_inv236 ( n4707, ex_wire111 );
dff g382_reg ( clk, reset, n2469, new_g11292_ );
not U_inv237 ( n4560, n2469 );
dff g456_reg ( clk, reset, n2433, new_g11340_ );
not U_inv238 ( n4700, n2433 );
dff g461_reg ( clk, reset, n2203, new_g11372_ );
not U_inv239 ( n4701, n2203 );
dff g466_reg ( clk, reset, n2262, new_g11376_ );
not U_inv240 ( n4702, n2262 );
dff g471_reg ( clk, reset, n2246, new_g11380_ );
not U_inv241 ( n4703, n2246 );
dff g481_reg ( clk, reset, n2310, n1234 );
not U_inv242 ( n4644, n2310 );
dff g486_reg ( clk, reset, n2283, n1239 );
not U_inv243 ( n4645, n2283 );
dff g491_reg ( clk, reset, n2232, n1244 );
not U_inv244 ( n4696, n2232 );
dff g354_reg ( clk, reset, n2361, new_g11483_ );
dff g1086_reg ( clk, reset, n2348, new_g6071_ );
dff g1003_reg ( clk, reset, n2300, new_g6902_ );
not U_inv245 ( n4503, n2300 );
dff g496_reg ( clk, reset, n2231, n1249 );
not U_inv246 ( n4646, n2231 );
dff g501_reg ( clk, reset, n2284, n1254 );
not U_inv247 ( n4647, n2284 );
dff g360_reg ( clk, reset, n2359, new_g11485_ );
dff g1092_reg ( clk, reset, n2346, new_g6088_ );
dff g1011_reg ( clk, reset, n2299, new_g6912_ );
not U_inv248 ( n4505, n2299 );
dff g506_reg ( clk, reset, n2215, n1259 );
dff g511_reg ( clk, reset, n2309, n1264 );
not U_inv249 ( n4642, n2309 );
dff g516_reg ( clk, reset, n2216, n1269 );
dff g476_reg ( clk, reset, n2275, n1274 );
not U_inv250 ( n4697, n2275 );
dff g339_reg ( clk, reset, n2364, new_g11478_ );
dff g1071_reg ( clk, reset, n2353, new_g5910_ );
dff g1023_reg ( clk, reset, ex_wire112, new_g7244_ );
not U_inv251 ( n4511, ex_wire112 );
dff g542_reg ( clk, reset, n2334, n1279 );
not U_inv252 ( n4643, n2334 );
dff g538_reg ( clk, reset, n2280, n1284 );
dff g534_reg ( clk, reset, n2236, n1289 );
dff g530_reg ( clk, reset, n2293, n1294 );
dff g525_reg ( clk, reset, n2315, n1299 );
not U_inv253 ( n4698, n2315 );
dff g521_reg ( clk, reset, n2329, n1304 );
not U_inv254 ( n4699, n2329 );
dff g345_reg ( clk, reset, n2355, new_g11625_ );
dff g1077_reg ( clk, reset, n2352, new_g5914_ );
dff g1032_reg ( clk, reset, n2432, new_g7257_ );
dff g1275_reg ( clk, reset, n2211, n2136 );
dff g1235_reg ( clk, reset, n2205, n2141 );
dff g1240_reg ( clk, reset, n2307, n2146 );
not U_inv255 ( n4539, n2307 );
dff g1245_reg ( clk, reset, n2209, n2151 );
dff g1250_reg ( clk, reset, n2272, n2156 );
not U_inv256 ( n4732, n2272 );
dff g1255_reg ( clk, reset, n2271, n2161 );
not U_inv257 ( n4540, n2271 );
dff g1260_reg ( clk, reset, n2243, n2166 );
dff g1265_reg ( clk, reset, n2210, n2171 );
dff g1270_reg ( clk, reset, n2255, n2176 );
not U_inv258 ( n4537, n2255 );
dff g108_reg ( clk, reset, g108, new_g11561_ );
dff g1336_reg ( clk, reset, n2219, new_g11636_ );
dff g1341_reg ( clk, reset, n2229, new_g11639_ );
not U_inv259 ( n4731, n2229 );
dff g1206_reg ( clk, reset, g3069, new_g4114_ );
dff g1361_reg ( clk, reset, ex_wire113, g3069 );
not U_inv260 ( n4528, ex_wire113 );
dff g1356_reg ( clk, reset, n2235, new_g5763_ );
dff g1317_reg ( clk, reset, g1317, n2235 );
dff g1346_reg ( clk, reset, n2311, new_g11640_ );
not U_inv261 ( n4612, n2311 );
dff g1351_reg ( clk, reset, n2266, new_g11641_ );
dff g1333_reg ( clk, reset, ex_wire114, new_g11610_ );
not U_inv262 ( n4625, ex_wire114 );
dff g1330_reg ( clk, reset, ex_wire115, new_g11609_ );
not U_inv263 ( n4566, ex_wire115 );
dff g1327_reg ( clk, reset, ex_wire116, new_g11608_ );
not U_inv264 ( n4593, ex_wire116 );
dff g1324_reg ( clk, reset, ex_wire117, new_g11607_ );
not U_inv265 ( n4604, ex_wire117 );
dff g1321_reg ( clk, reset, ex_wire118, new_g11606_ );
not U_inv266 ( n4615, ex_wire118 );
dff g1318_reg ( clk, reset, n2419, new_g11605_ );
dff g1314_reg ( clk, reset, n2404, new_g11604_ );
dff g1311_reg ( clk, reset, ex_wire119, new_g11603_ );
not U_inv267 ( n4574, ex_wire119 );
dff g1308_reg ( clk, reset, ex_wire120, new_g11602_ );
not U_inv268 ( n4622, ex_wire120 );
dff g39_reg ( clk, reset, ex_wire121, new_g10663_ );
not U_inv269 ( n4626, ex_wire121 );
dff g1654_reg ( clk, reset, n2392, new_g10765_ );
dff g569_reg ( clk, reset, n2395, new_g10717_ );
dff g261_reg ( clk, reset, g261, new_g6038_ );
dff g330_reg ( clk, reset, ex_wire122, g261 );
not U_inv270 ( n4519, ex_wire122 );
dff g363_reg ( clk, reset, n2358, new_g11486_ );
dff g1095_reg ( clk, reset, n2345, new_g6093_ );
dff g1007_reg ( clk, reset, ex_wire123, new_g6918_ );
not U_inv271 ( n4504, ex_wire123 );
dff g1857_reg ( clk, reset, n2282, new_g11294_ );
not U_inv272 ( n4720, n2282 );
dff g1814_reg ( clk, reset, n2220, new_g9266_ );
not U_inv273 ( n4717, n2220 );
dff g1828_reg ( clk, reset, n2253, new_g9272_ );
not U_inv274 ( n4718, n2253 );
dff g1822_reg ( clk, reset, n2202, new_g9269_ );
not U_inv275 ( n4550, n2202 );
dff g16_reg ( clk, reset, ex_wire124, new_g3524_ );
not U_inv276 ( n4599, ex_wire124 );
dff g1853_reg ( clk, reset, ex_wire125, new_g4904_ );
not U_inv277 ( n4479, ex_wire125 );
dff g1845_reg ( clk, reset, n2445, new_g4905_ );
not U_inv278 ( n4719, n2445 );
dff g1848_reg ( clk, reset, ex_wire126, new_g6755_ );
not U_inv279 ( n4481, ex_wire126 );
dff g1849_reg ( clk, reset, ex_wire127, new_g4902_ );
not U_inv280 ( n4480, ex_wire127 );
dff g1850_reg ( clk, reset, g1850, new_g4903_ );
dff g1864_reg ( clk, reset, ex_wire128, new_g6795_ );
not U_inv281 ( n4721, ex_wire128 );
dff g1861_reg ( clk, reset, ex_wire129, new_g6471_ );
not U_inv282 ( n4552, ex_wire129 );
dff g1868_reg ( clk, reset, ex_wire130, new_g6909_ );
not U_inv283 ( n4553, ex_wire130 );
dff g1878_reg ( clk, reset, n2326, new_g8559_ );
not U_inv284 ( n4551, n2326 );
dff g1887_reg ( clk, reset, n2248, n1810 );
dff g1896_reg ( clk, reset, n2287, n1815 );
dff g1905_reg ( clk, reset, n2337, n1820 );
not U_inv285 ( n4549, n2337 );
dff g1914_reg ( clk, reset, n2336, n1825 );
not U_inv286 ( n4548, n2336 );
dff g1923_reg ( clk, reset, n2286, n1830 );
dff g1932_reg ( clk, reset, n2335, n1835 );
not U_inv287 ( n4547, n2335 );
dff g1941_reg ( clk, reset, n2291, n1840 );
dff g1950_reg ( clk, reset, n2455, n1845 );
not U_inv288 ( n4729, n2455 );
dff g1840_reg ( clk, reset, n2303, new_g8384_ );
not U_inv289 ( n4716, n2303 );
dff g1834_reg ( clk, reset, ex_wire131, new_g9555_ );
not U_inv290 ( n4715, ex_wire131 );
dff g1872_reg ( clk, reset, n2204, new_g8921_ );
not U_inv291 ( n4722, n2204 );
dff g1882_reg ( clk, reset, n2269, new_g8943_ );
not U_inv292 ( n4723, n2269 );
dff g1891_reg ( clk, reset, n2194, new_g8937_ );
not U_inv293 ( n4724, n2194 );
dff g1900_reg ( clk, reset, n2237, new_g8938_ );
not U_inv294 ( n4725, n2237 );
dff g1909_reg ( clk, reset, n2304, new_g8939_ );
not U_inv295 ( n4726, n2304 );
dff g1918_reg ( clk, reset, n2242, new_g8940_ );
not U_inv296 ( n4434, n2242 );
dff g1927_reg ( clk, reset, ex_wire132, new_g8941_ );
not U_inv297 ( n4727, ex_wire132 );
dff g1936_reg ( clk, reset, n2297, new_g8944_ );
not U_inv298 ( n4433, n2297 );
dff g1945_reg ( clk, reset, n2453, new_g8945_ );
not U_inv299 ( n4728, n2453 );
dff g1854_reg ( clk, reset, g1854, new_g11293_ );
dff g7_reg ( clk, reset, ex_wire133, g1854 );
not U_inv300 ( n4596, ex_wire133 );
dff g37_reg ( clk, reset, ex_wire134, n7 );
not U_inv301 ( n4589, ex_wire134 );
dff g1684_reg ( clk, reset, n2365, new_g10866_ );
dff g563_reg ( clk, reset, n2379, new_g10798_ );
dff g259_reg ( clk, reset, g259, new_g6026_ );
dff g324_reg ( clk, reset, ex_wire135, g259 );
not U_inv302 ( n4517, ex_wire135 );
dff g357_reg ( clk, reset, n2360, new_g11484_ );
dff g1089_reg ( clk, reset, n2347, new_g6080_ );
dff g999_reg ( clk, reset, ex_wire136, new_g6908_ );
not U_inv303 ( n4510, ex_wire136 );
dff g174_reg ( clk, reset, ex_wire137, new_g8050_ );
not U_inv304 ( n4445, ex_wire137 );
dff g162_reg ( clk, reset, n2221, new_g8054_ );
dff g278_reg ( clk, reset, n2415, new_g6922_ );
dff g123_reg ( clk, reset, n2403, new_g7032_ );
dff g33_reg ( clk, reset, ex_wire138, new_g10719_ );
not U_inv305 ( n4583, ex_wire138 );
dff g1660_reg ( clk, reset, n2372, new_g10859_ );
dff g575_reg ( clk, reset, n2376, new_g10800_ );
dff g254_reg ( clk, reset, g254, new_g6045_ );
dff g309_reg ( clk, reset, ex_wire139, g254 );
not U_inv306 ( n4520, ex_wire139 );
dff g342_reg ( clk, reset, n2356, new_g11488_ );
dff g1074_reg ( clk, reset, n2343, new_g6099_ );
dff g1015_reg ( clk, reset, ex_wire140, new_g6930_ );
not U_inv307 ( n4506, ex_wire140 );
dff g135_reg ( clk, reset, n2260, new_g8053_ );
dff g293_reg ( clk, reset, n2429, new_g6911_ );
dff g1672_reg ( clk, reset, n2373, new_g10858_ );
dff g546_reg ( clk, reset, n2387, new_g10791_ );
dff g253_reg ( clk, reset, g253, new_g5996_ );
dff g305_reg ( clk, reset, n2258, g253 );
dff g426_reg ( clk, reset, n2214, n1379 );
dff g386_reg ( clk, reset, n2207, n1384 );
dff g391_reg ( clk, reset, n2308, n1389 );
not U_inv308 ( n4556, n2308 );
dff g396_reg ( clk, reset, n2212, n1394 );
dff g401_reg ( clk, reset, n2274, n1399 );
not U_inv309 ( n4704, n2274 );
dff g406_reg ( clk, reset, n2273, n1404 );
not U_inv310 ( n4557, n2273 );
dff g411_reg ( clk, reset, n2244, n1409 );
dff g416_reg ( clk, reset, n2213, n1414 );
dff g421_reg ( clk, reset, n2256, n1419 );
not U_inv311 ( n4554, n2256 );
dff g452_reg ( clk, reset, n2333, n1424 );
not U_inv312 ( n4555, n2333 );
dff g448_reg ( clk, reset, n2279, n1429 );
dff g444_reg ( clk, reset, n2234, n1434 );
dff g440_reg ( clk, reset, n2292, n1439 );
dff g435_reg ( clk, reset, n2314, n1444 );
not U_inv313 ( n4705, n2314 );
dff g431_reg ( clk, reset, n2327, n1449 );
not U_inv314 ( n4706, n2327 );
dff g148_reg ( clk, reset, n2306, new_g8048_ );
not U_inv315 ( n4462, n2306 );
dff g269_reg ( clk, reset, n2428, new_g6906_ );
dff g178_reg ( clk, reset, ex_wire141, new_g6759_ );
not U_inv316 ( n4448, ex_wire141 );
dff g266_reg ( clk, reset, n2420, new_g6900_ );
dff g34_reg ( clk, reset, ex_wire142, new_g10720_ );
not U_inv317 ( n4635, ex_wire142 );
dff g1675_reg ( clk, reset, n2371, new_g10860_ );
dff g554_reg ( clk, reset, n2385, new_g10793_ );
dff g256_reg ( clk, reset, g256, new_g6000_ );
dff g315_reg ( clk, reset, ex_wire143, g256 );
not U_inv318 ( n4516, ex_wire143 );
dff g348_reg ( clk, reset, n2363, new_g11481_ );
dff g1080_reg ( clk, reset, n2350, new_g6059_ );
dff g995_reg ( clk, reset, ex_wire144, new_g6895_ );
not U_inv319 ( n4509, ex_wire144 );
dff g757_reg ( clk, reset, g757, new_g10788_ );
dff g971_reg ( clk, reset, n2264, new_g11349_ );
not U_inv320 ( n4576, n2264 );
dff g976_reg ( clk, reset, n2322, new_g11391_ );
not U_inv321 ( n4665, n2322 );
dff g878_reg ( clk, reset, g3007, new_g3506_ );
dff g876_reg ( clk, reset, ex_wire145, g3007 );
not U_inv322 ( n4530, ex_wire145 );
dff g981_reg ( clk, reset, n2227, new_g11392_ );
not U_inv323 ( n4611, n2227 );
dff g986_reg ( clk, reset, ex_wire146, new_g11393_ );
not U_inv324 ( n4601, ex_wire146 );
dff g968_reg ( clk, reset, ex_wire147, new_g11314_ );
not U_inv325 ( n4621, ex_wire147 );
dff g965_reg ( clk, reset, ex_wire148, new_g11312_ );
not U_inv326 ( n4569, ex_wire148 );
dff g962_reg ( clk, reset, ex_wire149, new_g11310_ );
not U_inv327 ( n4598, ex_wire149 );
dff g959_reg ( clk, reset, n2412, new_g11308_ );
dff g956_reg ( clk, reset, n2425, new_g11306_ );
dff g35_reg ( clk, reset, ex_wire150, new_g10721_ );
not U_inv328 ( n4619, ex_wire150 );
dff g1666_reg ( clk, reset, n2368, new_g10863_ );
dff g1678_reg ( clk, reset, n2369, new_g10862_ );
dff g557_reg ( clk, reset, n2383, new_g10795_ );
dff g257_reg ( clk, reset, g257, new_g6002_ );
dff g318_reg ( clk, reset, ex_wire151, g257 );
not U_inv329 ( n4514, ex_wire151 );
dff g351_reg ( clk, reset, n2362, new_g11482_ );
dff g1083_reg ( clk, reset, n2349, new_g6068_ );
dff g991_reg ( clk, reset, ex_wire152, new_g6898_ );
not U_inv330 ( n4508, ex_wire152 );
dff g158_reg ( clk, reset, ex_wire153, new_g8060_ );
not U_inv331 ( n4447, ex_wire153 );
dff g275_reg ( clk, reset, ex_wire154, new_g6915_ );
not U_inv332 ( n4585, ex_wire154 );
dff g1727_reg ( clk, reset, n2424, new_g10773_ );
dff g953_reg ( clk, reset, ex_wire155, new_g11305_ );
not U_inv333 ( n4630, ex_wire155 );
dff g950_reg ( clk, reset, n2401, new_g11303_ );
dff g947_reg ( clk, reset, ex_wire156, new_g11300_ );
not U_inv334 ( n4573, ex_wire156 );
dff g40_reg ( clk, reset, g40, new_g10664_ );
dff g1657_reg ( clk, reset, n2391, new_g10767_ );
dff g572_reg ( clk, reset, n2393, new_g10718_ );
dff g262_reg ( clk, reset, g262, new_g6042_ );
dff g333_reg ( clk, reset, ex_wire157, g262 );
not U_inv335 ( n4518, ex_wire157 );
dff g336_reg ( clk, reset, n2354, new_g11647_ );
dff g1068_reg ( clk, reset, n2351, new_g6054_ );
dff g1027_reg ( clk, reset, n2298, new_g6894_ );
not U_inv336 ( n4544, n2298 );
dff g366_reg ( clk, reset, n2357, new_g11487_ );
dff g1098_reg ( clk, reset, n2344, new_g6096_ );
dff g1019_reg ( clk, reset, ex_wire158, new_g6924_ );
not U_inv337 ( n4507, ex_wire158 );
dff g105_reg ( clk, reset, n2342, new_g10898_ );
dff g131_reg ( clk, reset, n2261, new_g8059_ );
dff g127_reg ( clk, reset, n2223, new_g8044_ );
dff g170_reg ( clk, reset, ex_wire159, new_g8047_ );
not U_inv338 ( n4444, ex_wire159 );
dff g284_reg ( clk, reset, n2397, new_g6934_ );
dff g287_reg ( clk, reset, ex_wire160, new_g6901_ );
not U_inv339 ( n4584, ex_wire160 );
dff g290_reg ( clk, reset, ex_wire161, new_g6907_ );
not U_inv340 ( n4634, ex_wire161 );
dff g944_reg ( clk, reset, n2408, new_g11298_ );
dff g153_reg ( clk, reset, n2257, new_g7843_ );
not U_inv341 ( n4463, n2257 );
dff g272_reg ( clk, reset, n2413, new_g6910_ );
dff g32_reg ( clk, reset, ex_wire162, n3 );
not U_inv342 ( n4527, ex_wire162 );
dff g1663_reg ( clk, reset, n2370, new_g10861_ );
dff g1724_reg ( clk, reset, ex_wire163, new_g10771_ );
not U_inv343 ( n4631, ex_wire163 );
dff g182_reg ( clk, reset, ex_wire164, new_g6786_ );
not U_inv344 ( n4464, ex_wire164 );
dff g263_reg ( clk, reset, n2405, new_g6897_ );
dff g143_reg ( clk, reset, n2228, new_g6439_ );
not U_inv345 ( n4461, n2228 );
dff g302_reg ( clk, reset, ex_wire165, new_g6929_ );
not U_inv346 ( n4564, ex_wire165 );
dff g166_reg ( clk, reset, ex_wire166, new_g6757_ );
not U_inv347 ( n4446, ex_wire166 );
dff g299_reg ( clk, reset, ex_wire167, new_g6923_ );
not U_inv348 ( n4588, ex_wire167 );
dff g1721_reg ( clk, reset, n2402, new_g10770_ );
dff g281_reg ( clk, reset, ex_wire168, new_g6928_ );
not U_inv349 ( n4628, ex_wire168 );
dff g1733_reg ( clk, reset, ex_wire169, new_g10711_ );
not U_inv350 ( n4595, ex_wire169 );
dff g1304_reg ( clk, reset, n2332, n2181 );
not U_inv351 ( n4538, n2332 );
dff g1300_reg ( clk, reset, n2278, n2186 );
dff g1296_reg ( clk, reset, n2233, n2191 );
dff g1292_reg ( clk, reset, n2290, n2196 );
dff g1284_reg ( clk, reset, n2313, n2201 );
not U_inv352 ( n4733, n2313 );
dff g1280_reg ( clk, reset, n2325, n2206 );
not U_inv353 ( n4734, n2325 );
dff g1669_reg ( clk, reset, n2366, new_g10865_ );
dff g1730_reg ( clk, reset, n2411, new_g10707_ );
nor U2611 ( n3849, n2784, n3850 );
not U2612 ( n2784, g109 );
not U2613 ( n2775, n2774 );
nand U2614 ( n2774, n4546, n4708 );
nand U2615 ( n3107, g109, n3082 );
nor U2616 ( n3196, n2250, n4546 );
nor U2617 ( n3101, g4172, n4671 );
not U2618 ( n2472, g18 );
not U2619 ( n3389, n3391 );
nand U2620 ( n3391, n4017, n4018 );
nand U2621 ( g9961, n2470, n4639 );
nor U2622 ( n2470, n2471, g30 );
nor U2623 ( new_g9721_, n2472, n2473 );
xnor U2624 ( n2473, n2245, n2474 );
nor U2625 ( n2474, n2475, n2476 );
nor U2626 ( n2475, n2449, n2477 );
nand U2627 ( n2477, n2478, n2479 );
nand U2628 ( n2478, n2480, n2481 );
nor U2629 ( new_g9555_, n2482, n2472 );
nor U2630 ( n2482, n2483, n2484 );
nor U2631 ( n2483, n4715, n2485 );
nor U2632 ( n2485, n2486, n2487 );
nor U2633 ( n2486, n2488, n2303 );
nor U2634 ( n2488, n2489, n2490 );
nor U2635 ( new_g9272_, n2491, n2472 );
xnor U2636 ( n2491, n2492, n2253 );
nand U2637 ( n2492, n2493, n2494 );
nand U2638 ( n2494, n2489, n2495 );
nand U2639 ( n2495, n2496, n2497 );
nand U2640 ( n2497, n2498, n2202 );
nand U2641 ( n2498, n2499, n2500 );
nor U2642 ( new_g9269_, n2472, n2501 );
xnor U2643 ( n2501, n4550, n2502 );
nand U2644 ( n2502, n2503, n2489 );
nor U2645 ( n2503, n2504, n2505 );
nor U2646 ( n2505, n4550, n4718 );
not U2647 ( n2504, n2506 );
nor U2648 ( new_g9266_, n2472, n2507 );
xnor U2649 ( n2507, n4717, n2508 );
nand U2650 ( n2508, n2489, n2509 );
nand U2651 ( n2509, n2510, n2490 );
nor U2652 ( n2510, n2511, n2512 );
nor U2653 ( n2512, n2202, n2499 );
nor U2654 ( n2511, n4550, n2220 );
nor U2655 ( new_g9150_, n2513, n2472 );
xnor U2656 ( n2513, n4685, n2514 );
nor U2657 ( n2514, n2515, n2516 );
nand U2658 ( n2516, n2479, n2517 );
nor U2659 ( n2515, n2518, n2481 );
nor U2660 ( n2518, n2519, n2520 );
nor U2661 ( n2519, n4684, n2521 );
nor U2662 ( n2521, n2522, n2523 );
nor U2663 ( new_g9124_, n2472, n2524 );
xnor U2664 ( n2524, n2199, n2525 );
nor U2665 ( n2525, n2481, n2526 );
nand U2666 ( n2526, n2527, n2528 );
nand U2667 ( n2527, n2265, n2199 );
nor U2668 ( new_g9110_, n2472, n2529 );
xnor U2669 ( n2529, n2208, n2530 );
nor U2670 ( n2530, n2531, n2481 );
nor U2671 ( n2531, n2480, n2532 );
nand U2672 ( n2532, n2533, n2534 );
nand U2673 ( n2534, n4683, n2199 );
nand U2674 ( n2533, n2523, n4684 );
nand U2675 ( new_g8973_, n2535, n2536 );
nand U2676 ( n2536, n2537, n2538 );
xor U2677 ( n2537, n2539, n4689 );
nand U2678 ( n2539, n2540, n2541 );
nand U2679 ( n2541, n4652, n2542 );
nand U2680 ( new_g8945_, n2543, n2544 );
nand U2681 ( n2544, n2545, n2546 );
xnor U2682 ( n2545, n4728, n2547 );
nor U2683 ( n2547, n2548, n2549 );
nand U2684 ( n2549, n2550, n2551 );
nand U2685 ( n2551, n2552, n2553 );
nor U2686 ( n2552, n2554, n2555 );
nand U2687 ( n2550, n4729, n2556 );
nand U2688 ( new_g8944_, n2543, n2557 );
nand U2689 ( n2557, n2558, n2546 );
xnor U2690 ( n2558, n2559, n2297 );
nand U2691 ( n2559, n2560, n2561 );
nor U2692 ( n2561, n2548, n2562 );
and U2693 ( n2562, n2563, n2564 );
nor U2694 ( n2560, n2565, n2566 );
nor U2695 ( n2566, n2553, n2291 );
and U2696 ( n2565, n2567, n2568 );
nand U2697 ( new_g8943_, n2543, n2569 );
nand U2698 ( n2569, n2546, n2570 );
nand U2699 ( n2570, n2571, n2572 );
nand U2700 ( n2572, n2573, n2574 );
nand U2701 ( n2573, n2575, n2576 );
nand U2702 ( n2576, n4723, n2577 );
nand U2703 ( n2577, n2578, n2579 );
nand U2704 ( n2579, n2568, n2204 );
nand U2705 ( n2578, n2556, n2248 );
nand U2706 ( n2571, n2580, n2269 );
nand U2707 ( n2580, n2581, n2582 );
nor U2708 ( n2582, n2583, n2584 );
and U2709 ( n2584, n4722, n2568 );
and U2710 ( n2583, n2204, n2564 );
nor U2711 ( n2581, n2548, n2585 );
nor U2712 ( n2585, n2553, n2248 );
nand U2713 ( new_g8941_, n2543, n2586 );
nand U2714 ( n2586, n2587, n2546 );
xnor U2715 ( n2587, n4727, n2588 );
nor U2716 ( n2588, n2589, n2548 );
nor U2717 ( n2589, n2590, n2591 );
nand U2718 ( n2591, n2592, n2593 );
nand U2719 ( n2593, n2594, n2242 );
nand U2720 ( n2592, n2595, n4434 );
nor U2721 ( n2590, n4547, n2553 );
nand U2722 ( new_g8940_, n2543, n2596 );
nand U2723 ( n2596, n2597, n2546 );
xnor U2724 ( n2597, n2598, n2242 );
nand U2725 ( n2598, n2574, n2599 );
nand U2726 ( n2599, n2600, n2601 );
nand U2727 ( n2601, n2556, n2286 );
nor U2728 ( n2600, n2594, n2595 );
nor U2729 ( n2595, n2304, n2602 );
nor U2730 ( n2594, n4726, n2603 );
nand U2731 ( new_g8939_, n2543, n2604 );
nand U2732 ( n2604, n2605, n2546 );
xnor U2733 ( n2605, n4726, n2606 );
nor U2734 ( n2606, n2607, n2548 );
nor U2735 ( n2607, n2608, n2609 );
nand U2736 ( n2609, n2603, n2602 );
nand U2737 ( n2602, n2610, n2611 );
nor U2738 ( n2610, n2237, n2194 );
nand U2739 ( n2603, n2612, n2613 );
nor U2740 ( n2612, n4724, n4725 );
nor U2741 ( n2608, n4548, n2553 );
nand U2742 ( new_g8938_, n2543, n2614 );
nand U2743 ( n2614, n2615, n2546 );
xnor U2744 ( n2615, n4725, n2616 );
nor U2745 ( n2616, n2548, n2617 );
nor U2746 ( n2617, n2618, n2619 );
nand U2747 ( n2619, n2620, n2621 );
nand U2748 ( n2621, n2613, n2194 );
nand U2749 ( n2620, n2611, n4724 );
nor U2750 ( n2618, n4549, n2553 );
not U2751 ( n2548, n2574 );
nand U2752 ( new_g8937_, n2543, n2622 );
nand U2753 ( n2622, n2623, n2546 );
xnor U2754 ( n2623, n2624, n2194 );
nand U2755 ( n2624, n2574, n2625 );
nand U2756 ( n2625, n2626, n2627 );
nand U2757 ( n2627, n2556, n2287 );
nor U2758 ( n2626, n2613, n2611 );
not U2759 ( n2611, n2575 );
nand U2760 ( n2575, n2628, n2564 );
nor U2761 ( n2564, n2629, n2556 );
nor U2762 ( n2628, n2269, n2204 );
and U2763 ( n2613, n2630, n2568 );
and U2764 ( n2568, n2553, n2629 );
nor U2765 ( n2630, n4722, n4723 );
nand U2766 ( new_g8926_, n2535, n2631 );
nand U2767 ( n2631, n2632, n2538 );
xnor U2768 ( n2632, n4435, n2633 );
nor U2769 ( n2633, n2634, n2635 );
nand U2770 ( n2635, n2636, n2637 );
nand U2771 ( n2637, n2638, n2639 );
nor U2772 ( n2638, n2640, n2641 );
nand U2773 ( n2636, n4695, n2542 );
nand U2774 ( new_g8923_, n2535, n2642 );
nand U2775 ( n2642, n2643, n2538 );
xnor U2776 ( n2643, n4436, n2644 );
nor U2777 ( n2644, n2634, n2645 );
nand U2778 ( n2645, n2646, n2647 );
nand U2779 ( n2647, n2648, n2639 );
nor U2780 ( n2648, n2649, n2650 );
nor U2781 ( n2649, n2651, n2652 );
nand U2782 ( n2646, n4648, n2542 );
nand U2783 ( new_g8922_, n2535, n2653 );
nand U2784 ( n2653, n2538, n2654 );
nand U2785 ( n2654, n2655, n2656 );
nand U2786 ( n2656, n2657, n2540 );
nand U2787 ( n2657, n2658, n2659 );
nand U2788 ( n2659, n4690, n2660 );
nand U2789 ( n2660, n2661, n2662 );
nand U2790 ( n2662, n2542, n2249 );
nand U2791 ( n2655, n2663, n2305 );
nand U2792 ( n2663, n2664, n2540 );
nor U2793 ( n2664, n2665, n2666 );
nor U2794 ( n2666, n2639, n2249 );
nor U2795 ( n2665, n2542, n2667 );
xnor U2796 ( n2667, n2651, n4689 );
nand U2797 ( new_g8921_, n2543, n2668 );
nand U2798 ( n2668, n2669, n2546 );
xnor U2799 ( n2669, n2670, n2204 );
nand U2800 ( n2670, n2574, n2671 );
nand U2801 ( n2671, n4551, n2556 );
not U2802 ( n2556, n2553 );
nand U2803 ( n2574, n2672, n2553 );
nand U2804 ( n2553, n2673, n2674 );
nand U2805 ( n2674, n4716, n2675 );
nand U2806 ( n2543, n2676, n2677 );
nor U2807 ( n2677, n4718, n2546 );
nor U2808 ( n2546, n2678, n2489 );
nor U2809 ( n2489, n2679, n2672 );
nand U2810 ( n2672, n2673, n2680 );
nand U2811 ( n2680, n2681, n2490 );
nand U2812 ( n2681, n2282, n2682 );
nand U2813 ( n2682, n4550, n4718 );
or U2814 ( n2679, n2683, n2684 );
nor U2815 ( n2684, n4728, n2555 );
nor U2816 ( n2555, n2567, n2685 );
nand U2817 ( n2685, n2629, n2297 );
nand U2818 ( n2567, n2686, n2687 );
nor U2819 ( n2687, n2688, n2689 );
nand U2820 ( n2689, n2194, n2269 );
nand U2821 ( n2688, n2204, n2242 );
nor U2822 ( n2686, n4727, n2690 );
nand U2823 ( n2690, n2304, n2237 );
nor U2824 ( n2683, n2554, n2453 );
and U2825 ( n2554, n2691, n4433 );
nor U2826 ( n2691, n2563, n2629 );
nand U2827 ( n2629, n2500, n2202 );
nand U2828 ( n2500, n4717, n4718 );
nand U2829 ( n2563, n2692, n2693 );
nor U2830 ( n2693, n2694, n2695 );
nand U2831 ( n2695, n4724, n4725 );
nand U2832 ( n2694, n4726, n4727 );
nor U2833 ( n2692, n2242, n2696 );
nand U2834 ( n2696, n4722, n4723 );
and U2835 ( n2676, n2490, n2496 );
nand U2836 ( n2490, n2697, n4716 );
nor U2837 ( n2697, n4715, n4717 );
nand U2838 ( new_g8920_, n2535, n2698 );
nand U2839 ( n2698, n2699, n2538 );
xnor U2840 ( n2699, n4694, n2700 );
nor U2841 ( n2700, n2701, n2634 );
nor U2842 ( n2701, n2702, n2703 );
nand U2843 ( n2703, n2704, n2705 );
nand U2844 ( n2705, n2706, n2294 );
nand U2845 ( n2704, n2707, n4437 );
nor U2846 ( n2702, n4649, n2639 );
nand U2847 ( new_g8889_, n2535, n2708 );
nand U2848 ( n2708, n2709, n2538 );
xnor U2849 ( n2709, n2710, n2294 );
nand U2850 ( n2710, n2540, n2711 );
nand U2851 ( n2711, n2712, n2713 );
nand U2852 ( n2713, n2542, n2288 );
nor U2853 ( n2712, n2706, n2707 );
nor U2854 ( n2707, n2714, n2658 );
not U2855 ( n2658, n2715 );
nor U2856 ( n2706, n4693, n2716 );
nand U2857 ( new_g8887_, n2535, n2717 );
nand U2858 ( n2717, n2718, n2538 );
xnor U2859 ( n2718, n4693, n2719 );
nor U2860 ( n2719, n2720, n2634 );
nor U2861 ( n2720, n2721, n2722 );
nand U2862 ( n2722, n2723, n2716 );
nand U2863 ( n2716, n2724, n2725 );
nor U2864 ( n2724, n4691, n4692 );
nand U2865 ( n2723, n2726, n2715 );
nor U2866 ( n2726, n2230, n2195 );
nor U2867 ( n2721, n4650, n2639 );
nand U2868 ( new_g8885_, n2535, n2727 );
nand U2869 ( n2727, n2728, n2538 );
xnor U2870 ( n2728, n4692, n2729 );
nor U2871 ( n2729, n2634, n2730 );
nor U2872 ( n2730, n2731, n2732 );
nand U2873 ( n2732, n2733, n2734 );
nand U2874 ( n2734, n2725, n2195 );
nand U2875 ( n2733, n2715, n4691 );
nor U2876 ( n2731, n4651, n2639 );
nand U2877 ( new_g8883_, n2535, n2735 );
nand U2878 ( n2735, n2736, n2538 );
xnor U2879 ( n2736, n2737, n2195 );
nand U2880 ( n2737, n2540, n2738 );
nand U2881 ( n2738, n2739, n2740 );
nand U2882 ( n2740, n2542, n2289 );
nor U2883 ( n2739, n2725, n2715 );
nor U2884 ( n2715, n2741, n2542 );
nor U2885 ( n2725, n2661, n4690 );
nand U2886 ( n2661, n2742, n2639 );
nor U2887 ( n2742, n4689, n2651 );
not U2888 ( n2540, n2634 );
nor U2889 ( n2634, n2743, n2542 );
not U2890 ( n2542, n2639 );
nand U2891 ( n2639, n2744, n2745 );
nand U2892 ( n2745, n4682, n2746 );
nand U2893 ( n2535, n2747, n2748 );
nor U2894 ( n2748, n4685, n2538 );
not U2895 ( n2538, n2749 );
nor U2896 ( n2747, n2480, n2520 );
not U2897 ( n2480, n2750 );
nand U2898 ( new_g8820_, n2751, n2479 );
nand U2899 ( n2479, n2752, n4439 );
nor U2900 ( n2752, n2750, n2481 );
nand U2901 ( n2751, n2753, n2450 );
nand U2902 ( n2753, n2749, n2754 );
nand U2903 ( n2754, n2750, n2517 );
nand U2904 ( n2749, n2481, n2517 );
nand U2905 ( n2481, n2755, n2743 );
and U2906 ( n2743, n2744, n2756 );
nand U2907 ( n2756, n2757, n2750 );
nand U2908 ( n2750, n2758, n4682 );
nor U2909 ( n2758, n4681, n4683 );
nand U2910 ( n2757, n2281, n2759 );
nand U2911 ( n2759, n4684, n4685 );
nor U2912 ( n2755, n2760, n2761 );
nor U2913 ( n2761, n4435, n2641 );
nor U2914 ( n2641, n2762, n2652 );
nand U2915 ( n2652, n2763, n2764 );
nor U2916 ( n2764, n2765, n2766 );
nand U2917 ( n2766, n2195, n2305 );
or U2918 ( n2765, n4689, n4437 );
nor U2919 ( n2763, n4694, n2767 );
nand U2920 ( n2767, n2312, n2230 );
or U2921 ( n2762, n4436, n2651 );
nor U2922 ( n2760, n2640, n2454 );
and U2923 ( n2640, n4436, n2650 );
and U2924 ( n2650, n2768, n2769 );
nor U2925 ( n2769, n2741, n2714 );
nand U2926 ( n2714, n2770, n4691 );
nor U2927 ( n2770, n2312, n2230 );
nand U2928 ( n2741, n2771, n4689 );
and U2929 ( n2771, n2651, n4690 );
nor U2930 ( n2651, n2522, n4684 );
and U2931 ( n2768, n4694, n4437 );
nand U2932 ( new_g8779_, n2772, n2773 );
nand U2933 ( n2773, n2774, n2377 );
nand U2934 ( n2772, n2775, n2776 );
nand U2935 ( new_g8777_, n2777, n2778 );
nand U2936 ( n2778, n2774, n2394 );
nand U2937 ( n2777, n2775, n2779 );
nand U2938 ( new_g8776_, n2780, n2781 );
nand U2939 ( n2781, n2774, n2396 );
nand U2940 ( n2780, n2775, n2782 );
nor U2941 ( new_g8775_, n2783, n2784 );
xor U2942 ( n2783, n2785, n4458 );
nand U2943 ( new_g8774_, n2786, n2787 );
nand U2944 ( n2787, n2774, n2390 );
nand U2945 ( n2786, n2775, n2785 );
nand U2946 ( n2785, n2788, n2789 );
nand U2947 ( n2789, n2790, n2472 );
xor U2948 ( n2790, n2791, n4738 );
nand U2949 ( n2791, n2792, n2268 );
nand U2950 ( new_g8773_, n2793, n2794 );
nand U2951 ( n2794, n2774, n2380 );
nand U2952 ( n2793, n2775, n2795 );
nor U2953 ( new_g8772_, n2796, n2784 );
xor U2954 ( n2796, n2782, n4457 );
nand U2955 ( n2782, n2797, n2798 );
nand U2956 ( n2798, n2799, n2472 );
xor U2957 ( n2799, n2800, n4739 );
nand U2958 ( n2800, n2801, n2802 );
nor U2959 ( n2801, n4743, n4745 );
nand U2960 ( new_g8771_, n2803, n2804 );
nand U2961 ( n2804, n2774, n2382 );
nand U2962 ( n2803, n2775, n2805 );
nand U2963 ( new_g8770_, n2806, n2807 );
nand U2964 ( n2807, n2774, n2384 );
nand U2965 ( n2806, n2775, n2808 );
nor U2966 ( new_g8769_, n2809, n2784 );
xor U2967 ( n2809, n2808, n4454 );
nand U2968 ( n2808, n2810, n2811 );
nand U2969 ( n2811, n2812, n2472 );
xnor U2970 ( n2812, n2813, n2295 );
nand U2971 ( n2813, n2802, n2814 );
nor U2972 ( new_g8768_, n2815, n2784 );
xor U2973 ( n2815, n2779, n4456 );
nand U2974 ( n2779, n2816, n2817 );
nand U2975 ( n2817, n2818, n2472 );
xnor U2976 ( n2818, n4488, n2819 );
nor U2977 ( n2819, n2251, n2820 );
nor U2978 ( new_g8767_, n2821, n2784 );
xor U2979 ( n2821, n2805, n4460 );
nand U2980 ( n2805, n2822, n2823 );
nand U2981 ( n2823, n2824, n2472 );
xnor U2982 ( n2824, n4737, n2825 );
nor U2983 ( n2825, n2448, n2826 );
nor U2984 ( new_g8766_, n2827, n2784 );
xnor U2985 ( n2827, n2776, n2254 );
nand U2986 ( n2776, n2828, n2829 );
nand U2987 ( n2829, n2830, n2472 );
xor U2988 ( n2830, n2831, n4489 );
nand U2989 ( n2831, n2832, n4744 );
nor U2990 ( n2832, n4746, n2833 );
nor U2991 ( new_g8765_, n2834, n2784 );
xor U2992 ( n2834, n2795, n4459 );
nand U2993 ( n2795, n2835, n2836 );
nand U2994 ( n2836, n2837, n2472 );
xnor U2995 ( n2837, n4495, n2838 );
nor U2996 ( n2838, n4743, n2826 );
nand U2997 ( n2826, n2839, n4746 );
nor U2998 ( n2839, n4745, n2251 );
nand U2999 ( new_g8649_, n2840, n2841 );
nand U3000 ( n2841, n2842, n2331 );
nor U3001 ( n2840, n2843, n2844 );
nand U3002 ( new_g8631_, n2845, n2846 );
nand U3003 ( n2846, n2843, n2847 );
nand U3004 ( n2847, n2848, n2849 );
or U3005 ( n2849, n2850, n2851 );
nor U3006 ( n2848, n4440, n2852 );
nor U3007 ( n2852, n2853, n2854 );
nor U3008 ( n2854, n4678, n4443 );
nand U3009 ( n2845, n2855, n2517 );
nand U3010 ( n2855, n2856, n2857 );
nand U3011 ( n2857, n2858, g636 );
nand U3012 ( n2858, n2859, n68 );
nor U3013 ( n2859, n2860, n2861 );
xor U3014 ( n2861, n2862, n2863 );
nor U3015 ( n2863, n2864, n2865 );
nor U3016 ( n2865, n4687, n2208 );
nor U3017 ( n2864, n2866, n2281 );
nor U3018 ( n2866, n2523, n2245 );
nor U3019 ( n2862, n4439, n4438 );
nor U3020 ( n2860, n2867, n2868 );
nand U3021 ( n2868, n4681, n4684 );
nand U3022 ( n2867, n2746, n2869 );
not U3023 ( n2869, n2523 );
nand U3024 ( n2856, n2520, n4439 );
nand U3025 ( new_g8559_, n2870, n2871 );
nand U3026 ( n2871, n2872, n2326 );
nor U3027 ( n2870, n2678, n2873 );
nor U3028 ( new_g8505_, n2874, n2472 );
xnor U3029 ( n2874, n4682, n2875 );
nor U3030 ( n2875, n2844, n2876 );
nor U3031 ( n2876, n2476, n2746 );
nand U3032 ( n2746, n2877, n2878 );
nor U3033 ( n2878, n2265, n2879 );
nand U3034 ( n2879, n4682, n2208 );
nor U3035 ( n2844, n2842, n4695 );
nor U3036 ( new_g8384_, n2880, n2472 );
xnor U3037 ( n2880, n4716, n2881 );
nor U3038 ( n2881, n2873, n2882 );
nor U3039 ( n2882, n2487, n2675 );
nor U3040 ( n2873, n2872, n4729 );
nor U3041 ( new_g8260_, n4669, n2883 );
nor U3042 ( new_g8254_, n4668, n2883 );
nor U3043 ( new_g8250_, n4667, n2883 );
nor U3044 ( new_g8245_, n2884, n2885 );
xor U3045 ( n2885, n4440, n2886 );
nor U3046 ( n2886, n2887, n2888 );
not U3047 ( n2887, n2853 );
nor U3048 ( n2853, n4442, n4679 );
nor U3049 ( new_g8244_, n2889, n2890 );
xnor U3050 ( n2890, g4181, n2891 );
nand U3051 ( g8349, n4664, n2439 );
nand U3052 ( g8340, n4664, n2440 );
nand U3053 ( g8335, n4664, n2434 );
nand U3054 ( g8331, n4664, n2441 );
nand U3055 ( g8328, n4664, n2435 );
nand U3056 ( g8323, n4664, n2442 );
nand U3057 ( g8318, n4664, n2436 );
nand U3058 ( g8316, n4664, n2443 );
nand U3059 ( g8313, n4664, n2437 );
nand U3060 ( g8347, n4664, n2444 );
nand U3061 ( new_g8194_, n2892, n2893 );
nand U3062 ( n2893, n2774, n2375 );
nand U3063 ( n2892, n2894, n2775 );
xnor U3064 ( n2894, n4740, n2895 );
nor U3065 ( n2895, n4744, n2820 );
nand U3066 ( n2820, n2896, n4743 );
nor U3067 ( n2896, n4746, n2268 );
nand U3068 ( new_g8193_, n2897, n2898 );
nand U3069 ( n2898, n2774, n2386 );
nand U3070 ( n2897, n2899, n2775 );
xor U3071 ( n2899, n2900, n4494 );
nand U3072 ( n2900, n2792, n4745 );
and U3073 ( n2792, n2802, n4743 );
and U3074 ( n2802, n4746, n2251 );
nand U3075 ( g8352, n4664, n2438 );
nor U3076 ( new_g8173_, g1713, n2901 );
xnor U3077 ( n2901, n2263, n2902 );
nor U3078 ( n2902, n4714, n2903 );
nor U3079 ( new_g8147_, n4666, n2883 );
nand U3080 ( n2883, g109, n2904 );
nand U3081 ( n2904, n4441, n44 );
nor U3082 ( new_g8060_, n2905, n2784 );
xnor U3083 ( n2905, new_g6002_, n2221 );
nor U3084 ( new_g8059_, n2784, n2906 );
xnor U3085 ( n2906, new_g6042_, n2260 );
nor U3086 ( new_g8055_, n2907, n2784 );
xor U3087 ( n2907, n2908, n4751 );
nor U3088 ( new_g8054_, n2909, n2784 );
xor U3089 ( n2909, new_g6015_, n4445 );
nor U3090 ( new_g8053_, n2784, n2910 );
xnor U3091 ( n2910, new_g6045_, n2222 );
nor U3092 ( new_g8052_, n2911, n2784 );
xnor U3093 ( n2911, n2912, n2225 );
nor U3094 ( new_g8051_, n2784, n2913 );
xnor U3095 ( n2913, n2914, n4453 );
nor U3096 ( new_g8050_, n2915, n2784 );
xor U3097 ( n2915, new_g6026_, n4444 );
nor U3098 ( new_g8049_, n2784, n2916 );
xor U3099 ( n2916, new_g6049_, n4446 );
nor U3100 ( new_g8048_, n2917, n2784 );
xnor U3101 ( n2917, new_g5996_, n2257 );
nor U3102 ( new_g8047_, n2918, n2784 );
xnor U3103 ( n2918, new_g6035_, n2223 );
nor U3104 ( new_g8046_, n2919, n2784 );
xnor U3105 ( n2919, n2920, n2224 );
nor U3106 ( new_g8045_, n2784, n2921 );
xnor U3107 ( n2921, n2922, n4452 );
nor U3108 ( new_g8044_, n2923, n2784 );
xnor U3109 ( n2923, new_g6038_, n2261 );
nor U3110 ( new_g8043_, n2924, n2784 );
xor U3111 ( n2924, n2925, n4450 );
nor U3112 ( new_g8042_, n2784, n2926 );
xnor U3113 ( n2926, n2927, n4451 );
nor U3114 ( new_g8041_, n2928, n2784 );
xnor U3115 ( n2928, n2929, n2252 );
nor U3116 ( new_g8040_, n2930, n2784 );
xor U3117 ( n2930, n2931, n4455 );
nor U3118 ( new_g8039_, n2932, n2784 );
xor U3119 ( n2932, n2933, n4750 );
nor U3120 ( new_g8024_, n2884, n2934 );
xor U3121 ( n2934, n4679, n2935 );
nor U3122 ( n2935, n4442, n2888 );
nor U3123 ( new_g8019_, n2889, n2936 );
xnor U3124 ( n2936, n4533, n2937 );
nor U3125 ( new_g7930_, g1713, n2938 );
xnor U3126 ( n2938, n4714, n2903 );
nand U3127 ( n2903, n2939, n2200 );
nor U3128 ( new_g7843_, n2940, n2784 );
xor U3129 ( n2940, new_g6000_, n4447 );
nor U3130 ( new_g7709_, n2884, n2941 );
xnor U3131 ( n2941, n4442, n2888 );
nand U3132 ( n2888, n2942, g814 );
nor U3133 ( new_g7705_, n2889, n2943 );
xnor U3134 ( n2943, n4675, n2944 );
nand U3135 ( new_g7660_, n2945, n2946 );
or U3136 ( n2946, n2947, n4655 );
nor U3137 ( new_g7632_, n2948, n2949 );
xnor U3138 ( n2949, n2301, n2950 );
nand U3139 ( new_g7626_, n2951, n2517 );
nor U3140 ( n2951, n2952, n2953 );
nor U3141 ( n2953, n2281, n2954 );
nand U3142 ( n2954, n2744, n2528 );
nand U3143 ( n2528, n2955, n4684 );
nor U3144 ( n2955, n2523, n2520 );
and U3145 ( n2520, n2956, n4683 );
nor U3146 ( n2956, n4685, n2199 );
nor U3147 ( n2523, n4685, n4683 );
nor U3148 ( n2952, n4687, n2744 );
nor U3149 ( new_g7590_, n2957, n2948 );
nor U3150 ( n2957, n2958, n2467 );
nor U3151 ( n2958, n4543, n2959 );
nor U3152 ( new_g7586_, n2948, n2960 );
xnor U3153 ( n2960, n4543, n2959 );
or U3154 ( n2959, n2961, n4735 );
nor U3155 ( new_g7581_, n2948, n2962 );
xnor U3156 ( n2962, n4735, n2961 );
nand U3157 ( n2961, n2950, n2301 );
nor U3158 ( n2950, n2963, n2964 );
nand U3159 ( n2948, n4487, g109 );
nor U3160 ( new_g7541_, g1713, n2965 );
xnor U3161 ( n2965, n2200, n2939 );
nor U3162 ( n2939, n2966, n2967 );
nand U3163 ( new_g7441_, n2968, n2945 );
nor U3164 ( n2968, n2969, n2970 );
nor U3165 ( n2970, n4653, n2446 );
nand U3166 ( new_g7257_, n2971, n2972 );
nand U3167 ( n2972, n2775, n2352 );
nand U3168 ( n2971, n2774, n2432 );
nand U3169 ( new_g7244_, n2973, n2974 );
nand U3170 ( n2974, n2775, n2353 );
or U3171 ( n2973, n2775, n4511 );
nand U3172 ( new_g7219_, n2440, n2975 );
nand U3173 ( new_g7204_, n2441, n2975 );
nor U3174 ( new_g7202_, n2884, n2976 );
xnor U3175 ( n2976, g814, n2942 );
nor U3176 ( n2942, n2977, n4678 );
nor U3177 ( new_g7191_, n2889, n2978 );
xnor U3178 ( n2978, n4534, n2979 );
nand U3179 ( new_g7189_, n2442, n2975 );
nand U3180 ( new_g7183_, n2443, n2975 );
nand U3181 ( new_g7143_, n2444, n2975 );
nor U3182 ( new_g7137_, n2980, n2981 );
nor U3183 ( n2980, n2982, n2947 );
nor U3184 ( n2982, n4654, n2983 );
nor U3185 ( new_g7134_, n2984, n2981 );
not U3186 ( n2981, n2945 );
nor U3187 ( n2945, n2744, n2843 );
not U3188 ( n2744, n2476 );
nor U3189 ( n2984, n2985, n2983 );
nor U3190 ( n2985, n4688, n2969 );
nand U3191 ( new_g7133_, n4709, n2986 );
xnor U3192 ( n2986, n4500, n2987 );
nand U3193 ( new_g7032_, n2988, n2989 );
nand U3194 ( n2989, n2990, n2991 );
nor U3195 ( n2991, n2992, n2993 );
nand U3196 ( n2993, n2994, n2995 );
nor U3197 ( n2995, n2221, n2260 );
nor U3198 ( n2994, n2222, n2257 );
nand U3199 ( n2992, n2996, n2997 );
nor U3200 ( n2997, n4444, n4445 );
nor U3201 ( n2996, n4446, n4464 );
nor U3202 ( n2990, n2998, n2999 );
nand U3203 ( n2999, n3000, n3001 );
and U3204 ( n3001, new_g6786_, n4656 );
nor U3205 ( n3000, n2306, n2228 );
nand U3206 ( n2998, n3002, n3003 );
nor U3207 ( n3003, n2223, n2261 );
and U3208 ( n3002, n4447, n3004 );
nand U3209 ( n2988, g109, n2403 );
nor U3210 ( new_g6983_, g1713, n3005 );
xnor U3211 ( n3005, n2217, n3006 );
nor U3212 ( n3006, n4713, n2966 );
nand U3213 ( new_g6934_, n3007, n3008 );
nand U3214 ( n3008, n3009, n2397 );
or U3215 ( n3007, n3009, n4444 );
nand U3216 ( new_g6930_, n3010, n3011 );
nand U3217 ( n3011, n2775, n2343 );
or U3218 ( n3010, n2775, n4506 );
nand U3219 ( new_g6929_, n3012, n3013 );
or U3220 ( n3013, n3014, n4564 );
nand U3221 ( n3012, n3014, n2228 );
nand U3222 ( new_g6928_, n3015, n3016 );
or U3223 ( n3016, n3014, n4628 );
or U3224 ( n3015, n3009, n4445 );
nand U3225 ( new_g6924_, n3017, n3018 );
nand U3226 ( n3018, n2775, n2344 );
or U3227 ( n3017, n2775, n4507 );
nand U3228 ( new_g6923_, n3019, n3020 );
or U3229 ( n3020, n3014, n4588 );
or U3230 ( n3019, n3009, n4446 );
nand U3231 ( new_g6922_, n3021, n3022 );
nand U3232 ( n3022, n3009, n2415 );
nand U3233 ( n3021, n3014, n2221 );
nand U3234 ( new_g6918_, n3023, n3024 );
nand U3235 ( n3024, n2775, n2345 );
or U3236 ( n3023, n2775, n4504 );
nand U3237 ( new_g6916_, n3025, n3026 );
nand U3238 ( n3026, n3009, n2414 );
nand U3239 ( n3025, n3014, n2222 );
nand U3240 ( new_g6915_, n3027, n3028 );
or U3241 ( n3028, n3014, n4585 );
or U3242 ( n3027, n3009, n4447 );
nand U3243 ( new_g6912_, n3029, n3030 );
nand U3244 ( n3030, n2775, n2346 );
nand U3245 ( n3029, n2774, n2299 );
nand U3246 ( new_g6911_, n3031, n3032 );
nand U3247 ( n3032, n3009, n2429 );
nand U3248 ( n3031, n3014, n2260 );
nand U3249 ( new_g6910_, n3033, n3034 );
nand U3250 ( n3034, n3009, n2413 );
nand U3251 ( n3033, n3014, n2257 );
nand U3252 ( new_g6909_, n3035, n3036 );
or U3253 ( n3036, n3037, n4553 );
nand U3254 ( new_g6908_, n3038, n3039 );
nand U3255 ( n3039, n2775, n2347 );
or U3256 ( n3038, n2775, n4510 );
nand U3257 ( new_g6907_, n3040, n3041 );
or U3258 ( n3041, n3014, n4634 );
nand U3259 ( n3040, n3014, n2261 );
nand U3260 ( new_g6906_, n3042, n3043 );
nand U3261 ( n3043, n3009, n2428 );
nand U3262 ( n3042, n3014, n2306 );
nand U3263 ( new_g6902_, n3044, n3045 );
nand U3264 ( n3045, n2775, n2348 );
nand U3265 ( n3044, n2774, n2300 );
nand U3266 ( new_g6901_, n3046, n3047 );
or U3267 ( n3047, n3014, n4584 );
nand U3268 ( n3046, n3014, n2223 );
nand U3269 ( new_g6900_, n3048, n3049 );
nand U3270 ( n3049, n3009, n2420 );
or U3271 ( n3048, n3009, n4448 );
nand U3272 ( new_g6898_, n3050, n3051 );
nand U3273 ( n3051, n2775, n2349 );
or U3274 ( n3050, n2775, n4508 );
nand U3275 ( new_g6897_, n3052, n3053 );
nand U3276 ( n3053, n3009, n2405 );
or U3277 ( n3052, n3009, n4464 );
not U3278 ( n3009, n3014 );
nand U3279 ( n3014, g109, n3054 );
nand U3280 ( n3054, n4656, n3004 );
nand U3281 ( new_g6895_, n3055, n3056 );
nand U3282 ( n3056, n2775, n2350 );
or U3283 ( n3055, n2775, n4509 );
nand U3284 ( new_g6894_, n3057, n3058 );
nand U3285 ( n3058, n2775, n2351 );
nand U3286 ( n3057, n2774, n2298 );
nor U3287 ( new_g6841_, n4756, n2784 );
nor U3288 ( new_g6840_, n4512, n2784 );
nor U3289 ( new_g6839_, n4474, n2784 );
nor U3290 ( new_g6838_, n4755, n2784 );
nor U3291 ( new_g6834_, n4760, n2784 );
nor U3292 ( new_g6833_, n4771, n2784 );
nor U3293 ( new_g6832_, n4770, n2784 );
nor U3294 ( new_g6831_, n4769, n2784 );
nor U3295 ( new_g6830_, n4768, n2784 );
nor U3296 ( new_g6829_, n4767, n2784 );
nor U3297 ( new_g6828_, n4766, n2784 );
nor U3298 ( new_g6827_, n4765, n2784 );
nor U3299 ( new_g6826_, n4763, n2784 );
nor U3300 ( new_g6824_, n4764, n2784 );
nor U3301 ( new_g6823_, n4762, n2784 );
nor U3302 ( new_g6822_, n4761, n2784 );
nor U3303 ( new_g6821_, n4759, n2784 );
nor U3304 ( new_g6820_, n4758, n2784 );
nor U3305 ( new_g6819_, n4757, n2784 );
nor U3306 ( new_g6795_, n3059, n3060 );
nor U3307 ( n3059, n3061, n3037 );
nor U3308 ( n3061, n4721, n3062 );
nor U3309 ( new_g6786_, n2784, n4448 );
nor U3310 ( new_g6759_, n4462, n2784 );
nor U3311 ( new_g6757_, n4461, n2784 );
nand U3312 ( new_g6755_, n4719, n3063 );
nor U3313 ( new_g6747_, n2460, n3064 );
nand U3314 ( n3064, g109, n3065 );
nand U3315 ( n3065, n4449, n4470 );
nor U3316 ( new_g6733_, n2884, n3066 );
xnor U3317 ( n3066, n4678, n2977 );
nand U3318 ( n2977, n2851, n2850 );
nor U3319 ( n2850, n4676, n4677 );
nor U3320 ( new_g6728_, n2889, n3067 );
xnor U3321 ( n3067, n4535, n3068 );
nand U3322 ( new_g6679_, n3069, n3070 );
nand U3323 ( n3070, n3071, n3072 );
nor U3324 ( n3072, n3073, n3074 );
nand U3325 ( n3074, n3075, n4460 );
nor U3326 ( n3075, n4459, n4466 );
nand U3327 ( n3073, n3076, n3077 );
nor U3328 ( n3077, n4454, n4456 );
nor U3329 ( n3076, n4457, n4458 );
nor U3330 ( n3071, n3078, n3079 );
nand U3331 ( n3079, n3080, n4465 );
nor U3332 ( n3080, n2238, n2341 );
nand U3333 ( n3078, n3081, new_g6224_ );
nor U3334 ( n3081, n3082, n3083 );
nand U3335 ( n3069, g109, n2427 );
nand U3336 ( new_g6672_, n4686, n3084 );
nand U3337 ( new_g6656_, n3085, n3086 );
nand U3338 ( n3086, n3087, n3088 );
nor U3339 ( n3088, n3089, n3090 );
nand U3340 ( n3090, n3091, n3092 );
nor U3341 ( n3092, n4471, n4473 );
nor U3342 ( n3091, n4750, n4751 );
nand U3343 ( n3089, n3093, n3094 );
nor U3344 ( n3094, n4450, n4452 );
nor U3345 ( n3093, n4455, n4469 );
nor U3346 ( n3087, n3095, n3096 );
nand U3347 ( n3096, n3097, n4472 );
nor U3348 ( n3097, n3082, n3098 );
not U3349 ( n3098, new_g6180_ );
nand U3350 ( n3095, n3099, n3100 );
nor U3351 ( n3100, n2225, n2324 );
nor U3352 ( n3099, n2224, n2323 );
nand U3353 ( n3085, g109, n2418 );
nor U3354 ( new_g6653_, n3101, n2434 );
nor U3355 ( new_g6638_, n3101, n2435 );
nor U3356 ( new_g6627_, n3101, n2436 );
nor U3357 ( new_g6621_, n3101, n2437 );
nand U3358 ( new_g6551_, n3102, n3103 );
nand U3359 ( n3103, n3104, n2400 );
or U3360 ( n3102, n3104, n4450 );
nand U3361 ( new_g6546_, n3105, n3106 );
or U3362 ( n3106, n3107, n4565 );
nand U3363 ( n3105, n3107, n2452 );
nand U3364 ( new_g6545_, n3108, n3109 );
or U3365 ( n3109, n3107, n4627 );
nand U3366 ( n3108, n3107, n2224 );
nand U3367 ( new_g6542_, n3110, n3111 );
or U3368 ( n3111, n3107, n4587 );
nand U3369 ( n3110, n3107, n2323 );
nand U3370 ( new_g6541_, n3112, n3113 );
nand U3371 ( n3113, n3104, n2416 );
nand U3372 ( n3112, n3107, n2225 );
nand U3373 ( new_g6538_, n3114, n3115 );
or U3374 ( n3115, n3107, n4606 );
or U3375 ( n3114, n3104, n4452 );
nand U3376 ( new_g6537_, n3116, n3117 );
or U3377 ( n3117, n3107, n4591 );
or U3378 ( n3116, n3104, n4751 );
nand U3379 ( new_g6534_, n3118, n3119 );
or U3380 ( n3119, n3107, n4617 );
nand U3381 ( n3118, n3107, n2324 );
nand U3382 ( new_g6533_, n3120, n3121 );
or U3383 ( n3121, n3107, n4607 );
nand U3384 ( n3120, n3107, n2252 );
nor U3385 ( new_g6531_, n3101, n2438 );
nand U3386 ( new_g6529_, n3122, n3123 );
or U3387 ( n3123, n3107, n4637 );
or U3388 ( n3122, n3104, n4750 );
nand U3389 ( new_g6528_, n3124, n3125 );
or U3390 ( n3125, n3107, n4618 );
nand U3391 ( n3124, n3107, n2316 );
nor U3392 ( new_g6526_, n3101, n2439 );
nor U3393 ( new_g6525_, g1713, n3126 );
xnor U3394 ( n3126, n4713, n2966 );
nand U3395 ( n2966, n3127, n2198 );
nand U3396 ( new_g6524_, n3128, n3129 );
nand U3397 ( n3129, n3104, n2399 );
or U3398 ( n3128, n3104, n4454 );
nand U3399 ( new_g6523_, n3130, n3131 );
or U3400 ( n3131, n3107, n4579 );
or U3401 ( n3130, n3104, n4455 );
nand U3402 ( new_g6522_, n3132, n3133 );
nand U3403 ( n3133, n3104, n2422 );
or U3404 ( n3132, n3104, n4469 );
nor U3405 ( new_g6516_, g1713, n3134 );
xnor U3406 ( n3134, n2198, n3127 );
nor U3407 ( n3127, n3135, n4712 );
nand U3408 ( new_g6515_, n3136, n3137 );
or U3409 ( n3137, n3107, n4568 );
nand U3410 ( n3136, n3107, n2254 );
nand U3411 ( new_g6514_, n3138, n3139 );
nand U3412 ( n3139, n3104, n2409 );
nand U3413 ( n3138, n3107, n2341 );
nand U3414 ( new_g6513_, n3140, n3141 );
nand U3415 ( n3141, n3104, n2407 );
or U3416 ( n3140, n3104, n4473 );
nor U3417 ( new_g6508_, g1713, n3142 );
xnor U3418 ( n3142, n4712, n3135 );
nand U3419 ( n3135, n3143, n2241 );
nand U3420 ( new_g6507_, n3144, n3145 );
or U3421 ( n3145, n3107, n4597 );
or U3422 ( n3144, n3104, n4456 );
nand U3423 ( new_g6506_, n3146, n3147 );
or U3424 ( n3147, n3107, n4571 );
or U3425 ( n3146, n3104, n4466 );
nor U3426 ( new_g6502_, g1713, n3148 );
xnor U3427 ( n3148, n2241, n3143 );
nor U3428 ( n3143, n2987, n4500 );
nand U3429 ( new_g6501_, n3149, n3150 );
or U3430 ( n3150, n3107, n4605 );
or U3431 ( n3149, n3104, n4457 );
nand U3432 ( new_g6500_, n3151, n3152 );
or U3433 ( n3152, n3107, n4590 );
or U3434 ( n3151, n3104, n4465 );
nand U3435 ( new_g6481_, n3153, n3154 );
or U3436 ( n3154, n3107, n4616 );
or U3437 ( n3153, n3104, n4458 );
nand U3438 ( new_g6480_, n3155, n3156 );
or U3439 ( n3156, n3107, n4609 );
nand U3440 ( n3155, n3107, n2226 );
nand U3441 ( new_g6479_, n3157, n3158 );
or U3442 ( n3158, n3107, n4636 );
or U3443 ( n3157, n3104, n4459 );
nand U3444 ( new_g6478_, n3159, n3160 );
or U3445 ( n3160, n3107, n4620 );
nand U3446 ( n3159, n3107, n2277 );
nor U3447 ( new_g6471_, n3161, n3060 );
nor U3448 ( n3161, n3162, n3062 );
nor U3449 ( n3162, n4552, n2445 );
nand U3450 ( new_g6470_, n3163, n3164 );
or U3451 ( n3164, n3107, n4580 );
or U3452 ( n3163, n3104, n4460 );
nand U3453 ( new_g6469_, n3165, n3166 );
nand U3454 ( n3166, n3104, n2421 );
or U3455 ( n3165, n3104, n4467 );
nand U3456 ( new_g6468_, n3167, n3168 );
nand U3457 ( n3168, n3104, n2406 );
not U3458 ( n3104, n3107 );
nand U3459 ( n3167, n3107, n2238 );
nand U3460 ( n3082, n4773, n3004 );
nor U3461 ( new_g6439_, n3169, n2784 );
xor U3462 ( n3169, n3170, n3171 );
xnor U3463 ( n3171, n2228, n4462 );
xnor U3464 ( n3170, n4464, n4463 );
nor U3465 ( new_g6334_, n4754, n2784 );
nor U3466 ( new_g6332_, n4752, n2784 );
nor U3467 ( new_g6244_, n4465, n2784 );
nand U3468 ( new_g6243_, n3172, n3173 );
not U3469 ( n3173, n2884 );
xnor U3470 ( n3172, n4476, n4475 );
nor U3471 ( new_g6224_, n2784, n4467 );
nor U3472 ( new_g6216_, n4468, n2784 );
nor U3473 ( new_g6205_, n4748, n2784 );
nor U3474 ( new_g6193_, n4747, n2784 );
nor U3475 ( new_g6180_, n2784, n4749 );
nor U3476 ( new_g6179_, n4470, n3174 );
not U3477 ( n3174, new_g6163_ );
nor U3478 ( new_g6163_, n3175, n3176 );
nand U3479 ( new_g6155_, n3177, n3178 );
nand U3480 ( n3178, new_g4076_, n2197 );
nand U3481 ( n3177, n3179, n4730 );
nor U3482 ( n3179, n4486, n122 );
nand U3483 ( new_g6126_, n3180, n3181 );
nand U3484 ( n3181, n3182, g806 );
nor U3485 ( n3182, n3183, n2884 );
and U3486 ( n3183, g802, n2851 );
nand U3487 ( n3180, n3184, n4677 );
nor U3488 ( n3184, new_g5849_, n3185 );
or U3489 ( n3185, n4676, n4475 );
nand U3490 ( new_g6123_, n3186, n3187 );
nand U3491 ( n3187, n3188, g4176 );
nand U3492 ( n3188, n3189, n3190 );
nand U3493 ( n3190, n4536, n3191 );
not U3494 ( n3191, n2889 );
nand U3495 ( n3186, n3192, n4674 );
nor U3496 ( n3192, n3193, n2889 );
nand U3497 ( new_g6099_, n3194, n3195 );
nand U3498 ( n3195, n3196, n2356 );
nand U3499 ( n3194, n3197, n2343 );
nand U3500 ( new_g6096_, n3198, n3199 );
nand U3501 ( n3199, n3196, n2357 );
nand U3502 ( n3198, n3197, n2344 );
nand U3503 ( new_g6093_, n3200, n3201 );
nand U3504 ( n3201, n3196, n2358 );
nand U3505 ( n3200, n3197, n2345 );
nand U3506 ( new_g6088_, n3202, n3203 );
nand U3507 ( n3203, n3196, n2359 );
nand U3508 ( n3202, n3197, n2346 );
nand U3509 ( new_g6080_, n3204, n3205 );
nand U3510 ( n3205, n3196, n2360 );
nand U3511 ( n3204, n3197, n2347 );
nand U3512 ( new_g6071_, n3206, n3207 );
nand U3513 ( n3207, n3196, n2361 );
nand U3514 ( n3206, n3197, n2348 );
nand U3515 ( new_g6068_, n3208, n3209 );
nand U3516 ( n3209, n3196, n2362 );
nand U3517 ( n3208, n3197, n2349 );
nand U3518 ( new_g6059_, n3210, n3211 );
nand U3519 ( n3211, n3196, n2363 );
nand U3520 ( n3210, n3197, n2350 );
nand U3521 ( new_g6054_, n3212, n3213 );
nand U3522 ( n3213, n3196, n2354 );
nand U3523 ( n3212, n3197, n2351 );
nand U3524 ( new_g6049_, n3214, n3215 );
nand U3525 ( n3214, n2472, n2374 );
nand U3526 ( new_g6045_, n3216, n3217 );
nand U3527 ( n3216, n2472, n2376 );
nand U3528 ( new_g6042_, n3218, n3219 );
nand U3529 ( n3218, n2472, n2393 );
nand U3530 ( new_g6038_, n2828, n3220 );
nand U3531 ( n3220, n2472, n2395 );
nand U3532 ( new_g6035_, n2816, n3221 );
nand U3533 ( n3221, n2472, n2378 );
nand U3534 ( new_g6026_, n2797, n3222 );
nand U3535 ( n3222, n2472, n2379 );
nand U3536 ( new_g6015_, n2788, n3223 );
nand U3537 ( n3223, n2472, n2381 );
nand U3538 ( new_g6002_, n2835, n3224 );
nand U3539 ( n3224, n2472, n2383 );
nand U3540 ( new_g6000_, n2822, n3225 );
nand U3541 ( n3225, n2472, n2385 );
nand U3542 ( new_g5996_, n2810, n3226 );
nand U3543 ( n3226, n2472, n2387 );
nand U3544 ( new_g5914_, n3227, n3228 );
nand U3545 ( n3228, n3196, n2355 );
nand U3546 ( n3227, n3197, n2352 );
nand U3547 ( new_g5910_, n3229, n3230 );
nand U3548 ( n3230, n3196, n2364 );
nand U3549 ( n3229, n3197, n2353 );
nand U3550 ( new_g5770_, n3231, n3232 );
nand U3551 ( n3232, n3233, n3234 );
not U3552 ( n3234, n3235 );
nor U3553 ( n3233, n2784, n2316 );
nand U3554 ( n3231, new_g6198_, n3235 );
xor U3555 ( n3235, n4749, n3236 );
xnor U3556 ( n3236, n2252, n4473 );
nor U3557 ( new_g6198_, n2784, n4472 );
nor U3558 ( new_g5763_, n3237, n3238 );
nor U3559 ( n3238, n2784, n3239 );
nand U3560 ( new_g5755_, n3240, n3241 );
nand U3561 ( n3241, n4497, n3242 );
nor U3562 ( n3242, n3243, n3244 );
nor U3563 ( n3244, n3245, n3246 );
and U3564 ( n3245, g109, n4753 );
nor U3565 ( n3243, new_g6333_, n3247 );
nor U3566 ( n3240, n3248, n3249 );
nor U3567 ( n3249, n3247, n3250 );
nand U3568 ( n3250, new_g6331_, n4753 );
not U3569 ( new_g6331_, n3175 );
nand U3570 ( n3175, g109, n2247 );
nor U3571 ( n3248, n3246, n3251 );
nand U3572 ( n3251, new_g6333_, n2247 );
nor U3573 ( new_g6333_, n2784, n4753 );
not U3574 ( n3246, n3247 );
xor U3575 ( n3247, n4754, n3252 );
nor U3576 ( n3252, n3253, n2468 );
nor U3577 ( n3253, n3176, n2247 );
nand U3578 ( n3176, n3254, n3255 );
nor U3579 ( n3255, n3256, n3257 );
nand U3580 ( n3257, n3258, n3259 );
nor U3581 ( n3259, n2461, n3260 );
nand U3582 ( n3260, n4765, n4766 );
nor U3583 ( n3258, n2321, n3261 );
nand U3584 ( n3261, n4762, n4763 );
nand U3585 ( n3256, n3262, n3263 );
nor U3586 ( n3263, n2462, n3264 );
nand U3587 ( n3264, n4771, n4772 );
nor U3588 ( n3262, n2320, n3265 );
nand U3589 ( n3265, n4768, n4769 );
nor U3590 ( n3254, n3266, n3267 );
nand U3591 ( n3267, n3268, n3269 );
nor U3592 ( n3269, n2463, n3270 );
nand U3593 ( n3270, n4753, n4754 );
and U3594 ( n3268, n4512, n4474 );
nand U3595 ( n3266, n3271, n3272 );
nor U3596 ( n3272, n2464, n3273 );
nand U3597 ( n3273, n4759, n4760 );
nor U3598 ( n3271, n2319, n3274 );
nand U3599 ( n3274, n4756, n4757 );
nor U3600 ( new_g5556_, n3275, n3276 );
nand U3601 ( n3276, n3277, n3278 );
nor U3602 ( n3278, n4730, n2967 );
nor U3603 ( n3277, n2198, n3279 );
nand U3604 ( n3275, n3280, n3281 );
nor U3605 ( n3281, n4501, n3282 );
nand U3606 ( n3282, n2218, n2318 );
nor U3607 ( n3280, n4711, n4712 );
nand U3608 ( new_g5543_, n3283, n3284 );
nand U3609 ( n3284, n3285, g802 );
nor U3610 ( n3285, n2851, n2884 );
nor U3611 ( n2851, n4475, n4476 );
nand U3612 ( n3283, n3286, n4676 );
nor U3613 ( n3286, n4475, new_g5849_ );
or U3614 ( new_g5849_, n2884, n4476 );
nand U3615 ( n2884, n3287, g109 );
nor U3616 ( n3287, n4477, n4670 );
nand U3617 ( new_g5536_, n3288, n3289 );
or U3618 ( n3289, n3189, n4536 );
nor U3619 ( n3189, new_g4940_, n3290 );
nor U3620 ( n3290, g4174, n2889 );
nand U3621 ( n3288, n3291, n4536 );
nor U3622 ( n3291, n2889, n3292 );
nand U3623 ( n3292, g4174, g4173 );
nand U3624 ( new_g5529_, n3293, n3294 );
nand U3625 ( n3294, new_g4940_, g4174 );
nand U3626 ( n3293, n3295, n4673 );
nor U3627 ( n3295, n4672, n2889 );
nand U3628 ( new_g5445_, n3296, n3297 );
nand U3629 ( n3297, g109, n2328 );
nand U3630 ( new_g5421_, n3296, n3298 );
nand U3631 ( n3298, g109, n2426 );
nand U3632 ( new_g5404_, n3299, n3300 );
nand U3633 ( n3300, n2775, g1713 );
nand U3634 ( n3299, n2774, n2267 );
nand U3635 ( new_g5396_, n3301, n3302 );
nand U3636 ( n3302, n2775, g1710 );
nand U3637 ( n3301, n2774, g1713 );
nor U3638 ( new_g5390_, n4743, n3303 );
nor U3639 ( new_g5287_, new_g4089_, n2250 );
nor U3640 ( new_g5194_, n4529, n3304 );
nor U3641 ( new_g5173_, n4746, n3303 );
nor U3642 ( new_g5148_, n4745, n3303 );
nor U3643 ( new_g5126_, n4744, n3303 );
nand U3644 ( n3303, n4478, g109 );
nor U3645 ( new_g5083_, new_g4089_, n3305 );
nor U3646 ( n3305, n3304, n3196 );
nor U3647 ( new_g4940_, g4173, n2889 );
nand U3648 ( n2889, n4532, g109 );
nor U3649 ( new_g4905_, n4479, new_g3524_ );
not U3650 ( new_g4904_, n3306 );
nor U3651 ( new_g4903_, n4480, new_g3524_ );
nor U3652 ( new_g4902_, n4481, new_g3524_ );
nor U3653 ( new_g4893_, n4482, new_g4117_ );
nor U3654 ( new_g4891_, n4483, new_g4117_ );
nor U3655 ( new_g4890_, n4484, new_g4117_ );
nand U3656 ( new_g4556_, n4545, n4487 );
nor U3657 ( new_g4506_, n4740, n2784 );
nor U3658 ( new_g4500_, n4526, n2775 );
nor U3659 ( new_g4498_, n4489, n2784 );
nor U3660 ( new_g4490_, n4488, n2784 );
nor U3661 ( new_g4484_, n4739, n2784 );
nor U3662 ( new_g4480_, n4738, n2784 );
nor U3663 ( new_g4477_, n4495, n2784 );
nor U3664 ( new_g4473_, n4737, n2784 );
nor U3665 ( new_g4471_, n4736, n2784 );
nor U3666 ( new_g4465_, n4494, n2784 );
nor U3667 ( new_g4342_, n4742, n2784 );
nor U3668 ( new_g4340_, n4741, n2784 );
nor U3669 ( new_g4338_, n4492, n2784 );
nor U3670 ( new_g4334_, n4493, n2784 );
nor U3671 ( new_g4330_, n4490, n2784 );
nor U3672 ( new_g4325_, n4491, n2784 );
nand U3673 ( new_g4309_, n3307, n3308 );
nand U3674 ( n3308, n3309, n2263 );
or U3675 ( n3307, n3309, n4624 );
nand U3676 ( new_g4293_, n3310, n3311 );
nand U3677 ( n3311, n3309, n2276 );
or U3678 ( n3310, n3309, n4570 );
nand U3679 ( new_g4283_, n3312, n3313 );
nand U3680 ( n3313, n3309, n2200 );
or U3681 ( n3312, n3309, n4594 );
nand U3682 ( new_g4274_, n3314, n3315 );
nand U3683 ( n3315, n3309, n2217 );
nand U3684 ( n3314, n3316, n2410 );
nand U3685 ( new_g4264_, n3317, n3318 );
nand U3686 ( n3318, n3309, n2285 );
nand U3687 ( n3317, n3316, n2423 );
nand U3688 ( new_g4255_, n3319, n3320 );
nand U3689 ( n3320, n3309, n2198 );
nand U3690 ( n3319, n3316, n2417 );
nand U3691 ( new_g4239_, n3321, n3322 );
nand U3692 ( n3322, n3309, n2270 );
or U3693 ( n3321, n3309, n4577 );
nand U3694 ( new_g4238_, n3323, n3324 );
nand U3695 ( n3324, n3309, n2241 );
nand U3696 ( n3323, n3316, n2398 );
nand U3697 ( new_g4231_, n3325, n3326 );
nand U3698 ( n3326, n3309, n2218 );
or U3699 ( n3325, n3309, n4623 );
not U3700 ( n3309, n3316 );
nor U3701 ( new_g4114_, n3327, n3328 );
nand U3702 ( n3328, n2229, n2311 );
nand U3703 ( n3327, n2266, n2219 );
nand U3704 ( new_g4089_, n4485, n2451 );
nor U3705 ( new_g4076_, n2318, n122 );
nor U3706 ( new_g3506_, n3329, n3330 );
nand U3707 ( n3330, n2322, n2227 );
or U3708 ( n3329, n4601, n4576 );
nand U3709 ( new_g3462_, n3331, n3332 );
nand U3710 ( n3332, n3101, g746 );
nand U3711 ( n3331, new_g2791_, g4172 );
nand U3712 ( g6955, n3333, n3334 );
nand U3713 ( n3334, n4730, n2366 );
nand U3714 ( n3333, n2197, n2389 );
nand U3715 ( g6949, n3335, n3336 );
nand U3716 ( n3336, n4730, n2368 );
nand U3717 ( n3335, n2197, n2365 );
nand U3718 ( g6942, n3337, n3338 );
nand U3719 ( n3338, n4730, n2370 );
nand U3720 ( n3337, n2197, n2367 );
nand U3721 ( g6932, n3339, n3340 );
nand U3722 ( n3340, n4730, n2372 );
nand U3723 ( n3339, n2197, n2369 );
and U3724 ( g5659, n3341, g744 );
and U3725 ( n3341, g743, g109 );
nand U3726 ( g6926, n3342, n3343 );
nand U3727 ( n3343, n4730, n2391 );
nand U3728 ( n3342, n2197, n2371 );
and U3729 ( g5658, n3344, g742 );
and U3730 ( n3344, g741, g109 );
nand U3731 ( g6920, n3345, n3346 );
nand U3732 ( n3346, n4730, n2392 );
nand U3733 ( n3345, n2197, n2373 );
nor U3734 ( new_g3381_, n3347, n3348 );
or U3735 ( n3348, n4669, n4668 );
or U3736 ( n3347, n4667, n4666 );
and U3737 ( new_g2791_, n4671, g746 );
nor U3738 ( new_g2478_, n2259, g1737 );
nand U3739 ( new_g11647_, n3349, n3350 );
nand U3740 ( n3350, n2975, n2354 );
nand U3741 ( n3349, n3351, n3101 );
nand U3742 ( n3351, n3352, n3353 );
nand U3743 ( n3353, n3354, n3355 );
or U3744 ( n3352, n3355, n3356 );
nor U3745 ( new_g11641_, n3357, n3358 );
xnor U3746 ( n3358, n2266, n3359 );
nor U3747 ( n3359, n4612, n3360 );
nor U3748 ( new_g11640_, n3357, n3361 );
xnor U3749 ( n3361, n4612, n3360 );
nand U3750 ( n3360, n3362, n2229 );
nor U3751 ( new_g11639_, n3357, n3363 );
xnor U3752 ( n3363, n2229, n3362 );
and U3753 ( n3362, new_g11561_, n2219 );
nor U3754 ( new_g11636_, n3357, n3364 );
xnor U3755 ( n3364, n2219, new_g11561_ );
nand U3756 ( n3357, g109, n3365 );
nand U3757 ( n3365, n3366, n3239 );
nor U3758 ( n3366, n4487, n3237 );
not U3759 ( n3237, n3367 );
nand U3760 ( new_g11625_, n3368, n3369 );
nand U3761 ( n3369, n2975, n2355 );
nand U3762 ( n3368, n3370, n3101 );
xnor U3763 ( n3370, n3356, n3354 );
xor U3764 ( n3354, n3371, n3372 );
xor U3765 ( n3372, n3373, n3374 );
xor U3766 ( n3374, n3375, n3376 );
xor U3767 ( n3376, n3377, n3378 );
xor U3768 ( n3375, n3379, n3380 );
xor U3769 ( n3373, n3381, n3382 );
xor U3770 ( n3382, n3383, n3384 );
xor U3771 ( n3381, n3385, n3386 );
nand U3772 ( n3356, n3387, n3388 );
nand U3773 ( n3388, n3389, n2258 );
nand U3774 ( n3387, n3390, n3391 );
xnor U3775 ( n3390, n3392, n3393 );
or U3776 ( n3392, n2203, n3394 );
nand U3777 ( new_g11610_, n3395, n3396 );
nand U3778 ( n3396, n3397, n2263 );
or U3779 ( n3395, n3397, n4625 );
nand U3780 ( new_g11609_, n3398, n3399 );
nand U3781 ( n3399, n3397, n2276 );
or U3782 ( n3398, n3397, n4566 );
nand U3783 ( new_g11608_, n3400, n3401 );
nand U3784 ( n3401, n3397, n2200 );
or U3785 ( n3400, n3397, n4593 );
nand U3786 ( new_g11607_, n3402, n3403 );
nand U3787 ( n3403, n3397, n2217 );
or U3788 ( n3402, n3397, n4604 );
nand U3789 ( new_g11606_, n3404, n3405 );
nand U3790 ( n3405, n3397, n2285 );
or U3791 ( n3404, n3397, n4615 );
nand U3792 ( new_g11605_, n3406, n3407 );
nand U3793 ( n3407, n3397, n2198 );
nand U3794 ( n3406, n3408, n2419 );
nand U3795 ( new_g11604_, n3409, n3410 );
nand U3796 ( n3410, n3397, n2270 );
nand U3797 ( n3409, n3408, n2404 );
nand U3798 ( new_g11603_, n3411, n3412 );
nand U3799 ( n3412, n3397, n2241 );
or U3800 ( n3411, n3397, n4574 );
nand U3801 ( new_g11602_, n3413, n3414 );
nand U3802 ( n3414, n3397, n2218 );
or U3803 ( n3413, n3397, n4622 );
not U3804 ( n3397, n3408 );
nand U3805 ( n3408, new_g11561_, g1317 );
nand U3806 ( new_g11579_, n3415, n3416 );
nand U3807 ( n3416, n2774, n2388 );
nand U3808 ( n3415, n3417, n2775 );
xor U3809 ( n3417, n3418, n3419 );
xnor U3810 ( n3419, n3420, n2259 );
nand U3811 ( n3418, n3421, n3422 );
nand U3812 ( n3422, n3423, n2457 );
xnor U3813 ( n3423, n3424, n2296 );
nand U3814 ( n3421, n3425, n4742 );
xnor U3815 ( n3425, n3426, n3424 );
nand U3816 ( n3424, n3427, n4746 );
nor U3817 ( n3427, n2833, n2251 );
not U3818 ( n2833, n2814 );
nor U3819 ( n2814, n2268, n4743 );
nor U3820 ( n3426, n3428, n2296 );
nor U3821 ( n3428, n3429, n3430 );
nand U3822 ( n3430, n3431, n3432 );
nor U3823 ( n3432, n2465, n3433 );
nand U3824 ( n3433, n4494, n4740 );
nor U3825 ( n3431, n2466, n3434 );
nand U3826 ( n3434, n4491, n4492 );
nand U3827 ( n3429, n3435, n3436 );
nor U3828 ( n3436, n3437, n3438 );
nand U3829 ( n3438, n4738, n4739 );
nand U3830 ( n3437, n4488, n4489 );
nor U3831 ( n3435, n2295, n3439 );
nand U3832 ( n3439, n4737, n4495 );
and U3833 ( new_g11561_, n3440, n2964 );
nor U3834 ( n3440, n3441, n2963 );
nor U3835 ( n3441, n3442, n3443 );
nand U3836 ( n3443, n3444, n3445 );
nor U3837 ( n3445, n3446, n3447 );
nand U3838 ( n3447, n3448, n3449 );
xnor U3839 ( n3449, n4503, n4539 );
xnor U3840 ( n3448, n4504, n4540 );
xnor U3841 ( n3446, n4510, n2209 );
nor U3842 ( n3444, n3450, n3451 );
xnor U3843 ( n3451, n4511, n2255 );
xnor U3844 ( n3450, n4509, n2211 );
nand U3845 ( n3442, n3452, n3453 );
nor U3846 ( n3453, n3454, n3455 );
nand U3847 ( n3455, n3456, n3457 );
xnor U3848 ( n3457, n4505, n4732 );
xor U3849 ( n3456, n3458, n3459 );
xnor U3850 ( n3454, n4506, n2210 );
nor U3851 ( n3452, n3460, n3461 );
xnor U3852 ( n3461, n4507, n2243 );
xnor U3853 ( n3460, n4508, n2205 );
nor U3854 ( new_g11514_, n3462, n2784 );
xor U3855 ( n3462, n3420, n3463 );
xnor U3856 ( n3463, n4496, n3464 );
nor U3857 ( n3464, n3465, n3466 );
nand U3858 ( n3466, n3467, n3468 );
nand U3859 ( n3468, n3469, n2254 );
nor U3860 ( n3469, n2226, n2277 );
nand U3861 ( n3467, n3470, n4498 );
xnor U3862 ( n3470, n2226, n4748 );
not U3863 ( n3465, n3083 );
nand U3864 ( n3083, n3471, n2277 );
nor U3865 ( n3471, n4498, n4747 );
nand U3866 ( n3420, n3472, n3473 );
nand U3867 ( n3473, g18, n2247 );
nand U3868 ( n3472, n3474, n2472 );
nand U3869 ( n3474, n3475, n3476 );
or U3870 ( n3476, n3477, n2447 );
nand U3871 ( n3475, n3478, n3477 );
nand U3872 ( n3477, n3479, n3480 );
and U3873 ( n3480, n4525, n4524 );
and U3874 ( n3479, n4523, n4522 );
nand U3875 ( n3478, n3481, n3482 );
nand U3876 ( new_g11488_, n3483, n3484 );
nand U3877 ( n3484, n2975, n2356 );
nand U3878 ( n3483, n3378, n3101 );
nand U3879 ( n3378, n3485, n3486 );
or U3880 ( n3486, n3391, n4520 );
nand U3881 ( n3485, n3487, n3391 );
xnor U3882 ( n3487, n3488, n2216 );
nand U3883 ( n3488, n3489, n3490 );
nor U3884 ( n3490, n4700, n4703 );
nor U3885 ( n3489, n2262, n2203 );
nand U3886 ( new_g11487_, n3491, n3492 );
nand U3887 ( n3492, n2975, n2357 );
nand U3888 ( n3491, n3377, n3101 );
nand U3889 ( n3377, n3493, n3494 );
or U3890 ( n3494, n3391, n4518 );
nand U3891 ( n3493, n3495, n3391 );
xnor U3892 ( n3495, n4642, n3496 );
nor U3893 ( n3496, n2203, n3497 );
nand U3894 ( new_g11486_, n3498, n3499 );
nand U3895 ( n3499, n2975, n2358 );
nand U3896 ( n3498, n3380, n3101 );
nand U3897 ( n3380, n3500, n3501 );
or U3898 ( n3501, n3391, n4519 );
nand U3899 ( n3500, n3502, n3391 );
xnor U3900 ( n3502, n3503, n2215 );
nand U3901 ( new_g11485_, n3504, n3505 );
nand U3902 ( n3505, n2975, n2359 );
nand U3903 ( n3504, n3379, n3101 );
nand U3904 ( n3379, n3506, n3507 );
or U3905 ( n3507, n3391, n4513 );
nand U3906 ( n3506, n3508, n3391 );
xnor U3907 ( n3508, n4647, n3509 );
nor U3908 ( n3509, n4702, n3510 );
nand U3909 ( new_g11484_, n3511, n3512 );
nand U3910 ( n3512, n2975, n2360 );
nand U3911 ( n3511, n3384, n3101 );
nand U3912 ( n3384, n3513, n3514 );
or U3913 ( n3514, n3391, n4517 );
nand U3914 ( n3513, n3515, n3391 );
xnor U3915 ( n3515, n4646, n3516 );
nor U3916 ( n3516, n4700, n3517 );
nand U3917 ( new_g11483_, n3518, n3519 );
nand U3918 ( n3519, n2975, n2361 );
nand U3919 ( n3518, n3383, n3101 );
nand U3920 ( n3383, n3520, n3521 );
or U3921 ( n3521, n3391, n4515 );
nand U3922 ( n3520, n3522, n3391 );
xnor U3923 ( n3522, n4696, n3523 );
nor U3924 ( n3523, n2433, n3517 );
nand U3925 ( n3517, n3524, n4701 );
nand U3926 ( new_g11482_, n3525, n3526 );
nand U3927 ( n3526, n2975, n2362 );
nand U3928 ( n3525, n3386, n3101 );
nand U3929 ( n3386, n3527, n3528 );
or U3930 ( n3528, n3391, n4514 );
nand U3931 ( n3527, n3529, n3391 );
xnor U3932 ( n3529, n4645, n3530 );
nor U3933 ( n3530, n4701, n3394 );
nand U3934 ( n3394, n3531, n4702 );
nor U3935 ( n3531, n4700, n2246 );
nand U3936 ( new_g11481_, n3532, n3533 );
nand U3937 ( n3533, n2975, n2363 );
nand U3938 ( n3532, n3385, n3101 );
nand U3939 ( n3385, n3534, n3535 );
or U3940 ( n3535, n3391, n4516 );
nand U3941 ( n3534, n3536, n3391 );
xnor U3942 ( n3536, n4644, n3537 );
nor U3943 ( n3537, n2262, n3510 );
nand U3944 ( n3510, n3538, n4700 );
nor U3945 ( n3538, n4701, n2246 );
nand U3946 ( new_g11478_, n3539, n3540 );
nand U3947 ( n3540, n2975, n2364 );
not U3948 ( n2975, n3101 );
nand U3949 ( n3539, n3371, n3101 );
nand U3950 ( n3371, n3541, n3542 );
or U3951 ( n3542, n3391, n4521 );
nand U3952 ( n3541, n3543, n3391 );
xnor U3953 ( n3543, n4697, n3544 );
nor U3954 ( n3544, n4701, n3497 );
nand U3955 ( n3497, n3545, n4700 );
nor U3956 ( n3545, n4703, n2262 );
nor U3957 ( new_g11393_, n3546, n3547 );
xnor U3958 ( n3547, n4601, n3548 );
nand U3959 ( n3548, n3549, n2227 );
nor U3960 ( new_g11392_, n3546, n3550 );
xnor U3961 ( n3550, n2227, n3549 );
nor U3962 ( n3549, n3551, n4665 );
nor U3963 ( new_g11391_, n3546, n3552 );
xnor U3964 ( n3552, n4665, n3551 );
nand U3965 ( n3551, new_g10788_, n2264 );
nor U3966 ( new_g11380_, n3553, n3554 );
nor U3967 ( n3553, n3555, n2246 );
nor U3968 ( n3555, n3503, n3556 );
nand U3969 ( n3503, n3524, n3557 );
nor U3970 ( n3524, n4702, n2246 );
nor U3971 ( new_g11376_, n3554, n3558 );
xnor U3972 ( n3558, n4702, n3559 );
nand U3973 ( n3559, n3560, n2203 );
nor U3974 ( new_g11372_, n3554, n3561 );
xnor U3975 ( n3561, n2203, n3560 );
nor U3976 ( n3560, n3556, n4700 );
nor U3977 ( new_g11349_, n3546, n3562 );
xnor U3978 ( n3562, n2264, new_g10788_ );
nand U3979 ( n3546, g109, n3563 );
nand U3980 ( n3563, n3564, n3565 );
nor U3981 ( n3564, n4502, n3566 );
nor U3982 ( new_g11340_, n3554, n3567 );
xnor U3983 ( n3567, n4700, n3556 );
nand U3984 ( n3556, n3391, n3568 );
nand U3985 ( n3568, n3569, n3557 );
nor U3986 ( n3557, n4700, n4701 );
nor U3987 ( n3569, n4702, n4703 );
nand U3988 ( n3554, n4499, g109 );
nor U3989 ( new_g11320_, n3570, n3571 );
xnor U3990 ( n3571, n4559, n3572 );
nand U3991 ( new_g11314_, n3573, n3574 );
nand U3992 ( n3574, n3575, n2431 );
or U3993 ( n3573, n3575, n4621 );
nand U3994 ( new_g11312_, n3576, n3577 );
or U3995 ( n3577, n3578, n4563 );
or U3996 ( n3576, n3575, n4569 );
nand U3997 ( new_g11310_, n3579, n3580 );
or U3998 ( n3580, n3578, n4680 );
or U3999 ( n3579, n3575, n4598 );
nand U4000 ( new_g11308_, n3581, n3582 );
or U4001 ( n3582, n3578, n4562 );
nand U4002 ( n3581, n3578, n2412 );
nand U4003 ( new_g11306_, n3583, n3584 );
or U4004 ( n3584, n3578, n4561 );
nand U4005 ( n3583, n3578, n2425 );
nand U4006 ( new_g11305_, n3585, n3586 );
nand U4007 ( n3586, n3575, n2239 );
or U4008 ( n3585, n3575, n4630 );
nand U4009 ( new_g11303_, n3587, n3588 );
or U4010 ( n3588, n3578, n4641 );
nand U4011 ( n3587, n3578, n2401 );
nand U4012 ( new_g11300_, n3589, n3590 );
nand U4013 ( n3590, n3575, n2240 );
or U4014 ( n3589, n3575, n4573 );
nand U4015 ( new_g11298_, n3591, n3592 );
nand U4016 ( n3592, n3575, n2430 );
not U4017 ( n3575, n3578 );
nand U4018 ( n3591, n3578, n2408 );
nand U4019 ( n3578, n3593, new_g10788_ );
nor U4020 ( n3593, n3566, n3594 );
nor U4021 ( n3594, n2784, n3565 );
not U4022 ( n3566, n3595 );
nand U4023 ( new_g11294_, n3596, n3597 );
nand U4024 ( n3597, n3598, n2678 );
nor U4025 ( n3598, n3599, n3600 );
nor U4026 ( n3600, n2197, n3601 );
nand U4027 ( n3601, n3602, n3603 );
nand U4028 ( n3603, n3604, n3605 );
nand U4029 ( n3605, n2270, n2198 );
nand U4030 ( n3604, n2241, n2218 );
nand U4031 ( n3602, n3279, n2967 );
nand U4032 ( n2967, n2285, n2217 );
nand U4033 ( n3279, n2200, n2276 );
nor U4034 ( n3599, n4730, n3606 );
nand U4035 ( n3606, n3607, n3608 );
nand U4036 ( n3608, n3609, n3610 );
nand U4037 ( n3610, new_g10719_, new_g10720_ );
nand U4038 ( n3609, new_g10721_, new_g10722_ );
nand U4039 ( n3607, n3611, n3612 );
nand U4040 ( n3612, new_g10663_, new_g10664_ );
nor U4041 ( n3596, n3613, n3614 );
nor U4042 ( n3614, n2282, n3615 );
nand U4043 ( n3615, n2673, n2506 );
nand U4044 ( n2506, n3616, n4550 );
and U4045 ( n3616, n2499, n2496 );
nor U4046 ( n3613, n4720, n3060 );
not U4047 ( n3060, n3035 );
nor U4048 ( n3035, n2678, n2673 );
not U4049 ( n2673, n2487 );
nand U4050 ( new_g11293_, n3617, n3618 );
nand U4051 ( n3618, n3619, n2493 );
nand U4052 ( n3619, n2496, n3620 );
nand U4053 ( n3620, n3621, g1854 );
nand U4054 ( n3621, n3622, n3623 );
xnor U4055 ( n3623, n3624, n3625 );
nor U4056 ( n3625, n3626, n3627 );
nor U4057 ( n3627, n4720, n2220 );
nor U4058 ( n3626, n3628, n2282 );
and U4059 ( n3628, n2499, n4715 );
nor U4060 ( n3622, n3629, n3306 );
nand U4061 ( n3306, n3063, g1850 );
not U4062 ( n3063, new_g3524_ );
nand U4063 ( new_g3524_, n2493, n3630 );
or U4064 ( n3630, n2220, n4715 );
nor U4065 ( n3629, n3631, n3632 );
nand U4066 ( n3632, n4715, n4550 );
nand U4067 ( n3631, n2675, n2499 );
nand U4068 ( n2499, n2253, n2220 );
nand U4069 ( n2675, n3633, n3634 );
nor U4070 ( n3633, n4717, n2303 );
nand U4071 ( n2496, n3635, n4717 );
nor U4072 ( n3635, n4718, n2202 );
nand U4073 ( n3617, n3636, n2678 );
nand U4074 ( n3636, n3637, n3638 );
nand U4075 ( n3638, n3639, n2197 );
nand U4076 ( n3637, n4730, n4501 );
nor U4077 ( new_g11292_, n3640, n3570 );
nor U4078 ( n3640, n3641, n2469 );
nor U4079 ( n3641, n4707, n3642 );
nor U4080 ( new_g11291_, n3570, n3643 );
xnor U4081 ( n3643, n4707, n3642 );
nand U4082 ( n3642, n3644, n2302 );
nor U4083 ( new_g11290_, n3570, n3645 );
xnor U4084 ( n3645, n2302, n3644 );
nor U4085 ( n3644, n3572, n4559 );
nand U4086 ( n3572, n3391, n3646 );
nand U4087 ( n3570, n4502, g109 );
nand U4088 ( new_g10936_, n3647, n3648 );
nand U4089 ( n3648, n2987, n2447 );
nand U4090 ( n3647, n3304, n3649 );
nand U4091 ( n3649, n3650, n3651 );
nor U4092 ( n3651, new_g10719_, n3652 );
nand U4093 ( n3652, n3653, n3654 );
nor U4094 ( n3650, n3624, n3655 );
nand U4095 ( n3655, n3481, new_g10722_ );
nand U4096 ( new_g10898_, n3656, n3657 );
nand U4097 ( n3657, n2774, n2342 );
nand U4098 ( n3656, n2775, n3658 );
nand U4099 ( n3658, n3659, n3355 );
xor U4100 ( n3659, n3660, n3661 );
xor U4101 ( n3661, n3662, n3663 );
xor U4102 ( n3663, n3664, n3665 );
xor U4103 ( n3665, n4509, n4510 );
xor U4104 ( n3664, n4507, n4508 );
xor U4105 ( n3662, n3666, n3667 );
xnor U4106 ( n3667, n2299, n4506 );
xnor U4107 ( n3666, n2300, n4504 );
xnor U4108 ( n3660, n4544, n4511 );
nand U4109 ( new_g10866_, n3668, n3669 );
nand U4110 ( n3669, n2774, n2365 );
nand U4111 ( new_g10865_, n3670, n3671 );
nand U4112 ( n3671, n3197, n2366 );
nand U4113 ( n3670, n3672, n3196 );
nor U4114 ( n3672, n3673, n3674 );
nor U4115 ( n3673, new_g10722_, n2784 );
nand U4116 ( new_g10864_, n3675, n3676 );
nand U4117 ( n3676, n2774, n2367 );
nand U4118 ( new_g10863_, n3677, n3678 );
nand U4119 ( n3678, n3197, n2368 );
nand U4120 ( n3677, n3679, n3196 );
nor U4121 ( n3679, n3680, n3681 );
nor U4122 ( n3681, n3682, n2267 );
nor U4123 ( n3682, n3654, n2784 );
nand U4124 ( new_g10862_, n3683, n3684 );
nand U4125 ( n3684, n2774, n2369 );
nand U4126 ( new_g10861_, n3685, n3686 );
nand U4127 ( n3686, n3197, n2370 );
nand U4128 ( n3685, n3196, n3687 );
nand U4129 ( new_g10860_, n3688, n3689 );
nand U4130 ( n3689, n2774, n2371 );
nand U4131 ( new_g10859_, n3690, n3691 );
nand U4132 ( n3691, n3197, n2372 );
nand U4133 ( n3690, n3196, n3692 );
nand U4134 ( new_g10858_, n3693, n3694 );
nand U4135 ( n3694, n2774, n2373 );
nand U4136 ( new_g10855_, n3695, n3696 );
nand U4137 ( n3696, n2774, n2374 );
nand U4138 ( n3695, n2775, n3687 );
nand U4139 ( n3687, n3697, n4710 );
nor U4140 ( n3697, n3698, n3699 );
nor U4141 ( n3699, n3700, n2927 );
and U4142 ( n2927, n3701, n3215 );
nand U4143 ( n3215, g18, n2319 );
nand U4144 ( n3701, n2472, n2375 );
nor U4145 ( n3698, n3680, n3702 );
nand U4146 ( new_g10800_, n3703, n3704 );
nand U4147 ( n3704, n2774, n2376 );
nand U4148 ( n3703, n2775, n3692 );
nand U4149 ( n3692, n3705, n3706 );
not U4150 ( n3706, n3707 );
nor U4151 ( n3705, n3708, n3709 );
nor U4152 ( n3709, n3700, n2922 );
and U4153 ( n2922, n3710, n3217 );
nand U4154 ( n3217, g18, n2459 );
nand U4155 ( n3710, n2472, n2377 );
nor U4156 ( n3708, n3680, n3639 );
nand U4157 ( new_g10799_, n3711, n3712 );
nand U4158 ( n3712, n2774, n2378 );
nand U4159 ( new_g10798_, n3668, n3713 );
nand U4160 ( n3713, n2774, n2379 );
nand U4161 ( n3668, n2775, n3714 );
nand U4162 ( n3714, n3715, n3716 );
nand U4163 ( n3716, n3680, n2925 );
nand U4164 ( n2925, n2797, n3717 );
nand U4165 ( n3717, n2472, n2380 );
or U4166 ( n2797, n2472, n4763 );
nand U4167 ( n3715, n3718, n3624 );
nand U4168 ( new_g10797_, n3675, n3719 );
nand U4169 ( n3719, n2774, n2381 );
nand U4170 ( n3675, n3720, n3721 );
nor U4171 ( n3721, n3722, n3723 );
nor U4172 ( n3723, n3700, n2920 );
nand U4173 ( n2920, n2788, n3724 );
nand U4174 ( n3724, n2472, n2382 );
or U4175 ( n2788, n2472, n4765 );
nor U4176 ( n3722, new_g10722_, n3680 );
nand U4177 ( new_g10795_, n3683, n3725 );
nand U4178 ( n3725, n2774, n2383 );
nand U4179 ( n3683, n3720, n3726 );
nor U4180 ( n3726, n3727, n3728 );
nor U4181 ( n3728, n3700, n2912 );
nand U4182 ( n2912, n2835, n3729 );
nand U4183 ( n3729, n2472, n2384 );
nand U4184 ( n2835, g18, n2320 );
nor U4185 ( n3727, new_g10721_, n3680 );
nor U4186 ( n3720, n2774, n3707 );
nand U4187 ( n3707, n4710, n3730 );
nand U4188 ( n3730, n3700, n2784 );
nand U4189 ( new_g10793_, n3688, n3731 );
nand U4190 ( n3731, n2774, n2385 );
nand U4191 ( n3688, n3732, n2775 );
nor U4192 ( n3732, n3733, n3734 );
nor U4193 ( n3734, n2908, n3700 );
nand U4194 ( n2908, n2822, n3735 );
nand U4195 ( n3735, n2472, n2386 );
or U4196 ( n2822, n2472, n4769 );
nor U4197 ( n3733, n3674, n3736 );
nand U4198 ( n3736, g109, n3653 );
not U4199 ( n3674, n3718 );
nand U4200 ( new_g10791_, n3693, n3737 );
nand U4201 ( n3737, n2774, n2387 );
nand U4202 ( n3693, n2775, n3738 );
nand U4203 ( n3738, n3739, n3740 );
nand U4204 ( n3740, n3741, n3718 );
nand U4205 ( n3739, n3680, n2929 );
nand U4206 ( n2929, n2810, n3742 );
nand U4207 ( n3742, n2472, n2388 );
or U4208 ( n2810, n2472, n4771 );
and U4209 ( new_g10788_, n3743, n3744 );
nor U4210 ( n3743, n3389, n3745 );
nor U4211 ( n3745, n3746, n3747 );
nand U4212 ( n3747, n3748, n3749 );
nor U4213 ( n3749, n3750, n3751 );
nand U4214 ( n3751, n3752, n3753 );
xnor U4215 ( n3753, n4515, n4556 );
xnor U4216 ( n3752, n4519, n4557 );
xnor U4217 ( n3750, n4517, n2212 );
nor U4218 ( n3748, n3754, n3755 );
xnor U4219 ( n3755, n4521, n2256 );
xnor U4220 ( n3754, n4516, n2214 );
nand U4221 ( n3746, n3756, n3757 );
nor U4222 ( n3757, n3758, n3759 );
nand U4223 ( n3759, n3760, n3761 );
xnor U4224 ( n3761, n4513, n4704 );
xnor U4225 ( n3760, n3762, n2258 );
xnor U4226 ( n3758, n4520, n2213 );
nor U4227 ( n3756, n3763, n3764 );
xnor U4228 ( n3764, n4518, n2244 );
xnor U4229 ( n3763, n4514, n2207 );
nor U4230 ( new_g10785_, n4522, n3304 );
nor U4231 ( new_g10784_, n4523, n3304 );
nor U4232 ( new_g10782_, n4524, n3304 );
nor U4233 ( new_g10780_, n4525, n3304 );
not U4234 ( n3304, n2987 );
nand U4235 ( n2987, n4546, n2250 );
xnor U4236 ( g11163, n3765, n3 );
nand U4237 ( new_g10776_, n3711, n3766 );
nand U4238 ( n3766, n2774, n2389 );
nand U4239 ( n3711, n2775, n3767 );
nand U4240 ( n3767, n3768, n3769 );
nand U4241 ( n3769, n3680, n2931 );
nand U4242 ( n2931, n2816, n3770 );
nand U4243 ( n3770, n2472, n2390 );
nand U4244 ( n2816, g18, n2321 );
nand U4245 ( n3768, n3718, n3771 );
nand U4246 ( n3771, g109, n3482 );
nand U4247 ( new_g10773_, n3772, n3773 );
nand U4248 ( n3773, n3774, new_g10721_ );
nand U4249 ( n3772, n3775, n2424 );
nand U4250 ( new_g10771_, n3776, n3777 );
nand U4251 ( n3777, n3774, new_g10720_ );
or U4252 ( n3776, n3778, n4631 );
nand U4253 ( new_g10770_, n3779, n3780 );
nand U4254 ( n3780, n3774, new_g10719_ );
nand U4255 ( n3779, n3775, n2402 );
nand U4256 ( new_g10767_, n3781, n3782 );
nand U4257 ( n3782, n3197, n2391 );
nand U4258 ( n3781, n3196, n3783 );
nand U4259 ( new_g10765_, n3784, n3785 );
nand U4260 ( n3785, n3197, n2392 );
not U4261 ( n3197, n3196 );
nand U4262 ( n3784, n3196, n3786 );
nand U4263 ( new_g10718_, n3787, n3788 );
nand U4264 ( n3788, n2774, n2393 );
nand U4265 ( n3787, n2775, n3783 );
nand U4266 ( n3783, n3789, n4710 );
nor U4267 ( n3789, n3790, n3791 );
nor U4268 ( n3791, n3700, n2914 );
and U4269 ( n2914, n3792, n3219 );
nand U4270 ( n3219, g18, n2458 );
nand U4271 ( n3792, n2472, n2394 );
nor U4272 ( n3790, n3680, n3793 );
nand U4273 ( n3793, g109, new_g10664_ );
nand U4274 ( new_g10717_, n3794, n3795 );
nand U4275 ( n3795, n2774, n2395 );
nand U4276 ( n3794, n2775, n3786 );
nand U4277 ( n3786, n3796, n3797 );
nand U4278 ( n3797, n3718, n3798 );
nand U4279 ( n3798, g109, n3799 );
nor U4280 ( n3718, n2267, n3680 );
nand U4281 ( n3796, n3680, n2933 );
nand U4282 ( n2933, n2828, n3800 );
nand U4283 ( n3800, n2472, n2396 );
or U4284 ( n2828, n2472, n4759 );
not U4285 ( n3680, n3700 );
nand U4286 ( n3700, n4526, n4710 );
nand U4287 ( g10801, n3801, n3802 );
nand U4288 ( new_g10711_, n3803, n3804 );
nand U4289 ( n3804, n3778, n3624 );
nand U4290 ( n3624, g109, n3805 );
or U4291 ( n3803, n3778, n4595 );
nand U4292 ( new_g10707_, n3806, n3807 );
nand U4293 ( n3807, n3774, new_g10722_ );
nor U4294 ( n3774, n3775, n2784 );
nand U4295 ( n3806, n3775, n2411 );
not U4296 ( n3775, n3778 );
nor U4297 ( n3778, n4546, n4708 );
nor U4298 ( g11206, n3808, n3765 );
nand U4299 ( n3765, n3809, n3810 );
nand U4300 ( n3810, g109, n3811 );
nand U4301 ( n3811, n3812, n3813 );
or U4302 ( n3813, n3239, n3805 );
nand U4303 ( n3239, n4528, g3069 );
nand U4304 ( n3812, new_g10664_, g2648 );
and U4305 ( n3809, n3814, n3815 );
nand U4306 ( n3815, new_g5392_, new_g10663_ );
nor U4307 ( new_g5392_, n3316, n2784 );
nand U4308 ( n3316, n2259, g1765 );
nor U4309 ( n3814, n3816, n3817 );
nor U4310 ( n3817, n3818, n3367 );
nand U4311 ( n3367, g109, g108 );
nor U4312 ( n3816, n2342, n3819 );
nand U4313 ( n3819, g109, new_g10726_ );
not U4314 ( g10628, n3808 );
nand U4315 ( n3808, n3820, n3821 );
nor U4316 ( n3821, n3822, n3823 );
nand U4317 ( n3823, n3824, n3825 );
nand U4318 ( n3825, n3741, g877 );
nor U4319 ( n3741, n3639, n2784 );
nand U4320 ( n3824, n3826, n3827 );
not U4321 ( n3827, n3565 );
nand U4322 ( n3565, n4530, g3007 );
nor U4323 ( n3826, n3805, n2784 );
nor U4324 ( n3822, n3818, n3595 );
nand U4325 ( n3595, g109, g757 );
nor U4326 ( n3820, n3828, n3829 );
nor U4327 ( n3829, n3830, n3702 );
nand U4328 ( n3702, g109, new_g10720_ );
nor U4329 ( n3828, n3831, n3832 );
nand U4330 ( n3832, n4531, g109 );
nand U4331 ( n3831, new_g10721_, g2986 );
nand U4332 ( g10465, n3801, n3482 );
nand U4333 ( g10463, n3801, n3805 );
nand U4334 ( g10461, n3801, n3818 );
not U4335 ( n3818, new_g10722_ );
nand U4336 ( g10459, n3801, n3654 );
not U4337 ( n3654, new_g10721_ );
nand U4338 ( g10457, n3801, n3653 );
nand U4339 ( g10455, n3801, n3639 );
not U4340 ( n3639, new_g10719_ );
nand U4341 ( g10379, n3801, n3833 );
nand U4342 ( g10377, n3801, n3799 );
nor U4343 ( n3801, n3834, g30 );
and U4344 ( n68, n3084, g632 );
not U4345 ( n3084, new_g4117_ );
nand U4346 ( new_g4117_, n2517, n3835 );
nand U4347 ( n3835, n4683, n2245 );
nand U4348 ( n44, g109, n3836 );
nand U4349 ( n3836, n3830, n3837 );
nand U4350 ( n3837, n4531, g2986 );
not U4351 ( n3830, g881 );
not U4352 ( n3, n3802 );
xnor U4353 ( n3802, n3838, n3839 );
xor U4354 ( n3839, n3840, n3841 );
xnor U4355 ( n3841, n3799, n3842 );
nand U4356 ( n3842, n3611, n3843 );
nand U4357 ( n3843, n3805, n3482 );
not U4358 ( n3482, new_g10726_ );
not U4359 ( n3805, n7 );
nand U4360 ( n3611, new_g10726_, n7 );
xnor U4361 ( n3840, new_g10719_, n3833 );
not U4362 ( n3833, new_g10664_ );
xor U4363 ( n3838, n3844, n3845 );
xnor U4364 ( n3845, new_g10721_, n3653 );
not U4365 ( n3653, new_g10720_ );
xnor U4366 ( n3844, n3846, new_g10722_ );
nand U4367 ( n3846, n4527, n3834 );
nand U4368 ( n2206, n3847, n3848 );
nand U4369 ( n3848, n3849, n2325 );
nand U4370 ( n3847, n3850, n2313 );
nand U4371 ( n2201, n3851, n3852 );
nand U4372 ( n3852, n3849, n2313 );
nand U4373 ( n3851, n3850, n2290 );
nand U4374 ( n2196, n3853, n3854 );
nand U4375 ( n3854, n3849, n2290 );
nand U4376 ( n3853, n3850, n2233 );
xor U4377 ( n2192, n3855, n4532 );
nand U4378 ( n3855, n2891, g4181 );
nor U4379 ( n2891, n2937, n4533 );
or U4380 ( n2937, n2944, n4675 );
or U4381 ( n2944, n2979, n4534 );
or U4382 ( n2979, n3068, n4535 );
or U4383 ( n3068, n3193, n4674 );
nand U4384 ( n3193, n3856, g4174 );
nor U4385 ( n3856, n4536, n4672 );
nand U4386 ( n2191, n3857, n3858 );
nand U4387 ( n3858, n3849, n2233 );
nand U4388 ( n3857, n3850, n2278 );
nand U4389 ( n2190, n3859, n3860 );
nor U4390 ( n3859, n4640, g47 );
nand U4391 ( n2189, n3861, g46 );
nand U4392 ( n2188, n3862, n3860 );
and U4393 ( n3860, n3863, n3864 );
nor U4394 ( n3864, g45, n3865 );
nand U4395 ( n3865, n4663, n3866 );
nor U4396 ( n3863, g42, n3867 );
nand U4397 ( n3867, n4659, n4660 );
nor U4398 ( n3862, n4662, g46 );
nand U4399 ( n2187, n3868, n3869 );
nand U4400 ( n2186, n3870, n3871 );
nand U4401 ( n3871, n3849, n2278 );
nand U4402 ( n3870, n3850, n2332 );
nand U4403 ( n2181, n3872, n3873 );
nand U4404 ( n3873, n3849, n2332 );
nand U4405 ( n3872, n3850, n2255 );
nand U4406 ( n2176, n3874, n3875 );
nand U4407 ( n3875, n3849, n2255 );
nand U4408 ( n3874, n3850, n2210 );
nand U4409 ( n2171, n3876, n3877 );
nand U4410 ( n3877, n3849, n2210 );
nand U4411 ( n3876, n3850, n2243 );
nand U4412 ( n2166, n3878, n3879 );
nand U4413 ( n3879, n3849, n2243 );
nand U4414 ( n3878, n3850, n2271 );
nand U4415 ( n2161, n3880, n3881 );
nand U4416 ( n3881, n3849, n2271 );
nand U4417 ( n3880, n3850, n2272 );
nand U4418 ( n2156, n3882, n3883 );
nand U4419 ( n3883, n3849, n2272 );
nand U4420 ( n3882, n3850, n2209 );
nand U4421 ( n2151, n3884, n3885 );
nand U4422 ( n3885, n3849, n2209 );
nand U4423 ( n3884, n3850, n2307 );
nand U4424 ( n2146, n3886, n3887 );
nand U4425 ( n3887, n3849, n2307 );
nand U4426 ( n3886, n3850, n2205 );
nand U4427 ( n2141, n3888, n3889 );
nand U4428 ( n3889, n3849, n2205 );
nand U4429 ( n3888, n3850, n2211 );
nand U4430 ( n2136, n3890, n3891 );
nand U4431 ( n3891, n3849, n2211 );
nand U4432 ( n3890, n3850, n3458 );
nand U4433 ( n3458, n3892, n3893 );
or U4434 ( n3893, n3459, n2964 );
xor U4435 ( n3459, n3894, n2298 );
nand U4436 ( n3894, n2432, n3355 );
nand U4437 ( n3355, n3481, n3799 );
not U4438 ( n3799, new_g10663_ );
nand U4439 ( n3481, n3861, n4640 );
and U4440 ( n3861, n3895, n3868 );
and U4441 ( n3868, n3896, n3897 );
nor U4442 ( n3897, g48, g45 );
nor U4443 ( n3896, g43, n3898 );
nor U4444 ( n3895, n2471, g47 );
nand U4445 ( n3892, n3899, n2964 );
and U4446 ( n2964, n3900, n3901 );
nor U4447 ( n3901, n4541, n4542 );
nor U4448 ( n3900, n4543, n4735 );
nand U4449 ( n3899, n3902, n3903 );
nand U4450 ( n3903, n4733, n2325 );
nand U4451 ( n3902, n4734, n3904 );
nand U4452 ( n3904, n4733, n3905 );
nand U4453 ( n3905, n3906, n3907 );
nor U4454 ( n3907, n3908, n3909 );
nand U4455 ( n3909, n3910, n4539 );
nor U4456 ( n3910, n2271, n2209 );
nand U4457 ( n3908, n3911, n3912 );
nor U4458 ( n3912, n2272, n2210 );
nor U4459 ( n3911, n2205, n2243 );
nor U4460 ( n3906, n3913, n3914 );
nand U4461 ( n3914, n3915, n4537 );
nor U4462 ( n3915, n2278, n2211 );
nand U4463 ( n3913, n3916, n4538 );
nor U4464 ( n3916, n2233, n2290 );
not U4465 ( n3850, n2963 );
nand U4466 ( n2963, n3917, n4709 );
nor U4467 ( n3917, n4545, n2774 );
nor U4468 ( n192, n4469, n2784 );
nor U4469 ( n186, n4466, n2784 );
nand U4470 ( n1845, n3918, n3919 );
nand U4471 ( n3919, n3920, n2455 );
nand U4472 ( n3918, n2484, n2291 );
nand U4473 ( n1840, n3921, n3922 );
nand U4474 ( n3922, n3920, n2291 );
nand U4475 ( n3921, n2484, n2335 );
nand U4476 ( n1835, n3923, n3924 );
nand U4477 ( n3924, n3920, n2335 );
nand U4478 ( n3923, n2484, n2286 );
nand U4479 ( n1830, n3925, n3926 );
nand U4480 ( n3926, n3920, n2286 );
nand U4481 ( n3925, n2484, n2336 );
nand U4482 ( n1825, n3927, n3928 );
nand U4483 ( n3928, n3920, n2336 );
nand U4484 ( n3927, n2484, n2337 );
nand U4485 ( n1820, n3929, n3930 );
nand U4486 ( n3930, n3920, n2337 );
nand U4487 ( n3929, n2484, n2287 );
nand U4488 ( n1815, n3931, n3932 );
nand U4489 ( n3932, n3920, n2287 );
nand U4490 ( n3931, n2484, n2248 );
nand U4491 ( n1810, n3933, n3934 );
nand U4492 ( n3934, n3920, n2248 );
nor U4493 ( n3920, n2678, n2484 );
not U4494 ( n2678, n2493 );
nand U4495 ( n2493, n3634, n4717 );
and U4496 ( n3634, n3935, n4715 );
nor U4497 ( n3935, n2253, n2202 );
nand U4498 ( n3933, n2484, n2326 );
not U4499 ( n2484, n2872 );
nand U4500 ( n2872, n3936, n4715 );
nor U4501 ( n3936, n4716, n2487 );
nand U4502 ( n2487, n4553, n3037 );
and U4503 ( n3037, n4721, n3062 );
and U4504 ( n3062, n4552, n2445 );
nand U4505 ( n1449, n3937, n3938 );
nand U4506 ( n3938, n3389, n2327 );
nand U4507 ( n3937, n3391, n2314 );
nand U4508 ( n1444, n3939, n3940 );
nand U4509 ( n3940, n3389, n2314 );
nand U4510 ( n3939, n3391, n2292 );
nand U4511 ( n1439, n3941, n3942 );
nand U4512 ( n3942, n3389, n2292 );
nand U4513 ( n3941, n3391, n2234 );
nand U4514 ( n1434, n3943, n3944 );
nand U4515 ( n3944, n3389, n2234 );
nand U4516 ( n3943, n3391, n2279 );
nand U4517 ( n1429, n3945, n3946 );
nand U4518 ( n3946, n3389, n2279 );
nand U4519 ( n3945, n3391, n2333 );
nand U4520 ( n1424, n3947, n3948 );
nand U4521 ( n3948, n3389, n2333 );
nand U4522 ( n3947, n3391, n2256 );
nand U4523 ( n1419, n3949, n3950 );
nand U4524 ( n3950, n3389, n2256 );
nand U4525 ( n3949, n3391, n2213 );
nand U4526 ( n1414, n3951, n3952 );
nand U4527 ( n3952, n3389, n2213 );
nand U4528 ( n3951, n3391, n2244 );
nand U4529 ( n1409, n3953, n3954 );
nand U4530 ( n3954, n3389, n2244 );
nand U4531 ( n3953, n3391, n2273 );
nand U4532 ( n1404, n3955, n3956 );
nand U4533 ( n3956, n3389, n2273 );
nand U4534 ( n3955, n3391, n2274 );
nand U4535 ( n1399, n3957, n3958 );
nand U4536 ( n3958, n3389, n2274 );
nand U4537 ( n3957, n3391, n2212 );
nand U4538 ( n1394, n3959, n3960 );
nand U4539 ( n3960, n3389, n2212 );
nand U4540 ( n3959, n3391, n2308 );
nand U4541 ( n1389, n3961, n3962 );
nand U4542 ( n3962, n3389, n2308 );
nand U4543 ( n3961, n3391, n2207 );
nand U4544 ( n1384, n3963, n3964 );
nand U4545 ( n3964, n3389, n2207 );
nand U4546 ( n3963, n3391, n2214 );
nand U4547 ( n1379, n3965, n3966 );
nand U4548 ( n3966, n3389, n2214 );
nand U4549 ( n3965, n3762, n3391 );
nand U4550 ( n3762, n3967, n3968 );
nand U4551 ( n3968, n3646, n2258 );
nand U4552 ( n3967, n3969, n3744 );
not U4553 ( n3744, n3646 );
nand U4554 ( n3646, n3970, n3971 );
nor U4555 ( n3971, n4558, n4559 );
nor U4556 ( n3970, n4560, n4707 );
nand U4557 ( n3969, n3972, n3973 );
nand U4558 ( n3973, n4705, n2327 );
nand U4559 ( n3972, n4706, n3974 );
nand U4560 ( n3974, n4705, n3975 );
nand U4561 ( n3975, n3976, n3977 );
nor U4562 ( n3977, n3978, n3979 );
nand U4563 ( n3979, n3980, n4556 );
nor U4564 ( n3980, n2273, n2212 );
nand U4565 ( n3978, n3981, n3982 );
nor U4566 ( n3982, n2274, n2213 );
nor U4567 ( n3981, n2207, n2244 );
nor U4568 ( n3976, n3983, n3984 );
nand U4569 ( n3984, n3985, n4554 );
nor U4570 ( n3985, n2279, n2214 );
nand U4571 ( n3983, n3986, n4555 );
nor U4572 ( n3986, n2234, n2292 );
nand U4573 ( n1304, n3987, n3988 );
nand U4574 ( n3988, n3389, n2329 );
nand U4575 ( n3987, n3391, n2315 );
nand U4576 ( n1299, n3989, n3990 );
nand U4577 ( n3990, n3389, n2315 );
nand U4578 ( n3989, n3391, n2293 );
nand U4579 ( n1294, n3991, n3992 );
nand U4580 ( n3992, n3389, n2293 );
nand U4581 ( n3991, n3391, n2236 );
nand U4582 ( n1289, n3993, n3994 );
nand U4583 ( n3994, n3389, n2236 );
nand U4584 ( n3993, n3391, n2280 );
nand U4585 ( n1284, n3995, n3996 );
nand U4586 ( n3996, n3389, n2280 );
nand U4587 ( n3995, n3391, n2334 );
nand U4588 ( n1279, n3997, n3998 );
nand U4589 ( n3998, n3389, n2334 );
nand U4590 ( n3997, n3391, n2275 );
nand U4591 ( n1274, n3999, n4000 );
nand U4592 ( n4000, n3389, n2275 );
nand U4593 ( n3999, n3391, n2216 );
nand U4594 ( n1269, n4001, n4002 );
nand U4595 ( n4002, n3389, n2216 );
nand U4596 ( n4001, n3391, n2309 );
nand U4597 ( n1264, n4003, n4004 );
nand U4598 ( n4004, n3389, n2309 );
nand U4599 ( n4003, n3391, n2215 );
nand U4600 ( n1259, n4005, n4006 );
nand U4601 ( n4006, n3389, n2215 );
nand U4602 ( n4005, n3391, n2284 );
nand U4603 ( n1254, n4007, n4008 );
nand U4604 ( n4008, n3389, n2284 );
nand U4605 ( n4007, n3391, n2231 );
nand U4606 ( n1249, n4009, n4010 );
nand U4607 ( n4010, n3389, n2231 );
nand U4608 ( n4009, n3391, n2232 );
nand U4609 ( n1244, n4011, n4012 );
nand U4610 ( n4012, n3389, n2232 );
nand U4611 ( n4011, n3391, n2283 );
nand U4612 ( n1239, n4013, n4014 );
nand U4613 ( n4014, n3389, n2283 );
nand U4614 ( n4013, n3391, n2310 );
nand U4615 ( n1234, n4015, n4016 );
nand U4616 ( n4016, n3389, n2310 );
nand U4617 ( n4015, n3393, n3391 );
nor U4618 ( n4018, n4019, n4020 );
nand U4619 ( n4020, n4021, n4641 );
nor U4620 ( n4021, n2239, n2430 );
nand U4621 ( n4019, n4022, n4680 );
nor U4622 ( n4022, n4023, n2784 );
nor U4623 ( n4023, n4024, n4025 );
nand U4624 ( n4025, n4026, n4027 );
nor U4625 ( n4027, new_g10719_, new_g10664_ );
nand U4626 ( new_g10664_, n4028, n4029 );
nor U4627 ( n4029, n4030, n4031 );
nand U4628 ( n4031, n4032, n4033 );
nand U4629 ( n4033, n4034, g1191 );
nand U4630 ( n4032, n4035, n2397 );
nand U4631 ( n4030, n4036, n4037 );
nand U4632 ( n4037, n4038, n2398 );
nor U4633 ( n4036, n4039, n4040 );
nor U4634 ( n4040, n4573, n4041 );
nor U4635 ( n4039, n4575, n4042 );
nor U4636 ( n4028, n4043, n4044 );
nand U4637 ( n4044, n4045, n4046 );
nand U4638 ( n4046, n3834, g40 );
nor U4639 ( n4045, n4047, n4048 );
nor U4640 ( n4048, n4049, n4050 );
nand U4641 ( n4050, n4051, n4052 );
nor U4642 ( n4047, n4574, n4053 );
nand U4643 ( n4043, n4054, n4055 );
nand U4644 ( n4055, n4056, n2399 );
nand U4645 ( n4054, n4057, n2400 );
nand U4646 ( new_g10719_, n4058, n4059 );
nor U4647 ( n4059, n4060, n4061 );
nand U4648 ( n4061, n4062, n4063 );
nor U4649 ( n4063, n4064, n4065 );
nand U4650 ( n4065, n4066, n4067 );
nand U4651 ( n4067, n4068, n2401 );
nand U4652 ( n4066, n4069, n2264 );
nor U4653 ( n4064, n4577, n4070 );
nor U4654 ( n4062, n4071, n4072 );
nand U4655 ( n4072, n4073, n4074 );
nand U4656 ( n4074, n4038, n2402 );
nand U4657 ( n4073, n4075, g1194 );
nor U4658 ( n4071, n4578, n4076 );
nand U4659 ( n4060, n4077, n4078 );
nor U4660 ( n4078, n4079, n4080 );
nand U4661 ( n4080, n4081, n4052 );
nor U4662 ( n4079, n4581, n4082 );
not U4663 ( n4082, n4083 );
nor U4664 ( n4077, n4084, n4085 );
nand U4665 ( n4085, n4086, n4087 );
nand U4666 ( n4087, n4049, n2219 );
nand U4667 ( n4086, n4088, g886 );
nor U4668 ( n4084, n4582, n4042 );
nor U4669 ( n4058, n4089, n4090 );
nand U4670 ( n4090, n4091, n4092 );
nor U4671 ( n4092, n4093, n4094 );
nand U4672 ( n4094, n4095, n4096 );
nand U4673 ( n4096, n4097, n2317 );
nand U4674 ( n4095, n4098, n2403 );
nor U4675 ( n4093, n4580, n4099 );
nor U4676 ( n4091, n4100, n4101 );
nor U4677 ( n4101, n4583, n4102 );
nor U4678 ( n4100, n4579, n4103 );
nand U4679 ( n4089, n4104, n4105 );
nor U4680 ( n4105, n4106, n4107 );
nand U4681 ( n4107, n4108, n4109 );
nand U4682 ( n4109, n4110, n2404 );
nand U4683 ( n4108, n4035, n2405 );
nor U4684 ( n4106, n4584, n4111 );
nor U4685 ( n4104, n4112, n4113 );
nand U4686 ( n4113, n4114, n4115 );
nand U4687 ( n4115, n4056, n2406 );
nand U4688 ( n4114, n4057, n2407 );
nor U4689 ( n4112, n4666, n4116 );
nor U4690 ( n4026, new_g10663_, n7 );
nand U4691 ( n7, n4117, n4118 );
nor U4692 ( n4118, n4119, n4120 );
nand U4693 ( n4120, n4121, n4122 );
nor U4694 ( n4122, n4123, n4124 );
nor U4695 ( n4124, n4593, n4125 );
nor U4696 ( n4123, n4592, n4076 );
nor U4697 ( n4121, n4126, n4127 );
nor U4698 ( n4127, n4591, n4128 );
nor U4699 ( n4126, n4590, n4129 );
nand U4700 ( n4119, n4130, n4131 );
nor U4701 ( n4131, n4132, n4133 );
nor U4702 ( n4133, n4597, n4099 );
nor U4703 ( n4132, n4598, n4134 );
nor U4704 ( n4130, n4135, n4136 );
nor U4705 ( n4136, n4595, n4137 );
nor U4706 ( n4135, n4594, n4070 );
nor U4707 ( n4117, n4138, n4139 );
nand U4708 ( n4139, n4140, n4141 );
nor U4709 ( n4141, n4142, n4143 );
nor U4710 ( n4143, n4599, n4144 );
nor U4711 ( n4142, n4097, n4145 );
nand U4712 ( n4145, n4146, n4147 );
not U4713 ( n4147, n4148 );
nor U4714 ( n4146, n4098, n4149 );
nor U4715 ( n4140, n4150, n4151 );
nor U4716 ( n4151, n4596, n4152 );
nor U4717 ( n4150, n4585, n4153 );
nand U4718 ( n4138, n4154, n4155 );
nor U4719 ( n4155, n4156, n4157 );
nor U4720 ( n4157, n4588, n4111 );
nor U4721 ( n4156, n4589, n4102 );
nor U4722 ( n4154, n4158, n4159 );
nor U4723 ( n4159, n4586, n4042 );
nor U4724 ( n4158, n4587, n4103 );
nand U4725 ( new_g10663_, n4160, n4161 );
nor U4726 ( n4161, n4162, n4163 );
nand U4727 ( n4163, n4164, n4165 );
nand U4728 ( n4165, n4034, g1188 );
not U4729 ( n4034, n4076 );
nor U4730 ( n4164, n4166, n4167 );
nor U4731 ( n4167, n4623, n4137 );
nor U4732 ( n4166, n4624, n4070 );
nand U4733 ( n4162, n4168, n4169 );
nand U4734 ( n4169, n4069, n2408 );
nor U4735 ( n4168, n4170, n4171 );
nor U4736 ( n4171, n4621, n4134 );
nor U4737 ( n4170, n4629, n4042 );
nor U4738 ( n4160, n4172, n4173 );
nand U4739 ( n4173, n4174, n4175 );
nor U4740 ( n4175, n4176, n4177 );
nor U4741 ( n4177, n4049, n4148 );
nor U4742 ( n4176, n4622, n4053 );
nor U4743 ( n4174, n4178, n4179 );
nor U4744 ( n4179, n4626, n4102 );
nor U4745 ( n4178, n4627, n4128 );
nand U4746 ( n4172, n4180, n4181 );
nand U4747 ( n4181, n4056, n2409 );
nor U4748 ( n4180, n4182, n4183 );
nor U4749 ( n4183, n4628, n4153 );
nor U4750 ( n4182, n4625, n4125 );
nand U4751 ( n4024, n4184, n4185 );
nor U4752 ( n4185, new_g10726_, new_g10722_ );
nand U4753 ( new_g10722_, n4186, n4187 );
nor U4754 ( n4187, n4188, n4189 );
nand U4755 ( n4189, n4190, n4191 );
nor U4756 ( n4191, n4192, n4193 );
nand U4757 ( n4193, n4194, n4195 );
nand U4758 ( n4195, n4196, n2410 );
nand U4759 ( n4194, n4038, n2411 );
nor U4760 ( n4192, n4602, n4197 );
nor U4761 ( n4190, n4198, n4199 );
nor U4762 ( n4199, n4604, n4125 );
nor U4763 ( n4198, n4603, n4076 );
nand U4764 ( n4188, n4200, n4201 );
nor U4765 ( n4201, n4202, n4203 );
nand U4766 ( n4203, n4204, n4081 );
nand U4767 ( n4204, n4049, n2266 );
nor U4768 ( n4202, n4600, n4205 );
nor U4769 ( n4200, n4206, n4207 );
nand U4770 ( n4207, n4208, n4209 );
nand U4771 ( n4209, n4210, g907 );
nand U4772 ( n4208, n4068, n2412 );
nor U4773 ( n4206, n4601, n4041 );
nor U4774 ( n4186, n4211, n4212 );
nand U4775 ( n4212, n4213, n4214 );
nor U4776 ( n4214, n4215, n4216 );
nand U4777 ( n4216, n4217, n4218 );
nand U4778 ( n4218, n4097, g17 );
nand U4779 ( n4217, n4098, g8 );
nor U4780 ( n4215, n4605, n4099 );
nor U4781 ( n4213, n4219, n4220 );
nor U4782 ( n4220, n4608, n4102 );
nor U4783 ( n4219, n4606, n4103 );
nand U4784 ( n4211, n4221, n4222 );
nor U4785 ( n4222, n4223, n4224 );
nand U4786 ( n4224, n4225, n4226 );
nand U4787 ( n4226, n4035, n2413 );
nand U4788 ( n4225, n4227, n2414 );
nor U4789 ( n4223, n4609, n4129 );
nor U4790 ( n4221, n4228, n4229 );
nor U4791 ( n4229, n4669, n4116 );
nor U4792 ( n4228, n4607, n4128 );
nand U4793 ( new_g10726_, n4230, n4231 );
nor U4794 ( n4231, n4232, n4233 );
nand U4795 ( n4233, n4234, n4235 );
nand U4796 ( n4235, n4035, n2415 );
nor U4797 ( n4234, n4236, n4237 );
nor U4798 ( n4237, n4566, n4125 );
nor U4799 ( n4236, n4567, n4076 );
nand U4800 ( n4232, n4238, n4239 );
nor U4801 ( n4239, n4240, n4241 );
nor U4802 ( n4241, n4572, n4042 );
nor U4803 ( n4240, n4149, n4148 );
nor U4804 ( n4238, n4242, n4243 );
nor U4805 ( n4243, n4570, n4070 );
nor U4806 ( n4242, n4569, n4134 );
nor U4807 ( n4230, n4244, n4245 );
nand U4808 ( n4245, n4246, n4247 );
nand U4809 ( n4247, n3834, g38 );
nor U4810 ( n4246, n4248, n4249 );
nor U4811 ( n4249, n4565, n4103 );
nor U4812 ( n4248, n4568, n4099 );
nand U4813 ( n4244, n4250, n4251 );
nand U4814 ( n4251, n4057, n2416 );
nor U4815 ( n4250, n4252, n4253 );
nor U4816 ( n4253, n4571, n4129 );
nor U4817 ( n4252, n4564, n4111 );
nor U4818 ( n4184, new_g10721_, new_g10720_ );
nand U4819 ( new_g10720_, n4254, n4255 );
nor U4820 ( n4255, n4256, n4257 );
nand U4821 ( n4257, n4258, n4259 );
nor U4822 ( n4259, n4260, n4261 );
nand U4823 ( n4261, n4262, n4263 );
nand U4824 ( n4263, n4069, n2322 );
nand U4825 ( n4262, n4196, n2417 );
nor U4826 ( n4260, n4631, n4137 );
nor U4827 ( n4258, n4264, n4265 );
nor U4828 ( n4265, n4633, n4076 );
nor U4829 ( n4264, n4632, n4197 );
nand U4830 ( n4256, n4266, n4267 );
nor U4831 ( n4267, n4268, n4269 );
nand U4832 ( n4269, n4270, n4081 );
nand U4833 ( n4270, n4083, g925 );
nor U4834 ( n4268, n4731, n4053 );
nor U4835 ( n4266, n4271, n4272 );
nand U4836 ( n4272, n4273, n4274 );
nand U4837 ( n4274, n4088, g889 );
nand U4838 ( n4273, n4210, g901 );
nor U4839 ( n4271, n4630, n4134 );
nor U4840 ( n4254, n4275, n4276 );
nand U4841 ( n4276, n4277, n4278 );
nor U4842 ( n4278, n4279, n4280 );
nand U4843 ( n4280, n4281, n4282 );
nand U4844 ( n4282, n4097, n2328 );
nand U4845 ( n4281, n4098, n2418 );
nor U4846 ( n4279, n4636, n4099 );
nor U4847 ( n4277, n4283, n4284 );
nor U4848 ( n4284, n4635, n4102 );
nor U4849 ( n4283, n4637, n4103 );
nand U4850 ( n4275, n4285, n4286 );
nor U4851 ( n4286, n4287, n4288 );
nand U4852 ( n4288, n4289, n4290 );
nand U4853 ( n4290, n4110, n2419 );
nand U4854 ( n4289, n4035, n2420 );
nor U4855 ( n4287, n4634, n4111 );
nor U4856 ( n4285, n4291, n4292 );
nand U4857 ( n4292, n4293, n4294 );
nand U4858 ( n4294, n4056, n2421 );
not U4859 ( n4056, n4129 );
nand U4860 ( n4293, n4057, n2422 );
not U4861 ( n4057, n4128 );
nor U4862 ( n4291, n4667, n4116 );
nand U4863 ( new_g10721_, n4295, n4296 );
nor U4864 ( n4296, n4297, n4298 );
nand U4865 ( n4298, n4299, n4300 );
nor U4866 ( n4300, n4301, n4302 );
nand U4867 ( n4302, n4303, n4304 );
nand U4868 ( n4304, n4196, n2423 );
nand U4869 ( n4303, n4038, n2424 );
not U4870 ( n4038, n4137 );
nor U4871 ( n4301, n4613, n4197 );
nor U4872 ( n4299, n4305, n4306 );
nor U4873 ( n4306, n4615, n4125 );
nor U4874 ( n4305, n4614, n4076 );
nand U4875 ( n4297, n4307, n4308 );
nor U4876 ( n4308, n4309, n4310 );
nand U4877 ( n4310, n4311, n4081 );
nand U4878 ( n4081, n4312, n4313 );
nor U4879 ( n4313, n4149, n4314 );
nand U4880 ( n4314, n4197, n4152 );
not U4881 ( n4197, n4075 );
nor U4882 ( n4075, n4315, n4316 );
not U4883 ( n4149, n4052 );
nand U4884 ( n4052, n4317, n4318 );
nor U4885 ( n4318, n2471, n4319 );
nand U4886 ( n4319, g47, g46 );
nor U4887 ( n4317, n4320, n4315 );
nor U4888 ( n4312, n4148, n4321 );
nand U4889 ( n4321, n4053, n4144 );
nand U4890 ( n4148, n4322, n4051 );
and U4891 ( n4051, n4323, n4324 );
nor U4892 ( n4324, n4325, n4326 );
nand U4893 ( n4326, n4327, n4134 );
and U4894 ( n4327, n4099, n4076 );
nand U4895 ( n4076, n4328, n4329 );
nand U4896 ( n4325, n4330, n4331 );
nor U4897 ( n4331, n4088, n4332 );
not U4898 ( n4088, n4205 );
nor U4899 ( n4330, n4083, n4333 );
nor U4900 ( n4083, n4315, n4334 );
nor U4901 ( n4323, n4335, n4336 );
nand U4902 ( n4336, n4337, n4102 );
nor U4903 ( n4337, n4069, n4338 );
nor U4904 ( n4338, n4339, n4340 );
nor U4905 ( n4339, n4341, n4329 );
not U4906 ( n4069, n4041 );
nand U4907 ( n4335, n4342, n4137 );
nand U4908 ( n4137, n4343, g42 );
and U4909 ( n4342, n4042, n4116 );
nor U4910 ( n4322, n4110, n4196 );
not U4911 ( n4196, n4070 );
nand U4912 ( n4070, n4343, n4658 );
and U4913 ( n4343, n4344, n4345 );
nor U4914 ( n4345, n4659, n4660 );
nor U4915 ( n4344, n4661, n4316 );
not U4916 ( n4110, n4125 );
nand U4917 ( n4125, n4328, n4346 );
nand U4918 ( n4311, n4049, n2311 );
not U4919 ( n4049, n4053 );
nand U4920 ( n4053, n4328, n4341 );
not U4921 ( n4328, n4316 );
nand U4922 ( n4316, n3869, n4347 );
and U4923 ( n3869, n4348, n4640 );
nor U4924 ( n4348, n4662, n2471 );
nor U4925 ( n4309, n4610, n4205 );
nand U4926 ( n4205, n4349, n4350 );
nor U4927 ( n4350, n4659, n4661 );
nor U4928 ( n4349, n4334, n3898 );
nor U4929 ( n4307, n4351, n4352 );
nand U4930 ( n4352, n4353, n4354 );
nand U4931 ( n4354, n4210, g904 );
not U4932 ( n4210, n4042 );
nand U4933 ( n4042, n4355, n4329 );
nand U4934 ( n4353, n4068, n2425 );
not U4935 ( n4068, n4134 );
nand U4936 ( n4134, n4346, n4355 );
nor U4937 ( n4351, n4611, n4041 );
nand U4938 ( n4041, n4341, n4355 );
not U4939 ( n4355, n4334 );
nor U4940 ( n4295, n4356, n4357 );
nand U4941 ( n4357, n4358, n4359 );
nor U4942 ( n4359, n4360, n4361 );
nand U4943 ( n4361, n4362, n4363 );
nand U4944 ( n4363, n4097, n2426 );
not U4945 ( n4097, n4144 );
nand U4946 ( n4144, n4364, n4365 );
nor U4947 ( n4364, g44, n4340 );
nand U4948 ( n4362, n4098, n2427 );
not U4949 ( n4098, n4152 );
nand U4950 ( n4152, n4366, n4367 );
nor U4951 ( n4366, n3898, n4340 );
nor U4952 ( n4360, n4616, n4099 );
nand U4953 ( n4099, n4368, n4346 );
and U4954 ( n4346, n4369, n4370 );
nor U4955 ( n4370, n4661, g44 );
nor U4956 ( n4369, g43, g42 );
nor U4957 ( n4358, n4371, n4372 );
nor U4958 ( n4372, n4619, n4102 );
nor U4959 ( n4371, n4617, n4103 );
not U4960 ( n4103, n4333 );
nor U4961 ( n4333, n4315, n4340 );
nand U4962 ( n4315, n4365, g44 );
and U4963 ( n4365, n4367, n4658 );
nor U4964 ( n4367, n4659, g45 );
nand U4965 ( n4356, n4373, n4374 );
nor U4966 ( n4374, n4375, n4376 );
nand U4967 ( n4376, n4377, n4378 );
nand U4968 ( n4378, n4035, n2428 );
not U4969 ( n4035, n4153 );
nand U4970 ( n4153, n4332, n4111 );
nand U4971 ( n4377, n4227, n2429 );
not U4972 ( n4227, n4111 );
nand U4973 ( n4111, n4332, n4658 );
and U4974 ( n4332, n4379, n4380 );
nor U4975 ( n4379, g43, n4340 );
nor U4976 ( n4375, n4620, n4129 );
nand U4977 ( n4129, n4368, n4341 );
nor U4978 ( n4341, n4381, n3898 );
nand U4979 ( n3898, n4660, g42 );
nand U4980 ( n4381, g45, n4659 );
nor U4981 ( n4373, n4382, n4383 );
nor U4982 ( n4383, n4668, n4116 );
nand U4983 ( n4116, n4384, n4385 );
nor U4984 ( n4385, n4661, n4386 );
nand U4985 ( n4386, g44, g42 );
nor U4986 ( n4384, n4334, g43 );
nand U4987 ( n4334, n4387, n4388 );
nor U4988 ( n4388, n4640, n2471 );
nor U4989 ( n4387, n4320, g47 );
nor U4990 ( n4382, n4618, n4128 );
nand U4991 ( n4128, n4368, n4329 );
and U4992 ( n4329, n4380, n4389 );
nor U4993 ( n4389, n4658, n4659 );
nor U4994 ( n4380, n4660, g45 );
not U4995 ( n4368, n4340 );
nand U4996 ( n4340, n4390, n4391 );
nor U4997 ( n4391, n2471, n4320 );
not U4998 ( n2471, n3866 );
nand U4999 ( n3866, n4392, n4393 );
nand U5000 ( n4393, n4394, n4638 );
nor U5001 ( n4394, g48, g30 );
nand U5002 ( n4392, n4102, n4347 );
not U5003 ( n4347, n4320 );
nand U5004 ( n4320, n4638, g48 );
not U5005 ( n4102, n3834 );
nand U5006 ( n3834, n4639, g48 );
nor U5007 ( n4390, g47, g46 );
nor U5008 ( n4017, n4395, n4396 );
nand U5009 ( n4396, n4561, n4562 );
nand U5010 ( n4395, n4397, n4563 );
nor U5011 ( n4397, n2240, n2431 );
nand U5012 ( n3393, n4398, n4399 );
nand U5013 ( n4399, n4698, n2329 );
nand U5014 ( n4398, n4699, n4400 );
nand U5015 ( n4400, n4698, n4401 );
nand U5016 ( n4401, n4402, n4403 );
nor U5017 ( n4403, n4404, n4405 );
nand U5018 ( n4405, n4406, n4644 );
nor U5019 ( n4406, n2231, n2283 );
nand U5020 ( n4404, n4407, n4408 );
nor U5021 ( n4408, n2275, n2215 );
nor U5022 ( n4407, n2232, n2284 );
nor U5023 ( n4402, n4409, n4410 );
nand U5024 ( n4410, n4411, n4642 );
nor U5025 ( n4411, n2280, n2216 );
nand U5026 ( n4409, n4412, n4643 );
nor U5027 ( n4412, n2236, n2293 );
nand U5028 ( n1219, n4413, n4414 );
nand U5029 ( n4414, n4415, n2456 );
nand U5030 ( n4413, n4416, n2330 );
nand U5031 ( n1214, n4417, n4418 );
nand U5032 ( n4418, n4415, n2330 );
nand U5033 ( n4417, n4416, n2338 );
nand U5034 ( n1209, n4419, n4420 );
nand U5035 ( n4420, n4415, n2338 );
nand U5036 ( n4419, n4416, n2288 );
nand U5037 ( n1204, n4421, n4422 );
nand U5038 ( n4422, n4415, n2288 );
nand U5039 ( n4421, n4416, n2339 );
nand U5040 ( n1199, n4423, n4424 );
nand U5041 ( n4424, n4415, n2339 );
nand U5042 ( n4423, n4416, n2340 );
nand U5043 ( n1194, n4425, n4426 );
nand U5044 ( n4426, n4415, n2340 );
nand U5045 ( n4425, n4416, n2289 );
nand U5046 ( n1189, n4427, n4428 );
nand U5047 ( n4428, n4415, n2289 );
nand U5048 ( n4427, n4416, n2249 );
nand U5049 ( n1184, n4429, n4430 );
nand U5050 ( n4430, n4415, n2249 );
nor U5051 ( n4415, n4416, n2843 );
not U5052 ( n2843, n2517 );
nand U5053 ( n2517, n2877, n2522 );
nor U5054 ( n2522, n2208, n2265 );
nor U5055 ( n2877, n2199, n2245 );
nand U5056 ( n4429, n4416, n2331 );
not U5057 ( n4416, n2842 );
nand U5058 ( n2842, n4431, n4681 );
nor U5059 ( n4431, n4682, n2476 );
nand U5060 ( n2476, n4655, n2947 );
and U5061 ( n2947, n4654, n2983 );
and U5062 ( n2983, n4688, n2969 );
and U5063 ( n2969, n4653, n2446 );
nand U5064 ( N41, n3296, n4432 );
nand U5065 ( n4432, g109, n2317 );
nand U5066 ( n3296, n3004, g109 );
nor U5067 ( n3004, n2472, n4657 );
endmodule

