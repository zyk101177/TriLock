
module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule

module s5378_ori ( clk, reset, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat,
n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat,
n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat,
n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat,
n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat,
n3099gat, n3100gat, n3104gat, n3105gat, n3106gat, n3107gat, n3108gat,
n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat,
n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat,
n3123gat, n3124gat, n3125gat, n3126gat, n3127gat, n3128gat, n3129gat,
n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat,
n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat,
n3144gat, n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat,
n3151gat, n3152gat );
input clk, reset, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat,
n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat,
n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat,
n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat,
n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat,
n3100gat;
output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat;
wire n673gat, n398gat, n402gat, n919gat, n846gat, n394gat, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, n703gat,
n722gat, n726gat, n2510gat, n271gat, n160gat, n337gat, n842gat,
n341gat, n2522gat, n1821gat, n1825gat, n1829gat, n283gat, n165gat,
n279gat, n1026gat, n275gat, n2476gat, n1068gat, n957gat, n861gat,
n1294gat, n1241gat, n1298gat, n865gat, n1080gat, n1148gat, n2468gat,
n618gat, n491gat, n622gat, n626gat, n834gat, n707gat, n838gat,
n614gat, n2526gat, n680gat, n816gat, n580gat, n824gat, n820gat,
n883gat, n584gat, n684gat, n699gat, n2399gat, n2343gat, n2203gat,
n2562gat, n2207gat, n2626gat, n2490gat, n2622gat, n2630gat, n2543gat,
n2102gat, n1880gat, n495, n1763gat, new_n2989gat_, n2155gat, n1035gat,
n1121gat, n1072gat, n1282gat, n1226gat, n931gat, n1135gat, n1045gat,
n1197gat, n2518gat, n667gat, n659gat, n553gat, n777gat, n561gat,
n366gat, n322gat, n318gat, n314gat, n2599gat, n2588gat, n2640gat,
n2658gat, n2390gat, n2270gat, n2339gat, n2502gat, n2506gat, n1834gat,
n1767gat, n2084gat, n2143gat, n2061gat, n2139gat, n1899gat, n1850gat,
n2403gat, n2394gat, n2440gat, n2407gat, n2347gat, n1389gat, n2021gat,
n1394gat, n1496gat, n2091gat, n1740gat, n2179gat, n2190gat, n2135gat,
n2262gat, n2182gat, n1312gat, n1775gat, n1871gat, n1508gat, n1678gat,
n2169gat, n2454gat, n2040gat, n2099gat, new_n2194gat_, new_n2057gat_,
n2266gat, new_n2195gat_, new_n2556gat_, new_n2436gat_, new_n2387gat_,
new_n2330gat_, new_n2147gat_, new_n2396gat_, new_n2198gat_,
new_n2197gat_, new_n2196gat_, new_n1882gat_, n1975gat, n2644gat,
n156gat, n152gat, new_n2917gat_, new_n2892gat_, n388gat,
new_n2900gat_, new_n2929gat_, n463gat, n327gat, new_n2925gat_,
new_n2916gat_, n384gat, new_n2899gat_, n256gat, n470gat,
new_n2926gat_, new_n2924gat_, n148gat, new_n2923gat_, n665, n1771gat,
n625, n660, n1336gat, n1748gat, n1675gat, n1807gat, n1340gat,
n1456gat, n3142gat, n1525gat, n1596gat, n1588gat, n650, n560, n610,
n390, n440, n295, n344, n241, n211, n170, n300, n305, n310, n315,
n320, n329, n334, n339, n395, n400, n405, n425, n515, n520, n525,
n530, n535, n540, n545, n550, n555, n565, n570, n575, n580, n585,
n590, n595, n600, n605, n615, n790, n246, n256, n505, n730, n740,
n755, n810, n815, n825, n865, n875, n885, n995, n1000, n1005, n1020,
n1025, n1035, n1040, n1045, n2, n3, n4, n7, n8, n9, n10, n11, n12,
n13, n14, n15, n18, n19, n20, n21, n25, n41, n42, n45, n46, n48, n56,
n57, n58, n59, n68, n69, n70, n71, n72, n73, n92, n94, n95, n96, n97,
n98, n99, n100, n122, n123, n124, n125, n126, n127, n128, n129, n130,
n131, n132, n133, n134, n135, n136, n137, n139, n140, n141, n142,
n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
n165, n166, n167, n168, n169, n171, n172, n173, n174, n175, n176,
n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
n210, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
n233, n234, n235, n236, n237, n238, n239, n240, n242, n243, n244,
n245, n247, n248, n249, n250, n251, n252, n253, n254, n255, n257,
n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
n291, n292, n293, n294, n296, n297, n298, n299, n301, n302, n303,
n304, n306, n307, n308, n309, n311, n312, n313, n314, n316, n317,
n318, n319, n321, n322, n323, n324, n325, n326, n327, n328, n330,
n331, n332, n333, n335, n336, n337, n338, n340, n341, n342, n343,
n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
n389, n391, n392, n393, n394, n396, n397, n398, n399, n401, n402,
n403, n404, n406, n407, n408, n409, n410, n411, n412, n413, n414,
n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n426,
n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
n438, n439, n441, n442, n443, n444, n445, n446, n447, n448, n449,
n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
n494, n496, n497, n498, n499, n500, n501, n502, n503, n504, n506,
n507, n508, n509, n510, n511, n512, n513, n514, n516, n517, n518,
n519, n521, n522, n523, n524, n526, n527, n528, n529, n531, n532,
n533, n534, n536, n537, n538, n539, n541, n542, n543, n544, n546,
n547, n548, n549, n551, n552, n553, n554, n556, n557, n558, n559,
n561, n562, n563, n564, n566, n567, n568, n569, n571, n572, n573,
n574, n576, n577, n578, n579, n581, n582, n583, n584, n586, n587,
n588, n592, n593, n594, n596, n597, n598, n599, n601, n602, n603,
n604, n606, n607, n608, n611, n612, n613, n614, n616, n617, n618,
n619, n620, n621, n622, n623, n624, n626, n627, n628, n629, n630,
n631, n632, n633, n634, n636, n637, n638, n639, n640, n641, n642,
n643, n644, n645, n646, n647, n648, n649, n651, n652, n653, n654,
n655, n656, n657, n658, n659, n661, n662, n663, n664, n666, n667,
n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
n679, n680, n681, n683, n684, n685, n686, n687, n688, n689, n690,
n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
n724, n725, n726, n727, n728, n729, n731, n732, n733, n734, n735,
n736, n737, n738, n739, n741, n742, n743, n744, n745, n746, n747,
n748, n749, n750, n751, n752, n753, n754, n756, n757, n758, n759,
n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
n782, n783, n784, n785, n786, n787, n788, n789, n791, n792, n793,
n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
n805, n806, n807, n808, n809, n811, n812, n813, n814, n816, n817,
n818, n819, n820, n821, n822, n823, n824, n826, n827, n828, n829,
n830, n831, n833, n834, n835, n836, n837, n838, n839, n840, n841,
n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
n864, n866, n867, n868, n869, n870, n871, n872, n873, n874, n876,
n877, n878, n879, n880, n881, n882, n883, n884, n886, n887, n888,
n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
n911, n912, n913, n914, n915, n916, n917, n919, n920, n921, n922,
n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
n967, n968, n969, n3139gat, n971, n973, n974, n975, n976, n977, n978,
n980, n982, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n996, n997, n998, n999, n1001, n1002, n1004, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1021, n1023, n1024, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1036, n1037, n1038, n1039, n1041, n1042,
n1043, n1044, n1046, n1047, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074;
assign n3147gat = 1'b1;
assign n3141gat = n3142gat;
assign n3148gat = 1'b1;
assign n3140gat = n3139gat;
assign n3115gat = 1'b1;
assign n3112gat = 1'b1;
assign n3152gat = 1'b1;

dff n673gat_reg ( clk, reset, n673gat, n170 );
not U_inv0 ( n1034, n673gat );
dff n398gat_reg ( clk, reset, n398gat, n3069gat );
not U_inv1 ( n990, n398gat );
dff n402gat_reg ( clk, reset, n402gat, n3070gat );
dff n919gat_reg ( clk, reset, n919gat, n3072gat );
not U_inv2 ( n1030, n919gat );
dff n846gat_reg ( clk, reset, n846gat, n3071gat );
dff n394gat_reg ( clk, reset, n394gat, n3069gat );
not U_inv3 ( n1011, n394gat );
dff n703gat_reg ( clk, reset, n703gat, n3070gat );
not U_inv4 ( n1013, n703gat );
dff n726gat_reg ( clk, reset, n726gat, n3071gat );
dff n2510gat_reg ( clk, reset, n2510gat, n211 );
dff n271gat_reg ( clk, reset, n271gat, n3065gat );
dff n160gat_reg ( clk, reset, n160gat, n3067gat );
dff n337gat_reg ( clk, reset, n337gat, n3066gat );
dff n842gat_reg ( clk, reset, n842gat, n3073gat );
not U_inv5 ( n1033, n842gat );
dff n341gat_reg ( clk, reset, n341gat, n3068gat );
dff n2522gat_reg ( clk, reset, n2522gat, n241 );
dff n2472gat_reg ( clk, reset, ex_wire0, n246 );
not U_inv6 ( n1007, ex_wire0 );
dff n2319gat_reg ( clk, reset, ex_wire1, n1007 );
not U_inv7 ( n1058, ex_wire1 );
dff n1821gat_reg ( clk, reset, n1821gat, n256 );
dff n1825gat_reg ( clk, reset, n1825gat, n256 );
dff n2029gat_reg ( clk, reset, ex_wire2, n978 );
not U_inv8 ( n1068, ex_wire2 );
dff n1829gat_reg ( clk, reset, n1829gat, n1068 );
dff n283gat_reg ( clk, reset, n283gat, n3065gat );
dff n165gat_reg ( clk, reset, n165gat, n3067gat );
dff n279gat_reg ( clk, reset, n279gat, n3066gat );
not U_inv9 ( n1018, n279gat );
dff n1026gat_reg ( clk, reset, n1026gat, n3073gat );
dff n275gat_reg ( clk, reset, n275gat, n3068gat );
not U_inv10 ( n1015, n275gat );
dff n2476gat_reg ( clk, reset, n2476gat, n295 );
dff n1068gat_reg ( clk, reset, n1068gat, n300 );
dff n957gat_reg ( clk, reset, n957gat, n305 );
dff n861gat_reg ( clk, reset, n861gat, n310 );
not U_inv11 ( n1016, n861gat );
dff n1294gat_reg ( clk, reset, n1294gat, n315 );
dff n1241gat_reg ( clk, reset, n1241gat, n320 );
dff n1298gat_reg ( clk, reset, n1298gat, n170 );
dff n865gat_reg ( clk, reset, n865gat, n329 );
not U_inv12 ( n1017, n865gat );
dff n1080gat_reg ( clk, reset, n1080gat, n334 );
dff n1148gat_reg ( clk, reset, n1148gat, n339 );
dff n2468gat_reg ( clk, reset, n2468gat, n344 );
dff n618gat_reg ( clk, reset, n618gat, n3070gat );
dff n491gat_reg ( clk, reset, n491gat, n3069gat );
dff n622gat_reg ( clk, reset, n622gat, n3071gat );
dff n626gat_reg ( clk, reset, n626gat, n3072gat );
dff n148gat_reg ( clk, reset, n148gat, n1044 );
dff n834gat_reg ( clk, reset, n834gat, new_n2923gat_ );
not U_inv13 ( n1044, n834gat );
dff n2526gat_reg ( clk, reset, n2526gat, n390 );
dff n2588gat_reg ( clk, reset, n2588gat, n615 );
dff n1871gat_reg ( clk, reset, n1871gat, n815 );
not U_inv14 ( n3106gat, n1871gat );
dff n2095gat_reg ( clk, reset, ex_wire3, n982 );
not U_inv15 ( n1046, ex_wire3 );
dff n2176gat_reg ( clk, reset, ex_wire4, n1046 );
not U_inv16 ( n1001, ex_wire4 );
dff n2169gat_reg ( clk, reset, n2169gat, n1001 );
not U_inv17 ( n1057, n2169gat );
dff n2390gat_reg ( clk, reset, n2390gat, n18 );
not U_inv18 ( n3128gat, n2390gat );
dff n2262gat_reg ( clk, reset, n2262gat, n3128gat );
not U_inv19 ( n1056, n2262gat );
dff n2270gat_reg ( clk, reset, n2270gat, new_n2194gat_ );
not U_inv20 ( n3127gat, n2270gat );
dff n2190gat_reg ( clk, reset, n2190gat, n3127gat );
dff n2495gat_reg ( clk, reset, ex_wire5, n977 );
not U_inv21 ( n1039, ex_wire5 );
dff n2266gat_reg ( clk, reset, n2266gat, n1039 );
dff n2339gat_reg ( clk, reset, n2339gat, new_n2057gat_ );
not U_inv22 ( n3126gat, n2339gat );
dff n2135gat_reg ( clk, reset, n2135gat, n3126gat );
dff n2502gat_reg ( clk, reset, n2502gat, n650 );
dff n2626gat_reg ( clk, reset, n2626gat, new_n2195gat_ );
not U_inv23 ( n1036, n2626gat );
dff n1899gat_reg ( clk, reset, n1899gat, n1036 );
not U_inv24 ( n986, n1899gat );
dff n2490gat_reg ( clk, reset, n2490gat, new_n2330gat_ );
not U_inv25 ( n1038, n2490gat );
dff n2139gat_reg ( clk, reset, n2139gat, n1038 );
not U_inv26 ( n999, n2139gat );
dff n2622gat_reg ( clk, reset, n2622gat, new_n2387gat_ );
not U_inv27 ( n1027, n2622gat );
dff n2061gat_reg ( clk, reset, n2061gat, n1027 );
not U_inv28 ( n985, n2061gat );
dff n2543gat_reg ( clk, reset, n2543gat, new_n2436gat_ );
not U_inv29 ( n1037, n2543gat );
dff n2143gat_reg ( clk, reset, n2143gat, n1037 );
not U_inv30 ( n1004, n2143gat );
dff n2630gat_reg ( clk, reset, n2630gat, new_n2556gat_ );
not U_inv31 ( n993, n2630gat );
dff n1850gat_reg ( clk, reset, n1850gat, n993 );
not U_inv32 ( n1050, n1850gat );
dff n1678gat_reg ( clk, reset, n1678gat, n71 );
dff n2454gat_reg ( clk, reset, n2454gat, n865 );
dff n1767gat_reg ( clk, reset, n1767gat, n8 );
dff n1775gat_reg ( clk, reset, n1775gat, n810 );
not U_inv33 ( n1059, n1775gat );
dff n2592gat_reg ( clk, reset, ex_wire6, n1059 );
not U_inv34 ( n996, ex_wire6 );
dff n1834gat_reg ( clk, reset, n1834gat, n665 );
dff n2182gat_reg ( clk, reset, n2182gat, n969 );
dff n614gat_reg ( clk, reset, n614gat, new_n2892gat_ );
not U_inv35 ( n992, n614gat );
dff n156gat_reg ( clk, reset, n156gat, n992 );
not U_inv36 ( n1054, n156gat );
dff n707gat_reg ( clk, reset, n707gat, new_n2917gat_ );
not U_inv37 ( n1043, n707gat );
dff n152gat_reg ( clk, reset, n152gat, n1043 );
dff n838gat_reg ( clk, reset, n838gat, new_n2924gat_ );
not U_inv38 ( n991, n838gat );
dff n256gat_reg ( clk, reset, n256gat, n991 );
not U_inv39 ( n1055, n256gat );
dff n830gat_reg ( clk, reset, ex_wire7, new_n2926gat_ );
not U_inv40 ( n1026, ex_wire7 );
dff n470gat_reg ( clk, reset, n470gat, n1026 );
dff n2179gat_reg ( clk, reset, n2179gat, n974 );
dff n2091gat_reg ( clk, reset, n2091gat, n971 );
dff n2040gat_reg ( clk, reset, n2040gat, n9 );
dff n2021gat_reg ( clk, reset, n2021gat, n973 );
dff n2102gat_reg ( clk, reset, n2102gat, n495 );
dff n1763gat_reg ( clk, reset, n1763gat, n505 );
dff n2155gat_reg ( clk, reset, n2155gat, new_n2989gat_ );
dff n1508gat_reg ( clk, reset, n1508gat, n825 );
dff n2562gat_reg ( clk, reset, n2562gat, new_n2147gat_ );
not U_inv41 ( n1012, n2562gat );
dff n2440gat_reg ( clk, reset, n2440gat, n1012 );
not U_inv42 ( n997, n2440gat );
dff n2343gat_reg ( clk, reset, n2343gat, new_n2198gat_ );
not U_inv43 ( n988, n2343gat );
dff n2394gat_reg ( clk, reset, n2394gat, n988 );
not U_inv44 ( n1042, n2394gat );
dff n2399gat_reg ( clk, reset, n2399gat, new_n2396gat_ );
not U_inv45 ( n1014, n2399gat );
dff n2403gat_reg ( clk, reset, n2403gat, n1014 );
not U_inv46 ( n994, n2403gat );
dff n2203gat_reg ( clk, reset, n2203gat, new_n2196gat_ );
not U_inv47 ( n984, n2203gat );
dff n2347gat_reg ( clk, reset, n2347gat, n984 );
not U_inv48 ( n1053, n2347gat );
dff n2207gat_reg ( clk, reset, n2207gat, new_n2197gat_ );
not U_inv49 ( n989, n2207gat );
dff n2407gat_reg ( clk, reset, n2407gat, n989 );
not U_inv50 ( n1052, n2407gat );
dff n1394gat_reg ( clk, reset, n1394gat, n740 );
not U_inv51 ( n1031, n1394gat );
dff n1496gat_reg ( clk, reset, n1496gat, n1031 );
dff n1332gat_reg ( clk, reset, ex_wire8, n755 );
not U_inv52 ( n1067, ex_wire8 );
dff n1740gat_reg ( clk, reset, n1740gat, n1067 );
dff n1389gat_reg ( clk, reset, n1389gat, n730 );
dff n2640gat_reg ( clk, reset, n2640gat, n975 );
not U_inv53 ( n1041, n2640gat );
dff n2644gat_reg ( clk, reset, n2644gat, n1041 );
dff n2658gat_reg ( clk, reset, n2658gat, n625 );
dff n1433gat_reg ( clk, reset, ex_wire9, n790 );
not U_inv54 ( n1066, ex_wire9 );
dff n1316gat_reg ( clk, reset, ex_wire10, n1066 );
not U_inv55 ( n1010, ex_wire10 );
dff n1363gat_reg ( clk, reset, ex_wire11, n1010 );
not U_inv56 ( n1065, ex_wire11 );
dff n1312gat_reg ( clk, reset, n1312gat, n1065 );
not U_inv57 ( n1008, n1312gat );
dff n2044gat_reg ( clk, reset, ex_wire12, n875 );
not U_inv58 ( n1064, ex_wire12 );
dff n2037gat_reg ( clk, reset, ex_wire13, n1064 );
not U_inv59 ( n1002, ex_wire13 );
dff n2033gat_reg ( clk, reset, ex_wire14, n1002 );
not U_inv60 ( n1047, ex_wire14 );
dff n2110gat_reg ( clk, reset, ex_wire15, n1047 );
not U_inv61 ( n987, ex_wire15 );
dff n2125gat_reg ( clk, reset, ex_wire16, n987 );
not U_inv62 ( n1009, ex_wire16 );
dff n2121gat_reg ( clk, reset, ex_wire17, n1009 );
not U_inv63 ( n1063, ex_wire17 );
dff n2117gat_reg ( clk, reset, ex_wire18, n1063 );
not U_inv64 ( n1071, ex_wire18 );
dff n1880gat_reg ( clk, reset, n1880gat, new_n1882gat_ );
dff n2084gat_reg ( clk, reset, n2084gat, n3149gat );
dff n2025gat_reg ( clk, reset, ex_wire19, n885 );
not U_inv65 ( n1062, ex_wire19 );
dff n2099gat_reg ( clk, reset, n2099gat, n1062 );
dff n314gat_reg ( clk, reset, n314gat, n605 );
dff n318gat_reg ( clk, reset, n318gat, n600 );
dff n322gat_reg ( clk, reset, n322gat, n595 );
dff n366gat_reg ( clk, reset, n366gat, n590 );
dff n561gat_reg ( clk, reset, n561gat, n585 );
dff n777gat_reg ( clk, reset, n777gat, n580 );
dff n553gat_reg ( clk, reset, n553gat, n575 );
dff n659gat_reg ( clk, reset, n659gat, n570 );
dff n667gat_reg ( clk, reset, n667gat, n565 );
dff n2599gat_reg ( clk, reset, n2599gat, n610 );
dff n1197gat_reg ( clk, reset, n1197gat, n555 );
dff n1045gat_reg ( clk, reset, n1045gat, n550 );
dff n1135gat_reg ( clk, reset, n1135gat, n545 );
dff n931gat_reg ( clk, reset, n931gat, n540 );
dff n1226gat_reg ( clk, reset, n1226gat, n535 );
dff n1282gat_reg ( clk, reset, n1282gat, n530 );
dff n1072gat_reg ( clk, reset, n1072gat, n525 );
dff n1121gat_reg ( clk, reset, n1121gat, n520 );
dff n1035gat_reg ( clk, reset, n1035gat, n515 );
dff n2518gat_reg ( clk, reset, n2518gat, n560 );
dff n2634gat_reg ( clk, reset, ex_wire20, n976 );
not U_inv66 ( n1032, ex_wire20 );
dff n1975gat_reg ( clk, reset, n1975gat, n1032 );
dff n2506gat_reg ( clk, reset, n2506gat, n660 );
dff n584gat_reg ( clk, reset, n584gat, n425 );
dff n580gat_reg ( clk, reset, n580gat, n405 );
dff n816gat_reg ( clk, reset, n816gat, n400 );
dff n680gat_reg ( clk, reset, n680gat, n395 );
dff n883gat_reg ( clk, reset, n883gat, new_n2929gat_ );
not U_inv67 ( n1023, n883gat );
dff n388gat_reg ( clk, reset, n388gat, n1023 );
dff n824gat_reg ( clk, reset, n824gat, new_n2900gat_ );
not U_inv68 ( n1060, n824gat );
dff n331gat_reg ( clk, reset, ex_wire21, n1060 );
not U_inv69 ( n1006, ex_wire21 );
dff n684gat_reg ( clk, reset, n684gat, new_n2916gat_ );
not U_inv70 ( n1019, n684gat );
dff n327gat_reg ( clk, reset, n327gat, n1019 );
dff n820gat_reg ( clk, reset, n820gat, new_n2925gat_ );
not U_inv71 ( n1024, n820gat );
dff n463gat_reg ( clk, reset, n463gat, n1024 );
dff n699gat_reg ( clk, reset, n699gat, new_n2899gat_ );
not U_inv72 ( n1021, n699gat );
dff n384gat_reg ( clk, reset, n384gat, n1021 );
dff n2464gat_reg ( clk, reset, ex_wire22, n440 );
not U_inv73 ( n1072, ex_wire22 );
dff n2458gat_reg ( clk, reset, ex_wire23, n996 );
not U_inv74 ( n1061, ex_wire23 );
dff n2514gat_reg ( clk, reset, ex_wire24, n1061 );
not U_inv75 ( n998, ex_wire24 );
dff n1771gat_reg ( clk, reset, n1771gat, n995 );
dff n1336gat_reg ( clk, reset, n1336gat, n1000 );
dff n1748gat_reg ( clk, reset, n1748gat, n1005 );
dff n1675gat_reg ( clk, reset, n1675gat, n72 );
dff n1807gat_reg ( clk, reset, n1807gat, n68 );
dff n1340gat_reg ( clk, reset, n1340gat, n1020 );
not U_inv76 ( n1028, n1340gat );
dff n1456gat_reg ( clk, reset, n1456gat, n1025 );
dff n1525gat_reg ( clk, reset, n1525gat, n980 );
dff n1462gat_reg ( clk, reset, ex_wire25, n1035 );
not U_inv77 ( n1029, ex_wire25 );
dff n1596gat_reg ( clk, reset, n1596gat, n1040 );
dff n1588gat_reg ( clk, reset, n1588gat, n1045 );
dff n722gat_reg ( clk, reset, n722gat, n3072gat );
or U1053 ( n1051, n683, n684 );
not U1054 ( n130, n353 );
not U1055 ( n9, n151 );
not U1056 ( n69, n696 );
nor U1057 ( n353, n360, n135 );
not U1058 ( n133, n557 );
or U1059 ( n167, n370, n135 );
not U1060 ( n132, n163 );
nor U1061 ( n151, n156, n971 );
not U1062 ( n13, n974 );
not U1063 ( n41, n536 );
not U1064 ( n42, n528 );
nand U1065 ( n257, n95, n308 );
not U1066 ( n11, n156 );
nor U1067 ( n427, n46, n42 );
not U1068 ( n98, n308 );
not U1069 ( n129, n336 );
not U1070 ( n20, new_n2147gat_ );
nor U1071 ( new_n2396gat_, n564, n20 );
nor U1072 ( new_n2198gat_, n563, n20 );
not U1073 ( n19, new_n2195gat_ );
nor U1074 ( new_n2330gat_, n567, n19 );
nor U1075 ( new_n2387gat_, n19, n574 );
nor U1076 ( n995, n672, n7 );
not U1077 ( n12, n783 );
nor U1078 ( n940, n719, n59 );
nor U1079 ( n696, n70, n581 );
not U1080 ( n70, n656 );
nor U1081 ( n885, n686, n58 );
not U1082 ( n73, n704 );
not U1083 ( n2, n686 );
nor U1084 ( n1005, n69, n686 );
nand U1085 ( n973, n633, n7 );
nor U1086 ( n633, n9, n8 );
not U1087 ( n71, n657 );
not U1088 ( n72, n658 );
nand U1089 ( n360, n370, n361 );
nand U1090 ( n370, n133, n131 );
nor U1091 ( n557, n134, n139 );
nand U1092 ( n3122gat, n390, n380 );
nand U1093 ( n380, n128, n239 );
nand U1094 ( n3123gat, n610, n373 );
nand U1095 ( n373, n128, n195 );
nand U1096 ( n3121gat, n440, n387 );
nand U1097 ( n387, n128, n220 );
nand U1098 ( n3120gat, n295, n396 );
nand U1099 ( n396, n128, n168 );
nand U1100 ( n3119gat, n344, n404 );
nand U1101 ( n404, n128, n212 );
nand U1102 ( n3118gat, n241, n538 );
nand U1103 ( n538, n128, n228 );
nand U1104 ( n3117gat, n211, n547 );
nand U1105 ( n547, n128, n178 );
nand U1106 ( n3135gat, n229, n230 );
nand U1107 ( n230, n231, n160 );
nand U1108 ( n229, n239, n169 );
nand U1109 ( n231, n235, n236 );
nand U1110 ( n3136gat, n188, n189 );
nand U1111 ( n189, n190, n160 );
nand U1112 ( n188, n195, n169 );
nand U1113 ( n190, n191, n192 );
nand U1114 ( n3134gat, n213, n214 );
nand U1115 ( n214, n215, n160 );
nand U1116 ( n213, n220, n169 );
nand U1117 ( n215, n216, n217 );
nand U1118 ( n3133gat, n157, n158 );
nand U1119 ( n158, n159, n160 );
nand U1120 ( n157, n168, n169 );
nand U1121 ( n159, n161, n162 );
nand U1122 ( n3132gat, n204, n205 );
nand U1123 ( n205, n206, n160 );
nand U1124 ( n204, n212, n169 );
nand U1125 ( n206, n207, n208 );
nand U1126 ( n3131gat, n221, n222 );
nand U1127 ( n222, n223, n160 );
nand U1128 ( n221, n228, n169 );
nand U1129 ( n223, n224, n225 );
nand U1130 ( n3130gat, n171, n172 );
nand U1131 ( n172, n173, n160 );
nand U1132 ( n171, n178, n169 );
nand U1133 ( n173, n174, n175 );
nand U1134 ( n3124gat, n560, n362 );
nand U1135 ( n362, n128, n198 );
nand U1136 ( n3137gat, n196, n197 );
nand U1137 ( n196, n199, n160 );
nand U1138 ( n197, n198, n169 );
nand U1139 ( n199, n200, n201 );
or U1140 ( n166, n357, n360 );
nor U1141 ( n349, n166, n354 );
nand U1142 ( n187, n347, n348 );
nor U1143 ( n347, n355, n356 );
nor U1144 ( n348, n349, n350 );
nor U1145 ( n356, n357, n358 );
nand U1146 ( n3125gat, n650, n346 );
nand U1147 ( n346, n128, n187 );
nand U1148 ( n3129gat, n179, n180 );
nand U1149 ( n180, n181, n160 );
nand U1150 ( n179, n169, n187 );
nand U1151 ( n181, n182, n183 );
nor U1152 ( n163, n361, n135 );
not U1153 ( n135, n357 );
nand U1154 ( n358, n359, n360 );
nand U1155 ( n359, n361, n1034 );
not U1156 ( n127, n248 );
not U1157 ( n96, n341 );
nand U1158 ( n3104gat, n321, n322 );
nor U1159 ( n321, n323, n324 );
nor U1160 ( n324, n325, n326 );
nor U1161 ( n323, n327, n328 );
nand U1162 ( n3105gat, n330, n331 );
nor U1163 ( n330, n332, n333 );
nor U1164 ( n333, n100, n335 );
nor U1165 ( n332, n338, n340 );
not U1166 ( n100, n337 );
nand U1167 ( n3151gat, n566, n567 );
nor U1168 ( n566, n99, n568 );
nor U1169 ( n568, n341, n327 );
not U1170 ( n99, n326 );
nand U1171 ( n327, n569, n137 );
not U1172 ( n128, n233 );
nand U1173 ( n169, n240, n242 );
nand U1174 ( n240, n234, n137 );
nand U1175 ( n242, n243, n244 );
nor U1176 ( n244, n127, n245 );
nor U1177 ( n243, n247, n133 );
nand U1178 ( n340, n341, n137 );
nand U1179 ( n162, n163, n992 );
nand U1180 ( n208, n163, n1043 );
nand U1181 ( n225, n163, n991 );
nand U1182 ( n175, n163, n1044 );
nand U1183 ( n183, n163, n1026 );
nor U1184 ( n336, n131, n325 );
nand U1185 ( n335, n336, n134 );
nor U1186 ( n602, n606, n607 );
nor U1187 ( n607, n56, n608 );
nor U1188 ( n606, n611, n612 );
not U1189 ( n56, n420 );
nand U1190 ( n630, n9, n1028 );
nand U1191 ( n974, n259, n313 );
nand U1192 ( n971, n811, n534 );
and U1193 ( n811, n13, n598 );
not U1194 ( n15, n818 );
nor U1195 ( n536, n444, n1014 );
nor U1196 ( n516, n517, n45 );
not U1197 ( n45, n484 );
nor U1198 ( n517, n518, n519 );
nor U1199 ( n518, n59, n524 );
and U1200 ( n342, n412, n413 );
nor U1201 ( n413, n414, n415 );
and U1202 ( n412, n421, n422 );
nor U1203 ( n415, n3106gat, n416 );
nand U1204 ( n3143gat, n342, n660 );
nand U1205 ( n3144gat, n342, n625 );
nand U1206 ( n474, n3149gat, n1012 );
nand U1207 ( n456, n457, n458 );
nand U1208 ( n457, n483, n484 );
nand U1209 ( n458, n459, n460 );
nor U1210 ( n483, n485, n486 );
nor U1211 ( n486, n1014, n487 );
nor U1212 ( n487, n488, n489 );
nand U1213 ( n489, n490, n491 );
nand U1214 ( n488, n492, n493 );
nor U1215 ( n501, n988, n503 );
nor U1216 ( n503, n474, n1015 );
not U1217 ( n59, n3149gat );
nor U1218 ( n468, n59, n1012 );
nor U1219 ( n528, n445, n1014 );
nor U1220 ( n469, n3149gat, n1012 );
nor U1221 ( n455, n504, n506 );
nand U1222 ( n504, n988, n1014 );
nand U1223 ( n506, n460, n507 );
nand U1224 ( n507, n508, n509 );
nor U1225 ( n156, n1013, n634 );
nand U1226 ( n422, n156, n423 );
nand U1227 ( n423, n424, n426 );
nand U1228 ( n426, n427, n428 );
nand U1229 ( n424, n429, n430 );
not U1230 ( n95, n316 );
nor U1231 ( n296, n257, n298 );
xnor U1232 ( n298, n1006, n299 );
not U1233 ( n94, n266 );
nor U1234 ( n3145gat, n9, n631 );
nor U1235 ( n631, n632, n998 );
nand U1236 ( n537, n11, n534 );
and U1237 ( n514, n460, n529 );
nand U1238 ( n529, n531, n532 );
nand U1239 ( n532, n528, n533 );
nand U1240 ( n531, n536, n537 );
not U1241 ( n46, n597 );
nand U1242 ( n792, n801, n802 );
nand U1243 ( n802, n803, n337 );
nand U1244 ( n801, n806, n96 );
nor U1245 ( n803, n134, n129 );
nor U1246 ( n317, n129, n805 );
nand U1247 ( n308, n671, n134 );
nor U1248 ( n3138gat, n592, n593 );
nand U1249 ( n593, n594, n536 );
nand U1250 ( n592, n596, n597 );
nor U1251 ( n596, n1027, n13 );
not U1252 ( n57, new_n2989gat_ );
nor U1253 ( n460, n989, n984 );
nor U1254 ( n733, n1014, n734 );
nor U1255 ( n734, n484, n429 );
nand U1256 ( n581, n583, n985 );
not U1257 ( n58, n653 );
not U1258 ( n3116gat, n186 );
nand U1259 ( n741, n445, n742 );
nand U1260 ( n742, n988, n1012 );
not U1261 ( n92, n632 );
nor U1262 ( new_n2147gat_, n637, n587 );
nor U1263 ( new_n2195gat_, n587, n643 );
nor U1264 ( new_n2196gat_, n20, n343 );
nor U1265 ( new_n2197gat_, n20, n345 );
nor U1266 ( new_n2556gat_, n322, n19 );
nor U1267 ( new_n2436gat_, n19, n331 );
nand U1268 ( n416, n996, n1034 );
xnor U1269 ( n574, n985, n583 );
nor U1270 ( n563, n997, n1042 );
xnor U1271 ( n564, n994, n582 );
nor U1272 ( n567, n999, n986 );
nand U1273 ( n565, n780, n781 );
nor U1274 ( n780, n12, n782 );
nor U1275 ( n782, n139, n126 );
nand U1276 ( n585, n768, n769 );
nor U1277 ( n768, n12, n770 );
nor U1278 ( n770, n139, n124 );
nand U1279 ( n590, n765, n766 );
nor U1280 ( n765, n12, n767 );
nor U1281 ( n767, n139, n125 );
nand U1282 ( n600, n759, n760 );
nor U1283 ( n759, n12, n761 );
nor U1284 ( n761, n139, n123 );
nand U1285 ( n605, n756, n757 );
nor U1286 ( n756, n12, n758 );
nor U1287 ( n758, n139, n122 );
not U1288 ( n18, n587 );
nor U1289 ( new_n2194gat_, n573, n587 );
nor U1290 ( new_n2057gat_, n587, n572 );
nor U1291 ( n3107gat, n3106gat, n92 );
nor U1292 ( n667, n1046, n1001 );
nand U1293 ( n672, n833, n3100gat );
nor U1294 ( n833, n1007, n614 );
nor U1295 ( n505, n672, n21 );
not U1296 ( n21, n495 );
nor U1297 ( n810, n672, n687 );
nand U1298 ( n783, n807, n808 );
nor U1299 ( n807, n823, n824 );
nor U1300 ( n808, n629, n809 );
nor U1301 ( n823, n826, n827 );
nand U1302 ( n809, n971, n989 );
nand U1303 ( n686, n928, n929 );
nor U1304 ( n928, n941, n942 );
nor U1305 ( n929, n930, n931 );
nor U1306 ( n942, n943, n944 );
nor U1307 ( n656, n1004, n1050 );
nor U1308 ( n931, n4, n932 );
nand U1309 ( n932, n933, n934 );
nand U1310 ( n934, n935, n936 );
nand U1311 ( n935, n582, n1030 );
and U1312 ( n719, n959, n960 );
nand U1313 ( n959, n73, new_n2989gat_ );
nand U1314 ( n960, n696, n57 );
and U1315 ( n933, n955, n956 );
nor U1316 ( n956, n1053, n957 );
and U1317 ( n955, n892, n940 );
nand U1318 ( n957, n994, n1052 );
nand U1319 ( n704, n962, n963 );
nor U1320 ( n962, n999, n985 );
nor U1321 ( n963, n1004, n964 );
nand U1322 ( n964, n1050, n986 );
nor U1323 ( n1025, n920, n921 );
nand U1324 ( n920, new_n2989gat_, n710 );
nand U1325 ( n921, n2, n73 );
nor U1326 ( n930, n938, n939 );
nand U1327 ( n938, n563, n1053 );
nand U1328 ( n939, n940, n708 );
nand U1329 ( n292, n299, n1006 );
nand U1330 ( n643, n690, n691 );
nor U1331 ( n691, n692, n693 );
nor U1332 ( n690, n702, n703 );
nor U1333 ( n692, n697, n658 );
nor U1334 ( n702, n577, n698 );
nor U1335 ( n693, n694, n695 );
nand U1336 ( n694, n698, n699 );
nand U1337 ( n695, n696, n697 );
not U1338 ( n4, n949 );
nor U1339 ( n951, n1042, n4 );
nand U1340 ( n943, n946, n947 );
nor U1341 ( n947, n892, n948 );
nor U1342 ( n946, n951, n952 );
nor U1343 ( n948, n949, n950 );
nor U1344 ( n950, n990, n1042 );
nor U1345 ( n703, n704, n699 );
nand U1346 ( n283, n14, n1054 );
not U1347 ( n14, n313 );
nand U1348 ( n282, n278, n1055 );
nand U1349 ( n658, n700, n985 );
nand U1350 ( n637, n705, n706 );
nand U1351 ( n706, n707, n708 );
or U1352 ( n705, n710, n57 );
nor U1353 ( n707, new_n2989gat_, n709 );
nor U1354 ( n730, n719, n715 );
not U1355 ( n8, n687 );
nand U1356 ( n969, n10, n598 );
not U1357 ( n10, n537 );
nor U1358 ( n1035, n577, n917 );
nor U1359 ( n1040, n69, n917 );
not U1360 ( n68, n577 );
nand U1361 ( n657, n924, n656 );
and U1362 ( n924, n985, n567 );
nor U1363 ( n1020, n715, n657 );
not U1364 ( n7, n665 );
not U1365 ( n139, n3095gat );
nor U1366 ( n384, n703gat, n130 );
nand U1367 ( n239, n381, n382 );
nor U1368 ( n381, n385, n386 );
nor U1369 ( n382, n383, n384 );
nor U1370 ( n386, n684gat, n132 );
nor U1371 ( n377, n726gat, n130 );
nor U1372 ( n392, n394gat, n130 );
nor U1373 ( n401, n341gat, n130 );
nor U1374 ( n409, n160gat, n130 );
nor U1375 ( n543, n337gat, n130 );
nor U1376 ( n552, n271gat, n130 );
nand U1377 ( n195, n374, n375 );
nor U1378 ( n374, n378, n379 );
nor U1379 ( n375, n376, n377 );
nor U1380 ( n379, n824gat, n132 );
nand U1381 ( n220, n388, n389 );
nor U1382 ( n388, n393, n394 );
nor U1383 ( n389, n391, n392 );
nor U1384 ( n394, n699gat, n132 );
nand U1385 ( n168, n397, n398 );
nor U1386 ( n397, n402, n403 );
nor U1387 ( n398, n399, n401 );
nor U1388 ( n403, n584gat, n132 );
nand U1389 ( n212, n406, n407 );
nor U1390 ( n406, n410, n411 );
nor U1391 ( n407, n408, n409 );
nor U1392 ( n411, n816gat, n132 );
nand U1393 ( n228, n539, n541 );
nor U1394 ( n539, n544, n546 );
nor U1395 ( n541, n542, n543 );
nor U1396 ( n546, n580gat, n132 );
nand U1397 ( n178, n548, n549 );
nor U1398 ( n548, n553, n554 );
nor U1399 ( n549, n551, n552 );
nor U1400 ( n554, n680gat, n132 );
nor U1401 ( n365, n722gat, n130 );
nand U1402 ( n198, n363, n364 );
nor U1403 ( n363, n371, n372 );
nor U1404 ( n364, n365, n366 );
nor U1405 ( n372, n883gat, n132 );
nor U1406 ( n371, n366gat, n166 );
nor U1407 ( n378, n561gat, n166 );
nor U1408 ( n385, n318gat, n166 );
nor U1409 ( n393, n314gat, n166 );
nor U1410 ( n402, n322gat, n166 );
nor U1411 ( n410, n553gat, n166 );
nor U1412 ( n544, n777gat, n166 );
nor U1413 ( n553, n659gat, n166 );
nor U1414 ( n191, n193, n194 );
nor U1415 ( n193, n846gat, n167 );
nor U1416 ( n194, n1282gat, n166 );
nor U1417 ( n235, n237, n238 );
nor U1418 ( n237, n402gat, n167 );
nor U1419 ( n238, n1135gat, n166 );
nor U1420 ( n216, n218, n219 );
nor U1421 ( n218, n398gat, n167 );
nor U1422 ( n219, n1045gat, n166 );
nor U1423 ( n161, n164, n165 );
nor U1424 ( n164, n275gat, n167 );
nor U1425 ( n165, n931gat, n166 );
nor U1426 ( n207, n209, n210 );
nor U1427 ( n209, n165gat, n167 );
nor U1428 ( n210, n1121gat, n166 );
nor U1429 ( n224, n226, n227 );
nor U1430 ( n226, n279gat, n167 );
nor U1431 ( n227, n1072gat, n166 );
nor U1432 ( n174, n176, n177 );
nor U1433 ( n176, n283gat, n167 );
nor U1434 ( n177, n1035gat, n166 );
nor U1435 ( n200, n202, n203 );
nor U1436 ( n202, n919gat, n167 );
nor U1437 ( n203, n1226gat, n166 );
nor U1438 ( n182, n184, n185 );
nor U1439 ( n184, n1026gat, n167 );
nor U1440 ( n185, n166, n186 );
not U1441 ( n134, n3086gat );
nand U1442 ( n350, n351, n352 );
nand U1443 ( n351, n353, n1033 );
or U1444 ( n352, n167, n1241gat );
nand U1445 ( n366, n367, n368 );
nand U1446 ( n368, n369, n135 );
or U1447 ( n367, n167, n1298gat );
nor U1448 ( n369, n673gat, n370 );
nor U1449 ( n376, n1294gat, n167 );
nor U1450 ( n383, n1080gat, n167 );
nor U1451 ( n391, n1148gat, n167 );
nor U1452 ( n399, n865gat, n167 );
nor U1453 ( n408, n957gat, n167 );
nor U1454 ( n542, n861gat, n167 );
nor U1455 ( n551, n1068gat, n167 );
nand U1456 ( n357, n558, n247 );
nand U1457 ( n558, n3093gat, n3087gat );
nand U1458 ( n247, n3088gat, n3095gat );
nor U1459 ( n355, n820gat, n132 );
not U1460 ( n131, n3085gat );
nand U1461 ( n361, n556, n250 );
nand U1462 ( n556, n3095gat, n3087gat );
nand U1463 ( n250, n3093gat, n3086gat );
nand U1464 ( n341, n850, n3087gat );
nor U1465 ( n248, n3083gat, n3084gat );
nand U1466 ( n328, n96, n3094gat );
and U1467 ( n850, n851, n852 );
nor U1468 ( n852, n3085gat, n3106gat );
nor U1469 ( n851, n139, n127 );
nand U1470 ( n338, n3094gat, n97 );
not U1471 ( n97, n569 );
nand U1472 ( n569, n850, n3086gat );
or U1473 ( n192, n132, n622gat );
or U1474 ( n236, n132, n618gat );
or U1475 ( n217, n132, n491gat );
or U1476 ( n201, n132, n626gat );
nand U1477 ( n805, n854, n3093gat );
nor U1478 ( n854, n3106gat, n127 );
nor U1479 ( n337, n804, n805 );
nand U1480 ( n804, n136, n3088gat );
nand U1481 ( n326, n571, n337 );
nor U1482 ( n571, n3085gat, n134 );
nand U1483 ( n160, n232, n233 );
nand U1484 ( n232, n3088gat, n234 );
nand U1485 ( n233, n559, n248 );
nor U1486 ( n559, n3085gat, n561 );
nor U1487 ( n561, n562, n557 );
nor U1488 ( n562, n136, n139 );
not U1489 ( n136, n3087gat );
xnor U1490 ( n211, n905, n906 );
xnor U1491 ( n905, n3087gat, n913 );
xnor U1492 ( n906, n3086gat, n907 );
xnor U1493 ( n913, n3089gat, n137 );
nand U1494 ( n907, n908, n909 );
nand U1495 ( n909, n910, n131 );
nand U1496 ( n908, n3085gat, n911 );
xor U1497 ( n910, n3084gat, n3083gat );
nand U1498 ( n911, n127, n912 );
nand U1499 ( n912, n3083gat, n3084gat );
nand U1500 ( n245, n3087gat, n131 );
and U1501 ( n234, n248, n249 );
nand U1502 ( n249, n250, n251 );
nand U1503 ( n251, n3093gat, n3085gat );
not U1504 ( n137, n3088gat );
nor U1505 ( n325, n3091gat, n3092gat );
nand U1506 ( n612, n613, n25 );
not U1507 ( n25, n614 );
nand U1508 ( n613, n1825gat, n616 );
nand U1509 ( n616, n3097gat, n58 );
nand U1510 ( n3139gat, n599, n601 );
nor U1511 ( n599, n618, n619 );
and U1512 ( n601, n602, n603 );
nor U1513 ( n619, n1525gat, n143 );
nand U1514 ( n611, n617, n1871gat );
nor U1515 ( n617, n3098gat, n1775gat );
nand U1516 ( n259, n819, n722gat );
nor U1517 ( n819, n703gat, n818 );
nand U1518 ( n818, n820, n726gat );
nor U1519 ( n820, n2454gat, n1011 );
nor U1520 ( n618, n57, n621 );
nor U1521 ( n621, n622, n623 );
nor U1522 ( n623, n1678gat, n1029 );
nor U1523 ( n622, n1508gat, n624 );
nor U1524 ( n624, n626, n627 );
nor U1525 ( n627, n59, n628 );
nor U1526 ( n626, n629, n630 );
nand U1527 ( n628, n1394gat, n1029 );
nand U1528 ( n313, n817, n15 );
nor U1529 ( n817, n722gat, n703gat );
nor U1530 ( n149, n3149gat, n150 );
nor U1531 ( n150, n1340gat, n151 );
nor U1532 ( n145, n57, n146 );
nor U1533 ( n146, n147, n148 );
nor U1534 ( n148, n1807gat, n1028 );
nor U1535 ( n147, n1456gat, n149 );
nand U1536 ( n3142gat, n141, n142 );
or U1537 ( n142, n1675gat, n143 );
nor U1538 ( n141, n144, n145 );
and U1539 ( n144, n152, n153 );
nand U1540 ( n598, n816, n15 );
nor U1541 ( n816, n722gat, n1013 );
nand U1542 ( n444, n2343gat, n1012 );
nor U1543 ( n519, n3149gat, n521 );
nor U1544 ( n521, n522, n523 );
nor U1545 ( n523, n824gat, n42 );
nor U1546 ( n522, n883gat, n41 );
nand U1547 ( n421, n1389gat, n452 );
nand U1548 ( n452, n453, n454 );
nor U1549 ( n454, n455, n456 );
nor U1550 ( n453, n514, n516 );
nor U1551 ( n463, n464, n465 );
nand U1552 ( n465, n466, n467 );
nand U1553 ( n464, n470, n471 );
nand U1554 ( n466, n680gat, n469 );
nor U1555 ( n470, n2343gat, n473 );
nor U1556 ( n473, n474, n1016 );
nor U1557 ( n459, n461, n462 );
nor U1558 ( n461, n2399gat, n475 );
nor U1559 ( n462, n1014, n463 );
nor U1560 ( n475, n476, n477 );
nor U1561 ( n492, n2343gat, n494 );
nor U1562 ( n494, n474, n1018 );
nor U1563 ( n524, n526, n527 );
nor U1564 ( n527, n1294gat, n42 );
nor U1565 ( n526, n1298gat, n41 );
nand U1566 ( n3149gat, n958, n1880gat );
and U1567 ( n958, n1834gat, n1767gat );
nand U1568 ( n476, n480, n481 );
nand U1569 ( n481, n584gat, n472 );
nor U1570 ( n480, n988, n482 );
nor U1571 ( n482, n474, n1017 );
nand U1572 ( n534, n812, n813 );
nor U1573 ( n813, n394gat, n2454gat );
nor U1574 ( n812, n1013, n814 );
nor U1575 ( n485, n2399gat, n496 );
nor U1576 ( n496, n497, n498 );
nand U1577 ( n498, n499, n500 );
nand U1578 ( n497, n501, n502 );
nand U1579 ( n814, n722gat, n726gat );
nand U1580 ( n467, n1068gat, n468 );
nand U1581 ( n477, n478, n479 );
nand U1582 ( n478, n816gat, n469 );
nand U1583 ( n479, n957gat, n468 );
nand U1584 ( n491, n283gat, n468 );
nand U1585 ( n500, n165gat, n468 );
nand U1586 ( n490, n469, n834gat );
nand U1587 ( n499, n469, n707gat );
nor U1588 ( n508, n512, n513 );
and U1589 ( n513, n1021, n469 );
nor U1590 ( n512, n1148gat, n48 );
not U1591 ( n48, n468 );
nand U1592 ( n445, n2562gat, n2343gat );
nor U1593 ( n472, n3149gat, n2562gat );
nand U1594 ( n471, n580gat, n472 );
nand U1595 ( n634, n722, n394gat );
nor U1596 ( n722, n726gat, n2454gat );
nand U1597 ( n493, n472, n838gat );
nand U1598 ( n502, n472, n614gat );
nand U1599 ( n439, n441, n988 );
nand U1600 ( n441, n442, n443 );
or U1601 ( n443, n2562gat, n366gat );
or U1602 ( n442, n1012, n561gat );
nor U1603 ( n434, n2399gat, n435 );
nor U1604 ( n435, n436, n437 );
nor U1605 ( n436, n314gat, n445 );
nand U1606 ( n437, n438, n439 );
nand U1607 ( n430, n431, n432 );
nor U1608 ( n431, n450, n451 );
nor U1609 ( n432, n433, n434 );
nor U1610 ( n451, n659gat, n42 );
nor U1611 ( n316, n849, n338 );
nand U1612 ( n849, n341, n3088gat );
nor U1613 ( n303, n257, n306 );
xor U1614 ( n306, n384gat, n307 );
nor U1615 ( n307, n327gat, n292 );
nor U1616 ( n269, n257, n271 );
xor U1617 ( n271, n463gat, n272 );
nor U1618 ( n272, n273, n259 );
nor U1619 ( n273, n274, n388gat );
nor U1620 ( n289, n257, n291 );
xnor U1621 ( n291, n327gat, n292 );
nor U1622 ( n254, n257, n258 );
xnor U1623 ( n258, n388gat, n259 );
nand U1624 ( new_n2899gat_, n301, n302 );
nand U1625 ( n302, n3069gat, n98 );
nor U1626 ( n301, n303, n304 );
nor U1627 ( n304, n95, n122 );
nand U1628 ( new_n2925gat_, n267, n268 );
nand U1629 ( n268, n3073gat, n98 );
nor U1630 ( n267, n269, n270 );
nor U1631 ( n270, n95, n126 );
nand U1632 ( new_n2916gat_, n287, n288 );
nand U1633 ( n288, n3070gat, n98 );
nor U1634 ( n287, n289, n290 );
nor U1635 ( n290, n95, n123 );
nand U1636 ( new_n2900gat_, n293, n294 );
nand U1637 ( n294, n3071gat, n98 );
nor U1638 ( n293, n296, n297 );
nor U1639 ( n297, n95, n124 );
nand U1640 ( new_n2929gat_, n252, n253 );
nand U1641 ( n253, n3072gat, n98 );
nor U1642 ( n252, n254, n255 );
nor U1643 ( n255, n95, n125 );
or U1644 ( n438, n444, n318gat );
nor U1645 ( n509, n510, n511 );
and U1646 ( n511, n1019, n472 );
nor U1647 ( n510, n1080gat, n474 );
nand U1648 ( n153, n154, n155 );
nor U1649 ( n154, n3149gat, n156 );
nand U1650 ( n155, n1336gat, n971 );
nor U1651 ( n450, n777gat, n41 );
nand U1652 ( n143, n620, n971 );
nor U1653 ( n620, n1394gat, new_n2989gat_ );
nand U1654 ( n266, n314, n95 );
nand U1655 ( n314, n317, n318 );
nor U1656 ( n318, n137, n319 );
nand U1657 ( n319, n3087gat, n134 );
nand U1658 ( new_n2926gat_, n260, n261 );
nand U1659 ( n260, n3073gat, n266 );
nand U1660 ( n261, n262, n94 );
xor U1661 ( n262, n263, n470gat );
nand U1662 ( new_n2917gat_, n284, n285 );
nand U1663 ( n284, n3067gat, n266 );
nand U1664 ( n285, n286, n94 );
xor U1665 ( n286, n283, n152gat );
nand U1666 ( new_n2923gat_, n279, n280 );
nand U1667 ( n279, n3065gat, n266 );
nand U1668 ( n280, n281, n94 );
xor U1669 ( n281, n282, n148gat );
nand U1670 ( new_n2924gat_, n275, n276 );
nand U1671 ( n275, n3066gat, n266 );
nand U1672 ( n276, n277, n94 );
xnor U1673 ( n277, n278, n256gat );
nand U1674 ( new_n2892gat_, n309, n311 );
nand U1675 ( n309, n3068gat, n266 );
nand U1676 ( n311, n312, n94 );
xnor U1677 ( n312, n14, n156gat );
and U1678 ( n629, n821, n822 );
nor U1679 ( n821, n1012, n46 );
nor U1680 ( n822, n2343gat, n1014 );
nand U1681 ( n533, n2084gat, n534 );
nor U1682 ( n449, n553gat, n1012 );
nor U1683 ( n433, n446, n447 );
nand U1684 ( n447, n2399gat, n988 );
nor U1685 ( n446, n448, n449 );
nor U1686 ( n448, n322gat, n2562gat );
nor U1687 ( n597, n2203gat, n2207gat );
nor U1688 ( n806, n3088gat, n338 );
nand U1689 ( n515, n783, n800 );
nand U1690 ( n800, n3065gat, n792 );
nand U1691 ( n520, n783, n799 );
nand U1692 ( n799, n3067gat, n792 );
nand U1693 ( n525, n783, n798 );
nand U1694 ( n798, n3066gat, n792 );
nand U1695 ( n530, n783, n797 );
nand U1696 ( n797, n3071gat, n792 );
nand U1697 ( n535, n783, n796 );
nand U1698 ( n796, n3072gat, n792 );
nand U1699 ( n540, n783, n795 );
nand U1700 ( n795, n3068gat, n792 );
nand U1701 ( n545, n783, n794 );
nand U1702 ( n794, n3070gat, n792 );
nand U1703 ( n550, n783, n793 );
nand U1704 ( n793, n3069gat, n792 );
nand U1705 ( n555, n783, n791 );
nand U1706 ( n791, n3073gat, n792 );
xnor U1707 ( n354, n749, n750 );
xor U1708 ( n749, n753, n754 );
xor U1709 ( n750, n751, n752 );
xnor U1710 ( n753, n314gat, n318gat );
xor U1711 ( n751, n777gat, n659gat );
xor U1712 ( n428, n722gat, n354 );
xor U1713 ( n752, n561gat, n553gat );
and U1714 ( n671, n317, n853 );
nor U1715 ( n853, n3088gat, n136 );
xor U1716 ( n754, n366gat, n322gat );
or U1717 ( n608, n1069, n1596gat );
and U1718 ( n1069, n11, n1031 );
nand U1719 ( new_n2989gat_, n2102gat, n961 );
or U1720 ( n961, n1880gat, n1763gat );
nor U1721 ( n414, n417, n418 );
nand U1722 ( n418, n3149gat, n1031 );
nor U1723 ( n417, n419, n420 );
nor U1724 ( n419, n1508gat, n57 );
nand U1725 ( n395, n847, n848 );
nand U1726 ( n848, n3074gat, n316 );
nand U1727 ( n847, n3065gat, n98 );
nand U1728 ( n400, n845, n846 );
nand U1729 ( n846, n3076gat, n316 );
nand U1730 ( n845, n3067gat, n98 );
nand U1731 ( n405, n843, n844 );
nand U1732 ( n844, n3075gat, n316 );
nand U1733 ( n843, n3066gat, n98 );
nand U1734 ( n425, n841, n842 );
nand U1735 ( n842, n3077gat, n316 );
nand U1736 ( n841, n3068gat, n98 );
nor U1737 ( n484, n989, n2203gat );
xnor U1738 ( n186, n784, n785 );
xor U1739 ( n784, n788, n789 );
xor U1740 ( n785, n786, n787 );
xnor U1741 ( n788, n1035gat, n1045gat );
xor U1742 ( n786, n931gat, n1282gat );
xor U1743 ( n787, n1226gat, n1135gat );
xor U1744 ( n789, n1121gat, n1072gat );
nand U1745 ( n982, n668, n669 );
nand U1746 ( n668, n671, n3086gat );
nand U1747 ( n669, n670, n96 );
nor U1748 ( n670, n137, n338 );
xnor U1749 ( n625, n729, n731 );
nand U1750 ( n729, n736, n737 );
nor U1751 ( n731, n732, n733 );
nand U1752 ( n736, n741, n2640gat );
nor U1753 ( n732, n2399gat, n735 );
nor U1754 ( n735, n597, n460 );
nor U1755 ( n420, new_n2989gat_, n1678gat );
xnor U1756 ( n295, n879, n880 );
xor U1757 ( n880, n881, n882 );
xor U1758 ( n879, n883, n884 );
xnor U1759 ( n882, n283gat, n1018 );
nand U1760 ( n888, n402gat, n891 );
xnor U1761 ( n891, n990, n275gat );
nor U1762 ( n884, n886, n887 );
and U1763 ( n886, n275gat, n892 );
nand U1764 ( n887, n888, n889 );
nand U1765 ( n889, n890, n1015 );
nor U1766 ( n429, n984, n2207gat );
nor U1767 ( n892, n990, n402gat );
nand U1768 ( n577, n1850gat, n579 );
nor U1769 ( n579, n581, n2143gat );
nor U1770 ( n583, n1899gat, n2139gat );
and U1771 ( n322, n577, n578 );
or U1772 ( n578, n579, n1850gat );
xnor U1773 ( n241, n894, n895 );
xor U1774 ( n894, n903, n904 );
xor U1775 ( n895, n896, n897 );
xnor U1776 ( n903, n337gat, n341gat );
nand U1777 ( n900, n814, n901 );
or U1778 ( n901, n722gat, n726gat );
nand U1779 ( n896, n898, n899 );
nand U1780 ( n898, n842gat, n902 );
nand U1781 ( n899, n900, n1033 );
xor U1782 ( n902, n726gat, n722gat );
nor U1783 ( n890, n402gat, n398gat );
nand U1784 ( n737, n738, n1041 );
nand U1785 ( n738, n444, n739 );
nand U1786 ( n739, n2562gat, n988 );
xor U1787 ( n610, n354, n667gat );
xnor U1788 ( n904, n1013, n394gat );
nand U1789 ( n653, n2021gat, n1880gat );
xnor U1790 ( n560, n3116gat, n1197gat );
nand U1791 ( n632, n1771gat, n1775gat );
nor U1792 ( n662, n987, n663 );
nor U1793 ( n663, n998, n664 );
nand U1794 ( n664, n92, n1871gat );
nor U1795 ( n3146gat, n659, n661 );
nand U1796 ( n659, n666, n667 );
nand U1797 ( n661, n662, n2169gat );
nor U1798 ( n666, n1002, n1047 );
xnor U1799 ( n440, n834, n835 );
xnor U1800 ( n835, n1021, n684gat );
xor U1801 ( n834, n836, n837 );
xnor U1802 ( n836, n580gat, n840 );
xor U1803 ( n837, n838, n839 );
xnor U1804 ( n839, n1024, n816gat );
xnor U1805 ( n838, n1023, n824gat );
xor U1806 ( n866, n867, n868 );
xor U1807 ( n868, n1298gat, n1294gat );
xnor U1808 ( n867, n957gat, n1016 );
xnor U1809 ( n344, n862, n863 );
xnor U1810 ( n863, n1017, n1148gat );
xor U1811 ( n862, n864, n866 );
xnor U1812 ( n864, n1068gat, n869 );
nor U1813 ( n614, n1829gat, n978 );
nand U1814 ( n978, n1825gat, n1821gat );
xor U1815 ( n869, n1241gat, n1080gat );
xnor U1816 ( n390, n855, n856 );
xnor U1817 ( n856, n618gat, n992 );
xor U1818 ( n855, n857, n858 );
xnor U1819 ( n857, n491gat, n861 );
xor U1820 ( n858, n859, n860 );
xnor U1821 ( n860, n1026, n707gat );
xnor U1822 ( n859, n991, n834gat );
xor U1823 ( n840, n680gat, n584gat );
nand U1824 ( n652, n1051, n140 );
nand U1825 ( n684, n2658gat, n2588gat );
not U1826 ( n140, n3100gat );
nand U1827 ( n587, n648, n649 );
nor U1828 ( n649, n1046, n1002 );
and U1829 ( n648, n651, n652 );
nand U1830 ( n651, n2099gat, n653 );
nor U1831 ( n152, n1748gat, new_n2989gat_ );
xor U1832 ( n861, n626gat, n622gat );
nand U1833 ( n603, n604, n1596gat );
nor U1834 ( n604, n1588gat, new_n2989gat_ );
xnor U1835 ( n726, n1027, n2543gat );
xor U1836 ( n660, n723, n724 );
xnor U1837 ( n724, n1036, n725 );
xnor U1838 ( n723, n2490gat, n726 );
xnor U1839 ( n725, n1032, n2630gat );
xnor U1840 ( n345, n584, n2407gat );
nand U1841 ( n584, n641, n582 );
nor U1842 ( n641, n2403gat, n2347gat );
nand U1843 ( n3108gat, n1035gat, n345 );
xnor U1844 ( n331, n581, n2143gat );
xnor U1845 ( n881, n1030, n846gat );
xnor U1846 ( n897, n160gat, n271gat );
nor U1847 ( n582, n2394gat, n2440gat );
and U1848 ( n594, n967, n968 );
nor U1849 ( n968, n2626gat, n1038 );
nor U1850 ( n967, n993, n1037 );
xnor U1851 ( n883, n1026gat, n165gat );
nand U1852 ( n975, n636, new_n2147gat_ );
xor U1853 ( n636, n638, n2644gat );
nand U1854 ( n638, n639, n640 );
and U1855 ( n639, n997, n584 );
xnor U1856 ( n343, n586, n2347gat );
nand U1857 ( n586, n582, n994 );
nand U1858 ( n3109gat, n1072gat, n343 );
nand U1859 ( n976, n642, new_n2195gat_ );
xor U1860 ( n642, n644, n1975gat );
nand U1861 ( n644, n645, n646 );
nor U1862 ( n645, n1899gat, n579 );
nand U1863 ( n3150gat, n574, n576 );
or U1864 ( n576, n2454gat, n337gat );
nand U1865 ( n3111gat, n563, n931gat );
nand U1866 ( n3110gat, n1121gat, n564 );
nand U1867 ( n977, n647, n18 );
xor U1868 ( n647, n654, n2266gat );
nand U1869 ( n654, n2190gat, n1056 );
xor U1870 ( n572, n2135gat, n588 );
nor U1871 ( n588, n2262gat, n2190gat );
nand U1872 ( n3113gat, n1135gat, n572 );
xor U1873 ( n650, n727, n728 );
xnor U1874 ( n727, n2270gat, n2339gat );
xnor U1875 ( n728, n1039, n2390gat );
not U1876 ( n126, n3082gat );
not U1877 ( n124, n3080gat );
not U1878 ( n125, n3081gat );
not U1879 ( n123, n3079gat );
not U1880 ( n122, n3078gat );
nor U1881 ( n815, n3, n680 );
not U1882 ( n3, n885 );
nand U1883 ( n680, n681, n652 );
nand U1884 ( n681, n1775gat, n1008 );
nor U1885 ( n865, n674, n675 );
nand U1886 ( n675, n1312gat, n2 );
nand U1887 ( n674, n652, n1057 );
and U1888 ( n573, n2262gat, n2190gat );
nand U1889 ( n3114gat, n573, n1282gat );
nor U1890 ( new_n1882gat_, n1070, n1071 );
nand U1891 ( n1070, n1009, n3100gat );
nand U1892 ( n570, n777, n778 );
nor U1893 ( n777, n12, n779 );
and U1894 ( n779, n3095gat, n3074gat );
nand U1895 ( n575, n774, n775 );
nor U1896 ( n774, n12, n776 );
and U1897 ( n776, n3095gat, n3076gat );
nand U1898 ( n580, n771, n772 );
nor U1899 ( n771, n12, n773 );
and U1900 ( n773, n3095gat, n3075gat );
nand U1901 ( n595, n762, n763 );
nor U1902 ( n762, n12, n764 );
and U1903 ( n764, n3095gat, n3077gat );
or U1904 ( n745, n1072, n3090gat );
nand U1905 ( n615, n743, n744 );
nor U1906 ( n743, n747, n748 );
nor U1907 ( n744, n745, n746 );
nand U1908 ( n747, n2522gat, n2518gat );
nand U1909 ( n766, n3072gat, n3093gat );
nand U1910 ( n170, n914, n766 );
nand U1911 ( n914, n3081gat, n3095gat );
nand U1912 ( n757, n3069gat, n3093gat );
nand U1913 ( n760, n3070gat, n3093gat );
nand U1914 ( n763, n3068gat, n3093gat );
nand U1915 ( n781, n3073gat, n3093gat );
nand U1916 ( n769, n3071gat, n3093gat );
nand U1917 ( n772, n3066gat, n3093gat );
nand U1918 ( n775, n3067gat, n3093gat );
nand U1919 ( n778, n3065gat, n3093gat );
nand U1920 ( n339, n870, n757 );
nand U1921 ( n870, n3078gat, n3095gat );
nand U1922 ( n334, n871, n760 );
nand U1923 ( n871, n3079gat, n3095gat );
nand U1924 ( n329, n872, n763 );
nand U1925 ( n872, n3077gat, n3095gat );
nand U1926 ( n320, n873, n781 );
nand U1927 ( n873, n3082gat, n3095gat );
nand U1928 ( n315, n874, n769 );
nand U1929 ( n874, n3080gat, n3095gat );
nand U1930 ( n310, n876, n772 );
nand U1931 ( n876, n3075gat, n3095gat );
nand U1932 ( n305, n877, n775 );
nand U1933 ( n877, n3076gat, n3095gat );
nand U1934 ( n300, n878, n778 );
nand U1935 ( n878, n3074gat, n3095gat );
nor U1936 ( n256, n3099gat, n1058 );
nor U1937 ( n941, n953, n954 );
or U1938 ( n953, n952, n949 );
nand U1939 ( n954, n933, n2394gat );
nand U1940 ( n944, n945, n940 );
and U1941 ( n945, n2347gat, n708 );
nor U1942 ( n824, n2203gat, n41 );
nor U1943 ( n299, n259, n388gat );
nand U1944 ( n697, n701, n57 );
nor U1945 ( n701, n2091gat, n1496gat );
and U1946 ( n826, n2155gat, n1073 );
and U1947 ( n1073, n594, n1027 );
or U1948 ( n699, n57, n1740gat );
nor U1949 ( n949, n990, n846gat );
nor U1950 ( n278, n283, n152gat );
and U1951 ( n700, n916, n656 );
nor U1952 ( n916, n1899gat, n999 );
nor U1953 ( n827, n828, n829 );
nand U1954 ( n828, n831, n1038 );
nand U1955 ( n829, n830, n2630gat );
nor U1956 ( n831, n2622gat, n2543gat );
nor U1957 ( n830, n2155gat, n1036 );
xnor U1958 ( n952, n919gat, n997 );
nand U1959 ( n698, n1740gat, new_n2989gat_ );
nor U1960 ( n708, n994, n2407gat );
nor U1961 ( n790, n688, n689 );
and U1962 ( n688, n2182gat, n711 );
nand U1963 ( n689, n637, n643 );
nand U1964 ( n711, n712, n588 );
nand U1965 ( n936, n937, n2440gat );
nor U1966 ( n937, n2394gat, n1030 );
nand U1967 ( n640, n2403gat, n1042 );
nand U1968 ( n710, n922, n923 );
nor U1969 ( n923, n2407gat, n2347gat );
nor U1970 ( n922, n997, n640 );
nand U1971 ( n709, n919, n2394gat );
nor U1972 ( n919, n2440gat, n2347gat );
nand U1973 ( n683, n685, n2510gat );
and U1974 ( n685, n2506gat, n2502gat );
nand U1975 ( n263, n14, n264 );
nand U1976 ( n264, n1054, n265 );
or U1977 ( n265, n1055, n152gat );
nand U1978 ( n687, n720, n722gat );
nor U1979 ( n720, n703gat, n634 );
and U1980 ( n274, n1006, n327gat );
nand U1981 ( n715, n925, n926 );
nor U1982 ( n925, n1052, n997 );
nor U1983 ( n926, n2347gat, n927 );
nand U1984 ( n927, n1042, n994 );
nor U1985 ( n755, n713, n714 );
nand U1986 ( n713, n2061gat, n583 );
or U1987 ( n714, n715, n70 );
nor U1988 ( n740, n716, n717 );
nand U1989 ( n717, n708, n700 );
nand U1990 ( n716, n718, n2061gat );
and U1991 ( n718, n2347gat, n563 );
nor U1992 ( n1000, n965, n966 );
nand U1993 ( n966, n594, n429 );
nand U1994 ( n965, n528, n2622gat );
or U1995 ( n917, n1074, n709 );
or U1996 ( n1074, n2403gat, n1052 );
nor U1997 ( n665, n721, n634 );
or U1998 ( n721, n722gat, n703gat );
nor U1999 ( n1045, n1008, n915 );
nand U2000 ( n915, n700, n2061gat );
nand U2001 ( n646, n2061gat, n999 );
nor U2002 ( n980, n646, n655 );
nand U2003 ( n655, n656, n1899gat );
nor U2004 ( n825, n676, n677 );
nand U2005 ( n677, n678, n2061gat );
nand U2006 ( n676, n679, new_n2989gat_ );
nor U2007 ( n678, n1050, n999 );
nor U2008 ( n679, n2143gat, n1899gat );
nor U2009 ( n495, n2454gat, n271gat );
nor U2010 ( n712, n2179gat, n2135gat );
nor U2011 ( n246, n814, n893 );
nand U2012 ( n893, n703gat, n394gat );
and U2013 ( n875, n673, n1010 );
nor U2014 ( n673, n2040gat, n1775gat );
nand U2015 ( n746, n2476gat, n2468gat );
nand U2016 ( n748, n2599gat, n2526gat );
endmodule

