module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end
endmodule

module iir_ori ( clk, reset, inData_0, inData_1, inData_2, inData_3, inData_4, inData_5, inData_6, inData_7, inData_8, inData_9, inData_10, inData_11, inData_12, inData_13, inData_14, inData_15, inData_16, inData_17, inData_18, inData_19, inData_20, inData_21, inData_22, inData_23, inData_24, inData_25, inData_26, inData_27, inData_28, inData_29, inData_30, inData_31, outData_0, outData_1, outData_2, outData_3, outData_4, outData_5, outData_6, outData_7, outData_8, outData_9, outData_10, outData_11, outData_12, outData_13, outData_14, outData_15, outData_16, outData_17, outData_18, outData_19, outData_20, outData_21, outData_22, outData_23, outData_24, outData_25, outData_26, outData_27, outData_28, outData_29, outData_30, outData_31 );
input clk, reset, inData_0, inData_1, inData_2, inData_3, inData_4, inData_5, inData_6, inData_7, inData_8, inData_9, inData_10, inData_11, inData_12, inData_13, inData_14, inData_15, inData_16, inData_17, inData_18, inData_19, inData_20, inData_21, inData_22, inData_23, inData_24, inData_25, inData_26, inData_27, inData_28, inData_29, inData_30, inData_31;
output outData_0, outData_1, outData_2, outData_3, outData_4, outData_5, outData_6, outData_7, outData_8, outData_9, outData_10, outData_11, outData_12, outData_13, outData_14, outData_15, outData_16, outData_17, outData_18, outData_19, outData_20, outData_21, outData_22, outData_23, outData_24, outData_25, outData_26, outData_27, outData_28, outData_29, outData_30, outData_31;
wire my_IIR_filter_firBlock_left_N288, ex_wire0, ex_wire1, ex_wire2, ex_wire3, my_IIR_filter_firBlock_left_N287,
my_IIR_filter_firBlock_left_N286, my_IIR_filter_firBlock_left_N285,
my_IIR_filter_firBlock_left_N284, my_IIR_filter_firBlock_left_N283,
my_IIR_filter_firBlock_left_N282, my_IIR_filter_firBlock_left_N281,
my_IIR_filter_firBlock_left_N280, my_IIR_filter_firBlock_left_N279,
my_IIR_filter_firBlock_left_N278, my_IIR_filter_firBlock_left_N277,
my_IIR_filter_firBlock_left_N276, my_IIR_filter_firBlock_left_N275,
my_IIR_filter_firBlock_left_N274, my_IIR_filter_firBlock_left_N273,
my_IIR_filter_firBlock_left_N272, my_IIR_filter_firBlock_left_N271,
my_IIR_filter_firBlock_left_N270, my_IIR_filter_firBlock_left_N269,
my_IIR_filter_firBlock_left_N268, my_IIR_filter_firBlock_left_N267,
my_IIR_filter_firBlock_left_N266, my_IIR_filter_firBlock_left_N265,
my_IIR_filter_firBlock_left_N264, my_IIR_filter_firBlock_left_N263,
my_IIR_filter_firBlock_left_N262, my_IIR_filter_firBlock_left_N261,
my_IIR_filter_firBlock_left_N260, my_IIR_filter_firBlock_left_N259,
my_IIR_filter_firBlock_left_N258, my_IIR_filter_firBlock_left_N257,
my_IIR_filter_firBlock_left_N256, my_IIR_filter_firBlock_left_N255,
my_IIR_filter_firBlock_left_N254, my_IIR_filter_firBlock_left_N253,
my_IIR_filter_firBlock_left_N252, my_IIR_filter_firBlock_left_N251,
my_IIR_filter_firBlock_left_N250, my_IIR_filter_firBlock_left_N249,
my_IIR_filter_firBlock_left_N248, my_IIR_filter_firBlock_left_N247,
my_IIR_filter_firBlock_left_N246, my_IIR_filter_firBlock_left_N245,
my_IIR_filter_firBlock_left_N244, my_IIR_filter_firBlock_left_N243,
my_IIR_filter_firBlock_left_N242, my_IIR_filter_firBlock_left_N241,
my_IIR_filter_firBlock_left_N240, my_IIR_filter_firBlock_left_N239,
my_IIR_filter_firBlock_left_N238, my_IIR_filter_firBlock_left_N237,
my_IIR_filter_firBlock_left_N236, my_IIR_filter_firBlock_left_N235,
my_IIR_filter_firBlock_left_N234, my_IIR_filter_firBlock_left_N233,
my_IIR_filter_firBlock_left_N232, my_IIR_filter_firBlock_left_N231,
my_IIR_filter_firBlock_left_N230, my_IIR_filter_firBlock_left_N229,
my_IIR_filter_firBlock_left_N228, my_IIR_filter_firBlock_left_N227,
my_IIR_filter_firBlock_left_N226, my_IIR_filter_firBlock_left_N225,
my_IIR_filter_firBlock_left_N224, my_IIR_filter_firBlock_left_N223,
my_IIR_filter_firBlock_left_N222, my_IIR_filter_firBlock_left_N221,
my_IIR_filter_firBlock_left_N220, my_IIR_filter_firBlock_left_N219,
my_IIR_filter_firBlock_left_N218, my_IIR_filter_firBlock_left_N217,
my_IIR_filter_firBlock_left_N216, my_IIR_filter_firBlock_left_N215,
my_IIR_filter_firBlock_left_N214, my_IIR_filter_firBlock_left_N213,
my_IIR_filter_firBlock_left_N212, my_IIR_filter_firBlock_left_N211,
my_IIR_filter_firBlock_left_N210, my_IIR_filter_firBlock_left_N209,
my_IIR_filter_firBlock_left_N208, my_IIR_filter_firBlock_left_N207,
my_IIR_filter_firBlock_left_N206, my_IIR_filter_firBlock_left_N205,
my_IIR_filter_firBlock_left_N204, my_IIR_filter_firBlock_left_N203,
my_IIR_filter_firBlock_left_N202, my_IIR_filter_firBlock_left_N201,
my_IIR_filter_firBlock_left_N200, my_IIR_filter_firBlock_left_N199,
my_IIR_filter_firBlock_left_N198, my_IIR_filter_firBlock_left_N197,
my_IIR_filter_firBlock_left_N196, my_IIR_filter_firBlock_left_N195,
my_IIR_filter_firBlock_left_N194, my_IIR_filter_firBlock_left_N193,
my_IIR_filter_firBlock_left_N192, my_IIR_filter_firBlock_left_N191,
my_IIR_filter_firBlock_left_N190, my_IIR_filter_firBlock_left_N189,
my_IIR_filter_firBlock_left_N188, my_IIR_filter_firBlock_left_N187,
my_IIR_filter_firBlock_left_N186, my_IIR_filter_firBlock_left_N185,
my_IIR_filter_firBlock_left_N184, my_IIR_filter_firBlock_left_N183,
my_IIR_filter_firBlock_left_N182, my_IIR_filter_firBlock_left_N181,
my_IIR_filter_firBlock_left_N180, my_IIR_filter_firBlock_left_N179,
my_IIR_filter_firBlock_left_N178, my_IIR_filter_firBlock_left_N177,
my_IIR_filter_firBlock_left_N176, my_IIR_filter_firBlock_left_N175,
my_IIR_filter_firBlock_left_N174, my_IIR_filter_firBlock_left_N173,
my_IIR_filter_firBlock_left_N172, my_IIR_filter_firBlock_left_N171,
my_IIR_filter_firBlock_left_N170, my_IIR_filter_firBlock_left_N169,
my_IIR_filter_firBlock_left_N168, my_IIR_filter_firBlock_left_N167,
my_IIR_filter_firBlock_left_N166, my_IIR_filter_firBlock_left_N165,
my_IIR_filter_firBlock_left_N164, my_IIR_filter_firBlock_left_N163,
my_IIR_filter_firBlock_left_N162, my_IIR_filter_firBlock_left_N161,
my_IIR_filter_firBlock_left_N160, my_IIR_filter_firBlock_left_N159,
my_IIR_filter_firBlock_left_N158, my_IIR_filter_firBlock_left_N157,
my_IIR_filter_firBlock_left_N156, my_IIR_filter_firBlock_left_N155,
my_IIR_filter_firBlock_left_N154, my_IIR_filter_firBlock_left_N153,
my_IIR_filter_firBlock_left_N152, my_IIR_filter_firBlock_left_N151,
my_IIR_filter_firBlock_left_N150, my_IIR_filter_firBlock_left_N149,
my_IIR_filter_firBlock_left_N148, my_IIR_filter_firBlock_left_N147,
my_IIR_filter_firBlock_left_N146, my_IIR_filter_firBlock_left_N145,
my_IIR_filter_firBlock_left_N144, my_IIR_filter_firBlock_left_N143,
my_IIR_filter_firBlock_left_N142, my_IIR_filter_firBlock_left_N141,
my_IIR_filter_firBlock_left_N140, my_IIR_filter_firBlock_left_N139,
my_IIR_filter_firBlock_left_N138, my_IIR_filter_firBlock_left_N137,
my_IIR_filter_firBlock_left_N136, my_IIR_filter_firBlock_left_N135,
my_IIR_filter_firBlock_left_N134, my_IIR_filter_firBlock_left_N133,
my_IIR_filter_firBlock_left_N132, my_IIR_filter_firBlock_left_N131,
my_IIR_filter_firBlock_left_N130, my_IIR_filter_firBlock_left_N129,
my_IIR_filter_firBlock_left_N128, my_IIR_filter_firBlock_left_N127,
my_IIR_filter_firBlock_left_N126, my_IIR_filter_firBlock_left_N125,
my_IIR_filter_firBlock_left_N124, my_IIR_filter_firBlock_left_N123,
my_IIR_filter_firBlock_left_N122, my_IIR_filter_firBlock_left_N121,
my_IIR_filter_firBlock_left_N120, my_IIR_filter_firBlock_left_N119,
my_IIR_filter_firBlock_left_N118, my_IIR_filter_firBlock_left_N117,
my_IIR_filter_firBlock_left_N116, my_IIR_filter_firBlock_left_N115,
my_IIR_filter_firBlock_left_N114, my_IIR_filter_firBlock_left_N113,
my_IIR_filter_firBlock_left_N112, my_IIR_filter_firBlock_left_N111,
my_IIR_filter_firBlock_left_N110, my_IIR_filter_firBlock_left_N109,
my_IIR_filter_firBlock_left_N108, my_IIR_filter_firBlock_left_N107,
my_IIR_filter_firBlock_left_N106, my_IIR_filter_firBlock_left_N105,
my_IIR_filter_firBlock_left_N104, my_IIR_filter_firBlock_left_N103,
my_IIR_filter_firBlock_left_N102, my_IIR_filter_firBlock_left_N101,
my_IIR_filter_firBlock_left_N100, my_IIR_filter_firBlock_left_N99,
my_IIR_filter_firBlock_left_N98, my_IIR_filter_firBlock_left_N97,
my_IIR_filter_firBlock_left_N96, my_IIR_filter_firBlock_left_N95,
my_IIR_filter_firBlock_left_N94, my_IIR_filter_firBlock_left_N93,
my_IIR_filter_firBlock_left_N92, my_IIR_filter_firBlock_left_N91,
my_IIR_filter_firBlock_left_N90, my_IIR_filter_firBlock_left_N89,
my_IIR_filter_firBlock_left_N88, my_IIR_filter_firBlock_left_N87,
my_IIR_filter_firBlock_left_N86, my_IIR_filter_firBlock_left_N85,
my_IIR_filter_firBlock_left_N84, my_IIR_filter_firBlock_left_N83,
my_IIR_filter_firBlock_left_N82, my_IIR_filter_firBlock_left_N81,
my_IIR_filter_firBlock_left_N80, my_IIR_filter_firBlock_left_N79,
my_IIR_filter_firBlock_left_N78, my_IIR_filter_firBlock_left_N77,
my_IIR_filter_firBlock_left_N76, my_IIR_filter_firBlock_left_N75,
my_IIR_filter_firBlock_left_N74, my_IIR_filter_firBlock_left_N73,
my_IIR_filter_firBlock_left_N72, my_IIR_filter_firBlock_left_N71,
my_IIR_filter_firBlock_left_N70, my_IIR_filter_firBlock_left_N69,
my_IIR_filter_firBlock_left_N68, my_IIR_filter_firBlock_left_N67,
my_IIR_filter_firBlock_left_N66, my_IIR_filter_firBlock_left_N65,
my_IIR_filter_firBlock_left_N64, my_IIR_filter_firBlock_left_N63,
my_IIR_filter_firBlock_left_N62, my_IIR_filter_firBlock_left_N61,
my_IIR_filter_firBlock_left_N60, my_IIR_filter_firBlock_left_N59,
my_IIR_filter_firBlock_left_N58, my_IIR_filter_firBlock_left_N57,
my_IIR_filter_firBlock_left_N56, my_IIR_filter_firBlock_left_N55,
my_IIR_filter_firBlock_left_N54, my_IIR_filter_firBlock_left_N53,
my_IIR_filter_firBlock_left_N52, my_IIR_filter_firBlock_left_N51,
my_IIR_filter_firBlock_left_N50, my_IIR_filter_firBlock_left_N49,
my_IIR_filter_firBlock_left_N48, my_IIR_filter_firBlock_left_N47,
my_IIR_filter_firBlock_left_N46, my_IIR_filter_firBlock_left_N45,
my_IIR_filter_firBlock_left_N44, my_IIR_filter_firBlock_left_N43,
my_IIR_filter_firBlock_left_N42, my_IIR_filter_firBlock_left_N41,
my_IIR_filter_firBlock_left_N40, my_IIR_filter_firBlock_left_N39,
my_IIR_filter_firBlock_left_N38, my_IIR_filter_firBlock_left_N37,
my_IIR_filter_firBlock_left_N36, my_IIR_filter_firBlock_left_N35,
my_IIR_filter_firBlock_left_N34, my_IIR_filter_firBlock_left_N33,
my_IIR_filter_firBlock_left_N32, my_IIR_filter_firBlock_left_N31,
my_IIR_filter_firBlock_left_N30, my_IIR_filter_firBlock_left_N29,
my_IIR_filter_firBlock_left_N28, my_IIR_filter_firBlock_left_N27,
my_IIR_filter_firBlock_left_N26, my_IIR_filter_firBlock_left_N25,
my_IIR_filter_firBlock_left_N24, my_IIR_filter_firBlock_left_N23,
my_IIR_filter_firBlock_left_N22, my_IIR_filter_firBlock_left_N21,
my_IIR_filter_firBlock_left_N20, my_IIR_filter_firBlock_left_N19,
my_IIR_filter_firBlock_left_N18, my_IIR_filter_firBlock_left_N17,
my_IIR_filter_firBlock_left_N16, my_IIR_filter_firBlock_left_N15,
my_IIR_filter_firBlock_left_N14, my_IIR_filter_firBlock_left_N13,
my_IIR_filter_firBlock_left_N12, my_IIR_filter_firBlock_left_N11,
my_IIR_filter_firBlock_left_N10, my_IIR_filter_firBlock_left_N9,
my_IIR_filter_firBlock_left_N8, my_IIR_filter_firBlock_left_N7,
my_IIR_filter_firBlock_left_N6, my_IIR_filter_firBlock_left_N5,
my_IIR_filter_firBlock_left_N4, my_IIR_filter_firBlock_left_N3,
my_IIR_filter_firBlock_left_N2, my_IIR_filter_firBlock_left_N1,
my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_,
my_IIR_filter_firBlock_right_N192, my_IIR_filter_firBlock_right_N191,
my_IIR_filter_firBlock_right_N190, my_IIR_filter_firBlock_right_N189,
my_IIR_filter_firBlock_right_N188, my_IIR_filter_firBlock_right_N187,
my_IIR_filter_firBlock_right_N186, my_IIR_filter_firBlock_right_N185,
my_IIR_filter_firBlock_right_N184, my_IIR_filter_firBlock_right_N183,
my_IIR_filter_firBlock_right_N182, my_IIR_filter_firBlock_right_N181,
my_IIR_filter_firBlock_right_N180, my_IIR_filter_firBlock_right_N179,
my_IIR_filter_firBlock_right_N178, my_IIR_filter_firBlock_right_N177,
my_IIR_filter_firBlock_right_N176, my_IIR_filter_firBlock_right_N175,
my_IIR_filter_firBlock_right_N174, my_IIR_filter_firBlock_right_N173,
my_IIR_filter_firBlock_right_N172, my_IIR_filter_firBlock_right_N171,
my_IIR_filter_firBlock_right_N170, my_IIR_filter_firBlock_right_N169,
my_IIR_filter_firBlock_right_N168, my_IIR_filter_firBlock_right_N167,
my_IIR_filter_firBlock_right_N166, my_IIR_filter_firBlock_right_N165,
my_IIR_filter_firBlock_right_N164, my_IIR_filter_firBlock_right_N163,
my_IIR_filter_firBlock_right_N162, my_IIR_filter_firBlock_right_N161,
my_IIR_filter_firBlock_right_N160, my_IIR_filter_firBlock_right_N159,
my_IIR_filter_firBlock_right_N158, my_IIR_filter_firBlock_right_N157,
my_IIR_filter_firBlock_right_N156, my_IIR_filter_firBlock_right_N155,
my_IIR_filter_firBlock_right_N154, my_IIR_filter_firBlock_right_N153,
my_IIR_filter_firBlock_right_N152, my_IIR_filter_firBlock_right_N151,
my_IIR_filter_firBlock_right_N150, my_IIR_filter_firBlock_right_N149,
my_IIR_filter_firBlock_right_N148, my_IIR_filter_firBlock_right_N147,
my_IIR_filter_firBlock_right_N146, my_IIR_filter_firBlock_right_N145,
my_IIR_filter_firBlock_right_N144, my_IIR_filter_firBlock_right_N143,
my_IIR_filter_firBlock_right_N142, my_IIR_filter_firBlock_right_N141,
my_IIR_filter_firBlock_right_N140, my_IIR_filter_firBlock_right_N139,
my_IIR_filter_firBlock_right_N138, my_IIR_filter_firBlock_right_N137,
my_IIR_filter_firBlock_right_N136, my_IIR_filter_firBlock_right_N135,
my_IIR_filter_firBlock_right_N134, my_IIR_filter_firBlock_right_N133,
my_IIR_filter_firBlock_right_N132, my_IIR_filter_firBlock_right_N131,
my_IIR_filter_firBlock_right_N130, my_IIR_filter_firBlock_right_N129,
my_IIR_filter_firBlock_right_N128, my_IIR_filter_firBlock_right_N127,
my_IIR_filter_firBlock_right_N126, my_IIR_filter_firBlock_right_N125,
my_IIR_filter_firBlock_right_N124, my_IIR_filter_firBlock_right_N123,
my_IIR_filter_firBlock_right_N122, my_IIR_filter_firBlock_right_N121,
my_IIR_filter_firBlock_right_N120, my_IIR_filter_firBlock_right_N119,
my_IIR_filter_firBlock_right_N118, my_IIR_filter_firBlock_right_N117,
my_IIR_filter_firBlock_right_N116, my_IIR_filter_firBlock_right_N115,
my_IIR_filter_firBlock_right_N114, my_IIR_filter_firBlock_right_N113,
my_IIR_filter_firBlock_right_N112, my_IIR_filter_firBlock_right_N111,
my_IIR_filter_firBlock_right_N110, my_IIR_filter_firBlock_right_N109,
my_IIR_filter_firBlock_right_N108, my_IIR_filter_firBlock_right_N107,
my_IIR_filter_firBlock_right_N106, my_IIR_filter_firBlock_right_N105,
my_IIR_filter_firBlock_right_N104, my_IIR_filter_firBlock_right_N103,
my_IIR_filter_firBlock_right_N102, my_IIR_filter_firBlock_right_N101,
my_IIR_filter_firBlock_right_N100, my_IIR_filter_firBlock_right_N99,
my_IIR_filter_firBlock_right_N98, my_IIR_filter_firBlock_right_N97,
my_IIR_filter_firBlock_right_N96, my_IIR_filter_firBlock_right_N95,
my_IIR_filter_firBlock_right_N94, my_IIR_filter_firBlock_right_N93,
my_IIR_filter_firBlock_right_N92, my_IIR_filter_firBlock_right_N91,
my_IIR_filter_firBlock_right_N90, my_IIR_filter_firBlock_right_N89,
my_IIR_filter_firBlock_right_N88, my_IIR_filter_firBlock_right_N87,
my_IIR_filter_firBlock_right_N86, my_IIR_filter_firBlock_right_N85,
my_IIR_filter_firBlock_right_N84, my_IIR_filter_firBlock_right_N83,
my_IIR_filter_firBlock_right_N82, my_IIR_filter_firBlock_right_N81,
my_IIR_filter_firBlock_right_N80, my_IIR_filter_firBlock_right_N79,
my_IIR_filter_firBlock_right_N78, my_IIR_filter_firBlock_right_N77,
my_IIR_filter_firBlock_right_N76, my_IIR_filter_firBlock_right_N75,
my_IIR_filter_firBlock_right_N74, my_IIR_filter_firBlock_right_N73,
my_IIR_filter_firBlock_right_N72, my_IIR_filter_firBlock_right_N71,
my_IIR_filter_firBlock_right_N70, my_IIR_filter_firBlock_right_N69,
my_IIR_filter_firBlock_right_N68, my_IIR_filter_firBlock_right_N67,
my_IIR_filter_firBlock_right_N66, my_IIR_filter_firBlock_right_N65,
my_IIR_filter_firBlock_right_N64, my_IIR_filter_firBlock_right_N63,
my_IIR_filter_firBlock_right_N62, my_IIR_filter_firBlock_right_N61,
my_IIR_filter_firBlock_right_N60, my_IIR_filter_firBlock_right_N59,
my_IIR_filter_firBlock_right_N58, my_IIR_filter_firBlock_right_N57,
my_IIR_filter_firBlock_right_N56, my_IIR_filter_firBlock_right_N55,
my_IIR_filter_firBlock_right_N54, my_IIR_filter_firBlock_right_N53,
my_IIR_filter_firBlock_right_N52, my_IIR_filter_firBlock_right_N51,
my_IIR_filter_firBlock_right_N50, my_IIR_filter_firBlock_right_N49,
my_IIR_filter_firBlock_right_N48, my_IIR_filter_firBlock_right_N47,
my_IIR_filter_firBlock_right_N46, my_IIR_filter_firBlock_right_N45,
my_IIR_filter_firBlock_right_N44, my_IIR_filter_firBlock_right_N43,
my_IIR_filter_firBlock_right_N42, my_IIR_filter_firBlock_right_N41,
my_IIR_filter_firBlock_right_N40, my_IIR_filter_firBlock_right_N39,
my_IIR_filter_firBlock_right_N38, my_IIR_filter_firBlock_right_N37,
my_IIR_filter_firBlock_right_N36, my_IIR_filter_firBlock_right_N35,
my_IIR_filter_firBlock_right_N34, my_IIR_filter_firBlock_right_N33,
my_IIR_filter_firBlock_right_N32, my_IIR_filter_firBlock_right_N31,
my_IIR_filter_firBlock_right_N30, my_IIR_filter_firBlock_right_N29,
my_IIR_filter_firBlock_right_N28, my_IIR_filter_firBlock_right_N27,
my_IIR_filter_firBlock_right_N26, my_IIR_filter_firBlock_right_N25,
my_IIR_filter_firBlock_right_N24, my_IIR_filter_firBlock_right_N23,
my_IIR_filter_firBlock_right_N22, my_IIR_filter_firBlock_right_N21,
my_IIR_filter_firBlock_right_N20, my_IIR_filter_firBlock_right_N19,
my_IIR_filter_firBlock_right_N18, my_IIR_filter_firBlock_right_N17,
my_IIR_filter_firBlock_right_N16, my_IIR_filter_firBlock_right_N15,
my_IIR_filter_firBlock_right_N14, my_IIR_filter_firBlock_right_N13,
my_IIR_filter_firBlock_right_N12, my_IIR_filter_firBlock_right_N11,
my_IIR_filter_firBlock_right_N10, my_IIR_filter_firBlock_right_N9,
my_IIR_filter_firBlock_right_N8, my_IIR_filter_firBlock_right_N7,
my_IIR_filter_firBlock_right_N6, my_IIR_filter_firBlock_right_N5,
my_IIR_filter_firBlock_right_N4, my_IIR_filter_firBlock_right_N3,
my_IIR_filter_firBlock_right_N2, my_IIR_filter_firBlock_right_N1,
my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10_39,
n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746;
wire [5:1] inData_in;
wire [30:2] outData_in;
wire [31:0] leftOut;
wire [31:0] rightOut;
wire [287:0] my_IIR_filter_firBlock_left_firStep;
wire [114:0] my_IIR_filter_firBlock_left_multProducts;
wire [31:0] my_IIR_filter_firBlock_left_Y_in;
wire [38:6] my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192;
wire [93:0] my_IIR_filter_firBlock_right_firStep;
wire [117:0] my_IIR_filter_firBlock_right_multProducts;
wire [31:0] my_IIR_filter_firBlock_right_Y_in;
wire [38:7] my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192;
wire [38:1] my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189;
wire [34:1] my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10;

dff inData_in_reg_31_ ( clk, n606_r, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, inData_31 );
not U_inv0 ( n39, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv1 ( n606_r, n606 );
dff inData_in_reg_3_ ( clk, n604_r, inData_in[3], inData_3 );
not U_inv2 ( n43, inData_in[3] );
not U_inv3 ( n604_r, n604 );
dff inData_in_reg_2_ ( clk, n604_r, inData_in[2], inData_2 );
not U_inv4 ( n42, inData_in[2] );
not U_inv5 ( n604_r, n604 );
dff inData_in_reg_0_ ( clk, n604_r, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[6], inData_0 );
not U_inv6 ( n41, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[6] );
not U_inv7 ( n604_r, n604 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__0_ ( clk, n604_r, my_IIR_filter_firBlock_left_firStep[256], my_IIR_filter_firBlock_left_multProducts[90] );
not U_inv8 ( n604_r, n604 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__1_ ( clk, n604_r, my_IIR_filter_firBlock_left_firStep[257], my_IIR_filter_firBlock_left_multProducts[91] );
not U_inv9 ( n604_r, n604 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__2_ ( clk, n604_r, my_IIR_filter_firBlock_left_firStep[258], my_IIR_filter_firBlock_left_multProducts[92] );
not U_inv10 ( n604_r, n604 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__3_ ( clk, n604_r, my_IIR_filter_firBlock_left_firStep[259], my_IIR_filter_firBlock_left_multProducts[93] );
not U_inv11 ( n604_r, n604 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__4_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[260], my_IIR_filter_firBlock_left_multProducts[94] );
not U_inv12 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__5_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[261], my_IIR_filter_firBlock_left_multProducts[95] );
not U_inv13 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__6_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[262], my_IIR_filter_firBlock_left_multProducts[96] );
not U_inv14 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__7_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[263], my_IIR_filter_firBlock_left_multProducts[97] );
not U_inv15 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__8_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[264], my_IIR_filter_firBlock_left_multProducts[98] );
not U_inv16 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__9_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[265], my_IIR_filter_firBlock_left_multProducts[99] );
not U_inv17 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__10_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[266], my_IIR_filter_firBlock_left_multProducts[100] );
not U_inv18 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__11_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[267], my_IIR_filter_firBlock_left_multProducts[101] );
not U_inv19 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__12_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[268], my_IIR_filter_firBlock_left_multProducts[102] );
not U_inv20 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__13_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[269], my_IIR_filter_firBlock_left_multProducts[103] );
not U_inv21 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__14_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[270], my_IIR_filter_firBlock_left_multProducts[104] );
not U_inv22 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__15_ ( clk, n603_r, my_IIR_filter_firBlock_left_firStep[271], my_IIR_filter_firBlock_left_multProducts[105] );
not U_inv23 ( n603_r, n603 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__16_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[272], my_IIR_filter_firBlock_left_multProducts[106] );
not U_inv24 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__17_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[273], my_IIR_filter_firBlock_left_multProducts[107] );
not U_inv25 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__18_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[274], my_IIR_filter_firBlock_left_multProducts[108] );
not U_inv26 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__19_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[275], my_IIR_filter_firBlock_left_multProducts[109] );
not U_inv27 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__20_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[276], my_IIR_filter_firBlock_left_multProducts[110] );
not U_inv28 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__21_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[277], my_IIR_filter_firBlock_left_multProducts[111] );
not U_inv29 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__22_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[278], my_IIR_filter_firBlock_left_multProducts[112] );
not U_inv30 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__23_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[279], my_IIR_filter_firBlock_left_multProducts[113] );
not U_inv31 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__24_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[280], my_IIR_filter_firBlock_left_multProducts[114] );
not U_inv32 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__25_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[281], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv33 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__26_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[282], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv34 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__27_ ( clk, n602_r, my_IIR_filter_firBlock_left_firStep[283], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv35 ( n602_r, n602 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__28_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[284], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv36 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__29_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[285], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv37 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__30_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[286], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv38 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_0__31_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[287], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
not U_inv39 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__0_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[224], my_IIR_filter_firBlock_left_N1 );
not U_inv40 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__1_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[225], my_IIR_filter_firBlock_left_N2 );
not U_inv41 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__2_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[226], my_IIR_filter_firBlock_left_N3 );
not U_inv42 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__3_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[227], my_IIR_filter_firBlock_left_N4 );
not U_inv43 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__4_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[228], my_IIR_filter_firBlock_left_N5 );
not U_inv44 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__5_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[229], my_IIR_filter_firBlock_left_N6 );
not U_inv45 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__6_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[230], my_IIR_filter_firBlock_left_N7 );
not U_inv46 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__7_ ( clk, n601_r, my_IIR_filter_firBlock_left_firStep[231], my_IIR_filter_firBlock_left_N8 );
not U_inv47 ( n601_r, n601 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__8_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[232], my_IIR_filter_firBlock_left_N9 );
not U_inv48 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__9_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[233], my_IIR_filter_firBlock_left_N10 );
not U_inv49 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__10_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[234], my_IIR_filter_firBlock_left_N11 );
not U_inv50 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__11_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[235], my_IIR_filter_firBlock_left_N12 );
not U_inv51 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__12_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[236], my_IIR_filter_firBlock_left_N13 );
not U_inv52 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__13_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[237], my_IIR_filter_firBlock_left_N14 );
not U_inv53 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__14_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[238], my_IIR_filter_firBlock_left_N15 );
not U_inv54 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__15_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[239], my_IIR_filter_firBlock_left_N16 );
not U_inv55 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__16_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[240], my_IIR_filter_firBlock_left_N17 );
not U_inv56 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__17_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[241], my_IIR_filter_firBlock_left_N18 );
not U_inv57 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__18_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[242], my_IIR_filter_firBlock_left_N19 );
not U_inv58 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__19_ ( clk, n600_r, my_IIR_filter_firBlock_left_firStep[243], my_IIR_filter_firBlock_left_N20 );
not U_inv59 ( n600_r, n600 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__20_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[244], my_IIR_filter_firBlock_left_N21 );
not U_inv60 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__21_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[245], my_IIR_filter_firBlock_left_N22 );
not U_inv61 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__22_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[246], my_IIR_filter_firBlock_left_N23 );
not U_inv62 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__23_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[247], my_IIR_filter_firBlock_left_N24 );
not U_inv63 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__24_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[248], my_IIR_filter_firBlock_left_N25 );
not U_inv64 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__25_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[249], my_IIR_filter_firBlock_left_N26 );
not U_inv65 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__26_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[250], my_IIR_filter_firBlock_left_N27 );
not U_inv66 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__27_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[251], my_IIR_filter_firBlock_left_N28 );
not U_inv67 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__28_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[252], my_IIR_filter_firBlock_left_N29 );
not U_inv68 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__29_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[253], my_IIR_filter_firBlock_left_N30 );
not U_inv69 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__30_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[254], my_IIR_filter_firBlock_left_N31 );
not U_inv70 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_1__31_ ( clk, n599_r, my_IIR_filter_firBlock_left_firStep[255], my_IIR_filter_firBlock_left_N32 );
not U_inv71 ( n599_r, n599 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__0_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[192], my_IIR_filter_firBlock_left_N33 );
not U_inv72 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__1_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[193], my_IIR_filter_firBlock_left_N34 );
not U_inv73 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__2_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[194], my_IIR_filter_firBlock_left_N35 );
not U_inv74 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__3_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[195], my_IIR_filter_firBlock_left_N36 );
not U_inv75 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__4_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[196], my_IIR_filter_firBlock_left_N37 );
not U_inv76 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__5_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[197], my_IIR_filter_firBlock_left_N38 );
not U_inv77 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__6_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[198], my_IIR_filter_firBlock_left_N39 );
not U_inv78 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__7_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[199], my_IIR_filter_firBlock_left_N40 );
not U_inv79 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__8_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[200], my_IIR_filter_firBlock_left_N41 );
not U_inv80 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__9_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[201], my_IIR_filter_firBlock_left_N42 );
not U_inv81 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__10_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[202], my_IIR_filter_firBlock_left_N43 );
not U_inv82 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__11_ ( clk, n598_r, my_IIR_filter_firBlock_left_firStep[203], my_IIR_filter_firBlock_left_N44 );
not U_inv83 ( n598_r, n598 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__12_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[204], my_IIR_filter_firBlock_left_N45 );
not U_inv84 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__13_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[205], my_IIR_filter_firBlock_left_N46 );
not U_inv85 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__14_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[206], my_IIR_filter_firBlock_left_N47 );
not U_inv86 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__15_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[207], my_IIR_filter_firBlock_left_N48 );
not U_inv87 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__16_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[208], my_IIR_filter_firBlock_left_N49 );
not U_inv88 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__17_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[209], my_IIR_filter_firBlock_left_N50 );
not U_inv89 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__18_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[210], my_IIR_filter_firBlock_left_N51 );
not U_inv90 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__19_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[211], my_IIR_filter_firBlock_left_N52 );
not U_inv91 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__20_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[212], my_IIR_filter_firBlock_left_N53 );
not U_inv92 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__21_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[213], my_IIR_filter_firBlock_left_N54 );
not U_inv93 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__22_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[214], my_IIR_filter_firBlock_left_N55 );
not U_inv94 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__23_ ( clk, n597_r, my_IIR_filter_firBlock_left_firStep[215], my_IIR_filter_firBlock_left_N56 );
not U_inv95 ( n597_r, n597 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__24_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[216], my_IIR_filter_firBlock_left_N57 );
not U_inv96 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__25_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[217], my_IIR_filter_firBlock_left_N58 );
not U_inv97 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__26_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[218], my_IIR_filter_firBlock_left_N59 );
not U_inv98 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__27_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[219], my_IIR_filter_firBlock_left_N60 );
not U_inv99 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__28_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[220], my_IIR_filter_firBlock_left_N61 );
not U_inv100 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__29_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[221], my_IIR_filter_firBlock_left_N62 );
not U_inv101 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__30_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[222], my_IIR_filter_firBlock_left_N63 );
not U_inv102 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_2__31_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[223], my_IIR_filter_firBlock_left_N64 );
not U_inv103 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__0_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[160], my_IIR_filter_firBlock_left_N65 );
not U_inv104 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__1_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[161], my_IIR_filter_firBlock_left_N66 );
not U_inv105 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__2_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[162], my_IIR_filter_firBlock_left_N67 );
not U_inv106 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__3_ ( clk, n596_r, my_IIR_filter_firBlock_left_firStep[163], my_IIR_filter_firBlock_left_N68 );
not U_inv107 ( n596_r, n596 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__4_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[164], my_IIR_filter_firBlock_left_N69 );
not U_inv108 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__5_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[165], my_IIR_filter_firBlock_left_N70 );
not U_inv109 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__6_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[166], my_IIR_filter_firBlock_left_N71 );
not U_inv110 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__7_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[167], my_IIR_filter_firBlock_left_N72 );
not U_inv111 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__8_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[168], my_IIR_filter_firBlock_left_N73 );
not U_inv112 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__9_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[169], my_IIR_filter_firBlock_left_N74 );
not U_inv113 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__10_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[170], my_IIR_filter_firBlock_left_N75 );
not U_inv114 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__11_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[171], my_IIR_filter_firBlock_left_N76 );
not U_inv115 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__12_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[172], my_IIR_filter_firBlock_left_N77 );
not U_inv116 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__13_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[173], my_IIR_filter_firBlock_left_N78 );
not U_inv117 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__14_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[174], my_IIR_filter_firBlock_left_N79 );
not U_inv118 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__15_ ( clk, n595_r, my_IIR_filter_firBlock_left_firStep[175], my_IIR_filter_firBlock_left_N80 );
not U_inv119 ( n595_r, n595 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__16_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[176], my_IIR_filter_firBlock_left_N81 );
not U_inv120 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__17_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[177], my_IIR_filter_firBlock_left_N82 );
not U_inv121 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__18_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[178], my_IIR_filter_firBlock_left_N83 );
not U_inv122 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__19_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[179], my_IIR_filter_firBlock_left_N84 );
not U_inv123 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__20_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[180], my_IIR_filter_firBlock_left_N85 );
not U_inv124 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__21_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[181], my_IIR_filter_firBlock_left_N86 );
not U_inv125 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__22_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[182], my_IIR_filter_firBlock_left_N87 );
not U_inv126 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__23_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[183], my_IIR_filter_firBlock_left_N88 );
not U_inv127 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__24_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[184], my_IIR_filter_firBlock_left_N89 );
not U_inv128 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__25_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[185], my_IIR_filter_firBlock_left_N90 );
not U_inv129 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__26_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[186], my_IIR_filter_firBlock_left_N91 );
not U_inv130 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__27_ ( clk, n594_r, my_IIR_filter_firBlock_left_firStep[187], my_IIR_filter_firBlock_left_N92 );
not U_inv131 ( n594_r, n594 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__28_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[188], my_IIR_filter_firBlock_left_N93 );
not U_inv132 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__29_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[189], my_IIR_filter_firBlock_left_N94 );
not U_inv133 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__30_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[190], my_IIR_filter_firBlock_left_N95 );
not U_inv134 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_3__31_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[191], my_IIR_filter_firBlock_left_N96 );
not U_inv135 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__0_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[128], my_IIR_filter_firBlock_left_N97 );
not U_inv136 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__1_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[129], my_IIR_filter_firBlock_left_N98 );
not U_inv137 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__2_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[130], my_IIR_filter_firBlock_left_N99 );
not U_inv138 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__3_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[131], my_IIR_filter_firBlock_left_N100 );
not U_inv139 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__4_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[132], my_IIR_filter_firBlock_left_N101 );
not U_inv140 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__5_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[133], my_IIR_filter_firBlock_left_N102 );
not U_inv141 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__6_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[134], my_IIR_filter_firBlock_left_N103 );
not U_inv142 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__7_ ( clk, n593_r, my_IIR_filter_firBlock_left_firStep[135], my_IIR_filter_firBlock_left_N104 );
not U_inv143 ( n593_r, n593 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__8_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[136], my_IIR_filter_firBlock_left_N105 );
not U_inv144 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__9_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[137], my_IIR_filter_firBlock_left_N106 );
not U_inv145 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__10_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[138], my_IIR_filter_firBlock_left_N107 );
not U_inv146 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__11_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[139], my_IIR_filter_firBlock_left_N108 );
not U_inv147 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__12_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[140], my_IIR_filter_firBlock_left_N109 );
not U_inv148 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__13_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[141], my_IIR_filter_firBlock_left_N110 );
not U_inv149 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__14_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[142], my_IIR_filter_firBlock_left_N111 );
not U_inv150 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__15_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[143], my_IIR_filter_firBlock_left_N112 );
not U_inv151 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__16_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[144], my_IIR_filter_firBlock_left_N113 );
not U_inv152 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__17_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[145], my_IIR_filter_firBlock_left_N114 );
not U_inv153 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__18_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[146], my_IIR_filter_firBlock_left_N115 );
not U_inv154 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__19_ ( clk, n592_r, my_IIR_filter_firBlock_left_firStep[147], my_IIR_filter_firBlock_left_N116 );
not U_inv155 ( n592_r, n592 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__20_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[148], my_IIR_filter_firBlock_left_N117 );
not U_inv156 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__21_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[149], my_IIR_filter_firBlock_left_N118 );
not U_inv157 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__22_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[150], my_IIR_filter_firBlock_left_N119 );
not U_inv158 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__23_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[151], my_IIR_filter_firBlock_left_N120 );
not U_inv159 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__24_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[152], my_IIR_filter_firBlock_left_N121 );
not U_inv160 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__25_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[153], my_IIR_filter_firBlock_left_N122 );
not U_inv161 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__26_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[154], my_IIR_filter_firBlock_left_N123 );
not U_inv162 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__27_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[155], my_IIR_filter_firBlock_left_N124 );
not U_inv163 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__28_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[156], my_IIR_filter_firBlock_left_N125 );
not U_inv164 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__29_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[157], my_IIR_filter_firBlock_left_N126 );
not U_inv165 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__30_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[158], my_IIR_filter_firBlock_left_N127 );
not U_inv166 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_4__31_ ( clk, n591_r, my_IIR_filter_firBlock_left_firStep[159], my_IIR_filter_firBlock_left_N128 );
not U_inv167 ( n591_r, n591 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__0_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[96], my_IIR_filter_firBlock_left_N129 );
not U_inv168 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__1_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[97], my_IIR_filter_firBlock_left_N130 );
not U_inv169 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__2_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[98], my_IIR_filter_firBlock_left_N131 );
not U_inv170 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__3_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[99], my_IIR_filter_firBlock_left_N132 );
not U_inv171 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__4_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[100], my_IIR_filter_firBlock_left_N133 );
not U_inv172 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__5_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[101], my_IIR_filter_firBlock_left_N134 );
not U_inv173 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__6_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[102], my_IIR_filter_firBlock_left_N135 );
not U_inv174 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__7_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[103], my_IIR_filter_firBlock_left_N136 );
not U_inv175 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__8_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[104], my_IIR_filter_firBlock_left_N137 );
not U_inv176 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__9_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[105], my_IIR_filter_firBlock_left_N138 );
not U_inv177 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__10_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[106], my_IIR_filter_firBlock_left_N139 );
not U_inv178 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__11_ ( clk, n590_r, my_IIR_filter_firBlock_left_firStep[107], my_IIR_filter_firBlock_left_N140 );
not U_inv179 ( n590_r, n590 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__12_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[108], my_IIR_filter_firBlock_left_N141 );
not U_inv180 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__13_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[109], my_IIR_filter_firBlock_left_N142 );
not U_inv181 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__14_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[110], my_IIR_filter_firBlock_left_N143 );
not U_inv182 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__15_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[111], my_IIR_filter_firBlock_left_N144 );
not U_inv183 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__16_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[112], my_IIR_filter_firBlock_left_N145 );
not U_inv184 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__17_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[113], my_IIR_filter_firBlock_left_N146 );
not U_inv185 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__18_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[114], my_IIR_filter_firBlock_left_N147 );
not U_inv186 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__19_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[115], my_IIR_filter_firBlock_left_N148 );
not U_inv187 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__20_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[116], my_IIR_filter_firBlock_left_N149 );
not U_inv188 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__21_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[117], my_IIR_filter_firBlock_left_N150 );
not U_inv189 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__22_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[118], my_IIR_filter_firBlock_left_N151 );
not U_inv190 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__23_ ( clk, n589_r, my_IIR_filter_firBlock_left_firStep[119], my_IIR_filter_firBlock_left_N152 );
not U_inv191 ( n589_r, n589 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__24_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[120], my_IIR_filter_firBlock_left_N153 );
not U_inv192 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__25_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[121], my_IIR_filter_firBlock_left_N154 );
not U_inv193 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__26_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[122], my_IIR_filter_firBlock_left_N155 );
not U_inv194 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__27_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[123], my_IIR_filter_firBlock_left_N156 );
not U_inv195 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__28_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[124], my_IIR_filter_firBlock_left_N157 );
not U_inv196 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__29_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[125], my_IIR_filter_firBlock_left_N158 );
not U_inv197 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__30_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[126], my_IIR_filter_firBlock_left_N159 );
not U_inv198 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_5__31_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[127], my_IIR_filter_firBlock_left_N160 );
not U_inv199 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__0_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[64], my_IIR_filter_firBlock_left_N161 );
not U_inv200 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__1_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[65], my_IIR_filter_firBlock_left_N162 );
not U_inv201 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__2_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[66], my_IIR_filter_firBlock_left_N163 );
not U_inv202 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__3_ ( clk, n588_r, my_IIR_filter_firBlock_left_firStep[67], my_IIR_filter_firBlock_left_N164 );
not U_inv203 ( n588_r, n588 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__4_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[68], my_IIR_filter_firBlock_left_N165 );
not U_inv204 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__5_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[69], my_IIR_filter_firBlock_left_N166 );
not U_inv205 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__6_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[70], my_IIR_filter_firBlock_left_N167 );
not U_inv206 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__7_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[71], my_IIR_filter_firBlock_left_N168 );
not U_inv207 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__8_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[72], my_IIR_filter_firBlock_left_N169 );
not U_inv208 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__9_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[73], my_IIR_filter_firBlock_left_N170 );
not U_inv209 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__10_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[74], my_IIR_filter_firBlock_left_N171 );
not U_inv210 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__11_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[75], my_IIR_filter_firBlock_left_N172 );
not U_inv211 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__12_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[76], my_IIR_filter_firBlock_left_N173 );
not U_inv212 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__13_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[77], my_IIR_filter_firBlock_left_N174 );
not U_inv213 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__14_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[78], my_IIR_filter_firBlock_left_N175 );
not U_inv214 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__15_ ( clk, n587_r, my_IIR_filter_firBlock_left_firStep[79], my_IIR_filter_firBlock_left_N176 );
not U_inv215 ( n587_r, n587 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__16_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[80], my_IIR_filter_firBlock_left_N177 );
not U_inv216 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__17_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[81], my_IIR_filter_firBlock_left_N178 );
not U_inv217 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__18_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[82], my_IIR_filter_firBlock_left_N179 );
not U_inv218 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__19_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[83], my_IIR_filter_firBlock_left_N180 );
not U_inv219 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__20_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[84], my_IIR_filter_firBlock_left_N181 );
not U_inv220 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__21_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[85], my_IIR_filter_firBlock_left_N182 );
not U_inv221 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__22_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[86], my_IIR_filter_firBlock_left_N183 );
not U_inv222 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__23_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[87], my_IIR_filter_firBlock_left_N184 );
not U_inv223 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__24_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[88], my_IIR_filter_firBlock_left_N185 );
not U_inv224 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__25_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[89], my_IIR_filter_firBlock_left_N186 );
not U_inv225 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__26_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[90], my_IIR_filter_firBlock_left_N187 );
not U_inv226 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__27_ ( clk, n586_r, my_IIR_filter_firBlock_left_firStep[91], my_IIR_filter_firBlock_left_N188 );
not U_inv227 ( n586_r, n586 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__28_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[92], my_IIR_filter_firBlock_left_N189 );
not U_inv228 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__29_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[93], my_IIR_filter_firBlock_left_N190 );
not U_inv229 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__30_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[94], my_IIR_filter_firBlock_left_N191 );
not U_inv230 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_6__31_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[95], my_IIR_filter_firBlock_left_N192 );
not U_inv231 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__0_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[32], my_IIR_filter_firBlock_left_N193 );
not U_inv232 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__1_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[33], my_IIR_filter_firBlock_left_N194 );
not U_inv233 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__2_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[34], my_IIR_filter_firBlock_left_N195 );
not U_inv234 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__3_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[35], my_IIR_filter_firBlock_left_N196 );
not U_inv235 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__4_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[36], my_IIR_filter_firBlock_left_N197 );
not U_inv236 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__5_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[37], my_IIR_filter_firBlock_left_N198 );
not U_inv237 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__6_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[38], my_IIR_filter_firBlock_left_N199 );
not U_inv238 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__7_ ( clk, n585_r, my_IIR_filter_firBlock_left_firStep[39], my_IIR_filter_firBlock_left_N200 );
not U_inv239 ( n585_r, n585 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__8_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[40], my_IIR_filter_firBlock_left_N201 );
not U_inv240 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__9_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[41], my_IIR_filter_firBlock_left_N202 );
not U_inv241 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__10_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[42], my_IIR_filter_firBlock_left_N203 );
not U_inv242 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__11_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[43], my_IIR_filter_firBlock_left_N204 );
not U_inv243 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__12_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[44], my_IIR_filter_firBlock_left_N205 );
not U_inv244 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__13_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[45], my_IIR_filter_firBlock_left_N206 );
not U_inv245 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__14_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[46], my_IIR_filter_firBlock_left_N207 );
not U_inv246 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__15_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[47], my_IIR_filter_firBlock_left_N208 );
not U_inv247 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__16_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[48], my_IIR_filter_firBlock_left_N209 );
not U_inv248 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__17_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[49], my_IIR_filter_firBlock_left_N210 );
not U_inv249 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__18_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[50], my_IIR_filter_firBlock_left_N211 );
not U_inv250 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__19_ ( clk, n584_r, my_IIR_filter_firBlock_left_firStep[51], my_IIR_filter_firBlock_left_N212 );
not U_inv251 ( n584_r, n584 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__20_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[52], my_IIR_filter_firBlock_left_N213 );
not U_inv252 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__21_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[53], my_IIR_filter_firBlock_left_N214 );
not U_inv253 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__22_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[54], my_IIR_filter_firBlock_left_N215 );
not U_inv254 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__23_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[55], my_IIR_filter_firBlock_left_N216 );
not U_inv255 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__24_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[56], my_IIR_filter_firBlock_left_N217 );
not U_inv256 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__25_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[57], my_IIR_filter_firBlock_left_N218 );
not U_inv257 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__26_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[58], my_IIR_filter_firBlock_left_N219 );
not U_inv258 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__27_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[59], my_IIR_filter_firBlock_left_N220 );
not U_inv259 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__28_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[60], my_IIR_filter_firBlock_left_N221 );
not U_inv260 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__29_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[61], my_IIR_filter_firBlock_left_N222 );
not U_inv261 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__30_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[62], my_IIR_filter_firBlock_left_N223 );
not U_inv262 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_7__31_ ( clk, n583_r, my_IIR_filter_firBlock_left_firStep[63], my_IIR_filter_firBlock_left_N224 );
not U_inv263 ( n583_r, n583 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__0_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[0], my_IIR_filter_firBlock_left_N225 );
not U_inv264 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__1_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[1], my_IIR_filter_firBlock_left_N226 );
not U_inv265 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__2_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[2], my_IIR_filter_firBlock_left_N227 );
not U_inv266 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__3_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[3], my_IIR_filter_firBlock_left_N228 );
not U_inv267 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__4_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[4], my_IIR_filter_firBlock_left_N229 );
not U_inv268 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__5_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[5], my_IIR_filter_firBlock_left_N230 );
not U_inv269 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__6_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[6], my_IIR_filter_firBlock_left_N231 );
not U_inv270 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__7_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[7], my_IIR_filter_firBlock_left_N232 );
not U_inv271 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__8_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[8], my_IIR_filter_firBlock_left_N233 );
not U_inv272 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__9_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[9], my_IIR_filter_firBlock_left_N234 );
not U_inv273 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__10_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[10], my_IIR_filter_firBlock_left_N235 );
not U_inv274 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__11_ ( clk, n582_r, my_IIR_filter_firBlock_left_firStep[11], my_IIR_filter_firBlock_left_N236 );
not U_inv275 ( n582_r, n582 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__12_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[12], my_IIR_filter_firBlock_left_N237 );
not U_inv276 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__13_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[13], my_IIR_filter_firBlock_left_N238 );
not U_inv277 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__14_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[14], my_IIR_filter_firBlock_left_N239 );
not U_inv278 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__15_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[15], my_IIR_filter_firBlock_left_N240 );
not U_inv279 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__16_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[16], my_IIR_filter_firBlock_left_N241 );
not U_inv280 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__17_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[17], my_IIR_filter_firBlock_left_N242 );
not U_inv281 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__18_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[18], my_IIR_filter_firBlock_left_N243 );
not U_inv282 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__19_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[19], my_IIR_filter_firBlock_left_N244 );
not U_inv283 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__20_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[20], my_IIR_filter_firBlock_left_N245 );
not U_inv284 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__21_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[21], my_IIR_filter_firBlock_left_N246 );
not U_inv285 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__22_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[22], my_IIR_filter_firBlock_left_N247 );
not U_inv286 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__23_ ( clk, n581_r, my_IIR_filter_firBlock_left_firStep[23], my_IIR_filter_firBlock_left_N248 );
not U_inv287 ( n581_r, n581 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__24_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[24], my_IIR_filter_firBlock_left_N249 );
not U_inv288 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__25_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[25], my_IIR_filter_firBlock_left_N250 );
not U_inv289 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__26_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[26], my_IIR_filter_firBlock_left_N251 );
not U_inv290 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__27_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[27], my_IIR_filter_firBlock_left_N252 );
not U_inv291 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__28_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[28], my_IIR_filter_firBlock_left_N253 );
not U_inv292 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__29_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[29], my_IIR_filter_firBlock_left_N254 );
not U_inv293 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__30_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[30], my_IIR_filter_firBlock_left_N255 );
not U_inv294 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__0_ ( clk, n580_r, my_IIR_filter_firBlock_left_Y_in[0], my_IIR_filter_firBlock_left_N257 );
not U_inv295 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__1_ ( clk, n580_r, my_IIR_filter_firBlock_left_Y_in[1], my_IIR_filter_firBlock_left_N258 );
not U_inv296 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__2_ ( clk, n580_r, my_IIR_filter_firBlock_left_Y_in[2], my_IIR_filter_firBlock_left_N259 );
not U_inv297 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__3_ ( clk, n580_r, my_IIR_filter_firBlock_left_Y_in[3], my_IIR_filter_firBlock_left_N260 );
not U_inv298 ( n580_r, n580 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__4_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[4], my_IIR_filter_firBlock_left_N261 );
not U_inv299 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__5_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[5], my_IIR_filter_firBlock_left_N262 );
not U_inv300 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__6_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[6], my_IIR_filter_firBlock_left_N263 );
not U_inv301 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__7_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[7], my_IIR_filter_firBlock_left_N264 );
not U_inv302 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__8_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[8], my_IIR_filter_firBlock_left_N265 );
not U_inv303 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__9_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[9], my_IIR_filter_firBlock_left_N266 );
not U_inv304 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__10_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[10], my_IIR_filter_firBlock_left_N267 );
not U_inv305 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__11_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[11], my_IIR_filter_firBlock_left_N268 );
not U_inv306 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__12_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[12], my_IIR_filter_firBlock_left_N269 );
not U_inv307 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__13_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[13], my_IIR_filter_firBlock_left_N270 );
not U_inv308 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__14_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[14], my_IIR_filter_firBlock_left_N271 );
not U_inv309 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__15_ ( clk, n579_r, my_IIR_filter_firBlock_left_Y_in[15], my_IIR_filter_firBlock_left_N272 );
not U_inv310 ( n579_r, n579 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__16_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[16], my_IIR_filter_firBlock_left_N273 );
not U_inv311 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__17_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[17], my_IIR_filter_firBlock_left_N274 );
not U_inv312 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__18_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[18], my_IIR_filter_firBlock_left_N275 );
not U_inv313 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__19_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[19], my_IIR_filter_firBlock_left_N276 );
not U_inv314 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__20_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[20], my_IIR_filter_firBlock_left_N277 );
not U_inv315 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__21_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[21], my_IIR_filter_firBlock_left_N278 );
not U_inv316 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__22_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[22], my_IIR_filter_firBlock_left_N279 );
not U_inv317 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__23_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[23], my_IIR_filter_firBlock_left_N280 );
not U_inv318 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__24_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[24], my_IIR_filter_firBlock_left_N281 );
not U_inv319 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__25_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[25], my_IIR_filter_firBlock_left_N282 );
not U_inv320 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__26_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[26], my_IIR_filter_firBlock_left_N283 );
not U_inv321 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__27_ ( clk, n578_r, my_IIR_filter_firBlock_left_Y_in[27], my_IIR_filter_firBlock_left_N284 );
not U_inv322 ( n578_r, n578 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__28_ ( clk, n577_r, my_IIR_filter_firBlock_left_Y_in[28], my_IIR_filter_firBlock_left_N285 );
not U_inv323 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__29_ ( clk, n577_r, my_IIR_filter_firBlock_left_Y_in[29], my_IIR_filter_firBlock_left_N286 );
not U_inv324 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__30_ ( clk, n577_r, my_IIR_filter_firBlock_left_Y_in[30], my_IIR_filter_firBlock_left_N287 );
not U_inv325 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_firStep_reg_9__31_ ( clk, n577_r, my_IIR_filter_firBlock_left_Y_in[31], my_IIR_filter_firBlock_left_N288 );
not U_inv326 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_0_ ( clk, n577_r, leftOut[0], my_IIR_filter_firBlock_left_Y_in[0] );
not U_inv327 ( n208, leftOut[0] );
not U_inv328 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_1_ ( clk, n577_r, leftOut[1], my_IIR_filter_firBlock_left_Y_in[1] );
not U_inv329 ( n127, leftOut[1] );
not U_inv330 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_2_ ( clk, n577_r, leftOut[2], my_IIR_filter_firBlock_left_Y_in[2] );
not U_inv331 ( n263, leftOut[2] );
not U_inv332 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_3_ ( clk, n577_r, leftOut[3], my_IIR_filter_firBlock_left_Y_in[3] );
not U_inv333 ( n143, leftOut[3] );
not U_inv334 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_4_ ( clk, n577_r, leftOut[4], my_IIR_filter_firBlock_left_Y_in[4] );
not U_inv335 ( n279, leftOut[4] );
not U_inv336 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_5_ ( clk, n577_r, leftOut[5], my_IIR_filter_firBlock_left_Y_in[5] );
not U_inv337 ( n156, leftOut[5] );
not U_inv338 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_6_ ( clk, n577_r, leftOut[6], my_IIR_filter_firBlock_left_Y_in[6] );
not U_inv339 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_7_ ( clk, n577_r, leftOut[7], my_IIR_filter_firBlock_left_Y_in[7] );
not U_inv340 ( n577_r, n577 );
dff my_IIR_filter_firBlock_left_Y_reg_8_ ( clk, n576_r, leftOut[8], my_IIR_filter_firBlock_left_Y_in[8] );
not U_inv341 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_9_ ( clk, n576_r, leftOut[9], my_IIR_filter_firBlock_left_Y_in[9] );
not U_inv342 ( n146, leftOut[9] );
not U_inv343 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_10_ ( clk, n576_r, leftOut[10], my_IIR_filter_firBlock_left_Y_in[10] );
not U_inv344 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_11_ ( clk, n576_r, leftOut[11], my_IIR_filter_firBlock_left_Y_in[11] );
not U_inv345 ( n149, leftOut[11] );
not U_inv346 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_12_ ( clk, n576_r, leftOut[12], my_IIR_filter_firBlock_left_Y_in[12] );
not U_inv347 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_13_ ( clk, n576_r, leftOut[13], my_IIR_filter_firBlock_left_Y_in[13] );
not U_inv348 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_14_ ( clk, n576_r, leftOut[14], my_IIR_filter_firBlock_left_Y_in[14] );
not U_inv349 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_15_ ( clk, n576_r, leftOut[15], my_IIR_filter_firBlock_left_Y_in[15] );
not U_inv350 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_16_ ( clk, n576_r, leftOut[16], my_IIR_filter_firBlock_left_Y_in[16] );
not U_inv351 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_17_ ( clk, n576_r, leftOut[17], my_IIR_filter_firBlock_left_Y_in[17] );
not U_inv352 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_18_ ( clk, n576_r, leftOut[18], my_IIR_filter_firBlock_left_Y_in[18] );
not U_inv353 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_19_ ( clk, n576_r, leftOut[19], my_IIR_filter_firBlock_left_Y_in[19] );
not U_inv354 ( n576_r, n576 );
dff my_IIR_filter_firBlock_left_Y_reg_20_ ( clk, n575_r, leftOut[20], my_IIR_filter_firBlock_left_Y_in[20] );
not U_inv355 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_21_ ( clk, n575_r, leftOut[21], my_IIR_filter_firBlock_left_Y_in[21] );
not U_inv356 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_22_ ( clk, n575_r, leftOut[22], my_IIR_filter_firBlock_left_Y_in[22] );
not U_inv357 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_23_ ( clk, n575_r, leftOut[23], my_IIR_filter_firBlock_left_Y_in[23] );
not U_inv358 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_24_ ( clk, n575_r, leftOut[24], my_IIR_filter_firBlock_left_Y_in[24] );
not U_inv359 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_25_ ( clk, n575_r, leftOut[25], my_IIR_filter_firBlock_left_Y_in[25] );
not U_inv360 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_26_ ( clk, n575_r, leftOut[26], my_IIR_filter_firBlock_left_Y_in[26] );
not U_inv361 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_27_ ( clk, n575_r, leftOut[27], my_IIR_filter_firBlock_left_Y_in[27] );
not U_inv362 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_28_ ( clk, n575_r, leftOut[28], my_IIR_filter_firBlock_left_Y_in[28] );
not U_inv363 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_29_ ( clk, n575_r, leftOut[29], my_IIR_filter_firBlock_left_Y_in[29] );
not U_inv364 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_30_ ( clk, n575_r, leftOut[30], my_IIR_filter_firBlock_left_Y_in[30] );
not U_inv365 ( n575_r, n575 );
dff my_IIR_filter_firBlock_left_Y_reg_31_ ( clk, n575_r, leftOut[31], my_IIR_filter_firBlock_left_Y_in[31] );
not U_inv366 ( n575_r, n575 );
dff my_IIR_filter_firBlock_right_Y_reg_31_ ( clk, n574_r, rightOut[31], my_IIR_filter_firBlock_right_Y_in[31] );
not U_inv367 ( n574_r, n574 );
dff outData_reg_0_ ( clk, n574_r, outData_0, n498 );
not U_inv368 ( n574_r, n574 );
dff outData_reg_1_ ( clk, n574_r, outData_1, n501 );
not U_inv369 ( n574_r, n574 );
dff outData_reg_2_ ( clk, n574_r, outData_2, n522 );
not U_inv370 ( n574_r, n574 );
dff outData_reg_3_ ( clk, n574_r, outData_3, n503 );
not U_inv371 ( n574_r, n574 );
dff outData_reg_4_ ( clk, n574_r, outData_4, n517 );
not U_inv372 ( n574_r, n574 );
dff outData_reg_5_ ( clk, n574_r, outData_5, outData_in[5] );
not U_inv373 ( n574_r, n574 );
dff outData_reg_6_ ( clk, n574_r, outData_6, n520 );
not U_inv374 ( n574_r, n574 );
dff outData_reg_7_ ( clk, n574_r, outData_7, outData_in[7] );
not U_inv375 ( n574_r, n574 );
dff outData_reg_8_ ( clk, n574_r, outData_8, n506 );
not U_inv376 ( n574_r, n574 );
dff outData_reg_9_ ( clk, n574_r, outData_9, n519 );
not U_inv377 ( n574_r, n574 );
dff outData_reg_10_ ( clk, n574_r, outData_10, n509 );
not U_inv378 ( n574_r, n574 );
dff outData_reg_11_ ( clk, n573_r, outData_11, n487 );
not U_inv379 ( n573_r, n573 );
dff outData_reg_12_ ( clk, n573_r, outData_12, n510 );
not U_inv380 ( n573_r, n573 );
dff outData_reg_13_ ( clk, n573_r, outData_13, n499 );
not U_inv381 ( n573_r, n573 );
dff outData_reg_14_ ( clk, n573_r, outData_14, n485 );
not U_inv382 ( n573_r, n573 );
dff outData_reg_15_ ( clk, n573_r, outData_15, n495 );
not U_inv383 ( n573_r, n573 );
dff outData_reg_16_ ( clk, n573_r, outData_16, outData_in[16] );
not U_inv384 ( n573_r, n573 );
dff outData_reg_17_ ( clk, n573_r, outData_17, n512 );
not U_inv385 ( n573_r, n573 );
dff outData_reg_18_ ( clk, n573_r, outData_18, outData_in[18] );
not U_inv386 ( n573_r, n573 );
dff outData_reg_19_ ( clk, n573_r, outData_19, n493 );
not U_inv387 ( n573_r, n573 );
dff outData_reg_20_ ( clk, n573_r, outData_20, outData_in[20] );
not U_inv388 ( n573_r, n573 );
dff outData_reg_21_ ( clk, n573_r, outData_21, n154 );
not U_inv389 ( n573_r, n573 );
dff outData_reg_22_ ( clk, n573_r, outData_22, n489 );
not U_inv390 ( n573_r, n573 );
dff outData_reg_23_ ( clk, n572_r, outData_23, n529 );
not U_inv391 ( n572_r, n572 );
dff outData_reg_24_ ( clk, n572_r, outData_24, n157 );
not U_inv392 ( n572_r, n572 );
dff outData_reg_25_ ( clk, n572_r, outData_25, n504 );
not U_inv393 ( n572_r, n572 );
dff outData_reg_26_ ( clk, n572_r, outData_26, n158 );
not U_inv394 ( n572_r, n572 );
dff outData_reg_27_ ( clk, n572_r, outData_27, n491 );
not U_inv395 ( n572_r, n572 );
dff outData_reg_28_ ( clk, n572_r, outData_28, n209 );
not U_inv396 ( n572_r, n572 );
dff outData_reg_29_ ( clk, n572_r, outData_29, n514 );
not U_inv397 ( n572_r, n572 );
dff outData_reg_30_ ( clk, n572_r, outData_30, outData_in[30] );
not U_inv398 ( n572_r, n572 );
dff outData_reg_31_ ( clk, n572_r, outData_31, n525 );
not U_inv399 ( n572_r, n572 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__0_ ( clk, n572_r, my_IIR_filter_firBlock_right_N1, my_IIR_filter_firBlock_right_multProducts[92] );
not U_inv400 ( n572_r, n572 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__1_ ( clk, n572_r, my_IIR_filter_firBlock_right_N2, my_IIR_filter_firBlock_right_multProducts[93] );
not U_inv401 ( n572_r, n572 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__2_ ( clk, n572_r, my_IIR_filter_firBlock_right_N3, my_IIR_filter_firBlock_right_multProducts[94] );
not U_inv402 ( n572_r, n572 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__3_ ( clk, n571_r, my_IIR_filter_firBlock_right_N4, my_IIR_filter_firBlock_right_multProducts[95] );
not U_inv403 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__4_ ( clk, n571_r, my_IIR_filter_firBlock_right_N5, my_IIR_filter_firBlock_right_multProducts[96] );
not U_inv404 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__5_ ( clk, n571_r, my_IIR_filter_firBlock_right_N6, my_IIR_filter_firBlock_right_multProducts[97] );
not U_inv405 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__6_ ( clk, n571_r, my_IIR_filter_firBlock_right_N7, my_IIR_filter_firBlock_right_multProducts[98] );
not U_inv406 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__7_ ( clk, n571_r, my_IIR_filter_firBlock_right_N8, my_IIR_filter_firBlock_right_multProducts[99] );
not U_inv407 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__8_ ( clk, n571_r, my_IIR_filter_firBlock_right_N9, my_IIR_filter_firBlock_right_multProducts[100] );
not U_inv408 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__9_ ( clk, n571_r, my_IIR_filter_firBlock_right_N10, my_IIR_filter_firBlock_right_multProducts[101] );
not U_inv409 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__10_ ( clk, n571_r, my_IIR_filter_firBlock_right_N11, my_IIR_filter_firBlock_right_multProducts[102] );
not U_inv410 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__11_ ( clk, n571_r, my_IIR_filter_firBlock_right_N12, my_IIR_filter_firBlock_right_multProducts[103] );
not U_inv411 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__12_ ( clk, n571_r, my_IIR_filter_firBlock_right_N13, my_IIR_filter_firBlock_right_multProducts[104] );
not U_inv412 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__13_ ( clk, n571_r, my_IIR_filter_firBlock_right_N14, my_IIR_filter_firBlock_right_multProducts[105] );
not U_inv413 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__14_ ( clk, n571_r, my_IIR_filter_firBlock_right_N15, my_IIR_filter_firBlock_right_multProducts[106] );
not U_inv414 ( n571_r, n571 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__15_ ( clk, n570_r, my_IIR_filter_firBlock_right_N16, my_IIR_filter_firBlock_right_multProducts[107] );
not U_inv415 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__16_ ( clk, n570_r, my_IIR_filter_firBlock_right_N17, my_IIR_filter_firBlock_right_multProducts[108] );
not U_inv416 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__17_ ( clk, n570_r, my_IIR_filter_firBlock_right_N18, my_IIR_filter_firBlock_right_multProducts[109] );
not U_inv417 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__18_ ( clk, n570_r, my_IIR_filter_firBlock_right_N19, my_IIR_filter_firBlock_right_multProducts[110] );
not U_inv418 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__19_ ( clk, n570_r, my_IIR_filter_firBlock_right_N20, my_IIR_filter_firBlock_right_multProducts[111] );
not U_inv419 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__20_ ( clk, n570_r, my_IIR_filter_firBlock_right_N21, my_IIR_filter_firBlock_right_multProducts[112] );
not U_inv420 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__21_ ( clk, n570_r, my_IIR_filter_firBlock_right_N22, my_IIR_filter_firBlock_right_multProducts[113] );
not U_inv421 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__22_ ( clk, n570_r, my_IIR_filter_firBlock_right_N23, my_IIR_filter_firBlock_right_multProducts[114] );
not U_inv422 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__23_ ( clk, n570_r, my_IIR_filter_firBlock_right_N24, my_IIR_filter_firBlock_right_multProducts[115] );
not U_inv423 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__24_ ( clk, n570_r, my_IIR_filter_firBlock_right_N25, my_IIR_filter_firBlock_right_multProducts[116] );
not U_inv424 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__31_ ( clk, n570_r, my_IIR_filter_firBlock_right_N32, my_IIR_filter_firBlock_right_multProducts[117] );
not U_inv425 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__29_ ( clk, n570_r, my_IIR_filter_firBlock_right_N30, my_IIR_filter_firBlock_right_multProducts[117] );
not U_inv426 ( n570_r, n570 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__27_ ( clk, n569_r, my_IIR_filter_firBlock_right_N28, my_IIR_filter_firBlock_right_multProducts[117] );
not U_inv427 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__25_ ( clk, n569_r, my_IIR_filter_firBlock_right_N26, my_IIR_filter_firBlock_right_multProducts[117] );
not U_inv428 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__26_ ( clk, n569_r, my_IIR_filter_firBlock_right_N27, my_IIR_filter_firBlock_right_multProducts[117] );
not U_inv429 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__28_ ( clk, n569_r, my_IIR_filter_firBlock_right_N29, my_IIR_filter_firBlock_right_multProducts[117] );
not U_inv430 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_0__30_ ( clk, n569_r, my_IIR_filter_firBlock_right_N31, my_IIR_filter_firBlock_right_multProducts[117] );
not U_inv431 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__0_ ( clk, n569_r, my_IIR_filter_firBlock_right_firStep[62], my_IIR_filter_firBlock_right_N1 );
not U_inv432 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__1_ ( clk, n569_r, my_IIR_filter_firBlock_right_firStep[63], my_IIR_filter_firBlock_right_N2 );
not U_inv433 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__2_ ( clk, n569_r, my_IIR_filter_firBlock_right_firStep[64], my_IIR_filter_firBlock_right_N3 );
not U_inv434 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__3_ ( clk, n569_r, my_IIR_filter_firBlock_right_firStep[65], my_IIR_filter_firBlock_right_N4 );
not U_inv435 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__4_ ( clk, n569_r, my_IIR_filter_firBlock_right_firStep[66], my_IIR_filter_firBlock_right_N5 );
not U_inv436 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__5_ ( clk, n569_r, my_IIR_filter_firBlock_right_firStep[67], my_IIR_filter_firBlock_right_N6 );
not U_inv437 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__6_ ( clk, n569_r, my_IIR_filter_firBlock_right_firStep[68], my_IIR_filter_firBlock_right_N7 );
not U_inv438 ( n569_r, n569 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__7_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[69], my_IIR_filter_firBlock_right_N8 );
not U_inv439 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__8_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[70], my_IIR_filter_firBlock_right_N9 );
not U_inv440 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__9_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[71], my_IIR_filter_firBlock_right_N10 );
not U_inv441 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__10_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[72], my_IIR_filter_firBlock_right_N11 );
not U_inv442 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__11_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[73], my_IIR_filter_firBlock_right_N12 );
not U_inv443 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__12_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[74], my_IIR_filter_firBlock_right_N13 );
not U_inv444 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__13_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[75], my_IIR_filter_firBlock_right_N14 );
not U_inv445 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__14_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[76], my_IIR_filter_firBlock_right_N15 );
not U_inv446 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__15_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[77], my_IIR_filter_firBlock_right_N16 );
not U_inv447 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__16_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[78], my_IIR_filter_firBlock_right_N17 );
not U_inv448 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__17_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[79], my_IIR_filter_firBlock_right_N18 );
not U_inv449 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__18_ ( clk, n568_r, my_IIR_filter_firBlock_right_firStep[80], my_IIR_filter_firBlock_right_N19 );
not U_inv450 ( n568_r, n568 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__19_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[81], my_IIR_filter_firBlock_right_N20 );
not U_inv451 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__20_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[82], my_IIR_filter_firBlock_right_N21 );
not U_inv452 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__21_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[83], my_IIR_filter_firBlock_right_N22 );
not U_inv453 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__22_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[84], my_IIR_filter_firBlock_right_N23 );
not U_inv454 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__23_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[85], my_IIR_filter_firBlock_right_N24 );
not U_inv455 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__24_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[86], my_IIR_filter_firBlock_right_N25 );
not U_inv456 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__25_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[87], my_IIR_filter_firBlock_right_N26 );
not U_inv457 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__26_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[88], my_IIR_filter_firBlock_right_N27 );
not U_inv458 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__27_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[89], my_IIR_filter_firBlock_right_N28 );
not U_inv459 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__28_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[90], my_IIR_filter_firBlock_right_N29 );
not U_inv460 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__29_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[91], my_IIR_filter_firBlock_right_N30 );
not U_inv461 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__30_ ( clk, n567_r, my_IIR_filter_firBlock_right_firStep[92], my_IIR_filter_firBlock_right_N31 );
not U_inv462 ( n567_r, n567 );
dff my_IIR_filter_firBlock_right_firStep_reg_1__31_ ( clk, n566_r, my_IIR_filter_firBlock_right_firStep[93], my_IIR_filter_firBlock_right_N32 );
not U_inv463 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__0_ ( clk, n566_r, my_IIR_filter_firBlock_right_N65, my_IIR_filter_firBlock_right_N33 );
not U_inv464 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__1_ ( clk, n566_r, my_IIR_filter_firBlock_right_N66, my_IIR_filter_firBlock_right_N34 );
not U_inv465 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__2_ ( clk, n566_r, my_IIR_filter_firBlock_right_N67, my_IIR_filter_firBlock_right_N35 );
not U_inv466 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__3_ ( clk, n566_r, my_IIR_filter_firBlock_right_N68, my_IIR_filter_firBlock_right_N36 );
not U_inv467 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__4_ ( clk, n566_r, my_IIR_filter_firBlock_right_N69, my_IIR_filter_firBlock_right_N37 );
not U_inv468 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__5_ ( clk, n566_r, my_IIR_filter_firBlock_right_N70, my_IIR_filter_firBlock_right_N38 );
not U_inv469 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__6_ ( clk, n566_r, my_IIR_filter_firBlock_right_N71, my_IIR_filter_firBlock_right_N39 );
not U_inv470 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__7_ ( clk, n566_r, my_IIR_filter_firBlock_right_N72, my_IIR_filter_firBlock_right_N40 );
not U_inv471 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__8_ ( clk, n566_r, my_IIR_filter_firBlock_right_N73, my_IIR_filter_firBlock_right_N41 );
not U_inv472 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__9_ ( clk, n566_r, my_IIR_filter_firBlock_right_N74, my_IIR_filter_firBlock_right_N42 );
not U_inv473 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__10_ ( clk, n566_r, my_IIR_filter_firBlock_right_N75, my_IIR_filter_firBlock_right_N43 );
not U_inv474 ( n566_r, n566 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__11_ ( clk, n565_r, my_IIR_filter_firBlock_right_N76, my_IIR_filter_firBlock_right_N44 );
not U_inv475 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__12_ ( clk, n565_r, my_IIR_filter_firBlock_right_N77, my_IIR_filter_firBlock_right_N45 );
not U_inv476 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__13_ ( clk, n565_r, my_IIR_filter_firBlock_right_N78, my_IIR_filter_firBlock_right_N46 );
not U_inv477 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__14_ ( clk, n565_r, my_IIR_filter_firBlock_right_N79, my_IIR_filter_firBlock_right_N47 );
not U_inv478 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__15_ ( clk, n565_r, my_IIR_filter_firBlock_right_N80, my_IIR_filter_firBlock_right_N48 );
not U_inv479 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__16_ ( clk, n565_r, my_IIR_filter_firBlock_right_N81, my_IIR_filter_firBlock_right_N49 );
not U_inv480 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__17_ ( clk, n565_r, my_IIR_filter_firBlock_right_N82, my_IIR_filter_firBlock_right_N50 );
not U_inv481 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__18_ ( clk, n565_r, my_IIR_filter_firBlock_right_N83, my_IIR_filter_firBlock_right_N51 );
not U_inv482 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__19_ ( clk, n565_r, my_IIR_filter_firBlock_right_N84, my_IIR_filter_firBlock_right_N52 );
not U_inv483 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__20_ ( clk, n565_r, my_IIR_filter_firBlock_right_N85, my_IIR_filter_firBlock_right_N53 );
not U_inv484 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__21_ ( clk, n565_r, my_IIR_filter_firBlock_right_N86, my_IIR_filter_firBlock_right_N54 );
not U_inv485 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__22_ ( clk, n565_r, my_IIR_filter_firBlock_right_N87, my_IIR_filter_firBlock_right_N55 );
not U_inv486 ( n565_r, n565 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__23_ ( clk, n564_r, my_IIR_filter_firBlock_right_N88, my_IIR_filter_firBlock_right_N56 );
not U_inv487 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__24_ ( clk, n564_r, my_IIR_filter_firBlock_right_N89, my_IIR_filter_firBlock_right_N57 );
not U_inv488 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__25_ ( clk, n564_r, my_IIR_filter_firBlock_right_N90, my_IIR_filter_firBlock_right_N58 );
not U_inv489 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__26_ ( clk, n564_r, my_IIR_filter_firBlock_right_N91, my_IIR_filter_firBlock_right_N59 );
not U_inv490 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__27_ ( clk, n564_r, my_IIR_filter_firBlock_right_N92, my_IIR_filter_firBlock_right_N60 );
not U_inv491 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__28_ ( clk, n564_r, my_IIR_filter_firBlock_right_N93, my_IIR_filter_firBlock_right_N61 );
not U_inv492 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__29_ ( clk, n564_r, my_IIR_filter_firBlock_right_N94, my_IIR_filter_firBlock_right_N62 );
not U_inv493 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__30_ ( clk, n564_r, my_IIR_filter_firBlock_right_N95, my_IIR_filter_firBlock_right_N63 );
not U_inv494 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_2__31_ ( clk, n564_r, my_IIR_filter_firBlock_right_N96, my_IIR_filter_firBlock_right_N64 );
not U_inv495 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__0_ ( clk, n564_r, my_IIR_filter_firBlock_right_firStep[31], my_IIR_filter_firBlock_right_N65 );
not U_inv496 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__1_ ( clk, n564_r, my_IIR_filter_firBlock_right_firStep[32], my_IIR_filter_firBlock_right_N66 );
not U_inv497 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__2_ ( clk, n564_r, my_IIR_filter_firBlock_right_firStep[33], my_IIR_filter_firBlock_right_N67 );
not U_inv498 ( n564_r, n564 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__3_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[34], my_IIR_filter_firBlock_right_N68 );
not U_inv499 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__4_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[35], my_IIR_filter_firBlock_right_N69 );
not U_inv500 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__5_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[36], my_IIR_filter_firBlock_right_N70 );
not U_inv501 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__6_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[37], my_IIR_filter_firBlock_right_N71 );
not U_inv502 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__7_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[38], my_IIR_filter_firBlock_right_N72 );
not U_inv503 ( n90, my_IIR_filter_firBlock_right_firStep[38] );
not U_inv504 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__8_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[39], my_IIR_filter_firBlock_right_N73 );
not U_inv505 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__9_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[40], my_IIR_filter_firBlock_right_N74 );
not U_inv506 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__10_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[41], my_IIR_filter_firBlock_right_N75 );
not U_inv507 ( n87, my_IIR_filter_firBlock_right_firStep[41] );
not U_inv508 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__11_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[42], my_IIR_filter_firBlock_right_N76 );
not U_inv509 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__12_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[43], my_IIR_filter_firBlock_right_N77 );
not U_inv510 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__13_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[44], my_IIR_filter_firBlock_right_N78 );
not U_inv511 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__14_ ( clk, n563_r, my_IIR_filter_firBlock_right_firStep[45], my_IIR_filter_firBlock_right_N79 );
not U_inv512 ( n84, my_IIR_filter_firBlock_right_firStep[45] );
not U_inv513 ( n563_r, n563 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__15_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[46], my_IIR_filter_firBlock_right_N80 );
not U_inv514 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__16_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[47], my_IIR_filter_firBlock_right_N81 );
not U_inv515 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__17_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[48], my_IIR_filter_firBlock_right_N82 );
not U_inv516 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__18_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[49], my_IIR_filter_firBlock_right_N83 );
not U_inv517 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__19_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[50], my_IIR_filter_firBlock_right_N84 );
not U_inv518 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__20_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[51], my_IIR_filter_firBlock_right_N85 );
not U_inv519 ( n81, my_IIR_filter_firBlock_right_firStep[51] );
not U_inv520 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__21_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[52], my_IIR_filter_firBlock_right_N86 );
not U_inv521 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__22_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[53], my_IIR_filter_firBlock_right_N87 );
not U_inv522 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__23_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[54], my_IIR_filter_firBlock_right_N88 );
not U_inv523 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__24_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[55], my_IIR_filter_firBlock_right_N89 );
not U_inv524 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__25_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[56], my_IIR_filter_firBlock_right_N90 );
not U_inv525 ( n537, my_IIR_filter_firBlock_right_firStep[56] );
not U_inv526 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__26_ ( clk, n562_r, my_IIR_filter_firBlock_right_firStep[57], my_IIR_filter_firBlock_right_N91 );
not U_inv527 ( n78, my_IIR_filter_firBlock_right_firStep[57] );
not U_inv528 ( n562_r, n562 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__27_ ( clk, n561_r, my_IIR_filter_firBlock_right_firStep[58], my_IIR_filter_firBlock_right_N92 );
not U_inv529 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__28_ ( clk, n561_r, my_IIR_filter_firBlock_right_firStep[59], my_IIR_filter_firBlock_right_N93 );
not U_inv530 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__29_ ( clk, n561_r, my_IIR_filter_firBlock_right_firStep[60], my_IIR_filter_firBlock_right_N94 );
not U_inv531 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__30_ ( clk, n561_r, my_IIR_filter_firBlock_right_firStep[61], my_IIR_filter_firBlock_right_N95 );
not U_inv532 ( n72, my_IIR_filter_firBlock_right_firStep[61] );
not U_inv533 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_3__31_ ( clk, n561_r, ex_wire0, my_IIR_filter_firBlock_right_N96 );
not U_inv534 ( n180, ex_wire0 );
not U_inv535 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__0_ ( clk, n561_r, my_IIR_filter_firBlock_right_N129, my_IIR_filter_firBlock_right_N97 );
not U_inv536 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__1_ ( clk, n561_r, my_IIR_filter_firBlock_right_N130, my_IIR_filter_firBlock_right_N98 );
not U_inv537 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__2_ ( clk, n561_r, my_IIR_filter_firBlock_right_N131, my_IIR_filter_firBlock_right_N99 );
not U_inv538 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__3_ ( clk, n561_r, my_IIR_filter_firBlock_right_N132, my_IIR_filter_firBlock_right_N100 );
not U_inv539 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__4_ ( clk, n561_r, my_IIR_filter_firBlock_right_N133, my_IIR_filter_firBlock_right_N101 );
not U_inv540 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__5_ ( clk, n561_r, my_IIR_filter_firBlock_right_N134, my_IIR_filter_firBlock_right_N102 );
not U_inv541 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__6_ ( clk, n561_r, my_IIR_filter_firBlock_right_N135, my_IIR_filter_firBlock_right_N103 );
not U_inv542 ( n561_r, n561 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__7_ ( clk, n560_r, my_IIR_filter_firBlock_right_N136, my_IIR_filter_firBlock_right_N104 );
not U_inv543 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__8_ ( clk, n560_r, my_IIR_filter_firBlock_right_N137, my_IIR_filter_firBlock_right_N105 );
not U_inv544 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__9_ ( clk, n560_r, my_IIR_filter_firBlock_right_N138, my_IIR_filter_firBlock_right_N106 );
not U_inv545 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__10_ ( clk, n560_r, my_IIR_filter_firBlock_right_N139, my_IIR_filter_firBlock_right_N107 );
not U_inv546 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__11_ ( clk, n560_r, my_IIR_filter_firBlock_right_N140, my_IIR_filter_firBlock_right_N108 );
not U_inv547 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__12_ ( clk, n560_r, my_IIR_filter_firBlock_right_N141, my_IIR_filter_firBlock_right_N109 );
not U_inv548 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__13_ ( clk, n560_r, my_IIR_filter_firBlock_right_N142, my_IIR_filter_firBlock_right_N110 );
not U_inv549 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__14_ ( clk, n560_r, my_IIR_filter_firBlock_right_N143, my_IIR_filter_firBlock_right_N111 );
not U_inv550 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__15_ ( clk, n560_r, my_IIR_filter_firBlock_right_N144, my_IIR_filter_firBlock_right_N112 );
not U_inv551 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__16_ ( clk, n560_r, my_IIR_filter_firBlock_right_N145, my_IIR_filter_firBlock_right_N113 );
not U_inv552 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__17_ ( clk, n560_r, my_IIR_filter_firBlock_right_N146, my_IIR_filter_firBlock_right_N114 );
not U_inv553 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__18_ ( clk, n560_r, my_IIR_filter_firBlock_right_N147, my_IIR_filter_firBlock_right_N115 );
not U_inv554 ( n560_r, n560 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__19_ ( clk, n559_r, my_IIR_filter_firBlock_right_N148, my_IIR_filter_firBlock_right_N116 );
not U_inv555 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__20_ ( clk, n559_r, my_IIR_filter_firBlock_right_N149, my_IIR_filter_firBlock_right_N117 );
not U_inv556 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__21_ ( clk, n559_r, my_IIR_filter_firBlock_right_N150, my_IIR_filter_firBlock_right_N118 );
not U_inv557 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__22_ ( clk, n559_r, my_IIR_filter_firBlock_right_N151, my_IIR_filter_firBlock_right_N119 );
not U_inv558 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__23_ ( clk, n559_r, my_IIR_filter_firBlock_right_N152, my_IIR_filter_firBlock_right_N120 );
not U_inv559 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__24_ ( clk, n559_r, my_IIR_filter_firBlock_right_N153, my_IIR_filter_firBlock_right_N121 );
not U_inv560 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__25_ ( clk, n559_r, my_IIR_filter_firBlock_right_N154, my_IIR_filter_firBlock_right_N122 );
not U_inv561 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__26_ ( clk, n559_r, my_IIR_filter_firBlock_right_N155, my_IIR_filter_firBlock_right_N123 );
not U_inv562 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__27_ ( clk, n559_r, my_IIR_filter_firBlock_right_N156, my_IIR_filter_firBlock_right_N124 );
not U_inv563 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__28_ ( clk, n559_r, my_IIR_filter_firBlock_right_N157, my_IIR_filter_firBlock_right_N125 );
not U_inv564 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__29_ ( clk, n559_r, my_IIR_filter_firBlock_right_N158, my_IIR_filter_firBlock_right_N126 );
not U_inv565 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__30_ ( clk, n559_r, my_IIR_filter_firBlock_right_N159, my_IIR_filter_firBlock_right_N127 );
not U_inv566 ( n559_r, n559 );
dff my_IIR_filter_firBlock_right_firStep_reg_4__31_ ( clk, n558_r, my_IIR_filter_firBlock_right_N160, my_IIR_filter_firBlock_right_N128 );
not U_inv567 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__0_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[0], my_IIR_filter_firBlock_right_N129 );
not U_inv568 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__1_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[1], my_IIR_filter_firBlock_right_N130 );
not U_inv569 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__2_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[2], my_IIR_filter_firBlock_right_N131 );
not U_inv570 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__3_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[3], my_IIR_filter_firBlock_right_N132 );
not U_inv571 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__4_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[4], my_IIR_filter_firBlock_right_N133 );
not U_inv572 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__5_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[5], my_IIR_filter_firBlock_right_N134 );
not U_inv573 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__6_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[6], my_IIR_filter_firBlock_right_N135 );
not U_inv574 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__7_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[7], my_IIR_filter_firBlock_right_N136 );
not U_inv575 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__8_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[8], my_IIR_filter_firBlock_right_N137 );
not U_inv576 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__9_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[9], my_IIR_filter_firBlock_right_N138 );
not U_inv577 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__10_ ( clk, n558_r, my_IIR_filter_firBlock_right_firStep[10], my_IIR_filter_firBlock_right_N139 );
not U_inv578 ( n558_r, n558 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__11_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[11], my_IIR_filter_firBlock_right_N140 );
not U_inv579 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__12_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[12], my_IIR_filter_firBlock_right_N141 );
not U_inv580 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__13_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[13], my_IIR_filter_firBlock_right_N142 );
not U_inv581 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__14_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[14], my_IIR_filter_firBlock_right_N143 );
not U_inv582 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__15_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[15], my_IIR_filter_firBlock_right_N144 );
not U_inv583 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__16_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[16], my_IIR_filter_firBlock_right_N145 );
not U_inv584 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__17_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[17], my_IIR_filter_firBlock_right_N146 );
not U_inv585 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__18_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[18], my_IIR_filter_firBlock_right_N147 );
not U_inv586 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__19_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[19], my_IIR_filter_firBlock_right_N148 );
not U_inv587 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__20_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[20], my_IIR_filter_firBlock_right_N149 );
not U_inv588 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__21_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[21], my_IIR_filter_firBlock_right_N150 );
not U_inv589 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__22_ ( clk, n557_r, my_IIR_filter_firBlock_right_firStep[22], my_IIR_filter_firBlock_right_N151 );
not U_inv590 ( n557_r, n557 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__23_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[23], my_IIR_filter_firBlock_right_N152 );
not U_inv591 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__24_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[24], my_IIR_filter_firBlock_right_N153 );
not U_inv592 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__25_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[25], my_IIR_filter_firBlock_right_N154 );
not U_inv593 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__26_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[26], my_IIR_filter_firBlock_right_N155 );
not U_inv594 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__27_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[27], my_IIR_filter_firBlock_right_N156 );
not U_inv595 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__28_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[28], my_IIR_filter_firBlock_right_N157 );
not U_inv596 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__29_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[29], my_IIR_filter_firBlock_right_N158 );
not U_inv597 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__30_ ( clk, n556_r, my_IIR_filter_firBlock_right_firStep[30], my_IIR_filter_firBlock_right_N159 );
not U_inv598 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_5__31_ ( clk, n556_r, ex_wire1, my_IIR_filter_firBlock_right_N160 );
not U_inv599 ( n195, ex_wire1 );
not U_inv600 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__0_ ( clk, n556_r, my_IIR_filter_firBlock_right_Y_in[0], my_IIR_filter_firBlock_right_N161 );
not U_inv601 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__1_ ( clk, n556_r, my_IIR_filter_firBlock_right_Y_in[1], my_IIR_filter_firBlock_right_N162 );
not U_inv602 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__2_ ( clk, n556_r, my_IIR_filter_firBlock_right_Y_in[2], my_IIR_filter_firBlock_right_N163 );
not U_inv603 ( n556_r, n556 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__3_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[3], my_IIR_filter_firBlock_right_N164 );
not U_inv604 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__4_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[4], my_IIR_filter_firBlock_right_N165 );
not U_inv605 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__5_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[5], my_IIR_filter_firBlock_right_N166 );
not U_inv606 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__6_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[6], my_IIR_filter_firBlock_right_N167 );
not U_inv607 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__7_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[7], my_IIR_filter_firBlock_right_N168 );
not U_inv608 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__8_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[8], my_IIR_filter_firBlock_right_N169 );
not U_inv609 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__9_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[9], my_IIR_filter_firBlock_right_N170 );
not U_inv610 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__10_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[10], my_IIR_filter_firBlock_right_N171 );
not U_inv611 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__11_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[11], my_IIR_filter_firBlock_right_N172 );
not U_inv612 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__12_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[12], my_IIR_filter_firBlock_right_N173 );
not U_inv613 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__13_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[13], my_IIR_filter_firBlock_right_N174 );
not U_inv614 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__14_ ( clk, n555_r, my_IIR_filter_firBlock_right_Y_in[14], my_IIR_filter_firBlock_right_N175 );
not U_inv615 ( n555_r, n555 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__15_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[15], my_IIR_filter_firBlock_right_N176 );
not U_inv616 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__16_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[16], my_IIR_filter_firBlock_right_N177 );
not U_inv617 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__17_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[17], my_IIR_filter_firBlock_right_N178 );
not U_inv618 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__18_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[18], my_IIR_filter_firBlock_right_N179 );
not U_inv619 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__19_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[19], my_IIR_filter_firBlock_right_N180 );
not U_inv620 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__20_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[20], my_IIR_filter_firBlock_right_N181 );
not U_inv621 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__21_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[21], my_IIR_filter_firBlock_right_N182 );
not U_inv622 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__22_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[22], my_IIR_filter_firBlock_right_N183 );
not U_inv623 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__23_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[23], my_IIR_filter_firBlock_right_N184 );
not U_inv624 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__24_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[24], my_IIR_filter_firBlock_right_N185 );
not U_inv625 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__25_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[25], my_IIR_filter_firBlock_right_N186 );
not U_inv626 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__26_ ( clk, n554_r, my_IIR_filter_firBlock_right_Y_in[26], my_IIR_filter_firBlock_right_N187 );
not U_inv627 ( n554_r, n554 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__27_ ( clk, n553_r, my_IIR_filter_firBlock_right_Y_in[27], my_IIR_filter_firBlock_right_N188 );
not U_inv628 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__28_ ( clk, n553_r, my_IIR_filter_firBlock_right_Y_in[28], my_IIR_filter_firBlock_right_N189 );
not U_inv629 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__29_ ( clk, n553_r, my_IIR_filter_firBlock_right_Y_in[29], my_IIR_filter_firBlock_right_N190 );
not U_inv630 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__30_ ( clk, n553_r, my_IIR_filter_firBlock_right_Y_in[30], my_IIR_filter_firBlock_right_N191 );
not U_inv631 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_firStep_reg_6__31_ ( clk, n553_r, my_IIR_filter_firBlock_right_Y_in[31], my_IIR_filter_firBlock_right_N192 );
not U_inv632 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_0_ ( clk, n553_r, rightOut[0], my_IIR_filter_firBlock_right_Y_in[0] );
not U_inv633 ( n207, rightOut[0] );
not U_inv634 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_1_ ( clk, n553_r, rightOut[1], my_IIR_filter_firBlock_right_Y_in[1] );
not U_inv635 ( n126, rightOut[1] );
not U_inv636 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_2_ ( clk, n553_r, n121, my_IIR_filter_firBlock_right_Y_in[2] );
not U_inv637 ( n538, n121 );
not U_inv638 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_3_ ( clk, n553_r, rightOut[3], my_IIR_filter_firBlock_right_Y_in[3] );
not U_inv639 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_4_ ( clk, n553_r, ex_wire2, my_IIR_filter_firBlock_right_Y_in[4] );
not U_inv640 ( n539, ex_wire2 );
not U_inv641 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_5_ ( clk, n553_r, rightOut[5], my_IIR_filter_firBlock_right_Y_in[5] );
not U_inv642 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_6_ ( clk, n553_r, rightOut[6], my_IIR_filter_firBlock_right_Y_in[6] );
not U_inv643 ( n553_r, n553 );
dff my_IIR_filter_firBlock_right_Y_reg_7_ ( clk, n552_r, rightOut[7], my_IIR_filter_firBlock_right_Y_in[7] );
not U_inv644 ( n113, rightOut[7] );
not U_inv645 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_8_ ( clk, n552_r, rightOut[8], my_IIR_filter_firBlock_right_Y_in[8] );
not U_inv646 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_9_ ( clk, n552_r, rightOut[9], my_IIR_filter_firBlock_right_Y_in[9] );
not U_inv647 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_10_ ( clk, n552_r, rightOut[10], my_IIR_filter_firBlock_right_Y_in[10] );
not U_inv648 ( n129, rightOut[10] );
not U_inv649 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_11_ ( clk, n552_r, rightOut[11], my_IIR_filter_firBlock_right_Y_in[11] );
not U_inv650 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_12_ ( clk, n552_r, rightOut[12], my_IIR_filter_firBlock_right_Y_in[12] );
not U_inv651 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_13_ ( clk, n552_r, rightOut[13], my_IIR_filter_firBlock_right_Y_in[13] );
not U_inv652 ( n541, rightOut[13] );
not U_inv653 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_14_ ( clk, n552_r, rightOut[14], my_IIR_filter_firBlock_right_Y_in[14] );
not U_inv654 ( n104, rightOut[14] );
not U_inv655 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_15_ ( clk, n552_r, rightOut[15], my_IIR_filter_firBlock_right_Y_in[15] );
not U_inv656 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_16_ ( clk, n552_r, rightOut[16], my_IIR_filter_firBlock_right_Y_in[16] );
not U_inv657 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_17_ ( clk, n552_r, rightOut[17], my_IIR_filter_firBlock_right_Y_in[17] );
not U_inv658 ( n106, rightOut[17] );
not U_inv659 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_18_ ( clk, n552_r, rightOut[18], my_IIR_filter_firBlock_right_Y_in[18] );
not U_inv660 ( n552_r, n552 );
dff my_IIR_filter_firBlock_right_Y_reg_19_ ( clk, n551_r, rightOut[19], my_IIR_filter_firBlock_right_Y_in[19] );
not U_inv661 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_20_ ( clk, n551_r, rightOut[20], my_IIR_filter_firBlock_right_Y_in[20] );
not U_inv662 ( n108, rightOut[20] );
not U_inv663 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_21_ ( clk, n551_r, rightOut[21], my_IIR_filter_firBlock_right_Y_in[21] );
not U_inv664 ( n110, rightOut[21] );
not U_inv665 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_22_ ( clk, n551_r, rightOut[22], my_IIR_filter_firBlock_right_Y_in[22] );
not U_inv666 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_23_ ( clk, n551_r, rightOut[23], my_IIR_filter_firBlock_right_Y_in[23] );
not U_inv667 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_24_ ( clk, n551_r, rightOut[24], my_IIR_filter_firBlock_right_Y_in[24] );
not U_inv668 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_25_ ( clk, n551_r, rightOut[25], my_IIR_filter_firBlock_right_Y_in[25] );
not U_inv669 ( n543, rightOut[25] );
not U_inv670 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_26_ ( clk, n551_r, rightOut[26], my_IIR_filter_firBlock_right_Y_in[26] );
not U_inv671 ( n545, rightOut[26] );
not U_inv672 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_27_ ( clk, n551_r, rightOut[27], my_IIR_filter_firBlock_right_Y_in[27] );
not U_inv673 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_28_ ( clk, n551_r, rightOut[28], my_IIR_filter_firBlock_right_Y_in[28] );
not U_inv674 ( n530, rightOut[28] );
not U_inv675 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_29_ ( clk, n551_r, rightOut[29], my_IIR_filter_firBlock_right_Y_in[29] );
not U_inv676 ( n551_r, n551 );
dff my_IIR_filter_firBlock_right_Y_reg_30_ ( clk, n551_r, ex_wire3, my_IIR_filter_firBlock_right_Y_in[30] );
not U_inv677 ( n58, ex_wire3 );
not U_inv678 ( n551_r, n551 );
dff my_IIR_filter_firBlock_left_firStep_reg_8__31_ ( clk, n580_r, my_IIR_filter_firBlock_left_firStep[31], my_IIR_filter_firBlock_left_N256 );
not U_inv679 ( n580_r, n580 );
dff inData_in_reg_30_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[114], inData_30 );
not U_inv680 ( n61, my_IIR_filter_firBlock_left_multProducts[114] );
not U_inv681 ( n606_r, n606 );
dff inData_in_reg_29_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[113], inData_29 );
not U_inv682 ( n60, my_IIR_filter_firBlock_left_multProducts[113] );
not U_inv683 ( n606_r, n606 );
dff inData_in_reg_28_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[112], inData_28 );
not U_inv684 ( n59, my_IIR_filter_firBlock_left_multProducts[112] );
not U_inv685 ( n606_r, n606 );
dff inData_in_reg_27_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[111], inData_27 );
not U_inv686 ( n57, my_IIR_filter_firBlock_left_multProducts[111] );
not U_inv687 ( n606_r, n606 );
dff inData_in_reg_26_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[110], inData_26 );
not U_inv688 ( n56, my_IIR_filter_firBlock_left_multProducts[110] );
not U_inv689 ( n606_r, n606 );
dff inData_in_reg_25_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[109], inData_25 );
not U_inv690 ( n55, my_IIR_filter_firBlock_left_multProducts[109] );
not U_inv691 ( n606_r, n606 );
dff inData_in_reg_24_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[108], inData_24 );
not U_inv692 ( n54, my_IIR_filter_firBlock_left_multProducts[108] );
not U_inv693 ( n606_r, n606 );
dff inData_in_reg_23_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[107], inData_23 );
not U_inv694 ( n308, my_IIR_filter_firBlock_left_multProducts[107] );
not U_inv695 ( n606_r, n606 );
dff inData_in_reg_22_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[106], inData_22 );
not U_inv696 ( n53, my_IIR_filter_firBlock_left_multProducts[106] );
not U_inv697 ( n606_r, n606 );
dff inData_in_reg_21_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[105], inData_21 );
not U_inv698 ( n52, my_IIR_filter_firBlock_left_multProducts[105] );
not U_inv699 ( n606_r, n606 );
dff inData_in_reg_20_ ( clk, n606_r, my_IIR_filter_firBlock_left_multProducts[104], inData_20 );
not U_inv700 ( n51, my_IIR_filter_firBlock_left_multProducts[104] );
not U_inv701 ( n606_r, n606 );
dff inData_in_reg_19_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[103], inData_19 );
not U_inv702 ( n304, my_IIR_filter_firBlock_left_multProducts[103] );
not U_inv703 ( n605_r, n605 );
dff inData_in_reg_18_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[102], inData_18 );
not U_inv704 ( n296, my_IIR_filter_firBlock_left_multProducts[102] );
not U_inv705 ( n605_r, n605 );
dff inData_in_reg_17_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[101], inData_17 );
not U_inv706 ( n300, my_IIR_filter_firBlock_left_multProducts[101] );
not U_inv707 ( n605_r, n605 );
dff inData_in_reg_16_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[100], inData_16 );
not U_inv708 ( n298, my_IIR_filter_firBlock_left_multProducts[100] );
not U_inv709 ( n605_r, n605 );
dff inData_in_reg_15_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[99], inData_15 );
not U_inv710 ( n302, my_IIR_filter_firBlock_left_multProducts[99] );
not U_inv711 ( n605_r, n605 );
dff inData_in_reg_14_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[98], inData_14 );
not U_inv712 ( n294, my_IIR_filter_firBlock_left_multProducts[98] );
not U_inv713 ( n605_r, n605 );
dff inData_in_reg_13_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[97], inData_13 );
not U_inv714 ( n306, my_IIR_filter_firBlock_left_multProducts[97] );
not U_inv715 ( n605_r, n605 );
dff inData_in_reg_12_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[96], inData_12 );
not U_inv716 ( n50, my_IIR_filter_firBlock_left_multProducts[96] );
not U_inv717 ( n605_r, n605 );
dff inData_in_reg_11_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[95], inData_11 );
not U_inv718 ( n49, my_IIR_filter_firBlock_left_multProducts[95] );
not U_inv719 ( n605_r, n605 );
dff inData_in_reg_1_ ( clk, n604_r, inData_in[1], inData_1 );
not U_inv720 ( n40, inData_in[1] );
not U_inv721 ( n604_r, n604 );
dff inData_in_reg_10_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[94], inData_10 );
not U_inv722 ( n48, my_IIR_filter_firBlock_left_multProducts[94] );
not U_inv723 ( n605_r, n605 );
dff inData_in_reg_9_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[93], inData_9 );
not U_inv724 ( n343, my_IIR_filter_firBlock_left_multProducts[93] );
not U_inv725 ( n605_r, n605 );
dff inData_in_reg_8_ ( clk, n605_r, my_IIR_filter_firBlock_left_multProducts[92], inData_8 );
not U_inv726 ( n341, my_IIR_filter_firBlock_left_multProducts[92] );
not U_inv727 ( n605_r, n605 );
dff inData_in_reg_7_ ( clk, n604_r, my_IIR_filter_firBlock_left_multProducts[91], inData_7 );
not U_inv728 ( n47, my_IIR_filter_firBlock_left_multProducts[91] );
not U_inv729 ( n604_r, n604 );
dff inData_in_reg_6_ ( clk, n604_r, my_IIR_filter_firBlock_left_multProducts[90], inData_6 );
not U_inv730 ( n46, my_IIR_filter_firBlock_left_multProducts[90] );
not U_inv731 ( n604_r, n604 );
dff inData_in_reg_5_ ( clk, n604_r, inData_in[5], inData_5 );
not U_inv732 ( n45, inData_in[5] );
not U_inv733 ( n604_r, n604 );
dff inData_in_reg_4_ ( clk, n604_r, inData_in[4], inData_4 );
not U_inv734 ( n44, inData_in[4] );
not U_inv735 ( n604_r, n604 );
and U34 ( n3090, n3089, n3088 );
nand U35 ( n874, my_IIR_filter_firBlock_left_multProducts[102], n872 );
not U36 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[33], n128 );
not U37 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[13], n115 );
nand U38 ( n1272, n1271, n1270 );
nand U39 ( n1271, my_IIR_filter_firBlock_left_multProducts[98], n1269 );
nand U40 ( n1265, n1264, n1263 );
nand U41 ( n1264, my_IIR_filter_firBlock_left_multProducts[96], n1262 );
nand U42 ( n1258, n1257, n1256 );
nand U43 ( n1257, my_IIR_filter_firBlock_left_multProducts[94], n1255 );
or U44 ( n2944, n123, n520 );
xor U45 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[29], n3011, n3010 );
xnor U46 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[22], n2981, n120 );
nand U47 ( n766, leftOut[20], n764 );
nand U48 ( n872, n870, n869 );
nand U49 ( n870, my_IIR_filter_firBlock_left_multProducts[101], n868 );
nand U50 ( n832, n830, n48 );
nand U51 ( n823, inData_in[4], n940 );
not U52 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[17], n125 );
xnor U53 ( n128, n3184, n3183 );
not U54 ( n648, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[31] );
not U55 ( n643, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[25] );
not U56 ( n640, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[22] );
xor U57 ( n115, n3090, n116 );
buf U58 ( n518, outData_in[4] );
nand U59 ( n1293, n1291, n1290 );
nand U60 ( n1291, my_IIR_filter_firBlock_left_multProducts[103], n1289 );
nand U61 ( n1276, n1274, n1273 );
nand U62 ( n1274, my_IIR_filter_firBlock_left_multProducts[99], n1272 );
nand U63 ( n1269, n1267, n1266 );
nand U64 ( n1267, my_IIR_filter_firBlock_left_multProducts[97], n1265 );
nand U65 ( n1262, n1260, n1259 );
nand U66 ( n1260, my_IIR_filter_firBlock_left_multProducts[95], n1258 );
nand U67 ( n1255, n1253, n1252 );
nand U68 ( n1253, my_IIR_filter_firBlock_left_multProducts[93], n1251 );
xor U69 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[15], n946, n945 );
and U70 ( n3477, my_IIR_filter_firBlock_right_multProducts[0], my_IIR_filter_firBlock_right_firStep[0] );
not U71 ( n700, outData_in[9] );
nand U72 ( n795, leftOut[29], n793 );
xnor U73 ( n133, n134, n804 );
nand U74 ( n2614, n2482, n2481 );
nand U75 ( n2482, my_IIR_filter_firBlock_left_firStep[3], n2612 );
nand U76 ( n2612, n2480, n2479 );
nand U77 ( n2480, my_IIR_filter_firBlock_left_firStep[2], n2600 );
or U78 ( n1908, n1907, my_IIR_filter_firBlock_left_firStep[189] );
xor U79 ( my_IIR_filter_firBlock_left_multProducts[59], n1339, n1338 );
nand U80 ( my_IIR_filter_firBlock_left_multProducts[88], n1075, n1074 );
not U81 ( n209, n697 );
buf U82 ( n499, outData_in[13] );
buf U83 ( n498, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[1] );
not U84 ( outData_in[5], n133 );
buf U85 ( n547, n548 );
buf U86 ( n509, outData_in[10] );
xor U87 ( n3057, n502, n133 );
xnor U88 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[15], n3099, n62 );
xor U89 ( n62, n672, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[21] );
or U90 ( n3038, n497, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[2] );
or U91 ( n3606, n63, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[8] );
nor U92 ( n63, n3745, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[8] );
or U93 ( n3613, n64, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[10] );
nor U94 ( n64, n3612, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[10] );
xnor U95 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[24], n2989, n65 );
xnor U96 ( n65, n685, outData_in[18] );
xor U97 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[8], n3038, n172 );
xor U98 ( n66, n67, n807 );
not U99 ( outData_in[7], n66 );
xnor U100 ( n67, leftOut[7], rightOut[7] );
not U101 ( n68, n2958 );
nand U102 ( n2960, n2957, n69 );
nor U103 ( n69, n680, n68 );
nand U104 ( n70, n3338, my_IIR_filter_firBlock_right_multProducts[60] );
and U105 ( n3341, n70, n71 );
and U106 ( n71, n72, n3340 );
nand U107 ( n73, n2949, n701 );
nand U108 ( n2952, n73, n74 );
and U109 ( n74, n702, n2951 );
nand U110 ( n2946, n2944, n75 );
and U111 ( n75, n2945, n133 );
nand U112 ( n76, n3319, my_IIR_filter_firBlock_right_multProducts[56] );
nand U113 ( n3324, n76, n77 );
and U114 ( n77, n78, n3321 );
nand U115 ( n79, n3292, my_IIR_filter_firBlock_right_multProducts[50] );
nand U116 ( n3297, n79, n80 );
and U117 ( n80, n81, n3294 );
nand U118 ( n82, n3263, my_IIR_filter_firBlock_right_multProducts[44] );
nand U119 ( n3268, n82, n83 );
and U120 ( n83, n84, n3265 );
nand U121 ( n85, n3245, my_IIR_filter_firBlock_right_multProducts[40] );
nand U122 ( n3250, n85, n86 );
and U123 ( n86, n87, n3247 );
nand U124 ( n88, n3236, my_IIR_filter_firBlock_right_multProducts[37] );
nand U125 ( n3239, n88, n89 );
and U126 ( n89, n90, n3238 );
buf U127 ( n519, outData_in[9] );
or U128 ( n3115, n91, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[24] );
nor U129 ( n91, n3114, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[18] );
or U130 ( n3134, n92, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[28] );
nor U131 ( n92, n3133, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[22] );
or U132 ( n3138, n93, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[29] );
nor U133 ( n93, n3137, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[23] );
or U134 ( n3162, n94, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[34] );
nor U135 ( n94, n3161, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[28] );
or U136 ( n3171, n95, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[36] );
nor U137 ( n95, n3170, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[30] );
or U138 ( n3017, n96, outData_in[24] );
nor U139 ( n96, n3016, n489 );
or U140 ( n3031, n97, n491 );
nor U141 ( n97, n3030, n504 );
or U142 ( n3639, n98, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[16] );
nor U143 ( n98, n3638, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[16] );
or U144 ( n3675, n99, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[24] );
nor U145 ( n99, n3674, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[24] );
or U146 ( n3713, n100, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[32] );
nor U147 ( n100, n3712, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[32] );
or U148 ( n3722, n101, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[34] );
nor U149 ( n101, n3721, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[34] );
and U150 ( n3099, n3098, n3097 );
xnor U151 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[14], n3062, n102 );
xnor U152 ( n102, n703, outData_in[8] );
xnor U153 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[15], n3063, n103 );
xnor U154 ( n103, n702, outData_in[9] );
xor U155 ( n3219, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[15], n167 );
or U156 ( n745, n104, n105 );
nor U157 ( n105, n744, leftOut[14] );
or U158 ( n754, n106, n107 );
nor U159 ( n107, n753, leftOut[17] );
or U160 ( n765, n108, n109 );
nor U161 ( n109, n764, leftOut[20] );
or U162 ( n768, n110, n111 );
nor U163 ( n111, n767, leftOut[21] );
xnor U164 ( n3043, outData_in[30], outData_in[28] );
or U165 ( n112, n132, n523 );
or U166 ( n3054, n132, n523 );
or U167 ( n722, n113, n114 );
nor U168 ( n114, n807, leftOut[7] );
xor U169 ( n116, n674, n160 );
xor U170 ( my_IIR_filter_firBlock_right_multProducts[36], n3624, n117 );
xor U171 ( n117, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[13], n115 );
or U172 ( n2939, n118, n516 );
nor U173 ( n118, n3056, n522 );
nand U174 ( n763, leftOut[19], n761 );
or U175 ( n2982, n119, outData_in[16] );
nor U176 ( n119, n2981, n485 );
xnor U177 ( n120, n683, outData_in[16] );
nand U178 ( n761, n758, n757 );
nand U179 ( n711, n121, n122 );
nand U180 ( n122, n152, n153 );
nor U181 ( n123, n3059, n517 );
xor U182 ( n160, n2967, n161 );
xnor U183 ( outData_in[3], n124, n801 );
xnor U184 ( n124, leftOut[3], rightOut[3] );
xnor U185 ( n125, n3109, n3108 );
xor U186 ( n759, n126, n127 );
xor U187 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[31], n3020, n3019 );
xnor U188 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[25], n2993, n235 );
xnor U189 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[28], n3006, n237 );
xnor U190 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[35], n3039, n233 );
or U191 ( n730, n129, n130 );
nor U192 ( n130, n729, leftOut[10] );
xnor U193 ( my_IIR_filter_firBlock_right_multProducts[41], n3646, n131 );
xor U194 ( n131, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[18], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[18] );
and U195 ( n132, n677, n3038 );
xnor U196 ( n3611, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[10], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[10] );
xnor U197 ( outData_in[23], n193, n775 );
xor U198 ( n134, leftOut[5], rightOut[5] );
xnor U199 ( my_IIR_filter_firBlock_right_multProducts[35], n3620, n135 );
xnor U200 ( n135, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[12], n136 );
buf U201 ( n523, outData_in[2] );
xnor U202 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[16], n2955, n216 );
xor U203 ( n136, n3086, n218 );
xor U204 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[23], n3137, n3136 );
nand U205 ( n137, n2960, n519 );
nand U206 ( n2964, n137, n138 );
and U207 ( n138, n679, n2962 );
xnor U208 ( my_IIR_filter_firBlock_right_multProducts[61], n3743, n139 );
xnor U209 ( n139, n525, n3212 );
xnor U210 ( n140, n3166, n3164 );
nand U211 ( n141, n792, leftOut[2] );
nand U212 ( n713, n141, n142 );
and U213 ( n142, n143, n711 );
nand U214 ( n144, n184, rightOut[8] );
nand U215 ( n189, n144, n145 );
and U216 ( n145, n146, n725 );
xnor U217 ( n147, n3082, n3081 );
and U218 ( n3082, n3080, n3079 );
nand U219 ( n188, n731, n148 );
and U220 ( n148, n730, n149 );
nand U221 ( n150, n713, rightOut[3] );
and U222 ( n540, n150, n151 );
and U223 ( n151, n279, n715 );
buf U224 ( n157, outData_in[24] );
nand U225 ( n152, n708, rightOut[1] );
and U226 ( n153, n710, n263 );
not U227 ( n154, n690 );
xor U228 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[18], n2963, n164 );
buf U229 ( n158, outData_in[26] );
nand U230 ( n718, n716, n155 );
and U231 ( n155, n717, n156 );
xnor U232 ( outData_in[24], n778, n264 );
xnor U233 ( outData_in[26], n784, n267 );
xor U234 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[7], n3217, n159 );
xnor U235 ( n159, n674, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[7] );
xor U236 ( n161, n682, n488 );
xor U237 ( my_IIR_filter_firBlock_right_multProducts[44], n3660, n162 );
xor U238 ( n162, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[21], n639 );
xnor U239 ( n163, n2959, n219 );
xor U240 ( n164, n681, n509 );
xor U241 ( my_IIR_filter_firBlock_right_multProducts[52], n3697, n165 );
xnor U242 ( n165, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[29], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[29] );
xor U243 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[6], n3216, n166 );
xnor U244 ( n166, n675, n498 );
xnor U245 ( n167, n112, n224 );
xnor U246 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[10], n168, n2935 );
xnor U247 ( n168, outData_in[7], n519 );
xor U248 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[13], n2837, n169 );
xor U249 ( n169, n511, n509 );
xor U250 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[32], n3025, n3024 );
xor U251 ( n3029, n694, outData_in[27] );
xor U252 ( n3019, n692, outData_in[25] );
buf U253 ( n494, outData_in[19] );
xnor U254 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[26], n2997, n236 );
xor U255 ( n2971, n681, outData_in[14] );
buf U256 ( n496, outData_in[15] );
xor U257 ( n2976, n682, outData_in[15] );
xor U258 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[12], n3059, n170 );
xor U259 ( n170, n704, outData_in[6] );
xor U260 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[33], n2922, n171 );
xor U261 ( n171, n525, outData_in[30] );
xor U262 ( n172, outData_in[2], n498 );
xor U263 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[29], n2904, n173 );
xor U264 ( n173, outData_in[28], n158 );
xor U265 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[23], n2878, n174 );
xor U266 ( n174, n490, outData_in[20] );
xor U267 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[21], n2870, n175 );
xor U268 ( n175, outData_in[20], outData_in[18] );
xor U269 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[17], n2853, n176 );
xor U270 ( n176, outData_in[16], n486 );
nand U271 ( my_IIR_filter_firBlock_left_multProducts[89], n1078, n1077 );
and U272 ( n246, n177, n178 );
nand U273 ( n177, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[38], n1785 );
nand U274 ( n178, n1786, n527 );
nand U275 ( n762, n179, rightOut[19] );
or U276 ( n179, n761, leftOut[19] );
xnor U277 ( n251, my_IIR_filter_firBlock_right_multProducts[61], n180 );
nand U278 ( n748, rightOut[15], n181 );
or U279 ( n181, n747, leftOut[15] );
nand U280 ( n776, rightOut[23], n182 );
or U281 ( n182, n775, leftOut[23] );
nand U282 ( n788, rightOut[27], n183 );
or U283 ( n183, n787, leftOut[27] );
nand U284 ( n724, rightOut[8], n184 );
or U285 ( n184, n809, leftOut[8] );
nand U286 ( n737, n185, rightOut[12] );
or U287 ( n185, n736, leftOut[12] );
nand U288 ( n751, rightOut[16], n186 );
or U289 ( n186, n750, leftOut[16] );
nand U290 ( n779, rightOut[24], n187 );
or U291 ( n187, n778, leftOut[24] );
nand U292 ( n734, rightOut[11], n188 );
nand U293 ( n726, rightOut[9], n189 );
nand U294 ( n757, rightOut[18], n190 );
or U295 ( n190, n756, leftOut[18] );
nand U296 ( n794, rightOut[29], n191 );
or U297 ( n191, n793, leftOut[29] );
xnor U298 ( outData_in[21], n192, n767 );
xnor U299 ( n192, leftOut[21], rightOut[21] );
xnor U300 ( n193, leftOut[23], rightOut[23] );
xor U301 ( outData_in[12], n736, n194 );
xor U302 ( n194, rightOut[12], leftOut[12] );
xnor U303 ( n248, my_IIR_filter_firBlock_right_multProducts[30], n195 );
nand U304 ( n822, n196, n46 );
or U305 ( n196, n940, inData_in[4] );
nand U306 ( n869, n197, n304 );
or U307 ( n197, n868, my_IIR_filter_firBlock_left_multProducts[101] );
or U308 ( n868, n257, n258 );
nand U309 ( n830, n198, n199 );
nand U310 ( n198, my_IIR_filter_firBlock_left_multProducts[91], n946 );
nand U311 ( n199, n828, n343 );
nand U312 ( n1041, n200, n201 );
nand U313 ( n200, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[31], n1038 );
nand U314 ( n201, my_IIR_filter_firBlock_left_multProducts[106], n1039 );
nand U315 ( n1067, n202, n203 );
nand U316 ( n202, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[37], n1065 );
nand U317 ( n203, my_IIR_filter_firBlock_left_multProducts[112], n1066 );
nand U318 ( n873, n204, n51 );
or U319 ( n204, n872, my_IIR_filter_firBlock_left_multProducts[102] );
xnor U320 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[32], n900, n252 );
and U321 ( n2739, my_IIR_filter_firBlock_right_multProducts[62], my_IIR_filter_firBlock_right_firStep[62] );
or U322 ( n1634, n1633, n1632 );
nand U323 ( n1911, n205, n206 );
nand U324 ( n205, my_IIR_filter_firBlock_left_firStep[189], n1907 );
nand U325 ( n206, my_IIR_filter_firBlock_left_multProducts[29], n1908 );
buf U326 ( n626, reset );
buf U327 ( n627, reset );
buf U328 ( n628, reset );
nor U329 ( n760, n207, n208 );
xnor U330 ( outData_in[28], n790, n266 );
xor U331 ( n210, n3739, n211 );
xnor U332 ( n211, n654, n525 );
buf U333 ( n524, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10_39 );
xor U334 ( my_IIR_filter_firBlock_right_multProducts[3], n3362, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[10] );
nand U335 ( n3362, n3363, n655 );
buf U336 ( n525, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10_39 );
nand U337 ( n3366, n3364, n3363 );
nand U338 ( n3405, n3404, n653 );
xnor U339 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[38], n3208, n212 );
xor U340 ( n212, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[38], n524 );
not U341 ( n652, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[36] );
xor U342 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[10], n3077, n3076 );
not U343 ( n646, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[28] );
nand U344 ( n3660, n3659, n3658 );
nand U345 ( n3658, n3657, n638 );
nand U346 ( n3651, n3649, n3648 );
nand U347 ( n3648, n3647, n636 );
nand U348 ( n3629, n3627, n3626 );
nand U349 ( n3624, n3623, n3622 );
nand U350 ( n3622, n3621, n136 );
nand U351 ( n3633, n3632, n3631 );
nand U352 ( n3631, n3630, n633 );
not U353 ( n653, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[37] );
not U354 ( n644, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[26] );
not U355 ( n650, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[34] );
nand U356 ( n3620, n3619, n3618 );
xor U357 ( n3628, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[14], n633 );
not U358 ( n633, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[14] );
nand U359 ( n3612, n3610, n3609 );
nand U360 ( n3609, n3608, n655 );
nand U361 ( n3212, n3211, n3210 );
xnor U362 ( my_IIR_filter_firBlock_right_multProducts[32], n3746, n213 );
xnor U363 ( n213, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[9], n655 );
not U364 ( n637, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[19] );
xor U365 ( n3655, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[20], n638 );
nand U366 ( n3598, n3597, n3596 );
nand U367 ( n3745, n3605, n3604 );
nand U368 ( n3590, n3589, n3588 );
nand U369 ( n3589, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[3], n3586 );
nor U370 ( n3587, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[3], n3586 );
nand U371 ( n3594, n3593, n3592 );
or U372 ( n3592, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[4], n3591 );
xnor U373 ( my_IIR_filter_firBlock_right_multProducts[1], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[8], n3407 );
xnor U374 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[4], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[10], n3214 );
nand U375 ( n3079, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[10], n3078 );
nand U376 ( n3217, n3066, n675 );
nand U377 ( n3066, n677, n3216 );
nand U378 ( n3218, n3069, n3068 );
or U379 ( n3069, n678, n3217 );
nand U380 ( n3068, n3067, n674 );
nand U381 ( n3067, n3217, n678 );
nand U382 ( n3216, n3215, n676 );
nand U383 ( n3077, n3075, n3074 );
nand U384 ( n3074, n3073, n672 );
nor U385 ( n3363, n3361, n3406 );
xnor U386 ( my_IIR_filter_firBlock_right_multProducts[38], n3633, n214 );
xnor U387 ( n214, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[15], n634 );
not U388 ( n656, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[1] );
nor U389 ( n3215, n3065, n3213 );
xor U390 ( my_IIR_filter_firBlock_right_multProducts[12], n3378, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[19] );
nor U391 ( n3369, n3367, n3366 );
xor U392 ( my_IIR_filter_firBlock_right_multProducts[7], n3368, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[14] );
nand U393 ( n3368, n3369, n115 );
xnor U394 ( my_IIR_filter_firBlock_right_multProducts[10], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[17], n3375 );
nor U395 ( n3375, n3373, n3372 );
xor U396 ( my_IIR_filter_firBlock_right_multProducts[19], n3386, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[26] );
nand U397 ( n3386, n3387, n643 );
nor U398 ( n3377, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[19], n3378 );
nand U399 ( n3374, n3375, n125 );
nor U400 ( n3381, n3379, n3378 );
nor U401 ( n3387, n3385, n3384 );
xnor U402 ( my_IIR_filter_firBlock_right_multProducts[21], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[28], n3389 );
nor U403 ( n3383, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[23], n3384 );
nand U404 ( n3380, n3381, n639 );
nand U405 ( n3378, n3376, n3375 );
nand U406 ( n3372, n3370, n3369 );
nand U407 ( n3392, n3393, n140 );
nand U408 ( n3390, n3388, n3387 );
nor U409 ( n3393, n3391, n3390 );
nand U410 ( n3384, n3382, n3381 );
nand U411 ( n3396, n3394, n3393 );
nor U412 ( n3404, n3403, n3402 );
xor U413 ( n215, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[37], n3404 );
nor U414 ( n3399, n3397, n3396 );
xor U415 ( my_IIR_filter_firBlock_right_multProducts[27], n3398, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[34] );
xnor U416 ( my_IIR_filter_firBlock_right_multProducts[29], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[36], n3401 );
nand U417 ( n3402, n3400, n3399 );
not U418 ( n632, my_IIR_filter_firBlock_right_multProducts[91] );
xor U419 ( my_IIR_filter_firBlock_right_multProducts[108], n3571, n529 );
nand U420 ( n3406, n3360, n3359 );
nor U421 ( n3360, n498, n3356 );
and U422 ( n3359, n3358, n3357 );
nand U423 ( n3159, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[27], n3156 );
nand U424 ( n3154, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[26], n3151 );
not U425 ( n665, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[30] );
not U426 ( n660, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[22] );
not U427 ( n663, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[26] );
nand U428 ( n3139, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[23], n3137 );
not U429 ( n662, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[25] );
not U430 ( n671, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[38] );
not U431 ( n670, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[37] );
nand U432 ( n3172, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[30], n3170 );
not U433 ( n661, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[23] );
nand U434 ( n3104, n3102, n3101 );
nand U435 ( n3095, n3093, n3092 );
not U436 ( n666, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[31] );
nand U437 ( n3056, n2938, n2937 );
or U438 ( n2938, n707, n112 );
nand U439 ( n2936, n3054, n707 );
nand U440 ( n2955, n2954, n2953 );
nand U441 ( n2953, n2952, n700 );
nand U442 ( n3059, n2943, n2942 );
nand U443 ( n2967, n2966, n2965 );
nand U444 ( n2965, n2964, n681 );
nand U445 ( n3061, n2944, n2945 );
nand U446 ( n2969, n2968, n682 );
nand U447 ( n3058, n2939, n2940 );
nand U448 ( n2977, n2975, n2974 );
nand U449 ( n2974, n2973, n683 );
nand U450 ( n3020, n3018, n3017 );
xor U451 ( n3673, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[24], n642 );
xor U452 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[36], n3199, n3198 );
xnor U453 ( n216, n701, n508 );
xor U454 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[28], n3161, n3160 );
xnor U455 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[30], n3170, n217 );
xor U456 ( n217, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[30], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[36] );
nand U457 ( n3664, n3663, n3662 );
nand U458 ( n3646, n3645, n3644 );
xnor U459 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[12], n3086, n218 );
xor U460 ( n218, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[12], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[18] );
xor U461 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[26], n3151, n3150 );
xor U462 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[34], n3189, n3188 );
xnor U463 ( n219, n700, outData_in[11] );
xor U464 ( n3677, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[25], n643 );
xor U465 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[25], n3146, n3145 );
xnor U466 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[8], n3218, n220 );
xor U467 ( n220, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[8], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[14] );
nand U468 ( n3746, n3607, n3606 );
xor U469 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[27], n3156, n3155 );
not U470 ( n672, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[15] );
xor U471 ( n3650, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[19], n637 );
xor U472 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[19], n3118, n3117 );
nand U473 ( n2833, n2832, n2831 );
nand U474 ( n2849, n2848, n2847 );
nand U475 ( n2848, n511, n2845 );
or U476 ( n2846, n2845, n511 );
nand U477 ( n2932, n2819, n2818 );
nand U478 ( n2935, n2825, n2824 );
nand U479 ( n2841, n2840, n2839 );
nand U480 ( n2839, n511, n2838 );
nand U481 ( n2861, n2860, n2859 );
nand U482 ( n2859, n513, n2858 );
nand U483 ( n2853, n2852, n2851 );
nand U484 ( n2851, n495, n2850 );
nand U485 ( n2837, n2836, n2835 );
nand U486 ( n2870, n2869, n2868 );
nand U487 ( n2869, n512, n2866 );
or U488 ( n2867, n2866, n513 );
nand U489 ( n2829, n2828, n2827 );
nand U490 ( n2928, n2810, n2809 );
nand U491 ( n2913, n2912, n2911 );
nand U492 ( n2911, n515, n2910 );
nand U493 ( n2895, n2894, n2893 );
nand U494 ( n2894, n529, n2891 );
or U495 ( n2892, n2891, n529 );
nand U496 ( n2922, n2921, n2920 );
nand U497 ( n2921, n514, n2918 );
nand U498 ( n2920, n524, n2919 );
or U499 ( n2919, n2918, n515 );
nand U500 ( n2929, n2813, n2812 );
nand U501 ( n2812, n518, n2811 );
nand U502 ( n2845, n2844, n2843 );
nand U503 ( n2904, n2903, n2902 );
xnor U504 ( n3052, n699, n547 );
xor U505 ( n3641, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[17], n125 );
nand U506 ( n3586, n221, n222 );
or U507 ( n221, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[2], n3585 );
nand U508 ( n222, n656, n501 );
nand U509 ( n3602, n3601, n3600 );
nand U510 ( n3601, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[6], n3598 );
nor U511 ( n3599, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[6], n3598 );
xnor U512 ( n3132, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[22], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[28] );
xnor U513 ( my_IIR_filter_firBlock_right_multProducts[45], n3664, n223 );
xnor U514 ( n223, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[22], n640 );
xnor U515 ( n224, n503, n501 );
xnor U516 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[32], n2917, n2918 );
xor U517 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[10], n3056, n3055 );
nand U518 ( n3086, n3085, n3084 );
nand U519 ( n3220, n3072, n3071 );
nand U520 ( n3071, n3070, n673 );
not U521 ( n676, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[11] );
xor U522 ( n3744, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[8], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[8] );
xnor U523 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[5], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[11], n3215 );
xnor U524 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[1], n678, n498 );
not U525 ( n677, n497 );
nand U526 ( n3213, n3064, n677 );
xnor U527 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[30], n2908, n2909 );
not U528 ( n684, n496 );
nor U529 ( n2668, n498, n2625 );
not U530 ( n698, n515 );
xor U531 ( my_IIR_filter_firBlock_right_multProducts[63], n2669, n518 );
xnor U532 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[28], n2899, n2900 );
xnor U533 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[26], n2890, n2891 );
nand U534 ( n2628, n2626, n2668 );
not U535 ( n631, my_IIR_filter_firBlock_left_multProducts[89] );
xnor U536 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[4], n2926, n225 );
xnor U537 ( n225, n503, n501 );
nand U538 ( n1785, n1783, n1782 );
nand U539 ( n1782, n1781, n526 );
xor U540 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[5], n2928, n2927 );
xnor U541 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[20], n2865, n2866 );
xor U542 ( my_IIR_filter_firBlock_left_multProducts[29], n1780, n1779 );
xor U543 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[9], n2934, n2933 );
xor U544 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[18], n226, n2857 );
xor U545 ( n226, n495, n512 );
xor U546 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[7], n2931, n2930 );
xnor U547 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[11], n2829, n227 );
xnor U548 ( n227, n509, n507 );
xor U549 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[16], n228, n2849 );
xor U550 ( n228, n499, n496 );
xnor U551 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[15], n2845, n229 );
xnor U552 ( n229, n486, n511 );
xor U553 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[12], n230, n2833 );
xor U554 ( n230, n488, n519 );
nand U555 ( n2634, n2632, n2631 );
xor U556 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[14], n231, n2841 );
xor U557 ( n231, n487, n499 );
xor U558 ( my_IIR_filter_firBlock_right_multProducts[70], n680, n2637 );
nor U559 ( n2637, n2635, n2634 );
xor U560 ( my_IIR_filter_firBlock_right_multProducts[71], n2636, n510 );
nand U561 ( n2636, n2637, n680 );
nand U562 ( n2640, n2638, n2637 );
nand U563 ( my_IIR_filter_firBlock_right_multProducts[90], n632, n2667 );
nand U564 ( n2667, n524, n2666 );
xor U565 ( my_IIR_filter_firBlock_right_multProducts[76], n2646, n513 );
nor U566 ( n2643, n2641, n2640 );
xor U567 ( my_IIR_filter_firBlock_right_multProducts[80], n2652, n154 );
nor U568 ( n2651, n154, n2652 );
xor U569 ( my_IIR_filter_firBlock_right_multProducts[82], n692, n2655 );
nor U570 ( n2655, n2653, n2652 );
xor U571 ( my_IIR_filter_firBlock_right_multProducts[86], n696, n2661 );
xor U572 ( my_IIR_filter_firBlock_right_multProducts[88], n2664, n515 );
or U573 ( my_IIR_filter_firBlock_right_multProducts[116], my_IIR_filter_firBlock_right_multProducts[117], n232 );
and U574 ( n232, n524, n3582 );
xnor U575 ( my_IIR_filter_firBlock_right_multProducts[114], n515, n3580 );
nand U576 ( n3571, n3569, n3568 );
nand U577 ( n3567, n3568, n690 );
xnor U578 ( my_IIR_filter_firBlock_right_multProducts[106], n154, n3568 );
nand U579 ( n3559, n3557, n3556 );
nor U580 ( n3556, n3554, n3553 );
not U581 ( n549, n39 );
buf U582 ( n526, n550 );
nand U583 ( n3553, n3551, n3550 );
xnor U584 ( my_IIR_filter_firBlock_right_multProducts[102], n513, n3562 );
buf U585 ( n527, n550 );
nor U586 ( n3550, n3548, n3583 );
xor U587 ( my_IIR_filter_firBlock_right_multProducts[100], n3559, n496 );
nand U588 ( n3583, n3547, n3546 );
nor U589 ( n3547, n498, n3543 );
and U590 ( n3546, n3545, n3544 );
nand U591 ( n3555, n3556, n682 );
xnor U592 ( my_IIR_filter_firBlock_right_multProducts[97], n511, n3552 );
nand U593 ( n3549, n3550, n700 );
buf U594 ( n605, n607 );
buf U595 ( n606, n607 );
buf U596 ( n604, n607 );
buf U597 ( n580, n615 );
buf U598 ( n553, n624 );
buf U599 ( n554, n624 );
buf U600 ( n555, n624 );
buf U601 ( n556, n623 );
buf U602 ( n557, n623 );
buf U603 ( n558, n623 );
buf U604 ( n559, n622 );
buf U605 ( n560, n622 );
buf U606 ( n561, n622 );
buf U607 ( n562, n621 );
buf U608 ( n563, n621 );
buf U609 ( n564, n621 );
buf U610 ( n565, n620 );
buf U611 ( n566, n620 );
buf U612 ( n567, n620 );
buf U613 ( n568, n619 );
buf U614 ( n569, n619 );
buf U615 ( n570, n619 );
buf U616 ( n571, n618 );
buf U617 ( n572, n618 );
buf U618 ( n573, n618 );
buf U619 ( n574, n617 );
buf U620 ( n575, n617 );
buf U621 ( n576, n617 );
buf U622 ( n577, n616 );
buf U623 ( n578, n616 );
buf U624 ( n579, n616 );
buf U625 ( n581, n615 );
buf U626 ( n582, n615 );
buf U627 ( n583, n614 );
buf U628 ( n584, n614 );
buf U629 ( n585, n614 );
buf U630 ( n586, n613 );
buf U631 ( n587, n613 );
buf U632 ( n588, n613 );
buf U633 ( n589, n612 );
buf U634 ( n590, n612 );
buf U635 ( n591, n612 );
buf U636 ( n592, n611 );
buf U637 ( n593, n611 );
buf U638 ( n594, n611 );
buf U639 ( n595, n610 );
buf U640 ( n596, n610 );
buf U641 ( n597, n610 );
buf U642 ( n598, n609 );
buf U643 ( n599, n609 );
buf U644 ( n600, n609 );
buf U645 ( n601, n608 );
buf U646 ( n602, n608 );
buf U647 ( n603, n608 );
buf U648 ( n551, n625 );
buf U649 ( n552, n625 );
nand U650 ( n934, n812, n42 );
nand U651 ( n814, n813, n43 );
xor U652 ( n233, n492, outData_in[29] );
nand U653 ( n3011, n3009, n3008 );
nand U654 ( n3025, n3023, n3022 );
xnor U655 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[37], n3048, n234 );
xnor U656 ( n234, n698, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10_39 );
xor U657 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[34], n3034, n3033 );
nand U658 ( n1078, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, my_IIR_filter_firBlock_left_multProducts[88] );
nand U659 ( n1077, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n1076 );
or U660 ( n1076, my_IIR_filter_firBlock_left_multProducts[88], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
xnor U661 ( n235, n686, outData_in[19] );
nand U662 ( n2891, n2889, n2888 );
nand U663 ( n2866, n2864, n2863 );
nand U664 ( n2918, n2916, n2915 );
nand U665 ( n2882, n2881, n2880 );
nand U666 ( n2909, n2907, n2906 );
nand U667 ( n2874, n2873, n2872 );
nand U668 ( n2931, n2816, n2815 );
nand U669 ( n2934, n2822, n2821 );
buf U670 ( n522, outData_in[2] );
nand U671 ( n2878, n2877, n2876 );
nand U672 ( n2876, n154, n2875 );
nand U673 ( n2886, n2885, n2884 );
nand U674 ( n2885, n154, n2882 );
nand U675 ( n2884, outData_in[23], n2883 );
or U676 ( n2883, n2882, n154 );
nand U677 ( n2900, n2898, n2897 );
xnor U678 ( n3060, n133, n66 );
xnor U679 ( n236, n687, outData_in[20] );
xor U680 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[23], n2985, n2984 );
xor U681 ( n926, n60, n549 );
xnor U682 ( n237, n689, outData_in[22] );
buf U683 ( n503, outData_in[3] );
xor U684 ( my_IIR_filter_firBlock_left_multProducts[1], n1789, n1788 );
xor U685 ( n1788, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[9], n343 );
nand U686 ( n1789, n1640, n1639 );
nand U687 ( n1640, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[8], n1787 );
nand U688 ( n1639, n1638, n341 );
or U689 ( n1638, n1787, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[8] );
xor U690 ( my_IIR_filter_firBlock_left_multProducts[2], n1645, n1644 );
nand U691 ( n1645, n1643, n1642 );
nand U692 ( n1643, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[9], n1789 );
nand U693 ( n1642, n1641, n343 );
or U694 ( n1641, n1789, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[9] );
xor U695 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[11], n3058, n3057 );
xor U696 ( my_IIR_filter_firBlock_left_multProducts[3], n1650, n1649 );
xor U697 ( n1649, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[11], n49 );
nand U698 ( n1650, n1648, n1647 );
nand U699 ( n1647, n1646, n48 );
xor U700 ( my_IIR_filter_firBlock_left_multProducts[4], n1655, n1654 );
xor U701 ( n1654, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[12], n50 );
nand U702 ( n1655, n1653, n1652 );
nand U703 ( n1653, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[11], n1650 );
nand U704 ( n1652, n1651, n49 );
or U705 ( n1651, n1650, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[11] );
xor U706 ( my_IIR_filter_firBlock_left_multProducts[5], n1660, n1659 );
xor U707 ( n1659, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[13], n306 );
nand U708 ( n1660, n1658, n1657 );
nand U709 ( n1658, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[12], n1655 );
nand U710 ( n1657, n1656, n50 );
or U711 ( n1656, n1655, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[12] );
xor U712 ( my_IIR_filter_firBlock_left_multProducts[6], n1665, n1664 );
nand U713 ( n1665, n1663, n1662 );
nand U714 ( n1663, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[13], n1660 );
nand U715 ( n1662, n1661, n306 );
or U716 ( n1661, n1660, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[13] );
xnor U717 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[31], n2913, n238 );
xnor U718 ( n238, outData_in[30], n209 );
xor U719 ( my_IIR_filter_firBlock_left_multProducts[7], n1670, n1669 );
xor U720 ( n1669, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[15], n302 );
nand U721 ( n1670, n1668, n1667 );
nand U722 ( n1667, n1666, n294 );
xor U723 ( my_IIR_filter_firBlock_left_multProducts[8], n1675, n1674 );
xor U724 ( n1674, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[16], n298 );
nand U725 ( n1675, n1673, n1672 );
nand U726 ( n1673, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[15], n1670 );
nand U727 ( n1672, n1671, n302 );
or U728 ( n1671, n1670, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[15] );
xor U729 ( my_IIR_filter_firBlock_left_multProducts[9], n1680, n1679 );
nand U730 ( n1680, n1678, n1677 );
nand U731 ( n1678, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[16], n1675 );
nand U732 ( n1677, n1676, n298 );
or U733 ( n1676, n1675, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[16] );
nand U734 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[34], n2925, n2924 );
nand U735 ( n2924, n524, n2923 );
xor U736 ( my_IIR_filter_firBlock_left_multProducts[10], n1685, n1684 );
nand U737 ( n1685, n1683, n1682 );
nand U738 ( n1682, n1681, n300 );
xor U739 ( my_IIR_filter_firBlock_left_multProducts[11], n1690, n1689 );
nand U740 ( n1690, n1688, n1687 );
nand U741 ( n1687, n1686, n296 );
buf U742 ( n505, outData_in[25] );
not U743 ( n690, outData_in[21] );
xor U744 ( my_IIR_filter_firBlock_left_multProducts[12], n1695, n1694 );
nand U745 ( n1695, n1693, n1692 );
nand U746 ( n1692, n1691, n304 );
buf U747 ( n512, outData_in[17] );
buf U748 ( n515, outData_in[29] );
xor U749 ( my_IIR_filter_firBlock_left_multProducts[13], n1700, n1699 );
xor U750 ( n1699, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[21], n52 );
nand U751 ( n1700, n1698, n1697 );
nand U752 ( n1697, n1696, n51 );
buf U753 ( n491, outData_in[27] );
xor U754 ( my_IIR_filter_firBlock_left_multProducts[14], n1705, n1704 );
nand U755 ( n1705, n1703, n1702 );
nand U756 ( n1703, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[21], n1700 );
nand U757 ( n1702, n1701, n52 );
or U758 ( n1701, n1700, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[21] );
xnor U759 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[27], n2895, n239 );
xnor U760 ( n239, n158, n157 );
xor U761 ( my_IIR_filter_firBlock_left_multProducts[15], n1710, n1709 );
nand U762 ( n1710, n1708, n1707 );
nand U763 ( n1707, n1706, n53 );
xor U764 ( my_IIR_filter_firBlock_left_multProducts[16], n1715, n1714 );
nand U765 ( n1715, n1713, n1712 );
nand U766 ( n1712, n1711, n308 );
buf U767 ( n501, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[2] );
xor U768 ( my_IIR_filter_firBlock_left_multProducts[17], n1720, n1719 );
xor U769 ( n1719, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[25], n55 );
nand U770 ( n1720, n1718, n1717 );
nand U771 ( n1717, n1716, n54 );
xor U772 ( my_IIR_filter_firBlock_left_multProducts[18], n1725, n1724 );
xor U773 ( n1724, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[26], n56 );
nand U774 ( n1725, n1723, n1722 );
nand U775 ( n1723, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[25], n1720 );
nand U776 ( n1722, n1721, n55 );
or U777 ( n1721, n1720, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[25] );
xnor U778 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[25], n2886, n240 );
xnor U779 ( n240, n157, n490 );
nand U780 ( n1730, n1728, n1727 );
nand U781 ( n1728, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[26], n1725 );
nand U782 ( n1727, n1726, n56 );
or U783 ( n1726, n1725, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[26] );
xor U784 ( my_IIR_filter_firBlock_left_multProducts[19], n1730, n1729 );
xor U785 ( my_IIR_filter_firBlock_left_multProducts[20], n1735, n1734 );
nand U786 ( n1735, n1733, n1732 );
nand U787 ( n1732, n1731, n57 );
xor U788 ( my_IIR_filter_firBlock_left_multProducts[21], n1740, n1739 );
xor U789 ( n1739, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[29], n60 );
nand U790 ( n1740, n1738, n1737 );
nand U791 ( n1737, n1736, n59 );
xor U792 ( my_IIR_filter_firBlock_left_multProducts[22], n1745, n1744 );
nand U793 ( n1745, n1743, n1742 );
nand U794 ( n1743, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[29], n1740 );
nand U795 ( n1742, n1741, n60 );
or U796 ( n1741, n1740, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[29] );
xor U797 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[24], n241, n2882 );
xor U798 ( n241, n154, outData_in[23] );
xor U799 ( my_IIR_filter_firBlock_left_multProducts[23], n1750, n1749 );
nand U800 ( n1750, n1748, n1747 );
nand U801 ( n1747, n1746, n61 );
xor U802 ( my_IIR_filter_firBlock_left_multProducts[24], n1755, n1754 );
xor U803 ( n1754, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[32], n526 );
nand U804 ( n1755, n1753, n1752 );
nand U805 ( n1752, n1751, n527 );
xor U806 ( my_IIR_filter_firBlock_left_multProducts[25], n1760, n1759 );
nand U807 ( n1760, n1758, n1757 );
nand U808 ( n1758, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[32], n1755 );
nand U809 ( n1757, n1756, n527 );
or U810 ( n1756, n1755, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[32] );
xor U811 ( my_IIR_filter_firBlock_left_multProducts[26], n1765, n1764 );
nand U812 ( n1765, n1763, n1762 );
nand U813 ( n1762, n1761, n527 );
nor U814 ( n2631, n2629, n2628 );
xor U815 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[22], n242, n2874 );
xor U816 ( n242, n494, n154 );
xor U817 ( my_IIR_filter_firBlock_left_multProducts[27], n1770, n1769 );
xor U818 ( n1769, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[35], n526 );
nand U819 ( n1770, n1768, n1767 );
nand U820 ( n1767, n1766, n527 );
nand U821 ( n1775, n1773, n1772 );
nand U822 ( n1773, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[35], n1770 );
nand U823 ( n1772, n1771, n527 );
or U824 ( n1771, n1770, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[35] );
xnor U825 ( n243, n1785, n1784 );
nand U826 ( n1780, n1778, n1777 );
nand U827 ( n1777, n1776, n527 );
xor U828 ( my_IIR_filter_firBlock_left_multProducts[28], n1775, n1774 );
xnor U829 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[19], n2861, n244 );
xnor U830 ( n244, outData_in[18], outData_in[16] );
xor U831 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[6], n245, n2929 );
xor U832 ( n245, n503, outData_in[5] );
buf U833 ( n492, outData_in[27] );
xor U834 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[8], n247, n2932 );
xor U835 ( n247, outData_in[5], outData_in[7] );
not U836 ( n630, my_IIR_filter_firBlock_left_multProducts[60] );
nand U837 ( n2646, n2644, n2643 );
nor U838 ( n2645, n512, n2646 );
nor U839 ( n2649, n2647, n2646 );
nand U840 ( n2652, n2650, n2649 );
nand U841 ( n2654, n2655, n692 );
nand U842 ( n2658, n2656, n2655 );
nor U843 ( n2661, n2659, n2658 );
nand U844 ( n2660, n2661, n696 );
nor U845 ( n2666, n2665, n2664 );
nand U846 ( n2664, n2662, n2661 );
nor U847 ( n2663, n515, n2664 );
and U848 ( n3582, n3581, n3580 );
nor U849 ( n3580, n3578, n3577 );
nand U850 ( n3579, n3580, n698 );
nand U851 ( n3577, n3575, n3574 );
nor U852 ( n3574, n3572, n3571 );
nand U853 ( n3573, n3574, n694 );
nor U854 ( n3570, n529, n3571 );
nor U855 ( n3568, n3566, n3565 );
nand U856 ( n3565, n3563, n3562 );
nor U857 ( n3562, n3560, n3559 );
buf U858 ( n550, n39 );
nand U859 ( n3561, n3562, n686 );
nor U860 ( n3558, n495, n3559 );
buf U861 ( n624, n626 );
buf U862 ( n623, n626 );
buf U863 ( n622, n626 );
buf U864 ( n621, n626 );
buf U865 ( n620, n627 );
buf U866 ( n619, n627 );
buf U867 ( n618, n627 );
buf U868 ( n617, n627 );
buf U869 ( n616, n627 );
buf U870 ( n615, n628 );
buf U871 ( n614, n628 );
buf U872 ( n613, n628 );
buf U873 ( n612, n628 );
buf U874 ( n611, n628 );
buf U875 ( n610, n629 );
buf U876 ( n609, n629 );
buf U877 ( n608, n629 );
buf U878 ( n607, n629 );
buf U879 ( n625, n626 );
xnor U880 ( my_IIR_filter_firBlock_right_N192, n248, n3532 );
nand U881 ( n3474, my_IIR_filter_firBlock_right_multProducts[18], n3473 );
nor U882 ( n3528, my_IIR_filter_firBlock_right_firStep[30], n3529 );
nand U883 ( n3529, n3527, n3526 );
nand U884 ( n3496, n3495, n3494 );
nand U885 ( n3505, n3504, n3503 );
nand U886 ( n3503, my_IIR_filter_firBlock_right_multProducts[24], n3502 );
nand U887 ( n3514, n3513, n3512 );
nand U888 ( n3512, my_IIR_filter_firBlock_right_multProducts[26], n3511 );
nand U889 ( n3518, n3517, n3516 );
nand U890 ( n3492, n3490, n3489 );
nand U891 ( n3489, my_IIR_filter_firBlock_right_multProducts[21], n3488 );
nand U892 ( n3523, n3410, n3409 );
nand U893 ( n3410, my_IIR_filter_firBlock_right_firStep[1], n3477 );
nand U894 ( n3409, my_IIR_filter_firBlock_right_multProducts[1], n3408 );
or U895 ( n3408, my_IIR_filter_firBlock_right_firStep[1], n3477 );
xor U896 ( n805, rightOut[6], leftOut[6] );
nand U897 ( n3418, my_IIR_filter_firBlock_right_multProducts[4], n3417 );
nand U898 ( n3433, my_IIR_filter_firBlock_right_multProducts[9], n3432 );
nand U899 ( n3533, n3413, n3412 );
nand U900 ( n3412, my_IIR_filter_firBlock_right_multProducts[2], n3411 );
nand U901 ( n3458, n3457, n3456 );
nand U902 ( n3456, my_IIR_filter_firBlock_right_multProducts[14], n3455 );
nand U903 ( n3449, n3448, n3447 );
nand U904 ( n3440, n3439, n3438 );
nand U905 ( n3438, my_IIR_filter_firBlock_right_multProducts[10], n3437 );
nand U906 ( n3454, n3452, n3451 );
nand U907 ( n3451, my_IIR_filter_firBlock_right_multProducts[13], n3450 );
nand U908 ( n3538, n3422, n3421 );
nand U909 ( n3421, my_IIR_filter_firBlock_right_multProducts[5], n3420 );
nand U910 ( n3541, n3428, n3427 );
nand U911 ( n3427, my_IIR_filter_firBlock_right_multProducts[7], n3426 );
nand U912 ( n3535, n3416, n3415 );
nand U913 ( n3415, my_IIR_filter_firBlock_right_multProducts[3], n3414 );
or U914 ( n807, n249, n250 );
and U915 ( n249, leftOut[6], n806 );
and U916 ( n250, rightOut[6], n721 );
xnor U917 ( my_IIR_filter_firBlock_right_N128, n251, n3345 );
nor U918 ( n1206, my_IIR_filter_firBlock_left_firStep[286], n1207 );
nand U919 ( n1184, my_IIR_filter_firBlock_left_multProducts[86], n1183 );
nand U920 ( n1193, my_IIR_filter_firBlock_left_multProducts[88], n1192 );
xor U921 ( my_IIR_filter_firBlock_left_N32, n1211, n1210 );
xnor U922 ( n1211, my_IIR_filter_firBlock_left_multProducts[89], my_IIR_filter_firBlock_left_firStep[287] );
nor U923 ( n1210, n1209, n1208 );
nand U924 ( n1207, n1205, n1204 );
nand U925 ( n1204, my_IIR_filter_firBlock_left_multProducts[89], n1203 );
nand U926 ( n1182, n1181, n1180 );
nand U927 ( n1181, my_IIR_filter_firBlock_left_firStep[280], n1178 );
or U928 ( n1179, n1178, my_IIR_filter_firBlock_left_firStep[280] );
nand U929 ( n1191, n1190, n1189 );
nand U930 ( n1202, n1199, n1198 );
nand U931 ( n1198, my_IIR_filter_firBlock_left_multProducts[89], n1197 );
nand U932 ( n1178, n1176, n1175 );
nand U933 ( n1173, n1172, n1171 );
nand U934 ( n1171, my_IIR_filter_firBlock_left_multProducts[83], n1170 );
nand U935 ( n1164, n1163, n1162 );
nand U936 ( n1163, my_IIR_filter_firBlock_left_firStep[276], n1160 );
nand U937 ( n1162, my_IIR_filter_firBlock_left_multProducts[81], n1161 );
or U938 ( n1161, n1160, my_IIR_filter_firBlock_left_firStep[276] );
nand U939 ( n1169, n1167, n1166 );
nand U940 ( n1166, my_IIR_filter_firBlock_left_multProducts[82], n1165 );
xnor U941 ( n252, n54, my_IIR_filter_firBlock_left_multProducts[110] );
nand U942 ( n898, n897, n55 );
nand U943 ( n821, inData_in[3], n938 );
or U944 ( n819, n938, inData_in[3] );
or U945 ( n946, n253, n254 );
and U946 ( n253, my_IIR_filter_firBlock_left_multProducts[90], n944 );
and U947 ( n254, n827, n341 );
or U948 ( n850, n255, n256 );
and U949 ( n255, my_IIR_filter_firBlock_left_multProducts[96], n847 );
and U950 ( n256, n848, n294 );
and U951 ( n257, my_IIR_filter_firBlock_left_multProducts[100], n865 );
and U952 ( n258, n866, n296 );
nand U953 ( n886, n884, n883 );
nand U954 ( n883, n882, n53 );
nand U955 ( n938, n818, n817 );
nand U956 ( n817, n816, n44 );
or U957 ( n835, n343, n259 );
nor U958 ( n259, n49, n834 );
nand U959 ( n862, n861, n300 );
or U960 ( n831, n341, n260 );
nor U961 ( n260, n48, n830 );
nand U962 ( n855, n853, n852 );
nand U963 ( n853, my_IIR_filter_firBlock_left_multProducts[97], n850 );
nand U964 ( n852, n851, n302 );
or U965 ( n851, n850, my_IIR_filter_firBlock_left_multProducts[97] );
nand U966 ( n891, n889, n888 );
nand U967 ( n889, my_IIR_filter_firBlock_left_multProducts[105], n886 );
nand U968 ( n888, n887, n308 );
or U969 ( n887, n886, my_IIR_filter_firBlock_left_multProducts[105] );
nand U970 ( n842, n841, n840 );
nand U971 ( n840, n839, n50 );
nand U972 ( n881, n879, n878 );
nand U973 ( n878, n877, n52 );
nand U974 ( n860, n858, n857 );
nand U975 ( n858, my_IIR_filter_firBlock_left_multProducts[98], n855 );
nand U976 ( n857, n856, n298 );
or U977 ( n856, n855, my_IIR_filter_firBlock_left_multProducts[98] );
nand U978 ( n896, n894, n893 );
nand U979 ( n894, my_IIR_filter_firBlock_left_multProducts[106], n891 );
nand U980 ( n893, n892, n54 );
or U981 ( n892, n891, my_IIR_filter_firBlock_left_multProducts[106] );
nand U982 ( n944, n826, n825 );
nand U983 ( n825, n824, n47 );
nand U984 ( n844, n843, n306 );
nand U985 ( n1155, n1152, n1151 );
nand U986 ( n1152, my_IIR_filter_firBlock_left_firStep[274], n1149 );
nand U987 ( n1151, my_IIR_filter_firBlock_left_multProducts[79], n1150 );
or U988 ( n1150, n1149, my_IIR_filter_firBlock_left_firStep[274] );
nand U989 ( n1149, n1147, n1146 );
nand U990 ( n1146, my_IIR_filter_firBlock_left_multProducts[78], n1145 );
nand U991 ( n1144, n1143, n1142 );
nand U992 ( n1143, my_IIR_filter_firBlock_left_firStep[272], n1140 );
xnor U993 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[19], n842, n261 );
xnor U994 ( n261, n306, my_IIR_filter_firBlock_left_multProducts[95] );
xor U995 ( my_IIR_filter_firBlock_left_multProducts[67], n983, n982 );
nand U996 ( n1220, n1105, n1104 );
nand U997 ( n1104, my_IIR_filter_firBlock_left_multProducts[68], n1103 );
nand U998 ( n1113, n1111, n1110 );
nand U999 ( n1131, n1129, n1128 );
nand U1000 ( n1140, n1138, n1137 );
nand U1001 ( n1137, my_IIR_filter_firBlock_left_multProducts[76], n1136 );
nand U1002 ( n1135, n1134, n1133 );
nand U1003 ( n1134, my_IIR_filter_firBlock_left_firStep[270], n1131 );
nand U1004 ( n1133, my_IIR_filter_firBlock_left_multProducts[75], n1132 );
or U1005 ( n1132, n1131, my_IIR_filter_firBlock_left_firStep[270] );
nand U1006 ( n1122, n1120, n1119 );
nand U1007 ( n1119, my_IIR_filter_firBlock_left_multProducts[72], n1118 );
nand U1008 ( n1126, n1125, n1124 );
nand U1009 ( n1221, n1108, n1107 );
nand U1010 ( n1108, my_IIR_filter_firBlock_left_firStep[264], n1220 );
or U1011 ( n1106, n1220, my_IIR_filter_firBlock_left_firStep[264] );
nand U1012 ( n1117, n1116, n1115 );
nand U1013 ( n1116, my_IIR_filter_firBlock_left_firStep[266], n1113 );
nand U1014 ( n1115, my_IIR_filter_firBlock_left_multProducts[71], n1114 );
or U1015 ( n1114, n1113, my_IIR_filter_firBlock_left_firStep[266] );
nand U1016 ( n1218, n1102, n1101 );
nand U1017 ( n1102, my_IIR_filter_firBlock_left_firStep[262], n1217 );
nand U1018 ( n1101, my_IIR_filter_firBlock_left_multProducts[67], n1100 );
or U1019 ( n1100, n1217, my_IIR_filter_firBlock_left_firStep[262] );
xor U1020 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[26], n872, n871 );
xor U1021 ( n871, n296, my_IIR_filter_firBlock_left_multProducts[104] );
xor U1022 ( n890, n53, my_IIR_filter_firBlock_left_multProducts[108] );
xnor U1023 ( my_IIR_filter_firBlock_left_multProducts[78], n1033, n262 );
xnor U1024 ( n262, my_IIR_filter_firBlock_left_multProducts[105], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[30] );
xor U1025 ( n791, n538, n263 );
xnor U1026 ( n264, rightOut[24], leftOut[24] );
nand U1027 ( n746, leftOut[14], n744 );
nand U1028 ( n3333, my_IIR_filter_firBlock_right_multProducts[59], n3332 );
xor U1029 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[25], n868, n867 );
xor U1030 ( n867, n300, my_IIR_filter_firBlock_left_multProducts[103] );
xnor U1031 ( my_IIR_filter_firBlock_left_multProducts[73], n1009, n265 );
xnor U1032 ( n265, my_IIR_filter_firBlock_left_multProducts[100], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[25] );
xor U1033 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[16], n830, n829 );
xor U1034 ( n829, n341, my_IIR_filter_firBlock_left_multProducts[94] );
xor U1035 ( n968, my_IIR_filter_firBlock_left_multProducts[91], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[16] );
nand U1036 ( n1215, n1096, n1095 );
nand U1037 ( n1214, n1093, n1092 );
nand U1038 ( n1217, n1099, n1098 );
xor U1039 ( n728, rightOut[10], leftOut[10] );
nand U1040 ( n3255, my_IIR_filter_firBlock_right_multProducts[42], n3254 );
nand U1041 ( n3349, n3232, n3231 );
nand U1042 ( n3352, n3238, n3237 );
nand U1043 ( n3237, n3236, my_IIR_filter_firBlock_right_multProducts[37] );
nand U1044 ( n3346, n3226, n3225 );
nand U1045 ( n3226, my_IIR_filter_firBlock_right_firStep[33], n3336 );
nand U1046 ( n3225, my_IIR_filter_firBlock_right_multProducts[33], n3224 );
or U1047 ( n3224, n3336, my_IIR_filter_firBlock_right_firStep[33] );
nand U1048 ( n3354, n3241, n3240 );
nand U1049 ( n3351, n3235, n3234 );
nand U1050 ( n3348, n3229, n3228 );
xnor U1051 ( n266, rightOut[28], leftOut[28] );
xnor U1052 ( n267, rightOut[26], leftOut[26] );
xnor U1053 ( n739, leftOut[13], rightOut[13] );
xor U1054 ( n837, n50, my_IIR_filter_firBlock_left_multProducts[94] );
xnor U1055 ( my_IIR_filter_firBlock_left_multProducts[66], n978, n268 );
xnor U1056 ( n268, my_IIR_filter_firBlock_left_multProducts[93], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[18] );
xor U1057 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[21], n850, n849 );
xor U1058 ( n849, n306, my_IIR_filter_firBlock_left_multProducts[99] );
xnor U1059 ( my_IIR_filter_firBlock_left_multProducts[69], n991, n269 );
xnor U1060 ( n269, my_IIR_filter_firBlock_left_multProducts[96], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[21] );
xnor U1061 ( my_IIR_filter_firBlock_right_N127, n3342, n270 );
xor U1062 ( n270, n210, my_IIR_filter_firBlock_right_firStep[61] );
xor U1063 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[29], n886, n885 );
xor U1064 ( n885, n52, my_IIR_filter_firBlock_left_multProducts[107] );
nand U1065 ( n917, n913, n912 );
nand U1066 ( n912, n911, n59 );
nand U1067 ( n903, my_IIR_filter_firBlock_left_multProducts[108], n900 );
nand U1068 ( n902, n901, n56 );
or U1069 ( n901, n900, my_IIR_filter_firBlock_left_multProducts[108] );
nand U1070 ( n910, n908, n907 );
nand U1071 ( n907, n906, n57 );
xor U1072 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[36], n922, n921 );
xor U1073 ( n921, n61, my_IIR_filter_firBlock_left_multProducts[112] );
xnor U1074 ( my_IIR_filter_firBlock_left_multProducts[84], n1060, n271 );
xnor U1075 ( n271, my_IIR_filter_firBlock_left_multProducts[111], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[36] );
nand U1076 ( n922, n920, n919 );
nand U1077 ( n920, my_IIR_filter_firBlock_left_multProducts[111], n917 );
nand U1078 ( n919, n918, n60 );
or U1079 ( n918, n917, my_IIR_filter_firBlock_left_multProducts[111] );
xnor U1080 ( n732, leftOut[11], rightOut[11] );
xor U1081 ( n808, rightOut[8], leftOut[8] );
xor U1082 ( n859, n302, my_IIR_filter_firBlock_left_multProducts[101] );
xnor U1083 ( my_IIR_filter_firBlock_left_multProducts[71], n1000, n272 );
xnor U1084 ( n272, my_IIR_filter_firBlock_left_multProducts[98], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[23] );
xor U1085 ( n931, n61, n549 );
nand U1086 ( n932, n930, n929 );
nand U1087 ( n930, my_IIR_filter_firBlock_left_multProducts[113], n927 );
xnor U1088 ( my_IIR_filter_firBlock_left_multProducts[86], n1067, n273 );
xnor U1089 ( n273, my_IIR_filter_firBlock_left_multProducts[113], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[38] );
nand U1090 ( n927, n925, n924 );
nand U1091 ( n925, my_IIR_filter_firBlock_left_multProducts[112], n922 );
nand U1092 ( n924, n923, n61 );
or U1093 ( n923, n922, my_IIR_filter_firBlock_left_multProducts[112] );
nand U1094 ( n929, n928, n527 );
or U1095 ( n928, n927, my_IIR_filter_firBlock_left_multProducts[113] );
xor U1096 ( my_IIR_filter_firBlock_left_multProducts[87], n1072, n1071 );
xor U1097 ( n1071, my_IIR_filter_firBlock_left_multProducts[114], n549 );
nand U1098 ( n1072, n1070, n1069 );
nand U1099 ( n1069, my_IIR_filter_firBlock_left_multProducts[113], n1068 );
xor U1100 ( n935, n42, inData_in[4] );
nand U1101 ( n954, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[11], n951 );
nand U1102 ( n953, inData_in[2], n952 );
or U1103 ( n952, n951, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[11] );
nand U1104 ( n967, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[15], n1084 );
nand U1105 ( n966, my_IIR_filter_firBlock_left_multProducts[90], n965 );
or U1106 ( n965, n1084, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[15] );
nand U1107 ( n974, n972, n971 );
nand U1108 ( n971, my_IIR_filter_firBlock_left_multProducts[91], n970 );
nand U1109 ( n978, n977, n976 );
nand U1110 ( n976, my_IIR_filter_firBlock_left_multProducts[92], n975 );
nand U1111 ( n1084, n964, n963 );
nand U1112 ( n963, inData_in[5], n962 );
nand U1113 ( n1046, n1044, n1043 );
nand U1114 ( n1043, my_IIR_filter_firBlock_left_multProducts[107], n1042 );
nand U1115 ( n983, n981, n980 );
nand U1116 ( n980, my_IIR_filter_firBlock_left_multProducts[93], n979 );
nand U1117 ( n1024, n1022, n1021 );
nand U1118 ( n1021, my_IIR_filter_firBlock_left_multProducts[102], n1020 );
nand U1119 ( n1051, n1049, n1048 );
nand U1120 ( n1048, my_IIR_filter_firBlock_left_multProducts[108], n1047 );
nand U1121 ( n1000, n999, n998 );
nand U1122 ( n998, my_IIR_filter_firBlock_left_multProducts[97], n997 );
nand U1123 ( n1033, n1032, n1031 );
nand U1124 ( n1031, my_IIR_filter_firBlock_left_multProducts[104], n1030 );
nand U1125 ( n1060, n1059, n1058 );
nand U1126 ( n1058, my_IIR_filter_firBlock_left_multProducts[110], n1057 );
nand U1127 ( n1082, n961, n960 );
nand U1128 ( n960, inData_in[4], n959 );
nand U1129 ( n1014, n1012, n1011 );
nand U1130 ( n1011, my_IIR_filter_firBlock_left_multProducts[100], n1010 );
nand U1131 ( n951, n950, n949 );
and U1132 ( n948, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[9], n947 );
nand U1133 ( n1019, n1017, n1016 );
nand U1134 ( n1017, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[26], n1014 );
nand U1135 ( n1080, n958, n957 );
nand U1136 ( n958, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[12], n955 );
nand U1137 ( n957, inData_in[3], n956 );
or U1138 ( n956, n955, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[12] );
nand U1139 ( n1038, n1036, n1035 );
nand U1140 ( n1035, my_IIR_filter_firBlock_left_multProducts[105], n1034 );
nand U1141 ( n1029, n1027, n1026 );
nand U1142 ( n1026, my_IIR_filter_firBlock_left_multProducts[103], n1025 );
nand U1143 ( n1056, n1054, n1053 );
nand U1144 ( n1053, my_IIR_filter_firBlock_left_multProducts[109], n1052 );
nand U1145 ( n1009, n1008, n1007 );
nand U1146 ( n1007, my_IIR_filter_firBlock_left_multProducts[99], n1006 );
nand U1147 ( n1005, n1003, n1002 );
nand U1148 ( n1002, my_IIR_filter_firBlock_left_multProducts[98], n1001 );
nand U1149 ( n991, n990, n989 );
nand U1150 ( n989, my_IIR_filter_firBlock_left_multProducts[95], n988 );
nand U1151 ( n987, n986, n985 );
nand U1152 ( n985, my_IIR_filter_firBlock_left_multProducts[94], n984 );
nand U1153 ( n996, n994, n993 );
nand U1154 ( n993, my_IIR_filter_firBlock_left_multProducts[96], n992 );
nand U1155 ( n1065, n1063, n1062 );
nand U1156 ( n1062, my_IIR_filter_firBlock_left_multProducts[111], n1061 );
nand U1157 ( n1075, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n1072 );
nand U1158 ( n1074, my_IIR_filter_firBlock_left_multProducts[114], n1073 );
or U1159 ( n1073, n1072, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_ );
xor U1160 ( n875, n304, my_IIR_filter_firBlock_left_multProducts[105] );
xor U1161 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[35], n917, n914 );
xor U1162 ( n914, n57, my_IIR_filter_firBlock_left_multProducts[113] );
xor U1163 ( n880, n51, my_IIR_filter_firBlock_left_multProducts[106] );
xor U1164 ( my_IIR_filter_firBlock_left_multProducts[76], n1024, n1023 );
xnor U1165 ( n811, leftOut[9], rightOut[9] );
nand U1166 ( n3336, n3223, n3222 );
nand U1167 ( n3223, my_IIR_filter_firBlock_right_firStep[32], n3290 );
or U1168 ( n3221, my_IIR_filter_firBlock_right_firStep[32], n3290 );
xor U1169 ( n945, n47, my_IIR_filter_firBlock_left_multProducts[93] );
nand U1170 ( n1212, n1090, n1089 );
nand U1171 ( n1090, my_IIR_filter_firBlock_left_firStep[258], n1201 );
nand U1172 ( n1089, my_IIR_filter_firBlock_left_multProducts[63], n1088 );
or U1173 ( n1088, n1201, my_IIR_filter_firBlock_left_firStep[258] );
xor U1174 ( n895, n308, my_IIR_filter_firBlock_left_multProducts[109] );
xnor U1175 ( my_IIR_filter_firBlock_left_multProducts[68], n987, n274 );
xnor U1176 ( n274, my_IIR_filter_firBlock_left_multProducts[95], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[20] );
xor U1177 ( n846, n50, my_IIR_filter_firBlock_left_multProducts[98] );
xor U1178 ( n833, n343, my_IIR_filter_firBlock_left_multProducts[95] );
xnor U1179 ( outData_in[20], n764, n275 );
xnor U1180 ( n275, rightOut[20], leftOut[20] );
xor U1181 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[12], n940, n939 );
xor U1182 ( n939, n44, my_IIR_filter_firBlock_left_multProducts[90] );
xor U1183 ( n909, n56, my_IIR_filter_firBlock_left_multProducts[112] );
xor U1184 ( my_IIR_filter_firBlock_left_multProducts[82], n1051, n1050 );
xnor U1185 ( n2465, my_IIR_filter_firBlock_left_multProducts[89], my_IIR_filter_firBlock_left_firStep[63] );
nand U1186 ( n2450, n2448, n2447 );
nand U1187 ( n2447, my_IIR_filter_firBlock_left_multProducts[88], n2446 );
nand U1188 ( n2445, n2444, n2443 );
nand U1189 ( n2444, my_IIR_filter_firBlock_left_firStep[58], n2441 );
or U1190 ( n2442, n2441, my_IIR_filter_firBlock_left_firStep[58] );
nand U1191 ( n2456, n2453, n2452 );
nand U1192 ( n2453, my_IIR_filter_firBlock_left_firStep[60], n2450 );
nand U1193 ( n2452, my_IIR_filter_firBlock_left_multProducts[89], n2451 );
or U1194 ( n2451, n2450, my_IIR_filter_firBlock_left_firStep[60] );
nand U1195 ( n2461, n2459, n2458 );
nand U1196 ( n2458, my_IIR_filter_firBlock_left_multProducts[89], n2457 );
xnor U1197 ( outData_in[30], n797, n276 );
xor U1198 ( n276, n58, leftOut[30] );
or U1199 ( n793, n277, n278 );
nor U1200 ( n277, n531, n530 );
and U1201 ( n278, leftOut[28], n790 );
xor U1202 ( n904, n55, my_IIR_filter_firBlock_left_multProducts[111] );
xor U1203 ( n854, n294, my_IIR_filter_firBlock_left_multProducts[100] );
xor U1204 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[13], n942, n941 );
xor U1205 ( n941, n45, my_IIR_filter_firBlock_left_multProducts[91] );
xor U1206 ( n1079, inData_in[4], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[13] );
nand U1207 ( n1201, n1087, n1086 );
nand U1208 ( n1087, my_IIR_filter_firBlock_left_firStep[257], n1154 );
or U1209 ( n1085, my_IIR_filter_firBlock_left_firStep[257], n1154 );
and U1210 ( n1154, my_IIR_filter_firBlock_left_multProducts[61], my_IIR_filter_firBlock_left_firStep[256] );
xor U1211 ( n802, n539, n279 );
xor U1212 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[11], n938, n937 );
xor U1213 ( n937, n43, inData_in[5] );
xor U1214 ( n943, n46, my_IIR_filter_firBlock_left_multProducts[92] );
xor U1215 ( my_IIR_filter_firBlock_left_multProducts[62], n1082, n1081 );
nand U1216 ( n2049, n2046, n2045 );
nand U1217 ( n2046, my_IIR_filter_firBlock_left_firStep[157], n2043 );
nand U1218 ( n2045, my_IIR_filter_firBlock_left_multProducts[29], n2044 );
or U1219 ( n2044, n2043, my_IIR_filter_firBlock_left_firStep[157] );
nand U1220 ( n2032, n2031, n2030 );
nand U1221 ( n2031, my_IIR_filter_firBlock_left_firStep[154], n2028 );
nand U1222 ( n2030, my_IIR_filter_firBlock_left_multProducts[26], n2029 );
or U1223 ( n2029, n2028, my_IIR_filter_firBlock_left_firStep[154] );
nand U1224 ( n1896, n1895, n1894 );
nand U1225 ( n1895, my_IIR_filter_firBlock_left_firStep[186], n1892 );
nand U1226 ( n1894, my_IIR_filter_firBlock_left_multProducts[26], n1893 );
or U1227 ( n1893, n1892, my_IIR_filter_firBlock_left_firStep[186] );
nand U1228 ( n2023, n2022, n2021 );
nand U1229 ( n2022, my_IIR_filter_firBlock_left_firStep[152], n2019 );
nand U1230 ( n2021, my_IIR_filter_firBlock_left_multProducts[24], n2020 );
or U1231 ( n2020, n2019, my_IIR_filter_firBlock_left_firStep[152] );
nand U1232 ( n1887, n1886, n1885 );
nand U1233 ( n1886, my_IIR_filter_firBlock_left_firStep[184], n1883 );
nand U1234 ( n1885, my_IIR_filter_firBlock_left_multProducts[24], n1884 );
or U1235 ( n1884, n1883, my_IIR_filter_firBlock_left_firStep[184] );
nand U1236 ( n2043, n2040, n2039 );
nand U1237 ( n2040, my_IIR_filter_firBlock_left_firStep[156], n2037 );
nand U1238 ( n2039, my_IIR_filter_firBlock_left_multProducts[28], n2038 );
or U1239 ( n2038, n2037, my_IIR_filter_firBlock_left_firStep[156] );
nand U1240 ( n1907, n1904, n1903 );
nand U1241 ( n1904, my_IIR_filter_firBlock_left_firStep[188], n1901 );
nand U1242 ( n1903, my_IIR_filter_firBlock_left_multProducts[28], n1902 );
or U1243 ( n1902, n1901, my_IIR_filter_firBlock_left_firStep[188] );
nand U1244 ( n2014, n2013, n2012 );
nand U1245 ( n2013, my_IIR_filter_firBlock_left_firStep[150], n2010 );
nand U1246 ( n2012, my_IIR_filter_firBlock_left_multProducts[22], n2011 );
or U1247 ( n2011, n2010, my_IIR_filter_firBlock_left_firStep[150] );
nand U1248 ( n1878, n1877, n1876 );
nand U1249 ( n1877, my_IIR_filter_firBlock_left_firStep[182], n1874 );
nand U1250 ( n1876, my_IIR_filter_firBlock_left_multProducts[22], n1875 );
or U1251 ( n1875, n1874, my_IIR_filter_firBlock_left_firStep[182] );
nand U1252 ( n1985, n1984, n1983 );
nand U1253 ( n1984, my_IIR_filter_firBlock_left_firStep[144], n1981 );
nand U1254 ( n1983, my_IIR_filter_firBlock_left_multProducts[16], n1982 );
or U1255 ( n1982, n1981, my_IIR_filter_firBlock_left_firStep[144] );
nand U1256 ( n1849, n1848, n1847 );
nand U1257 ( n1848, my_IIR_filter_firBlock_left_firStep[176], n1845 );
nand U1258 ( n1847, my_IIR_filter_firBlock_left_multProducts[16], n1846 );
or U1259 ( n1846, n1845, my_IIR_filter_firBlock_left_firStep[176] );
nand U1260 ( n1976, n1975, n1974 );
nand U1261 ( n1975, my_IIR_filter_firBlock_left_firStep[142], n1972 );
nand U1262 ( n1974, my_IIR_filter_firBlock_left_multProducts[14], n1973 );
or U1263 ( n1973, n1972, my_IIR_filter_firBlock_left_firStep[142] );
nand U1264 ( n1840, n1839, n1838 );
nand U1265 ( n1839, my_IIR_filter_firBlock_left_firStep[174], n1836 );
nand U1266 ( n1838, my_IIR_filter_firBlock_left_multProducts[14], n1837 );
or U1267 ( n1837, n1836, my_IIR_filter_firBlock_left_firStep[174] );
nand U1268 ( n1967, n1966, n1965 );
nand U1269 ( n1966, my_IIR_filter_firBlock_left_firStep[140], n1963 );
nand U1270 ( n1965, my_IIR_filter_firBlock_left_multProducts[12], n1964 );
or U1271 ( n1964, n1963, my_IIR_filter_firBlock_left_firStep[140] );
nand U1272 ( n1831, n1830, n1829 );
nand U1273 ( n1830, my_IIR_filter_firBlock_left_firStep[172], n1827 );
nand U1274 ( n1829, my_IIR_filter_firBlock_left_multProducts[12], n1828 );
or U1275 ( n1828, n1827, my_IIR_filter_firBlock_left_firStep[172] );
nand U1276 ( n1958, n1957, n1956 );
nand U1277 ( n1957, my_IIR_filter_firBlock_left_firStep[138], n1954 );
nand U1278 ( n1956, my_IIR_filter_firBlock_left_multProducts[10], n1955 );
or U1279 ( n1955, n1954, my_IIR_filter_firBlock_left_firStep[138] );
nand U1280 ( n1822, n1821, n1820 );
nand U1281 ( n1821, my_IIR_filter_firBlock_left_firStep[170], n1818 );
nand U1282 ( n1820, my_IIR_filter_firBlock_left_multProducts[10], n1819 );
or U1283 ( n1819, n1818, my_IIR_filter_firBlock_left_firStep[170] );
nand U1284 ( n2063, n1949, n1948 );
nand U1285 ( n1949, my_IIR_filter_firBlock_left_firStep[136], n2062 );
nand U1286 ( n1948, my_IIR_filter_firBlock_left_multProducts[8], n1947 );
or U1287 ( n1947, n2062, my_IIR_filter_firBlock_left_firStep[136] );
nand U1288 ( n1925, n1813, n1812 );
nand U1289 ( n1813, my_IIR_filter_firBlock_left_firStep[168], n1924 );
nand U1290 ( n1812, my_IIR_filter_firBlock_left_multProducts[8], n1811 );
or U1291 ( n1811, n1924, my_IIR_filter_firBlock_left_firStep[168] );
nand U1292 ( n2060, n1943, n1942 );
nand U1293 ( n1943, my_IIR_filter_firBlock_left_firStep[134], n2059 );
nand U1294 ( n1942, my_IIR_filter_firBlock_left_multProducts[6], n1941 );
or U1295 ( n1941, n2059, my_IIR_filter_firBlock_left_firStep[134] );
nand U1296 ( n1922, n1807, n1806 );
nand U1297 ( n1807, my_IIR_filter_firBlock_left_firStep[166], n1921 );
nand U1298 ( n1806, my_IIR_filter_firBlock_left_multProducts[6], n1805 );
or U1299 ( n1805, n1921, my_IIR_filter_firBlock_left_firStep[166] );
nand U1300 ( n2057, n1937, n1936 );
nand U1301 ( n1937, my_IIR_filter_firBlock_left_firStep[132], n2056 );
nand U1302 ( n1936, my_IIR_filter_firBlock_left_multProducts[4], n1935 );
or U1303 ( n1935, n2056, my_IIR_filter_firBlock_left_firStep[132] );
nand U1304 ( n1919, n1801, n1800 );
nand U1305 ( n1801, my_IIR_filter_firBlock_left_firStep[164], n1918 );
nand U1306 ( n1800, my_IIR_filter_firBlock_left_multProducts[4], n1799 );
or U1307 ( n1799, n1918, my_IIR_filter_firBlock_left_firStep[164] );
nand U1308 ( n2054, n1931, n1930 );
nand U1309 ( n1931, my_IIR_filter_firBlock_left_firStep[130], n2042 );
nand U1310 ( n1930, my_IIR_filter_firBlock_left_multProducts[2], n1929 );
or U1311 ( n1929, n2042, my_IIR_filter_firBlock_left_firStep[130] );
nand U1312 ( n1916, n1795, n1794 );
nand U1313 ( n1795, my_IIR_filter_firBlock_left_firStep[162], n1906 );
nand U1314 ( n1794, my_IIR_filter_firBlock_left_multProducts[2], n1793 );
or U1315 ( n1793, n1906, my_IIR_filter_firBlock_left_firStep[162] );
nand U1316 ( n2037, n2035, n2034 );
nand U1317 ( n2035, my_IIR_filter_firBlock_left_firStep[155], n2032 );
nand U1318 ( n2034, my_IIR_filter_firBlock_left_multProducts[27], n2033 );
or U1319 ( n2033, n2032, my_IIR_filter_firBlock_left_firStep[155] );
nand U1320 ( n1901, n1899, n1898 );
nand U1321 ( n1899, my_IIR_filter_firBlock_left_firStep[187], n1896 );
nand U1322 ( n1898, my_IIR_filter_firBlock_left_multProducts[27], n1897 );
or U1323 ( n1897, n1896, my_IIR_filter_firBlock_left_firStep[187] );
nand U1324 ( n2028, n2026, n2025 );
nand U1325 ( n2026, my_IIR_filter_firBlock_left_firStep[153], n2023 );
nand U1326 ( n2025, my_IIR_filter_firBlock_left_multProducts[25], n2024 );
or U1327 ( n2024, n2023, my_IIR_filter_firBlock_left_firStep[153] );
nand U1328 ( n1892, n1890, n1889 );
nand U1329 ( n1890, my_IIR_filter_firBlock_left_firStep[185], n1887 );
nand U1330 ( n1889, my_IIR_filter_firBlock_left_multProducts[25], n1888 );
or U1331 ( n1888, n1887, my_IIR_filter_firBlock_left_firStep[185] );
nand U1332 ( n2019, n2017, n2016 );
nand U1333 ( n2017, my_IIR_filter_firBlock_left_firStep[151], n2014 );
nand U1334 ( n2016, my_IIR_filter_firBlock_left_multProducts[23], n2015 );
or U1335 ( n2015, n2014, my_IIR_filter_firBlock_left_firStep[151] );
nand U1336 ( n1883, n1881, n1880 );
nand U1337 ( n1881, my_IIR_filter_firBlock_left_firStep[183], n1878 );
nand U1338 ( n1880, my_IIR_filter_firBlock_left_multProducts[23], n1879 );
or U1339 ( n1879, n1878, my_IIR_filter_firBlock_left_firStep[183] );
nand U1340 ( n1990, n1988, n1987 );
nand U1341 ( n1988, my_IIR_filter_firBlock_left_firStep[145], n1985 );
nand U1342 ( n1987, my_IIR_filter_firBlock_left_multProducts[17], n1986 );
or U1343 ( n1986, n1985, my_IIR_filter_firBlock_left_firStep[145] );
nand U1344 ( n1854, n1852, n1851 );
nand U1345 ( n1852, my_IIR_filter_firBlock_left_firStep[177], n1849 );
nand U1346 ( n1851, my_IIR_filter_firBlock_left_multProducts[17], n1850 );
or U1347 ( n1850, n1849, my_IIR_filter_firBlock_left_firStep[177] );
nand U1348 ( n1981, n1979, n1978 );
nand U1349 ( n1979, my_IIR_filter_firBlock_left_firStep[143], n1976 );
nand U1350 ( n1978, my_IIR_filter_firBlock_left_multProducts[15], n1977 );
or U1351 ( n1977, n1976, my_IIR_filter_firBlock_left_firStep[143] );
nand U1352 ( n1845, n1843, n1842 );
nand U1353 ( n1843, my_IIR_filter_firBlock_left_firStep[175], n1840 );
nand U1354 ( n1842, my_IIR_filter_firBlock_left_multProducts[15], n1841 );
or U1355 ( n1841, n1840, my_IIR_filter_firBlock_left_firStep[175] );
nand U1356 ( n1972, n1970, n1969 );
nand U1357 ( n1970, my_IIR_filter_firBlock_left_firStep[141], n1967 );
nand U1358 ( n1969, my_IIR_filter_firBlock_left_multProducts[13], n1968 );
or U1359 ( n1968, n1967, my_IIR_filter_firBlock_left_firStep[141] );
nand U1360 ( n1836, n1834, n1833 );
nand U1361 ( n1834, my_IIR_filter_firBlock_left_firStep[173], n1831 );
nand U1362 ( n1833, my_IIR_filter_firBlock_left_multProducts[13], n1832 );
or U1363 ( n1832, n1831, my_IIR_filter_firBlock_left_firStep[173] );
nand U1364 ( n1963, n1961, n1960 );
nand U1365 ( n1961, my_IIR_filter_firBlock_left_firStep[139], n1958 );
nand U1366 ( n1960, my_IIR_filter_firBlock_left_multProducts[11], n1959 );
or U1367 ( n1959, n1958, my_IIR_filter_firBlock_left_firStep[139] );
nand U1368 ( n1827, n1825, n1824 );
nand U1369 ( n1825, my_IIR_filter_firBlock_left_firStep[171], n1822 );
nand U1370 ( n1824, my_IIR_filter_firBlock_left_multProducts[11], n1823 );
or U1371 ( n1823, n1822, my_IIR_filter_firBlock_left_firStep[171] );
nand U1372 ( n1954, n1952, n1951 );
nand U1373 ( n1952, my_IIR_filter_firBlock_left_firStep[137], n2063 );
nand U1374 ( n1951, my_IIR_filter_firBlock_left_multProducts[9], n1950 );
or U1375 ( n1950, n2063, my_IIR_filter_firBlock_left_firStep[137] );
nand U1376 ( n1818, n1816, n1815 );
nand U1377 ( n1816, my_IIR_filter_firBlock_left_firStep[169], n1925 );
nand U1378 ( n1815, my_IIR_filter_firBlock_left_multProducts[9], n1814 );
or U1379 ( n1814, n1925, my_IIR_filter_firBlock_left_firStep[169] );
nand U1380 ( n2062, n1946, n1945 );
nand U1381 ( n1946, my_IIR_filter_firBlock_left_firStep[135], n2060 );
nand U1382 ( n1945, my_IIR_filter_firBlock_left_multProducts[7], n1944 );
or U1383 ( n1944, n2060, my_IIR_filter_firBlock_left_firStep[135] );
nand U1384 ( n1924, n1810, n1809 );
nand U1385 ( n1810, my_IIR_filter_firBlock_left_firStep[167], n1922 );
nand U1386 ( n1809, my_IIR_filter_firBlock_left_multProducts[7], n1808 );
or U1387 ( n1808, n1922, my_IIR_filter_firBlock_left_firStep[167] );
nand U1388 ( n2059, n1940, n1939 );
nand U1389 ( n1940, my_IIR_filter_firBlock_left_firStep[133], n2057 );
nand U1390 ( n1939, my_IIR_filter_firBlock_left_multProducts[5], n1938 );
or U1391 ( n1938, n2057, my_IIR_filter_firBlock_left_firStep[133] );
nand U1392 ( n1921, n1804, n1803 );
nand U1393 ( n1804, my_IIR_filter_firBlock_left_firStep[165], n1919 );
nand U1394 ( n1803, my_IIR_filter_firBlock_left_multProducts[5], n1802 );
or U1395 ( n1802, n1919, my_IIR_filter_firBlock_left_firStep[165] );
nand U1396 ( n2056, n1934, n1933 );
nand U1397 ( n1934, my_IIR_filter_firBlock_left_firStep[131], n2054 );
nand U1398 ( n1933, my_IIR_filter_firBlock_left_multProducts[3], n1932 );
or U1399 ( n1932, n2054, my_IIR_filter_firBlock_left_firStep[131] );
nand U1400 ( n1918, n1798, n1797 );
nand U1401 ( n1798, my_IIR_filter_firBlock_left_firStep[163], n1916 );
nand U1402 ( n1797, my_IIR_filter_firBlock_left_multProducts[3], n1796 );
or U1403 ( n1796, n1916, my_IIR_filter_firBlock_left_firStep[163] );
nand U1404 ( n1787, n1637, n1636 );
nand U1405 ( n1637, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[7], n1634 );
or U1406 ( n1636, my_IIR_filter_firBlock_left_multProducts[91], n1635 );
nor U1407 ( n1635, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[7], n1634 );
xor U1408 ( my_IIR_filter_firBlock_left_N160, n2053, n2052 );
xnor U1409 ( n2053, n246, my_IIR_filter_firBlock_left_firStep[159] );
nor U1410 ( n2052, n2051, n2050 );
and U1411 ( n2050, n2049, my_IIR_filter_firBlock_left_firStep[158] );
xor U1412 ( my_IIR_filter_firBlock_left_N128, n1915, n1914 );
xnor U1413 ( n1915, n246, my_IIR_filter_firBlock_left_firStep[191] );
nor U1414 ( n1914, n1913, n1912 );
and U1415 ( n1912, n1911, my_IIR_filter_firBlock_left_firStep[190] );
nor U1416 ( n2051, n2048, n243 );
nor U1417 ( n2048, my_IIR_filter_firBlock_left_firStep[158], n2049 );
nor U1418 ( n1913, n1910, n243 );
nor U1419 ( n1910, my_IIR_filter_firBlock_left_firStep[190], n1911 );
nand U1420 ( n1996, n1993, n1992 );
nand U1421 ( n1993, my_IIR_filter_firBlock_left_firStep[146], n1990 );
nand U1422 ( n1992, my_IIR_filter_firBlock_left_multProducts[18], n1991 );
or U1423 ( n1991, n1990, my_IIR_filter_firBlock_left_firStep[146] );
nand U1424 ( n1860, n1857, n1856 );
nand U1425 ( n1857, my_IIR_filter_firBlock_left_firStep[178], n1854 );
nand U1426 ( n1856, my_IIR_filter_firBlock_left_multProducts[18], n1855 );
or U1427 ( n1855, n1854, my_IIR_filter_firBlock_left_firStep[178] );
nand U1428 ( n2042, n1928, n1927 );
nand U1429 ( n1928, my_IIR_filter_firBlock_left_firStep[129], n1995 );
nand U1430 ( n1927, my_IIR_filter_firBlock_left_multProducts[1], n1926 );
or U1431 ( n1926, my_IIR_filter_firBlock_left_firStep[129], n1995 );
nand U1432 ( n1906, n1792, n1791 );
nand U1433 ( n1792, my_IIR_filter_firBlock_left_firStep[161], n1859 );
nand U1434 ( n1791, my_IIR_filter_firBlock_left_multProducts[1], n1790 );
or U1435 ( n1790, my_IIR_filter_firBlock_left_firStep[161], n1859 );
nand U1436 ( n1631, n1627, n1626 );
nor U1437 ( n1626, inData_in[5], inData_in[4] );
nor U1438 ( n1627, inData_in[3], inData_in[2] );
nor U1439 ( n1633, n1631, n1630 );
nand U1440 ( n1630, n1629, n1628 );
nand U1441 ( n2005, n2004, n2003 );
nand U1442 ( n2004, my_IIR_filter_firBlock_left_firStep[148], n2001 );
nand U1443 ( n2003, my_IIR_filter_firBlock_left_multProducts[20], n2002 );
or U1444 ( n2002, n2001, my_IIR_filter_firBlock_left_firStep[148] );
nand U1445 ( n1869, n1868, n1867 );
nand U1446 ( n1868, my_IIR_filter_firBlock_left_firStep[180], n1865 );
nand U1447 ( n1867, my_IIR_filter_firBlock_left_multProducts[20], n1866 );
or U1448 ( n1866, n1865, my_IIR_filter_firBlock_left_firStep[180] );
nand U1449 ( n2010, n2008, n2007 );
nand U1450 ( n2008, my_IIR_filter_firBlock_left_firStep[149], n2005 );
nand U1451 ( n2007, my_IIR_filter_firBlock_left_multProducts[21], n2006 );
or U1452 ( n2006, n2005, my_IIR_filter_firBlock_left_firStep[149] );
nand U1453 ( n1874, n1872, n1871 );
nand U1454 ( n1872, my_IIR_filter_firBlock_left_firStep[181], n1869 );
nand U1455 ( n1871, my_IIR_filter_firBlock_left_multProducts[21], n1870 );
or U1456 ( n1870, n1869, my_IIR_filter_firBlock_left_firStep[181] );
nand U1457 ( n2001, n1999, n1998 );
nand U1458 ( n1999, my_IIR_filter_firBlock_left_firStep[147], n1996 );
nand U1459 ( n1998, my_IIR_filter_firBlock_left_multProducts[19], n1997 );
or U1460 ( n1997, n1996, my_IIR_filter_firBlock_left_firStep[147] );
nand U1461 ( n1865, n1863, n1862 );
nand U1462 ( n1863, my_IIR_filter_firBlock_left_firStep[179], n1860 );
nand U1463 ( n1862, my_IIR_filter_firBlock_left_multProducts[19], n1861 );
or U1464 ( n1861, n1860, my_IIR_filter_firBlock_left_firStep[179] );
xor U1465 ( n864, n298, my_IIR_filter_firBlock_left_multProducts[102] );
xnor U1466 ( outData_in[16], n750, n280 );
xnor U1467 ( n280, rightOut[16], leftOut[16] );
xnor U1468 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10_39, n281, n800 );
xor U1469 ( n281, rightOut[31], leftOut[31] );
xor U1470 ( outData_in[19], n282, n761 );
xor U1471 ( n282, leftOut[19], rightOut[19] );
nand U1472 ( n2436, n2435, n2434 );
nand U1473 ( n2435, my_IIR_filter_firBlock_left_firStep[56], n2432 );
nand U1474 ( n2432, n2430, n2429 );
xnor U1475 ( outData_in[18], n756, n283 );
xnor U1476 ( n283, rightOut[18], leftOut[18] );
xor U1477 ( outData_in[25], n284, n781 );
xor U1478 ( n284, leftOut[25], rightOut[25] );
nand U1479 ( n2427, n2426, n2425 );
nand U1480 ( n2418, n2417, n2416 );
nand U1481 ( n2417, my_IIR_filter_firBlock_left_firStep[52], n2414 );
nand U1482 ( n2423, n2421, n2420 );
nand U1483 ( n2420, my_IIR_filter_firBlock_left_multProducts[82], n2419 );
nand U1484 ( n2414, n2412, n2411 );
nand U1485 ( n2409, n2406, n2405 );
nand U1486 ( n2406, my_IIR_filter_firBlock_left_firStep[50], n2403 );
nand U1487 ( n2405, my_IIR_filter_firBlock_left_multProducts[79], n2404 );
or U1488 ( n2404, n2403, my_IIR_filter_firBlock_left_firStep[50] );
nand U1489 ( n2398, n2397, n2396 );
nand U1490 ( n2397, my_IIR_filter_firBlock_left_firStep[48], n2394 );
nand U1491 ( n2359, my_IIR_filter_firBlock_left_firStep[39], n2472 );
nand U1492 ( n2466, n2344, n2343 );
nand U1493 ( n2344, my_IIR_filter_firBlock_left_firStep[34], n2455 );
nand U1494 ( n2343, my_IIR_filter_firBlock_left_multProducts[63], n2342 );
or U1495 ( n2342, n2455, my_IIR_filter_firBlock_left_firStep[34] );
nand U1496 ( n2469, n2350, n2349 );
nand U1497 ( n2350, my_IIR_filter_firBlock_left_firStep[36], n2468 );
or U1498 ( n2348, n2468, my_IIR_filter_firBlock_left_firStep[36] );
nand U1499 ( n2468, n2347, n2346 );
nand U1500 ( n2347, my_IIR_filter_firBlock_left_firStep[35], n2466 );
or U1501 ( n2345, n2466, my_IIR_filter_firBlock_left_firStep[35] );
nand U1502 ( n2471, n2353, n2352 );
nand U1503 ( n2353, my_IIR_filter_firBlock_left_firStep[37], n2469 );
or U1504 ( n2351, n2469, my_IIR_filter_firBlock_left_firStep[37] );
nand U1505 ( n2385, n2383, n2382 );
nand U1506 ( n2472, n2356, n2355 );
nand U1507 ( n2356, my_IIR_filter_firBlock_left_firStep[38], n2471 );
nand U1508 ( n2355, my_IIR_filter_firBlock_left_multProducts[67], n2354 );
or U1509 ( n2354, n2471, my_IIR_filter_firBlock_left_firStep[38] );
nand U1510 ( n2376, n2374, n2373 );
nand U1511 ( n2475, n2362, n2361 );
nand U1512 ( n2362, my_IIR_filter_firBlock_left_firStep[40], n2474 );
or U1513 ( n2360, n2474, my_IIR_filter_firBlock_left_firStep[40] );
nand U1514 ( n2380, n2379, n2378 );
nand U1515 ( n2371, n2370, n2369 );
nand U1516 ( n2370, my_IIR_filter_firBlock_left_firStep[42], n2367 );
nand U1517 ( n2369, my_IIR_filter_firBlock_left_multProducts[71], n2368 );
or U1518 ( n2368, n2367, my_IIR_filter_firBlock_left_firStep[42] );
nand U1519 ( n2394, n2392, n2391 );
nand U1520 ( n2391, my_IIR_filter_firBlock_left_multProducts[76], n2390 );
nand U1521 ( n2389, n2388, n2387 );
nand U1522 ( n2388, my_IIR_filter_firBlock_left_firStep[46], n2385 );
nand U1523 ( n2387, my_IIR_filter_firBlock_left_multProducts[75], n2386 );
or U1524 ( n2386, n2385, my_IIR_filter_firBlock_left_firStep[46] );
nand U1525 ( n2455, n2341, n2340 );
nand U1526 ( n2341, my_IIR_filter_firBlock_left_firStep[33], n2408 );
or U1527 ( n2339, my_IIR_filter_firBlock_left_firStep[33], n2408 );
xor U1528 ( n743, rightOut[14], leftOut[14] );
and U1529 ( n3290, my_IIR_filter_firBlock_right_multProducts[31], my_IIR_filter_firBlock_right_firStep[31] );
xor U1530 ( n770, rightOut[22], leftOut[22] );
xor U1531 ( my_IIR_filter_firBlock_left_multProducts[0], n1787, n285 );
xnor U1532 ( n285, my_IIR_filter_firBlock_left_multProducts[92], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[8] );
and U1533 ( n1995, my_IIR_filter_firBlock_left_multProducts[0], my_IIR_filter_firBlock_left_firStep[128] );
and U1534 ( n1859, my_IIR_filter_firBlock_left_multProducts[0], my_IIR_filter_firBlock_left_firStep[160] );
xor U1535 ( outData_in[17], n286, n753 );
xor U1536 ( n286, leftOut[17], rightOut[17] );
xor U1537 ( outData_in[15], n287, n747 );
xor U1538 ( n287, leftOut[15], rightOut[15] );
xor U1539 ( outData_in[27], n288, n787 );
xor U1540 ( n288, leftOut[27], rightOut[27] );
xor U1541 ( outData_in[29], n289, n793 );
xor U1542 ( n289, leftOut[29], rightOut[29] );
xnor U1543 ( my_IIR_filter_firBlock_right_N191, n3529, n290 );
xor U1544 ( n290, n215, my_IIR_filter_firBlock_right_firStep[30] );
xor U1545 ( my_IIR_filter_firBlock_right_N126, n291, n3337 );
xor U1546 ( n291, my_IIR_filter_firBlock_right_firStep[60], my_IIR_filter_firBlock_right_multProducts[60] );
xnor U1547 ( my_IIR_filter_firBlock_left_N255, n2461, n292 );
xor U1548 ( n292, n631, my_IIR_filter_firBlock_left_firStep[62] );
nand U1549 ( n2793, n2790, n2789 );
nand U1550 ( n2790, my_IIR_filter_firBlock_right_firStep[91], n2787 );
nand U1551 ( n2789, my_IIR_filter_firBlock_right_multProducts[91], n2788 );
or U1552 ( n2788, n2787, my_IIR_filter_firBlock_right_firStep[91] );
nand U1553 ( n2804, n2687, n2686 );
nand U1554 ( n2687, my_IIR_filter_firBlock_right_firStep[68], n2803 );
nand U1555 ( n2686, my_IIR_filter_firBlock_right_multProducts[68], n2685 );
or U1556 ( n2685, n2803, my_IIR_filter_firBlock_right_firStep[68] );
nand U1557 ( n2729, n2728, n2727 );
nand U1558 ( n2728, my_IIR_filter_firBlock_right_firStep[78], n2725 );
nand U1559 ( n2727, my_IIR_filter_firBlock_right_multProducts[78], n2726 );
or U1560 ( n2726, n2725, my_IIR_filter_firBlock_right_firStep[78] );
nand U1561 ( n2801, n2681, n2680 );
nand U1562 ( n2681, my_IIR_filter_firBlock_right_firStep[66], n2800 );
nand U1563 ( n2680, my_IIR_filter_firBlock_right_multProducts[66], n2679 );
or U1564 ( n2679, n2800, my_IIR_filter_firBlock_right_firStep[66] );
nand U1565 ( n2758, n2757, n2756 );
nand U1566 ( n2757, my_IIR_filter_firBlock_right_firStep[84], n2754 );
nand U1567 ( n2756, my_IIR_filter_firBlock_right_multProducts[84], n2755 );
or U1568 ( n2755, n2754, my_IIR_filter_firBlock_right_firStep[84] );
nand U1569 ( n2798, n2675, n2674 );
nand U1570 ( n2675, my_IIR_filter_firBlock_right_firStep[64], n2786 );
nand U1571 ( n2674, my_IIR_filter_firBlock_right_multProducts[64], n2673 );
or U1572 ( n2673, n2786, my_IIR_filter_firBlock_right_firStep[64] );
nand U1573 ( n2711, n2710, n2709 );
nand U1574 ( n2710, my_IIR_filter_firBlock_right_firStep[74], n2707 );
nand U1575 ( n2709, my_IIR_filter_firBlock_right_multProducts[74], n2708 );
or U1576 ( n2708, n2707, my_IIR_filter_firBlock_right_firStep[74] );
nand U1577 ( n2702, n2701, n2700 );
nand U1578 ( n2701, my_IIR_filter_firBlock_right_firStep[72], n2698 );
nand U1579 ( n2700, my_IIR_filter_firBlock_right_multProducts[72], n2699 );
or U1580 ( n2699, n2698, my_IIR_filter_firBlock_right_firStep[72] );
nand U1581 ( n2720, n2719, n2718 );
nand U1582 ( n2719, my_IIR_filter_firBlock_right_firStep[76], n2716 );
nand U1583 ( n2718, my_IIR_filter_firBlock_right_multProducts[76], n2717 );
or U1584 ( n2717, n2716, my_IIR_filter_firBlock_right_firStep[76] );
nand U1585 ( n2749, n2748, n2747 );
nand U1586 ( n2748, my_IIR_filter_firBlock_right_firStep[82], n2745 );
nand U1587 ( n2747, my_IIR_filter_firBlock_right_multProducts[82], n2746 );
or U1588 ( n2746, n2745, my_IIR_filter_firBlock_right_firStep[82] );
nand U1589 ( n2767, n2766, n2765 );
nand U1590 ( n2766, my_IIR_filter_firBlock_right_firStep[86], n2763 );
nand U1591 ( n2765, my_IIR_filter_firBlock_right_multProducts[86], n2764 );
or U1592 ( n2764, n2763, my_IIR_filter_firBlock_right_firStep[86] );
nand U1593 ( n2776, n2775, n2774 );
nand U1594 ( n2775, my_IIR_filter_firBlock_right_firStep[88], n2772 );
nand U1595 ( n2774, my_IIR_filter_firBlock_right_multProducts[88], n2773 );
or U1596 ( n2773, n2772, my_IIR_filter_firBlock_right_firStep[88] );
nand U1597 ( n2740, n2737, n2736 );
nand U1598 ( n2737, my_IIR_filter_firBlock_right_firStep[80], n2734 );
nand U1599 ( n2736, my_IIR_filter_firBlock_right_multProducts[80], n2735 );
or U1600 ( n2735, n2734, my_IIR_filter_firBlock_right_firStep[80] );
nand U1601 ( n2807, n2693, n2692 );
nand U1602 ( n2693, my_IIR_filter_firBlock_right_firStep[70], n2806 );
nand U1603 ( n2692, my_IIR_filter_firBlock_right_multProducts[70], n2691 );
or U1604 ( n2691, n2806, my_IIR_filter_firBlock_right_firStep[70] );
nand U1605 ( n2787, n2784, n2783 );
nand U1606 ( n2784, my_IIR_filter_firBlock_right_firStep[90], n2781 );
nand U1607 ( n2783, my_IIR_filter_firBlock_right_multProducts[90], n2782 );
or U1608 ( n2782, n2781, my_IIR_filter_firBlock_right_firStep[90] );
nand U1609 ( n2803, n2684, n2683 );
nand U1610 ( n2684, my_IIR_filter_firBlock_right_firStep[67], n2801 );
nand U1611 ( n2683, my_IIR_filter_firBlock_right_multProducts[67], n2682 );
or U1612 ( n2682, n2801, my_IIR_filter_firBlock_right_firStep[67] );
nand U1613 ( n2725, n2723, n2722 );
nand U1614 ( n2723, my_IIR_filter_firBlock_right_firStep[77], n2720 );
nand U1615 ( n2722, my_IIR_filter_firBlock_right_multProducts[77], n2721 );
or U1616 ( n2721, n2720, my_IIR_filter_firBlock_right_firStep[77] );
nand U1617 ( n2745, n2743, n2742 );
nand U1618 ( n2743, my_IIR_filter_firBlock_right_firStep[81], n2740 );
nand U1619 ( n2742, my_IIR_filter_firBlock_right_multProducts[81], n2741 );
or U1620 ( n2741, n2740, my_IIR_filter_firBlock_right_firStep[81] );
nand U1621 ( n2763, n2761, n2760 );
nand U1622 ( n2761, my_IIR_filter_firBlock_right_firStep[85], n2758 );
nand U1623 ( n2760, my_IIR_filter_firBlock_right_multProducts[85], n2759 );
or U1624 ( n2759, n2758, my_IIR_filter_firBlock_right_firStep[85] );
nand U1625 ( n2772, n2770, n2769 );
nand U1626 ( n2770, my_IIR_filter_firBlock_right_firStep[87], n2767 );
nand U1627 ( n2769, my_IIR_filter_firBlock_right_multProducts[87], n2768 );
or U1628 ( n2768, n2767, my_IIR_filter_firBlock_right_firStep[87] );
nand U1629 ( n2781, n2779, n2778 );
nand U1630 ( n2779, my_IIR_filter_firBlock_right_firStep[89], n2776 );
nand U1631 ( n2778, my_IIR_filter_firBlock_right_multProducts[89], n2777 );
or U1632 ( n2777, n2776, my_IIR_filter_firBlock_right_firStep[89] );
nand U1633 ( n2800, n2678, n2677 );
nand U1634 ( n2678, my_IIR_filter_firBlock_right_firStep[65], n2798 );
nand U1635 ( n2677, my_IIR_filter_firBlock_right_multProducts[65], n2676 );
or U1636 ( n2676, n2798, my_IIR_filter_firBlock_right_firStep[65] );
nand U1637 ( n2716, n2714, n2713 );
nand U1638 ( n2714, my_IIR_filter_firBlock_right_firStep[75], n2711 );
nand U1639 ( n2713, my_IIR_filter_firBlock_right_multProducts[75], n2712 );
or U1640 ( n2712, n2711, my_IIR_filter_firBlock_right_firStep[75] );
nand U1641 ( n2734, n2732, n2731 );
nand U1642 ( n2732, my_IIR_filter_firBlock_right_firStep[79], n2729 );
nand U1643 ( n2731, my_IIR_filter_firBlock_right_multProducts[79], n2730 );
or U1644 ( n2730, n2729, my_IIR_filter_firBlock_right_firStep[79] );
nand U1645 ( n2707, n2705, n2704 );
nand U1646 ( n2705, my_IIR_filter_firBlock_right_firStep[73], n2702 );
nand U1647 ( n2704, my_IIR_filter_firBlock_right_multProducts[73], n2703 );
or U1648 ( n2703, n2702, my_IIR_filter_firBlock_right_firStep[73] );
nand U1649 ( n2806, n2690, n2689 );
nand U1650 ( n2690, my_IIR_filter_firBlock_right_firStep[69], n2804 );
nand U1651 ( n2689, my_IIR_filter_firBlock_right_multProducts[69], n2688 );
or U1652 ( n2688, n2804, my_IIR_filter_firBlock_right_firStep[69] );
nand U1653 ( n2786, n2672, n2671 );
nand U1654 ( n2672, my_IIR_filter_firBlock_right_firStep[63], n2739 );
nand U1655 ( n2671, my_IIR_filter_firBlock_right_multProducts[63], n2670 );
or U1656 ( n2670, my_IIR_filter_firBlock_right_firStep[63], n2739 );
nand U1657 ( n2698, n2696, n2695 );
nand U1658 ( n2696, my_IIR_filter_firBlock_right_firStep[71], n2807 );
nand U1659 ( n2695, my_IIR_filter_firBlock_right_multProducts[71], n2694 );
or U1660 ( n2694, n2807, my_IIR_filter_firBlock_right_firStep[71] );
nor U1661 ( n2795, n2792, n632 );
nor U1662 ( n2792, my_IIR_filter_firBlock_right_firStep[92], n2793 );
xor U1663 ( my_IIR_filter_firBlock_right_N64, n2797, n2796 );
xnor U1664 ( n2797, my_IIR_filter_firBlock_right_multProducts[91], my_IIR_filter_firBlock_right_firStep[93] );
nor U1665 ( n2796, n2795, n2794 );
and U1666 ( n2794, n2793, my_IIR_filter_firBlock_right_firStep[92] );
nand U1667 ( n2754, n2752, n2751 );
nand U1668 ( n2752, my_IIR_filter_firBlock_right_firStep[83], n2749 );
nand U1669 ( n2751, my_IIR_filter_firBlock_right_multProducts[83], n2750 );
or U1670 ( n2750, n2749, my_IIR_filter_firBlock_right_firStep[83] );
xnor U1671 ( my_IIR_filter_firBlock_left_N31, n1207, n293 );
xor U1672 ( n293, n631, my_IIR_filter_firBlock_left_firStep[286] );
nand U1673 ( n1347, n1227, n1226 );
nand U1674 ( n1227, my_IIR_filter_firBlock_left_multProducts[90], n1346 );
nand U1675 ( n1226, inData_in[2], n1225 );
or U1676 ( n1225, n1346, my_IIR_filter_firBlock_left_multProducts[90] );
nand U1677 ( n1242, n1241, n1240 );
nand U1678 ( n1241, my_IIR_filter_firBlock_left_multProducts[90], n1238 );
nand U1679 ( n1240, my_IIR_filter_firBlock_left_multProducts[94], n1239 );
or U1680 ( n1239, n1238, my_IIR_filter_firBlock_left_multProducts[90] );
or U1681 ( n1256, n294, n295 );
nor U1682 ( n295, n1255, my_IIR_filter_firBlock_left_multProducts[94] );
or U1683 ( n1270, n296, n297 );
nor U1684 ( n297, n1269, my_IIR_filter_firBlock_left_multProducts[98] );
or U1685 ( n1263, n298, n299 );
nor U1686 ( n299, n1262, my_IIR_filter_firBlock_left_multProducts[96] );
nand U1687 ( n1280, n1279, n1278 );
nand U1688 ( n1279, my_IIR_filter_firBlock_left_multProducts[100], n1276 );
nand U1689 ( n1278, my_IIR_filter_firBlock_left_multProducts[104], n1277 );
or U1690 ( n1277, n1276, my_IIR_filter_firBlock_left_multProducts[100] );
nand U1691 ( n1251, n1250, n1249 );
nand U1692 ( n1250, my_IIR_filter_firBlock_left_multProducts[92], n1247 );
nand U1693 ( n1249, my_IIR_filter_firBlock_left_multProducts[96], n1248 );
or U1694 ( n1248, n1247, my_IIR_filter_firBlock_left_multProducts[92] );
nand U1695 ( n1350, n1233, n1232 );
nand U1696 ( n1233, my_IIR_filter_firBlock_left_multProducts[92], n1349 );
nand U1697 ( n1232, inData_in[4], n1231 );
or U1698 ( n1231, n1349, my_IIR_filter_firBlock_left_multProducts[92] );
nand U1699 ( n1349, n1230, n1229 );
nand U1700 ( n1230, my_IIR_filter_firBlock_left_multProducts[91], n1347 );
nand U1701 ( n1229, inData_in[3], n1228 );
or U1702 ( n1228, n1347, my_IIR_filter_firBlock_left_multProducts[91] );
nand U1703 ( n1247, n1245, n1244 );
nand U1704 ( n1245, my_IIR_filter_firBlock_left_multProducts[91], n1242 );
nand U1705 ( n1244, my_IIR_filter_firBlock_left_multProducts[95], n1243 );
or U1706 ( n1243, n1242, my_IIR_filter_firBlock_left_multProducts[91] );
or U1707 ( n1266, n300, n301 );
nor U1708 ( n301, n1265, my_IIR_filter_firBlock_left_multProducts[97] );
or U1709 ( n1259, n302, n303 );
nor U1710 ( n303, n1258, my_IIR_filter_firBlock_left_multProducts[95] );
or U1711 ( n1273, n304, n305 );
nor U1712 ( n305, n1272, my_IIR_filter_firBlock_left_multProducts[99] );
or U1713 ( n1252, n306, n307 );
nor U1714 ( n307, n1251, my_IIR_filter_firBlock_left_multProducts[93] );
nand U1715 ( n1238, n1236, n1235 );
nand U1716 ( n1236, my_IIR_filter_firBlock_left_multProducts[93], n1350 );
nand U1717 ( n1235, inData_in[5], n1234 );
or U1718 ( n1234, n1350, my_IIR_filter_firBlock_left_multProducts[93] );
nand U1719 ( n1346, n1224, n1223 );
nand U1720 ( n1223, inData_in[5], n1222 );
nand U1721 ( n1285, n1283, n1282 );
nand U1722 ( n1283, my_IIR_filter_firBlock_left_multProducts[101], n1280 );
nand U1723 ( n1282, my_IIR_filter_firBlock_left_multProducts[105], n1281 );
or U1724 ( n1281, n1280, my_IIR_filter_firBlock_left_multProducts[101] );
nand U1725 ( n1315, n1314, n1313 );
nand U1726 ( n1314, my_IIR_filter_firBlock_left_multProducts[108], n1311 );
nand U1727 ( n1313, my_IIR_filter_firBlock_left_multProducts[112], n1312 );
or U1728 ( n1312, n1311, my_IIR_filter_firBlock_left_multProducts[108] );
nand U1729 ( n1289, n1288, n1287 );
nand U1730 ( n1288, my_IIR_filter_firBlock_left_multProducts[102], n1285 );
nand U1731 ( n1287, my_IIR_filter_firBlock_left_multProducts[106], n1286 );
or U1732 ( n1286, n1285, my_IIR_filter_firBlock_left_multProducts[102] );
nand U1733 ( n1297, n1296, n1295 );
nand U1734 ( n1296, my_IIR_filter_firBlock_left_multProducts[104], n1293 );
nand U1735 ( n1295, my_IIR_filter_firBlock_left_multProducts[108], n1294 );
or U1736 ( n1294, n1293, my_IIR_filter_firBlock_left_multProducts[104] );
nand U1737 ( n1306, n1305, n1304 );
nand U1738 ( n1305, my_IIR_filter_firBlock_left_multProducts[106], n1302 );
nand U1739 ( n1304, my_IIR_filter_firBlock_left_multProducts[110], n1303 );
or U1740 ( n1303, n1302, my_IIR_filter_firBlock_left_multProducts[106] );
nand U1741 ( n1311, n1309, n1308 );
nand U1742 ( n1309, my_IIR_filter_firBlock_left_multProducts[107], n1306 );
nand U1743 ( n1308, my_IIR_filter_firBlock_left_multProducts[111], n1307 );
or U1744 ( n1307, n1306, my_IIR_filter_firBlock_left_multProducts[107] );
or U1745 ( n1290, n308, n309 );
nor U1746 ( n309, n1289, my_IIR_filter_firBlock_left_multProducts[103] );
nand U1747 ( n1302, n1300, n1299 );
nand U1748 ( n1300, my_IIR_filter_firBlock_left_multProducts[105], n1297 );
nand U1749 ( n1299, my_IIR_filter_firBlock_left_multProducts[109], n1298 );
or U1750 ( n1298, n1297, my_IIR_filter_firBlock_left_multProducts[105] );
nand U1751 ( n1320, n1318, n1317 );
nand U1752 ( n1318, my_IIR_filter_firBlock_left_multProducts[109], n1315 );
nand U1753 ( n1317, my_IIR_filter_firBlock_left_multProducts[113], n1316 );
or U1754 ( n1316, n1315, my_IIR_filter_firBlock_left_multProducts[109] );
nand U1755 ( n1324, n1323, n1322 );
nand U1756 ( n1323, my_IIR_filter_firBlock_left_multProducts[110], n1320 );
nand U1757 ( n1322, my_IIR_filter_firBlock_left_multProducts[114], n1321 );
or U1758 ( n1321, n1320, my_IIR_filter_firBlock_left_multProducts[110] );
nand U1759 ( n1329, n1327, n1326 );
nand U1760 ( n1327, my_IIR_filter_firBlock_left_multProducts[111], n1324 );
nand U1761 ( n1326, n549, n1325 );
or U1762 ( n1325, n1324, my_IIR_filter_firBlock_left_multProducts[111] );
nand U1763 ( n1334, n1332, n1331 );
nand U1764 ( n1332, my_IIR_filter_firBlock_left_multProducts[112], n1329 );
nand U1765 ( n1331, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n1330 );
or U1766 ( n1330, n1329, my_IIR_filter_firBlock_left_multProducts[112] );
xnor U1767 ( my_IIR_filter_firBlock_left_multProducts[58], n1333, n1334 );
xnor U1768 ( n1333, my_IIR_filter_firBlock_left_multProducts[113], n549 );
nand U1769 ( n2324, n2322, n2321 );
nand U1770 ( n2322, my_IIR_filter_firBlock_left_firStep[93], n2319 );
nand U1771 ( n2321, my_IIR_filter_firBlock_left_multProducts[60], n2320 );
or U1772 ( n2320, n2319, my_IIR_filter_firBlock_left_firStep[93] );
nand U1773 ( n1473, n1471, n1470 );
nand U1774 ( n1471, my_IIR_filter_firBlock_left_firStep[253], n1468 );
nand U1775 ( n1470, my_IIR_filter_firBlock_left_multProducts[60], n1469 );
or U1776 ( n1469, n1468, my_IIR_filter_firBlock_left_firStep[253] );
nand U1777 ( n2319, n2316, n2315 );
nand U1778 ( n2316, my_IIR_filter_firBlock_left_firStep[92], n2313 );
nand U1779 ( n2315, my_IIR_filter_firBlock_left_multProducts[59], n2314 );
or U1780 ( n2314, n2313, my_IIR_filter_firBlock_left_firStep[92] );
nand U1781 ( n1468, n1465, n1464 );
nand U1782 ( n1465, my_IIR_filter_firBlock_left_firStep[252], n1462 );
nand U1783 ( n1464, my_IIR_filter_firBlock_left_multProducts[59], n1463 );
or U1784 ( n1463, n1462, my_IIR_filter_firBlock_left_firStep[252] );
nand U1785 ( n2313, n2311, n2310 );
nand U1786 ( n2311, my_IIR_filter_firBlock_left_firStep[91], n2308 );
nand U1787 ( n2310, my_IIR_filter_firBlock_left_multProducts[58], n2309 );
or U1788 ( n2309, n2308, my_IIR_filter_firBlock_left_firStep[91] );
nand U1789 ( n1462, n1460, n1459 );
nand U1790 ( n1460, my_IIR_filter_firBlock_left_firStep[251], n1457 );
nand U1791 ( n1459, my_IIR_filter_firBlock_left_multProducts[58], n1458 );
or U1792 ( n1458, n1457, my_IIR_filter_firBlock_left_firStep[251] );
xor U1793 ( my_IIR_filter_firBlock_left_N224, n2328, n2327 );
xnor U1794 ( n2328, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, my_IIR_filter_firBlock_left_firStep[95] );
nor U1795 ( n2327, n2326, n2325 );
and U1796 ( n2325, n2324, my_IIR_filter_firBlock_left_firStep[94] );
xor U1797 ( my_IIR_filter_firBlock_left_N64, n1477, n1476 );
xnor U1798 ( n1477, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, my_IIR_filter_firBlock_left_firStep[255] );
nor U1799 ( n1476, n1475, n1474 );
and U1800 ( n1474, n1473, my_IIR_filter_firBlock_left_firStep[254] );
nor U1801 ( n2326, n2323, n526 );
nor U1802 ( n2323, my_IIR_filter_firBlock_left_firStep[94], n2324 );
nor U1803 ( n1475, n1472, n526 );
nor U1804 ( n1472, my_IIR_filter_firBlock_left_firStep[254], n1473 );
nand U1805 ( n1339, n1337, n1336 );
nand U1806 ( n1337, my_IIR_filter_firBlock_left_multProducts[113], n1334 );
nand U1807 ( n1336, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n1335 );
or U1808 ( n1335, n1334, my_IIR_filter_firBlock_left_multProducts[113] );
xor U1809 ( n1338, n549, my_IIR_filter_firBlock_left_multProducts[114] );
xor U1810 ( my_IIR_filter_firBlock_left_multProducts[32], n310, n1347 );
xor U1811 ( n310, inData_in[3], my_IIR_filter_firBlock_left_multProducts[91] );
nand U1812 ( n2329, n2207, n2206 );
nand U1813 ( n2207, my_IIR_filter_firBlock_left_firStep[66], n2318 );
nand U1814 ( n2206, my_IIR_filter_firBlock_left_multProducts[33], n2205 );
or U1815 ( n2205, n2318, my_IIR_filter_firBlock_left_firStep[66] );
nand U1816 ( n1478, n1356, n1355 );
nand U1817 ( n1356, my_IIR_filter_firBlock_left_firStep[226], n1467 );
nand U1818 ( n1355, my_IIR_filter_firBlock_left_multProducts[33], n1354 );
or U1819 ( n1354, n1467, my_IIR_filter_firBlock_left_firStep[226] );
nand U1820 ( n2334, n2216, n2215 );
nand U1821 ( n2216, my_IIR_filter_firBlock_left_firStep[69], n2332 );
nand U1822 ( n2215, my_IIR_filter_firBlock_left_multProducts[36], n2214 );
or U1823 ( n2214, n2332, my_IIR_filter_firBlock_left_firStep[69] );
nand U1824 ( n1483, n1365, n1364 );
nand U1825 ( n1365, my_IIR_filter_firBlock_left_firStep[229], n1481 );
nand U1826 ( n1364, my_IIR_filter_firBlock_left_multProducts[36], n1363 );
or U1827 ( n1363, n1481, my_IIR_filter_firBlock_left_firStep[229] );
nand U1828 ( n2318, n2204, n2203 );
nand U1829 ( n2204, my_IIR_filter_firBlock_left_firStep[65], n2271 );
nand U1830 ( n2203, my_IIR_filter_firBlock_left_multProducts[32], n2202 );
or U1831 ( n2202, my_IIR_filter_firBlock_left_firStep[65], n2271 );
nand U1832 ( n1467, n1353, n1352 );
nand U1833 ( n1353, my_IIR_filter_firBlock_left_firStep[225], n1420 );
nand U1834 ( n1352, my_IIR_filter_firBlock_left_multProducts[32], n1351 );
or U1835 ( n1351, my_IIR_filter_firBlock_left_firStep[225], n1420 );
nand U1836 ( n2331, n2210, n2209 );
nand U1837 ( n2210, my_IIR_filter_firBlock_left_firStep[67], n2329 );
nand U1838 ( n2209, my_IIR_filter_firBlock_left_multProducts[34], n2208 );
or U1839 ( n2208, n2329, my_IIR_filter_firBlock_left_firStep[67] );
nand U1840 ( n1480, n1359, n1358 );
nand U1841 ( n1359, my_IIR_filter_firBlock_left_firStep[227], n1478 );
nand U1842 ( n1358, my_IIR_filter_firBlock_left_multProducts[34], n1357 );
or U1843 ( n1357, n1478, my_IIR_filter_firBlock_left_firStep[227] );
nand U1844 ( n2332, n2213, n2212 );
nand U1845 ( n2213, my_IIR_filter_firBlock_left_firStep[68], n2331 );
nand U1846 ( n2212, my_IIR_filter_firBlock_left_multProducts[35], n2211 );
or U1847 ( n2211, n2331, my_IIR_filter_firBlock_left_firStep[68] );
nand U1848 ( n1481, n1362, n1361 );
nand U1849 ( n1362, my_IIR_filter_firBlock_left_firStep[228], n1480 );
nand U1850 ( n1361, my_IIR_filter_firBlock_left_multProducts[35], n1360 );
or U1851 ( n1360, n1480, my_IIR_filter_firBlock_left_firStep[228] );
nand U1852 ( n2335, n2219, n2218 );
nand U1853 ( n2219, my_IIR_filter_firBlock_left_firStep[70], n2334 );
nand U1854 ( n2218, my_IIR_filter_firBlock_left_multProducts[37], n2217 );
or U1855 ( n2217, n2334, my_IIR_filter_firBlock_left_firStep[70] );
nand U1856 ( n1484, n1368, n1367 );
nand U1857 ( n1368, my_IIR_filter_firBlock_left_firStep[230], n1483 );
nand U1858 ( n1367, my_IIR_filter_firBlock_left_multProducts[37], n1366 );
or U1859 ( n1366, n1483, my_IIR_filter_firBlock_left_firStep[230] );
nand U1860 ( n2337, n2222, n2221 );
nand U1861 ( n2222, my_IIR_filter_firBlock_left_firStep[71], n2335 );
nand U1862 ( n2221, my_IIR_filter_firBlock_left_multProducts[38], n2220 );
or U1863 ( n2220, n2335, my_IIR_filter_firBlock_left_firStep[71] );
nand U1864 ( n1486, n1371, n1370 );
nand U1865 ( n1371, my_IIR_filter_firBlock_left_firStep[231], n1484 );
nand U1866 ( n1370, my_IIR_filter_firBlock_left_multProducts[38], n1369 );
or U1867 ( n1369, n1484, my_IIR_filter_firBlock_left_firStep[231] );
nand U1868 ( n2338, n2225, n2224 );
nand U1869 ( n2225, my_IIR_filter_firBlock_left_firStep[72], n2337 );
nand U1870 ( n2224, my_IIR_filter_firBlock_left_multProducts[39], n2223 );
or U1871 ( n2223, n2337, my_IIR_filter_firBlock_left_firStep[72] );
nand U1872 ( n1487, n1374, n1373 );
nand U1873 ( n1374, my_IIR_filter_firBlock_left_firStep[232], n1486 );
nand U1874 ( n1373, my_IIR_filter_firBlock_left_multProducts[39], n1372 );
or U1875 ( n1372, n1486, my_IIR_filter_firBlock_left_firStep[232] );
nand U1876 ( n2230, n2228, n2227 );
nand U1877 ( n2228, my_IIR_filter_firBlock_left_firStep[73], n2338 );
nand U1878 ( n2227, my_IIR_filter_firBlock_left_multProducts[40], n2226 );
or U1879 ( n2226, n2338, my_IIR_filter_firBlock_left_firStep[73] );
nand U1880 ( n1379, n1377, n1376 );
nand U1881 ( n1377, my_IIR_filter_firBlock_left_firStep[233], n1487 );
nand U1882 ( n1376, my_IIR_filter_firBlock_left_multProducts[40], n1375 );
or U1883 ( n1375, n1487, my_IIR_filter_firBlock_left_firStep[233] );
nand U1884 ( n2234, n2233, n2232 );
nand U1885 ( n2233, my_IIR_filter_firBlock_left_firStep[74], n2230 );
nand U1886 ( n2232, my_IIR_filter_firBlock_left_multProducts[41], n2231 );
or U1887 ( n2231, n2230, my_IIR_filter_firBlock_left_firStep[74] );
nand U1888 ( n1383, n1382, n1381 );
nand U1889 ( n1382, my_IIR_filter_firBlock_left_firStep[234], n1379 );
nand U1890 ( n1381, my_IIR_filter_firBlock_left_multProducts[41], n1380 );
or U1891 ( n1380, n1379, my_IIR_filter_firBlock_left_firStep[234] );
nand U1892 ( n2239, n2237, n2236 );
nand U1893 ( n2237, my_IIR_filter_firBlock_left_firStep[75], n2234 );
nand U1894 ( n2236, my_IIR_filter_firBlock_left_multProducts[42], n2235 );
or U1895 ( n2235, n2234, my_IIR_filter_firBlock_left_firStep[75] );
nand U1896 ( n1388, n1386, n1385 );
nand U1897 ( n1386, my_IIR_filter_firBlock_left_firStep[235], n1383 );
nand U1898 ( n1385, my_IIR_filter_firBlock_left_multProducts[42], n1384 );
or U1899 ( n1384, n1383, my_IIR_filter_firBlock_left_firStep[235] );
nand U1900 ( n2243, n2242, n2241 );
nand U1901 ( n2242, my_IIR_filter_firBlock_left_firStep[76], n2239 );
nand U1902 ( n2241, my_IIR_filter_firBlock_left_multProducts[43], n2240 );
or U1903 ( n2240, n2239, my_IIR_filter_firBlock_left_firStep[76] );
nand U1904 ( n1392, n1391, n1390 );
nand U1905 ( n1391, my_IIR_filter_firBlock_left_firStep[236], n1388 );
nand U1906 ( n1390, my_IIR_filter_firBlock_left_multProducts[43], n1389 );
or U1907 ( n1389, n1388, my_IIR_filter_firBlock_left_firStep[236] );
nand U1908 ( n2248, n2246, n2245 );
nand U1909 ( n2246, my_IIR_filter_firBlock_left_firStep[77], n2243 );
nand U1910 ( n2245, my_IIR_filter_firBlock_left_multProducts[44], n2244 );
or U1911 ( n2244, n2243, my_IIR_filter_firBlock_left_firStep[77] );
nand U1912 ( n1397, n1395, n1394 );
nand U1913 ( n1395, my_IIR_filter_firBlock_left_firStep[237], n1392 );
nand U1914 ( n1394, my_IIR_filter_firBlock_left_multProducts[44], n1393 );
or U1915 ( n1393, n1392, my_IIR_filter_firBlock_left_firStep[237] );
nand U1916 ( n2252, n2251, n2250 );
nand U1917 ( n2251, my_IIR_filter_firBlock_left_firStep[78], n2248 );
nand U1918 ( n2250, my_IIR_filter_firBlock_left_multProducts[45], n2249 );
or U1919 ( n2249, n2248, my_IIR_filter_firBlock_left_firStep[78] );
nand U1920 ( n1401, n1400, n1399 );
nand U1921 ( n1400, my_IIR_filter_firBlock_left_firStep[238], n1397 );
nand U1922 ( n1399, my_IIR_filter_firBlock_left_multProducts[45], n1398 );
or U1923 ( n1398, n1397, my_IIR_filter_firBlock_left_firStep[238] );
nand U1924 ( n2261, n2260, n2259 );
nand U1925 ( n2260, my_IIR_filter_firBlock_left_firStep[80], n2257 );
nand U1926 ( n2259, my_IIR_filter_firBlock_left_multProducts[47], n2258 );
or U1927 ( n2258, n2257, my_IIR_filter_firBlock_left_firStep[80] );
nand U1928 ( n1410, n1409, n1408 );
nand U1929 ( n1409, my_IIR_filter_firBlock_left_firStep[240], n1406 );
nand U1930 ( n1408, my_IIR_filter_firBlock_left_multProducts[47], n1407 );
or U1931 ( n1407, n1406, my_IIR_filter_firBlock_left_firStep[240] );
nand U1932 ( n2257, n2255, n2254 );
nand U1933 ( n2255, my_IIR_filter_firBlock_left_firStep[79], n2252 );
nand U1934 ( n2254, my_IIR_filter_firBlock_left_multProducts[46], n2253 );
or U1935 ( n2253, n2252, my_IIR_filter_firBlock_left_firStep[79] );
nand U1936 ( n1406, n1404, n1403 );
nand U1937 ( n1404, my_IIR_filter_firBlock_left_firStep[239], n1401 );
nand U1938 ( n1403, my_IIR_filter_firBlock_left_multProducts[46], n1402 );
or U1939 ( n1402, n1401, my_IIR_filter_firBlock_left_firStep[239] );
nand U1940 ( n2266, n2264, n2263 );
nand U1941 ( n2264, my_IIR_filter_firBlock_left_firStep[81], n2261 );
nand U1942 ( n2263, my_IIR_filter_firBlock_left_multProducts[48], n2262 );
or U1943 ( n2262, n2261, my_IIR_filter_firBlock_left_firStep[81] );
nand U1944 ( n1415, n1413, n1412 );
nand U1945 ( n1413, my_IIR_filter_firBlock_left_firStep[241], n1410 );
nand U1946 ( n1412, my_IIR_filter_firBlock_left_multProducts[48], n1411 );
or U1947 ( n1411, n1410, my_IIR_filter_firBlock_left_firStep[241] );
nand U1948 ( n2272, n2269, n2268 );
nand U1949 ( n2269, my_IIR_filter_firBlock_left_firStep[82], n2266 );
nand U1950 ( n2268, my_IIR_filter_firBlock_left_multProducts[49], n2267 );
or U1951 ( n2267, n2266, my_IIR_filter_firBlock_left_firStep[82] );
nand U1952 ( n1421, n1418, n1417 );
nand U1953 ( n1418, my_IIR_filter_firBlock_left_firStep[242], n1415 );
nand U1954 ( n1417, my_IIR_filter_firBlock_left_multProducts[49], n1416 );
or U1955 ( n1416, n1415, my_IIR_filter_firBlock_left_firStep[242] );
nand U1956 ( n2277, n2275, n2274 );
nand U1957 ( n2275, my_IIR_filter_firBlock_left_firStep[83], n2272 );
nand U1958 ( n2274, my_IIR_filter_firBlock_left_multProducts[50], n2273 );
or U1959 ( n2273, n2272, my_IIR_filter_firBlock_left_firStep[83] );
nand U1960 ( n1426, n1424, n1423 );
nand U1961 ( n1424, my_IIR_filter_firBlock_left_firStep[243], n1421 );
nand U1962 ( n1423, my_IIR_filter_firBlock_left_multProducts[50], n1422 );
or U1963 ( n1422, n1421, my_IIR_filter_firBlock_left_firStep[243] );
nand U1964 ( n2281, n2280, n2279 );
nand U1965 ( n2280, my_IIR_filter_firBlock_left_firStep[84], n2277 );
nand U1966 ( n2279, my_IIR_filter_firBlock_left_multProducts[51], n2278 );
or U1967 ( n2278, n2277, my_IIR_filter_firBlock_left_firStep[84] );
nand U1968 ( n1430, n1429, n1428 );
nand U1969 ( n1429, my_IIR_filter_firBlock_left_firStep[244], n1426 );
nand U1970 ( n1428, my_IIR_filter_firBlock_left_multProducts[51], n1427 );
or U1971 ( n1427, n1426, my_IIR_filter_firBlock_left_firStep[244] );
nand U1972 ( n2286, n2284, n2283 );
nand U1973 ( n2284, my_IIR_filter_firBlock_left_firStep[85], n2281 );
nand U1974 ( n2283, my_IIR_filter_firBlock_left_multProducts[52], n2282 );
or U1975 ( n2282, n2281, my_IIR_filter_firBlock_left_firStep[85] );
nand U1976 ( n1435, n1433, n1432 );
nand U1977 ( n1433, my_IIR_filter_firBlock_left_firStep[245], n1430 );
nand U1978 ( n1432, my_IIR_filter_firBlock_left_multProducts[52], n1431 );
or U1979 ( n1431, n1430, my_IIR_filter_firBlock_left_firStep[245] );
nand U1980 ( n2290, n2289, n2288 );
nand U1981 ( n2289, my_IIR_filter_firBlock_left_firStep[86], n2286 );
nand U1982 ( n2288, my_IIR_filter_firBlock_left_multProducts[53], n2287 );
or U1983 ( n2287, n2286, my_IIR_filter_firBlock_left_firStep[86] );
nand U1984 ( n1439, n1438, n1437 );
nand U1985 ( n1438, my_IIR_filter_firBlock_left_firStep[246], n1435 );
nand U1986 ( n1437, my_IIR_filter_firBlock_left_multProducts[53], n1436 );
or U1987 ( n1436, n1435, my_IIR_filter_firBlock_left_firStep[246] );
nand U1988 ( n2299, n2298, n2297 );
nand U1989 ( n2298, my_IIR_filter_firBlock_left_firStep[88], n2295 );
nand U1990 ( n2297, my_IIR_filter_firBlock_left_multProducts[55], n2296 );
or U1991 ( n2296, n2295, my_IIR_filter_firBlock_left_firStep[88] );
nand U1992 ( n1448, n1447, n1446 );
nand U1993 ( n1447, my_IIR_filter_firBlock_left_firStep[248], n1444 );
nand U1994 ( n1446, my_IIR_filter_firBlock_left_multProducts[55], n1445 );
or U1995 ( n1445, n1444, my_IIR_filter_firBlock_left_firStep[248] );
nand U1996 ( n2295, n2293, n2292 );
nand U1997 ( n2293, my_IIR_filter_firBlock_left_firStep[87], n2290 );
nand U1998 ( n2292, my_IIR_filter_firBlock_left_multProducts[54], n2291 );
or U1999 ( n2291, n2290, my_IIR_filter_firBlock_left_firStep[87] );
nand U2000 ( n1444, n1442, n1441 );
nand U2001 ( n1442, my_IIR_filter_firBlock_left_firStep[247], n1439 );
nand U2002 ( n1441, my_IIR_filter_firBlock_left_multProducts[54], n1440 );
or U2003 ( n1440, n1439, my_IIR_filter_firBlock_left_firStep[247] );
nand U2004 ( n2308, n2307, n2306 );
nand U2005 ( n2307, my_IIR_filter_firBlock_left_firStep[90], n2304 );
nand U2006 ( n2306, my_IIR_filter_firBlock_left_multProducts[57], n2305 );
or U2007 ( n2305, n2304, my_IIR_filter_firBlock_left_firStep[90] );
nand U2008 ( n1457, n1456, n1455 );
nand U2009 ( n1456, my_IIR_filter_firBlock_left_firStep[250], n1453 );
nand U2010 ( n1455, my_IIR_filter_firBlock_left_multProducts[57], n1454 );
or U2011 ( n1454, n1453, my_IIR_filter_firBlock_left_firStep[250] );
nand U2012 ( n2304, n2302, n2301 );
nand U2013 ( n2302, my_IIR_filter_firBlock_left_firStep[89], n2299 );
nand U2014 ( n2301, my_IIR_filter_firBlock_left_multProducts[56], n2300 );
or U2015 ( n2300, n2299, my_IIR_filter_firBlock_left_firStep[89] );
nand U2016 ( n1453, n1451, n1450 );
nand U2017 ( n1451, my_IIR_filter_firBlock_left_firStep[249], n1448 );
nand U2018 ( n1450, my_IIR_filter_firBlock_left_multProducts[56], n1449 );
or U2019 ( n1449, n1448, my_IIR_filter_firBlock_left_firStep[249] );
xor U2020 ( my_IIR_filter_firBlock_left_multProducts[56], n311, n1324 );
xor U2021 ( n311, my_IIR_filter_firBlock_left_multProducts[111], n549 );
xor U2022 ( my_IIR_filter_firBlock_left_multProducts[57], n1329, n1328 );
xor U2023 ( n1328, n549, my_IIR_filter_firBlock_left_multProducts[112] );
xor U2024 ( my_IIR_filter_firBlock_left_N159, n2049, n2047 );
xnor U2025 ( n2047, n243, my_IIR_filter_firBlock_left_firStep[158] );
xor U2026 ( my_IIR_filter_firBlock_left_N127, n1911, n1909 );
xnor U2027 ( n1909, n243, my_IIR_filter_firBlock_left_firStep[190] );
xor U2028 ( my_IIR_filter_firBlock_left_multProducts[33], n1349, n1348 );
xor U2029 ( n1348, inData_in[4], my_IIR_filter_firBlock_left_multProducts[92] );
xor U2030 ( my_IIR_filter_firBlock_left_multProducts[54], n312, n1315 );
xor U2031 ( n312, my_IIR_filter_firBlock_left_multProducts[109], my_IIR_filter_firBlock_left_multProducts[113] );
xor U2032 ( my_IIR_filter_firBlock_left_multProducts[34], n313, n1350 );
xor U2033 ( n313, inData_in[5], my_IIR_filter_firBlock_left_multProducts[93] );
xor U2034 ( my_IIR_filter_firBlock_left_multProducts[55], n1320, n1319 );
xor U2035 ( n1319, my_IIR_filter_firBlock_left_multProducts[114], my_IIR_filter_firBlock_left_multProducts[110] );
xnor U2036 ( my_IIR_filter_firBlock_right_N125, n3331, n314 );
xnor U2037 ( n314, my_IIR_filter_firBlock_right_multProducts[59], my_IIR_filter_firBlock_right_firStep[59] );
xor U2038 ( my_IIR_filter_firBlock_left_multProducts[35], n1238, n1237 );
xor U2039 ( n1237, my_IIR_filter_firBlock_left_multProducts[94], my_IIR_filter_firBlock_left_multProducts[90] );
xor U2040 ( my_IIR_filter_firBlock_left_multProducts[37], n1247, n1246 );
xor U2041 ( n1246, my_IIR_filter_firBlock_left_multProducts[96], my_IIR_filter_firBlock_left_multProducts[92] );
xor U2042 ( my_IIR_filter_firBlock_left_multProducts[39], n1255, n1254 );
xor U2043 ( n1254, my_IIR_filter_firBlock_left_multProducts[98], my_IIR_filter_firBlock_left_multProducts[94] );
xor U2044 ( my_IIR_filter_firBlock_left_multProducts[41], n1262, n1261 );
xor U2045 ( n1261, my_IIR_filter_firBlock_left_multProducts[100], my_IIR_filter_firBlock_left_multProducts[96] );
xor U2046 ( my_IIR_filter_firBlock_left_multProducts[43], n1269, n1268 );
xor U2047 ( n1268, my_IIR_filter_firBlock_left_multProducts[102], my_IIR_filter_firBlock_left_multProducts[98] );
xor U2048 ( my_IIR_filter_firBlock_left_multProducts[52], n315, n1306 );
xor U2049 ( n315, my_IIR_filter_firBlock_left_multProducts[107], my_IIR_filter_firBlock_left_multProducts[111] );
xor U2050 ( my_IIR_filter_firBlock_left_multProducts[31], n1346, n1345 );
xor U2051 ( n1345, inData_in[2], my_IIR_filter_firBlock_left_multProducts[90] );
and U2052 ( n2271, my_IIR_filter_firBlock_left_multProducts[31], my_IIR_filter_firBlock_left_firStep[64] );
and U2053 ( n1420, my_IIR_filter_firBlock_left_multProducts[31], my_IIR_filter_firBlock_left_firStep[224] );
xor U2054 ( my_IIR_filter_firBlock_left_multProducts[45], n1276, n1275 );
xor U2055 ( n1275, my_IIR_filter_firBlock_left_multProducts[104], my_IIR_filter_firBlock_left_multProducts[100] );
xor U2056 ( my_IIR_filter_firBlock_left_multProducts[36], n316, n1242 );
xor U2057 ( n316, my_IIR_filter_firBlock_left_multProducts[95], my_IIR_filter_firBlock_left_multProducts[91] );
xor U2058 ( my_IIR_filter_firBlock_left_multProducts[47], n1285, n1284 );
xor U2059 ( n1284, my_IIR_filter_firBlock_left_multProducts[106], my_IIR_filter_firBlock_left_multProducts[102] );
xor U2060 ( my_IIR_filter_firBlock_left_multProducts[38], n317, n1251 );
xor U2061 ( n317, my_IIR_filter_firBlock_left_multProducts[97], my_IIR_filter_firBlock_left_multProducts[93] );
xor U2062 ( my_IIR_filter_firBlock_left_multProducts[49], n1293, n1292 );
xor U2063 ( n1292, my_IIR_filter_firBlock_left_multProducts[108], my_IIR_filter_firBlock_left_multProducts[104] );
xor U2064 ( my_IIR_filter_firBlock_left_multProducts[53], n1311, n1310 );
xor U2065 ( n1310, my_IIR_filter_firBlock_left_multProducts[112], my_IIR_filter_firBlock_left_multProducts[108] );
xor U2066 ( my_IIR_filter_firBlock_left_multProducts[40], n318, n1258 );
xor U2067 ( n318, my_IIR_filter_firBlock_left_multProducts[95], my_IIR_filter_firBlock_left_multProducts[99] );
xor U2068 ( my_IIR_filter_firBlock_left_multProducts[51], n1302, n1301 );
xor U2069 ( n1301, my_IIR_filter_firBlock_left_multProducts[110], my_IIR_filter_firBlock_left_multProducts[106] );
xor U2070 ( my_IIR_filter_firBlock_left_multProducts[42], n319, n1265 );
xor U2071 ( n319, my_IIR_filter_firBlock_left_multProducts[97], my_IIR_filter_firBlock_left_multProducts[101] );
xor U2072 ( my_IIR_filter_firBlock_left_multProducts[44], n320, n1272 );
xor U2073 ( n320, my_IIR_filter_firBlock_left_multProducts[99], my_IIR_filter_firBlock_left_multProducts[103] );
xor U2074 ( my_IIR_filter_firBlock_left_multProducts[46], n321, n1280 );
xor U2075 ( n321, my_IIR_filter_firBlock_left_multProducts[101], my_IIR_filter_firBlock_left_multProducts[105] );
xor U2076 ( my_IIR_filter_firBlock_left_multProducts[48], n322, n1289 );
xor U2077 ( n322, my_IIR_filter_firBlock_left_multProducts[103], my_IIR_filter_firBlock_left_multProducts[107] );
xor U2078 ( my_IIR_filter_firBlock_left_multProducts[50], n323, n1297 );
xor U2079 ( n323, my_IIR_filter_firBlock_left_multProducts[105], my_IIR_filter_firBlock_left_multProducts[109] );
xor U2080 ( my_IIR_filter_firBlock_left_N253, n2450, n2449 );
xnor U2081 ( n2449, n631, my_IIR_filter_firBlock_left_firStep[60] );
xnor U2082 ( n1195, n631, my_IIR_filter_firBlock_left_firStep[284] );
xor U2083 ( my_IIR_filter_firBlock_right_N190, n324, n3524 );
xor U2084 ( n324, my_IIR_filter_firBlock_right_firStep[29], my_IIR_filter_firBlock_right_multProducts[29] );
xor U2085 ( my_IIR_filter_firBlock_left_N254, n325, n2456 );
xor U2086 ( n325, my_IIR_filter_firBlock_left_firStep[61], my_IIR_filter_firBlock_left_multProducts[89] );
xor U2087 ( my_IIR_filter_firBlock_left_N30, n326, n1202 );
xor U2088 ( n326, my_IIR_filter_firBlock_left_firStep[285], my_IIR_filter_firBlock_left_multProducts[89] );
xor U2089 ( my_IIR_filter_firBlock_right_N63, n2793, n2791 );
xnor U2090 ( n2791, n632, my_IIR_filter_firBlock_right_firStep[92] );
nand U2091 ( n2187, n2184, n2183 );
nand U2092 ( n2184, my_IIR_filter_firBlock_left_firStep[125], n2181 );
nand U2093 ( n2183, my_IIR_filter_firBlock_left_multProducts[59], n2182 );
or U2094 ( n2182, n2181, my_IIR_filter_firBlock_left_firStep[125] );
nand U2095 ( n1611, n1608, n1607 );
nand U2096 ( n1608, my_IIR_filter_firBlock_left_firStep[221], n1605 );
nand U2097 ( n1607, my_IIR_filter_firBlock_left_multProducts[59], n1606 );
or U2098 ( n1606, n1605, my_IIR_filter_firBlock_left_firStep[221] );
nand U2099 ( n2181, n2178, n2177 );
nand U2100 ( n2178, my_IIR_filter_firBlock_left_firStep[124], n2175 );
nand U2101 ( n2177, my_IIR_filter_firBlock_left_multProducts[58], n2176 );
or U2102 ( n2176, n2175, my_IIR_filter_firBlock_left_firStep[124] );
nand U2103 ( n1605, n1602, n1601 );
nand U2104 ( n1602, my_IIR_filter_firBlock_left_firStep[220], n1599 );
nand U2105 ( n1601, my_IIR_filter_firBlock_left_multProducts[58], n1600 );
or U2106 ( n1600, n1599, my_IIR_filter_firBlock_left_firStep[220] );
xor U2107 ( my_IIR_filter_firBlock_left_N192, n2191, n2190 );
xnor U2108 ( n2191, n549, my_IIR_filter_firBlock_left_firStep[127] );
nor U2109 ( n2190, n2189, n2188 );
and U2110 ( n2188, n2187, my_IIR_filter_firBlock_left_firStep[126] );
xor U2111 ( my_IIR_filter_firBlock_left_N96, n1615, n1614 );
xnor U2112 ( n1615, n549, my_IIR_filter_firBlock_left_firStep[223] );
nor U2113 ( n1614, n1613, n1612 );
and U2114 ( n1612, n1611, my_IIR_filter_firBlock_left_firStep[222] );
nor U2115 ( n2189, n2186, n630 );
nor U2116 ( n2186, my_IIR_filter_firBlock_left_firStep[126], n2187 );
nor U2117 ( n1613, n1610, n630 );
nor U2118 ( n1610, my_IIR_filter_firBlock_left_firStep[222], n1611 );
nand U2119 ( n2170, n2169, n2168 );
nand U2120 ( n2169, my_IIR_filter_firBlock_left_firStep[122], n2166 );
nand U2121 ( n2168, my_IIR_filter_firBlock_left_multProducts[56], n2167 );
or U2122 ( n2167, n2166, my_IIR_filter_firBlock_left_firStep[122] );
nand U2123 ( n1594, n1593, n1592 );
nand U2124 ( n1593, my_IIR_filter_firBlock_left_firStep[218], n1590 );
nand U2125 ( n1592, my_IIR_filter_firBlock_left_multProducts[56], n1591 );
or U2126 ( n1591, n1590, my_IIR_filter_firBlock_left_firStep[218] );
nand U2127 ( n2175, n2173, n2172 );
nand U2128 ( n2173, my_IIR_filter_firBlock_left_firStep[123], n2170 );
nand U2129 ( n2172, my_IIR_filter_firBlock_left_multProducts[57], n2171 );
or U2130 ( n2171, n2170, my_IIR_filter_firBlock_left_firStep[123] );
nand U2131 ( n1599, n1597, n1596 );
nand U2132 ( n1597, my_IIR_filter_firBlock_left_firStep[219], n1594 );
nand U2133 ( n1596, my_IIR_filter_firBlock_left_multProducts[57], n1595 );
or U2134 ( n1595, n1594, my_IIR_filter_firBlock_left_firStep[219] );
nand U2135 ( my_IIR_filter_firBlock_left_multProducts[60], n1342, n1341 );
nand U2136 ( n1342, my_IIR_filter_firBlock_left_multProducts[114], n1339 );
nand U2137 ( n1341, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n1340 );
or U2138 ( n1340, n1339, my_IIR_filter_firBlock_left_multProducts[114] );
nand U2139 ( n2194, n2072, n2071 );
nand U2140 ( n2072, my_IIR_filter_firBlock_left_firStep[99], n2192 );
nand U2141 ( n2071, my_IIR_filter_firBlock_left_multProducts[33], n2070 );
or U2142 ( n2070, n2192, my_IIR_filter_firBlock_left_firStep[99] );
nand U2143 ( n1618, n1496, n1495 );
nand U2144 ( n1496, my_IIR_filter_firBlock_left_firStep[195], n1616 );
nand U2145 ( n1495, my_IIR_filter_firBlock_left_multProducts[33], n1494 );
or U2146 ( n1494, n1616, my_IIR_filter_firBlock_left_firStep[195] );
nand U2147 ( n2197, n2078, n2077 );
nand U2148 ( n2078, my_IIR_filter_firBlock_left_firStep[101], n2195 );
nand U2149 ( n2077, my_IIR_filter_firBlock_left_multProducts[35], n2076 );
or U2150 ( n2076, n2195, my_IIR_filter_firBlock_left_firStep[101] );
nand U2151 ( n1621, n1502, n1501 );
nand U2152 ( n1502, my_IIR_filter_firBlock_left_firStep[197], n1619 );
nand U2153 ( n1501, my_IIR_filter_firBlock_left_multProducts[35], n1500 );
or U2154 ( n1500, n1619, my_IIR_filter_firBlock_left_firStep[197] );
nand U2155 ( n2198, n2081, n2080 );
nand U2156 ( n2081, my_IIR_filter_firBlock_left_firStep[102], n2197 );
nand U2157 ( n2080, my_IIR_filter_firBlock_left_multProducts[36], n2079 );
or U2158 ( n2079, n2197, my_IIR_filter_firBlock_left_firStep[102] );
nand U2159 ( n1622, n1505, n1504 );
nand U2160 ( n1505, my_IIR_filter_firBlock_left_firStep[198], n1621 );
nand U2161 ( n1504, my_IIR_filter_firBlock_left_multProducts[36], n1503 );
or U2162 ( n1503, n1621, my_IIR_filter_firBlock_left_firStep[198] );
nand U2163 ( n2192, n2069, n2068 );
nand U2164 ( n2069, my_IIR_filter_firBlock_left_firStep[98], n2180 );
nand U2165 ( n2068, my_IIR_filter_firBlock_left_multProducts[32], n2067 );
or U2166 ( n2067, n2180, my_IIR_filter_firBlock_left_firStep[98] );
nand U2167 ( n1616, n1493, n1492 );
nand U2168 ( n1493, my_IIR_filter_firBlock_left_firStep[194], n1604 );
nand U2169 ( n1492, my_IIR_filter_firBlock_left_multProducts[32], n1491 );
or U2170 ( n1491, n1604, my_IIR_filter_firBlock_left_firStep[194] );
nand U2171 ( n2195, n2075, n2074 );
nand U2172 ( n2075, my_IIR_filter_firBlock_left_firStep[100], n2194 );
nand U2173 ( n2074, my_IIR_filter_firBlock_left_multProducts[34], n2073 );
or U2174 ( n2073, n2194, my_IIR_filter_firBlock_left_firStep[100] );
nand U2175 ( n1619, n1499, n1498 );
nand U2176 ( n1499, my_IIR_filter_firBlock_left_firStep[196], n1618 );
nand U2177 ( n1498, my_IIR_filter_firBlock_left_multProducts[34], n1497 );
or U2178 ( n1497, n1618, my_IIR_filter_firBlock_left_firStep[196] );
nand U2179 ( n2200, n2084, n2083 );
nand U2180 ( n2084, my_IIR_filter_firBlock_left_firStep[103], n2198 );
nand U2181 ( n2083, my_IIR_filter_firBlock_left_multProducts[37], n2082 );
or U2182 ( n2082, n2198, my_IIR_filter_firBlock_left_firStep[103] );
nand U2183 ( n1624, n1508, n1507 );
nand U2184 ( n1508, my_IIR_filter_firBlock_left_firStep[199], n1622 );
nand U2185 ( n1507, my_IIR_filter_firBlock_left_multProducts[37], n1506 );
or U2186 ( n1506, n1622, my_IIR_filter_firBlock_left_firStep[199] );
nand U2187 ( n2092, n2090, n2089 );
nand U2188 ( n2090, my_IIR_filter_firBlock_left_firStep[105], n2201 );
nand U2189 ( n2089, my_IIR_filter_firBlock_left_multProducts[39], n2088 );
or U2190 ( n2088, n2201, my_IIR_filter_firBlock_left_firStep[105] );
nand U2191 ( n1516, n1514, n1513 );
nand U2192 ( n1514, my_IIR_filter_firBlock_left_firStep[201], n1625 );
nand U2193 ( n1513, my_IIR_filter_firBlock_left_multProducts[39], n1512 );
or U2194 ( n1512, n1625, my_IIR_filter_firBlock_left_firStep[201] );
nand U2195 ( n2201, n2087, n2086 );
nand U2196 ( n2087, my_IIR_filter_firBlock_left_firStep[104], n2200 );
nand U2197 ( n2086, my_IIR_filter_firBlock_left_multProducts[38], n2085 );
or U2198 ( n2085, n2200, my_IIR_filter_firBlock_left_firStep[104] );
nand U2199 ( n1625, n1511, n1510 );
nand U2200 ( n1511, my_IIR_filter_firBlock_left_firStep[200], n1624 );
nand U2201 ( n1510, my_IIR_filter_firBlock_left_multProducts[38], n1509 );
or U2202 ( n1509, n1624, my_IIR_filter_firBlock_left_firStep[200] );
nand U2203 ( n2101, n2099, n2098 );
nand U2204 ( n2099, my_IIR_filter_firBlock_left_firStep[107], n2096 );
nand U2205 ( n2098, my_IIR_filter_firBlock_left_multProducts[41], n2097 );
or U2206 ( n2097, n2096, my_IIR_filter_firBlock_left_firStep[107] );
nand U2207 ( n1525, n1523, n1522 );
nand U2208 ( n1523, my_IIR_filter_firBlock_left_firStep[203], n1520 );
nand U2209 ( n1522, my_IIR_filter_firBlock_left_multProducts[41], n1521 );
or U2210 ( n1521, n1520, my_IIR_filter_firBlock_left_firStep[203] );
nand U2211 ( n2096, n2095, n2094 );
nand U2212 ( n2095, my_IIR_filter_firBlock_left_firStep[106], n2092 );
nand U2213 ( n2094, my_IIR_filter_firBlock_left_multProducts[40], n2093 );
or U2214 ( n2093, n2092, my_IIR_filter_firBlock_left_firStep[106] );
nand U2215 ( n1520, n1519, n1518 );
nand U2216 ( n1519, my_IIR_filter_firBlock_left_firStep[202], n1516 );
nand U2217 ( n1518, my_IIR_filter_firBlock_left_multProducts[40], n1517 );
or U2218 ( n1517, n1516, my_IIR_filter_firBlock_left_firStep[202] );
nand U2219 ( n2105, n2104, n2103 );
nand U2220 ( n2104, my_IIR_filter_firBlock_left_firStep[108], n2101 );
nand U2221 ( n2103, my_IIR_filter_firBlock_left_multProducts[42], n2102 );
or U2222 ( n2102, n2101, my_IIR_filter_firBlock_left_firStep[108] );
nand U2223 ( n1529, n1528, n1527 );
nand U2224 ( n1528, my_IIR_filter_firBlock_left_firStep[204], n1525 );
nand U2225 ( n1527, my_IIR_filter_firBlock_left_multProducts[42], n1526 );
or U2226 ( n1526, n1525, my_IIR_filter_firBlock_left_firStep[204] );
nand U2227 ( n2110, n2108, n2107 );
nand U2228 ( n2108, my_IIR_filter_firBlock_left_firStep[109], n2105 );
nand U2229 ( n2107, my_IIR_filter_firBlock_left_multProducts[43], n2106 );
or U2230 ( n2106, n2105, my_IIR_filter_firBlock_left_firStep[109] );
nand U2231 ( n1534, n1532, n1531 );
nand U2232 ( n1532, my_IIR_filter_firBlock_left_firStep[205], n1529 );
nand U2233 ( n1531, my_IIR_filter_firBlock_left_multProducts[43], n1530 );
or U2234 ( n1530, n1529, my_IIR_filter_firBlock_left_firStep[205] );
nand U2235 ( n2119, n2117, n2116 );
nand U2236 ( n2117, my_IIR_filter_firBlock_left_firStep[111], n2114 );
nand U2237 ( n2116, my_IIR_filter_firBlock_left_multProducts[45], n2115 );
or U2238 ( n2115, n2114, my_IIR_filter_firBlock_left_firStep[111] );
nand U2239 ( n1543, n1541, n1540 );
nand U2240 ( n1541, my_IIR_filter_firBlock_left_firStep[207], n1538 );
nand U2241 ( n1540, my_IIR_filter_firBlock_left_multProducts[45], n1539 );
or U2242 ( n1539, n1538, my_IIR_filter_firBlock_left_firStep[207] );
nand U2243 ( n2114, n2113, n2112 );
nand U2244 ( n2113, my_IIR_filter_firBlock_left_firStep[110], n2110 );
nand U2245 ( n2112, my_IIR_filter_firBlock_left_multProducts[44], n2111 );
or U2246 ( n2111, n2110, my_IIR_filter_firBlock_left_firStep[110] );
nand U2247 ( n1538, n1537, n1536 );
nand U2248 ( n1537, my_IIR_filter_firBlock_left_firStep[206], n1534 );
nand U2249 ( n1536, my_IIR_filter_firBlock_left_multProducts[44], n1535 );
or U2250 ( n1535, n1534, my_IIR_filter_firBlock_left_firStep[206] );
nand U2251 ( n2123, n2122, n2121 );
nand U2252 ( n2122, my_IIR_filter_firBlock_left_firStep[112], n2119 );
nand U2253 ( n2121, my_IIR_filter_firBlock_left_multProducts[46], n2120 );
or U2254 ( n2120, n2119, my_IIR_filter_firBlock_left_firStep[112] );
nand U2255 ( n1547, n1546, n1545 );
nand U2256 ( n1546, my_IIR_filter_firBlock_left_firStep[208], n1543 );
nand U2257 ( n1545, my_IIR_filter_firBlock_left_multProducts[46], n1544 );
or U2258 ( n1544, n1543, my_IIR_filter_firBlock_left_firStep[208] );
nand U2259 ( n2128, n2126, n2125 );
nand U2260 ( n2126, my_IIR_filter_firBlock_left_firStep[113], n2123 );
nand U2261 ( n2125, my_IIR_filter_firBlock_left_multProducts[47], n2124 );
or U2262 ( n2124, n2123, my_IIR_filter_firBlock_left_firStep[113] );
nand U2263 ( n1552, n1550, n1549 );
nand U2264 ( n1550, my_IIR_filter_firBlock_left_firStep[209], n1547 );
nand U2265 ( n1549, my_IIR_filter_firBlock_left_multProducts[47], n1548 );
or U2266 ( n1548, n1547, my_IIR_filter_firBlock_left_firStep[209] );
nand U2267 ( n2134, n2131, n2130 );
nand U2268 ( n2131, my_IIR_filter_firBlock_left_firStep[114], n2128 );
nand U2269 ( n2130, my_IIR_filter_firBlock_left_multProducts[48], n2129 );
or U2270 ( n2129, n2128, my_IIR_filter_firBlock_left_firStep[114] );
nand U2271 ( n1558, n1555, n1554 );
nand U2272 ( n1555, my_IIR_filter_firBlock_left_firStep[210], n1552 );
nand U2273 ( n1554, my_IIR_filter_firBlock_left_multProducts[48], n1553 );
or U2274 ( n1553, n1552, my_IIR_filter_firBlock_left_firStep[210] );
nand U2275 ( n2139, n2137, n2136 );
nand U2276 ( n2137, my_IIR_filter_firBlock_left_firStep[115], n2134 );
nand U2277 ( n2136, my_IIR_filter_firBlock_left_multProducts[49], n2135 );
or U2278 ( n2135, n2134, my_IIR_filter_firBlock_left_firStep[115] );
nand U2279 ( n1563, n1561, n1560 );
nand U2280 ( n1561, my_IIR_filter_firBlock_left_firStep[211], n1558 );
nand U2281 ( n1560, my_IIR_filter_firBlock_left_multProducts[49], n1559 );
or U2282 ( n1559, n1558, my_IIR_filter_firBlock_left_firStep[211] );
nand U2283 ( n2143, n2142, n2141 );
nand U2284 ( n2142, my_IIR_filter_firBlock_left_firStep[116], n2139 );
nand U2285 ( n2141, my_IIR_filter_firBlock_left_multProducts[50], n2140 );
or U2286 ( n2140, n2139, my_IIR_filter_firBlock_left_firStep[116] );
nand U2287 ( n1567, n1566, n1565 );
nand U2288 ( n1566, my_IIR_filter_firBlock_left_firStep[212], n1563 );
nand U2289 ( n1565, my_IIR_filter_firBlock_left_multProducts[50], n1564 );
or U2290 ( n1564, n1563, my_IIR_filter_firBlock_left_firStep[212] );
nand U2291 ( n2148, n2146, n2145 );
nand U2292 ( n2146, my_IIR_filter_firBlock_left_firStep[117], n2143 );
nand U2293 ( n2145, my_IIR_filter_firBlock_left_multProducts[51], n2144 );
or U2294 ( n2144, n2143, my_IIR_filter_firBlock_left_firStep[117] );
nand U2295 ( n1572, n1570, n1569 );
nand U2296 ( n1570, my_IIR_filter_firBlock_left_firStep[213], n1567 );
nand U2297 ( n1569, my_IIR_filter_firBlock_left_multProducts[51], n1568 );
or U2298 ( n1568, n1567, my_IIR_filter_firBlock_left_firStep[213] );
nand U2299 ( n2152, n2151, n2150 );
nand U2300 ( n2151, my_IIR_filter_firBlock_left_firStep[118], n2148 );
nand U2301 ( n2150, my_IIR_filter_firBlock_left_multProducts[52], n2149 );
or U2302 ( n2149, n2148, my_IIR_filter_firBlock_left_firStep[118] );
nand U2303 ( n1576, n1575, n1574 );
nand U2304 ( n1575, my_IIR_filter_firBlock_left_firStep[214], n1572 );
nand U2305 ( n1574, my_IIR_filter_firBlock_left_multProducts[52], n1573 );
or U2306 ( n1573, n1572, my_IIR_filter_firBlock_left_firStep[214] );
nand U2307 ( n2157, n2155, n2154 );
nand U2308 ( n2155, my_IIR_filter_firBlock_left_firStep[119], n2152 );
nand U2309 ( n2154, my_IIR_filter_firBlock_left_multProducts[53], n2153 );
or U2310 ( n2153, n2152, my_IIR_filter_firBlock_left_firStep[119] );
nand U2311 ( n1581, n1579, n1578 );
nand U2312 ( n1579, my_IIR_filter_firBlock_left_firStep[215], n1576 );
nand U2313 ( n1578, my_IIR_filter_firBlock_left_multProducts[53], n1577 );
or U2314 ( n1577, n1576, my_IIR_filter_firBlock_left_firStep[215] );
nand U2315 ( n2166, n2164, n2163 );
nand U2316 ( n2164, my_IIR_filter_firBlock_left_firStep[121], n2161 );
nand U2317 ( n2163, my_IIR_filter_firBlock_left_multProducts[55], n2162 );
or U2318 ( n2162, n2161, my_IIR_filter_firBlock_left_firStep[121] );
nand U2319 ( n1590, n1588, n1587 );
nand U2320 ( n1588, my_IIR_filter_firBlock_left_firStep[217], n1585 );
nand U2321 ( n1587, my_IIR_filter_firBlock_left_multProducts[55], n1586 );
or U2322 ( n1586, n1585, my_IIR_filter_firBlock_left_firStep[217] );
nand U2323 ( n2161, n2160, n2159 );
nand U2324 ( n2160, my_IIR_filter_firBlock_left_firStep[120], n2157 );
nand U2325 ( n2159, my_IIR_filter_firBlock_left_multProducts[54], n2158 );
or U2326 ( n2158, n2157, my_IIR_filter_firBlock_left_firStep[120] );
nand U2327 ( n1585, n1584, n1583 );
nand U2328 ( n1584, my_IIR_filter_firBlock_left_firStep[216], n1581 );
nand U2329 ( n1583, my_IIR_filter_firBlock_left_multProducts[54], n1582 );
or U2330 ( n1582, n1581, my_IIR_filter_firBlock_left_firStep[216] );
nand U2331 ( n2180, n2066, n2065 );
nand U2332 ( n2066, my_IIR_filter_firBlock_left_firStep[97], n2133 );
nand U2333 ( n2065, my_IIR_filter_firBlock_left_multProducts[31], n2064 );
or U2334 ( n2064, my_IIR_filter_firBlock_left_firStep[97], n2133 );
nand U2335 ( n1604, n1490, n1489 );
nand U2336 ( n1490, my_IIR_filter_firBlock_left_firStep[193], n1557 );
nand U2337 ( n1489, my_IIR_filter_firBlock_left_multProducts[31], n1488 );
or U2338 ( n1488, my_IIR_filter_firBlock_left_firStep[193], n1557 );
xnor U2339 ( my_IIR_filter_firBlock_right_N189, n3518, n327 );
xnor U2340 ( n327, my_IIR_filter_firBlock_right_multProducts[28], my_IIR_filter_firBlock_right_firStep[28] );
xnor U2341 ( my_IIR_filter_firBlock_left_N223, n2324, n328 );
xor U2342 ( n328, n526, my_IIR_filter_firBlock_left_firStep[94] );
xnor U2343 ( my_IIR_filter_firBlock_left_N63, n1473, n329 );
xor U2344 ( n329, n526, my_IIR_filter_firBlock_left_firStep[254] );
xor U2345 ( my_IIR_filter_firBlock_right_N124, n330, n3327 );
xor U2346 ( n330, my_IIR_filter_firBlock_right_firStep[58], my_IIR_filter_firBlock_right_multProducts[58] );
xor U2347 ( my_IIR_filter_firBlock_left_multProducts[30], n1344, n1343 );
and U2348 ( n2133, my_IIR_filter_firBlock_left_multProducts[30], my_IIR_filter_firBlock_left_firStep[96] );
and U2349 ( n1557, my_IIR_filter_firBlock_left_multProducts[30], my_IIR_filter_firBlock_left_firStep[192] );
xor U2350 ( my_IIR_filter_firBlock_left_N158, n331, n2043 );
xor U2351 ( n331, my_IIR_filter_firBlock_left_firStep[157], my_IIR_filter_firBlock_left_multProducts[29] );
xor U2352 ( my_IIR_filter_firBlock_left_N126, n332, n1907 );
xor U2353 ( n332, my_IIR_filter_firBlock_left_firStep[189], my_IIR_filter_firBlock_left_multProducts[29] );
xor U2354 ( n3322, my_IIR_filter_firBlock_right_multProducts[57], my_IIR_filter_firBlock_right_firStep[57] );
xor U2355 ( my_IIR_filter_firBlock_right_N62, n333, n2787 );
xor U2356 ( n333, my_IIR_filter_firBlock_right_firStep[91], my_IIR_filter_firBlock_right_multProducts[91] );
xor U2357 ( my_IIR_filter_firBlock_left_N191, n2187, n2185 );
xnor U2358 ( n2185, n630, my_IIR_filter_firBlock_left_firStep[126] );
xor U2359 ( my_IIR_filter_firBlock_left_N95, n1611, n1609 );
xnor U2360 ( n1609, n630, my_IIR_filter_firBlock_left_firStep[222] );
xor U2361 ( my_IIR_filter_firBlock_right_N188, n334, n3514 );
xor U2362 ( n334, my_IIR_filter_firBlock_right_firStep[27], my_IIR_filter_firBlock_right_multProducts[27] );
xor U2363 ( my_IIR_filter_firBlock_left_N252, n335, n2445 );
xor U2364 ( n335, my_IIR_filter_firBlock_left_firStep[59], my_IIR_filter_firBlock_left_multProducts[88] );
xor U2365 ( my_IIR_filter_firBlock_left_N28, n336, n1191 );
xor U2366 ( n336, my_IIR_filter_firBlock_left_firStep[283], my_IIR_filter_firBlock_left_multProducts[88] );
xor U2367 ( my_IIR_filter_firBlock_left_N157, n2037, n2036 );
xor U2368 ( n2036, my_IIR_filter_firBlock_left_multProducts[28], my_IIR_filter_firBlock_left_firStep[156] );
xor U2369 ( my_IIR_filter_firBlock_left_N125, n1901, n1900 );
xor U2370 ( n1900, my_IIR_filter_firBlock_left_multProducts[28], my_IIR_filter_firBlock_left_firStep[188] );
xor U2371 ( my_IIR_filter_firBlock_left_N222, n337, n2319 );
xor U2372 ( n337, my_IIR_filter_firBlock_left_firStep[93], my_IIR_filter_firBlock_left_multProducts[60] );
xor U2373 ( my_IIR_filter_firBlock_left_N62, n338, n1468 );
xor U2374 ( n338, my_IIR_filter_firBlock_left_firStep[253], my_IIR_filter_firBlock_left_multProducts[60] );
xor U2375 ( my_IIR_filter_firBlock_left_N221, n2313, n2312 );
xor U2376 ( n2312, my_IIR_filter_firBlock_left_multProducts[59], my_IIR_filter_firBlock_left_firStep[92] );
xor U2377 ( my_IIR_filter_firBlock_left_N61, n1462, n1461 );
xor U2378 ( n1461, my_IIR_filter_firBlock_left_multProducts[59], my_IIR_filter_firBlock_left_firStep[252] );
xor U2379 ( my_IIR_filter_firBlock_left_N251, n2441, n2440 );
xor U2380 ( my_IIR_filter_firBlock_left_N190, n339, n2181 );
xor U2381 ( n339, my_IIR_filter_firBlock_left_firStep[125], my_IIR_filter_firBlock_left_multProducts[59] );
xor U2382 ( my_IIR_filter_firBlock_left_N94, n340, n1605 );
xor U2383 ( n340, my_IIR_filter_firBlock_left_firStep[221], my_IIR_filter_firBlock_left_multProducts[59] );
nand U2384 ( n2607, n2604, n2603 );
nand U2385 ( n2604, my_IIR_filter_firBlock_left_firStep[29], n2601 );
nand U2386 ( n2603, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2602 );
or U2387 ( n2602, n2601, my_IIR_filter_firBlock_left_firStep[29] );
or U2388 ( n2479, n341, n342 );
nor U2389 ( n342, n2600, my_IIR_filter_firBlock_left_firStep[2] );
nand U2390 ( n2615, n2485, n2484 );
nand U2391 ( n2485, my_IIR_filter_firBlock_left_firStep[4], n2614 );
nand U2392 ( n2484, my_IIR_filter_firBlock_left_multProducts[94], n2483 );
or U2393 ( n2483, n2614, my_IIR_filter_firBlock_left_firStep[4] );
nand U2394 ( n2517, n2515, n2514 );
nand U2395 ( n2515, my_IIR_filter_firBlock_left_firStep[12], n2512 );
nand U2396 ( n2514, my_IIR_filter_firBlock_left_multProducts[102], n2513 );
or U2397 ( n2513, n2512, my_IIR_filter_firBlock_left_firStep[12] );
nand U2398 ( n2537, n2535, n2534 );
nand U2399 ( n2535, my_IIR_filter_firBlock_left_firStep[16], n2532 );
nand U2400 ( n2534, my_IIR_filter_firBlock_left_multProducts[106], n2533 );
or U2401 ( n2533, n2532, my_IIR_filter_firBlock_left_firStep[16] );
nand U2402 ( n2549, n2545, n2544 );
nand U2403 ( n2545, my_IIR_filter_firBlock_left_firStep[18], n2542 );
nand U2404 ( n2544, my_IIR_filter_firBlock_left_multProducts[108], n2543 );
or U2405 ( n2543, n2542, my_IIR_filter_firBlock_left_firStep[18] );
nand U2406 ( n2507, n2505, n2504 );
nand U2407 ( n2505, my_IIR_filter_firBlock_left_firStep[10], n2502 );
nand U2408 ( n2504, my_IIR_filter_firBlock_left_multProducts[100], n2503 );
or U2409 ( n2503, n2502, my_IIR_filter_firBlock_left_firStep[10] );
nand U2410 ( n2527, n2525, n2524 );
nand U2411 ( n2525, my_IIR_filter_firBlock_left_firStep[14], n2522 );
nand U2412 ( n2524, my_IIR_filter_firBlock_left_multProducts[104], n2523 );
or U2413 ( n2523, n2522, my_IIR_filter_firBlock_left_firStep[14] );
nand U2414 ( n2559, n2557, n2556 );
nand U2415 ( n2557, my_IIR_filter_firBlock_left_firStep[20], n2554 );
nand U2416 ( n2556, my_IIR_filter_firBlock_left_multProducts[110], n2555 );
or U2417 ( n2555, n2554, my_IIR_filter_firBlock_left_firStep[20] );
nand U2418 ( n2579, n2577, n2576 );
nand U2419 ( n2577, my_IIR_filter_firBlock_left_firStep[24], n2574 );
nand U2420 ( n2576, my_IIR_filter_firBlock_left_multProducts[114], n2575 );
or U2421 ( n2575, n2574, my_IIR_filter_firBlock_left_firStep[24] );
nand U2422 ( n2589, n2587, n2586 );
nand U2423 ( n2587, my_IIR_filter_firBlock_left_firStep[26], n2584 );
nand U2424 ( n2586, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2585 );
or U2425 ( n2585, n2584, my_IIR_filter_firBlock_left_firStep[26] );
nand U2426 ( n2601, n2597, n2596 );
nand U2427 ( n2597, my_IIR_filter_firBlock_left_firStep[28], n2594 );
nand U2428 ( n2596, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2595 );
or U2429 ( n2595, n2594, my_IIR_filter_firBlock_left_firStep[28] );
nand U2430 ( n2600, n2478, n2477 );
nand U2431 ( n2478, my_IIR_filter_firBlock_left_firStep[1], n2548 );
nand U2432 ( n2477, my_IIR_filter_firBlock_left_multProducts[91], n2476 );
or U2433 ( n2476, my_IIR_filter_firBlock_left_firStep[1], n2548 );
or U2434 ( n2481, n343, n344 );
nor U2435 ( n344, n2612, my_IIR_filter_firBlock_left_firStep[3] );
nand U2436 ( n2618, n2488, n2487 );
nand U2437 ( n2488, my_IIR_filter_firBlock_left_firStep[5], n2615 );
nand U2438 ( n2487, my_IIR_filter_firBlock_left_multProducts[95], n2486 );
or U2439 ( n2486, n2615, my_IIR_filter_firBlock_left_firStep[5] );
nand U2440 ( n2532, n2530, n2529 );
nand U2441 ( n2530, my_IIR_filter_firBlock_left_firStep[15], n2527 );
nand U2442 ( n2529, my_IIR_filter_firBlock_left_multProducts[105], n2528 );
or U2443 ( n2528, n2527, my_IIR_filter_firBlock_left_firStep[15] );
nand U2444 ( n2564, n2562, n2561 );
nand U2445 ( n2562, my_IIR_filter_firBlock_left_firStep[21], n2559 );
nand U2446 ( n2561, my_IIR_filter_firBlock_left_multProducts[111], n2560 );
or U2447 ( n2560, n2559, my_IIR_filter_firBlock_left_firStep[21] );
nand U2448 ( n2574, n2572, n2571 );
nand U2449 ( n2572, my_IIR_filter_firBlock_left_firStep[23], n2569 );
nand U2450 ( n2571, my_IIR_filter_firBlock_left_multProducts[113], n2570 );
or U2451 ( n2570, n2569, my_IIR_filter_firBlock_left_firStep[23] );
nand U2452 ( n2512, n2510, n2509 );
nand U2453 ( n2510, my_IIR_filter_firBlock_left_firStep[11], n2507 );
nand U2454 ( n2509, my_IIR_filter_firBlock_left_multProducts[101], n2508 );
or U2455 ( n2508, n2507, my_IIR_filter_firBlock_left_firStep[11] );
nand U2456 ( n2622, n2494, n2493 );
nand U2457 ( n2494, my_IIR_filter_firBlock_left_firStep[7], n2619 );
nand U2458 ( n2493, my_IIR_filter_firBlock_left_multProducts[97], n2492 );
or U2459 ( n2492, n2619, my_IIR_filter_firBlock_left_firStep[7] );
nand U2460 ( n2502, n2500, n2499 );
nand U2461 ( n2500, my_IIR_filter_firBlock_left_firStep[9], n2623 );
nand U2462 ( n2499, my_IIR_filter_firBlock_left_multProducts[99], n2498 );
or U2463 ( n2498, n2623, my_IIR_filter_firBlock_left_firStep[9] );
nand U2464 ( n2522, n2520, n2519 );
nand U2465 ( n2520, my_IIR_filter_firBlock_left_firStep[13], n2517 );
nand U2466 ( n2519, my_IIR_filter_firBlock_left_multProducts[103], n2518 );
or U2467 ( n2518, n2517, my_IIR_filter_firBlock_left_firStep[13] );
nand U2468 ( n2542, n2540, n2539 );
nand U2469 ( n2540, my_IIR_filter_firBlock_left_firStep[17], n2537 );
nand U2470 ( n2539, my_IIR_filter_firBlock_left_multProducts[107], n2538 );
or U2471 ( n2538, n2537, my_IIR_filter_firBlock_left_firStep[17] );
nand U2472 ( n2554, n2552, n2551 );
nand U2473 ( n2552, my_IIR_filter_firBlock_left_firStep[19], n2549 );
nand U2474 ( n2551, my_IIR_filter_firBlock_left_multProducts[109], n2550 );
or U2475 ( n2550, n2549, my_IIR_filter_firBlock_left_firStep[19] );
nand U2476 ( n2584, n2582, n2581 );
nand U2477 ( n2582, my_IIR_filter_firBlock_left_firStep[25], n2579 );
nand U2478 ( n2581, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2580 );
or U2479 ( n2580, n2579, my_IIR_filter_firBlock_left_firStep[25] );
nand U2480 ( n2594, n2592, n2591 );
nand U2481 ( n2592, my_IIR_filter_firBlock_left_firStep[27], n2589 );
nand U2482 ( n2591, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w3_38_, n2590 );
or U2483 ( n2590, n2589, my_IIR_filter_firBlock_left_firStep[27] );
nand U2484 ( n2569, n2567, n2566 );
nand U2485 ( n2567, my_IIR_filter_firBlock_left_firStep[22], n2564 );
nand U2486 ( n2566, my_IIR_filter_firBlock_left_multProducts[112], n2565 );
or U2487 ( n2565, n2564, my_IIR_filter_firBlock_left_firStep[22] );
nand U2488 ( n2623, n2497, n2496 );
nand U2489 ( n2497, my_IIR_filter_firBlock_left_firStep[8], n2622 );
nand U2490 ( n2496, my_IIR_filter_firBlock_left_multProducts[98], n2495 );
or U2491 ( n2495, n2622, my_IIR_filter_firBlock_left_firStep[8] );
nor U2492 ( n2609, n2606, n526 );
nor U2493 ( n2606, my_IIR_filter_firBlock_left_firStep[30], n2607 );
and U2494 ( n2548, my_IIR_filter_firBlock_left_multProducts[90], my_IIR_filter_firBlock_left_firStep[0] );
nand U2495 ( n2619, n2491, n2490 );
nand U2496 ( n2491, my_IIR_filter_firBlock_left_firStep[6], n2618 );
nand U2497 ( n2490, my_IIR_filter_firBlock_left_multProducts[96], n2489 );
or U2498 ( n2489, n2618, my_IIR_filter_firBlock_left_firStep[6] );
xor U2499 ( my_IIR_filter_firBlock_left_N288, n2611, n2610 );
xnor U2500 ( n2611, n549, my_IIR_filter_firBlock_left_firStep[31] );
nor U2501 ( n2610, n2609, n2608 );
and U2502 ( n2608, n2607, my_IIR_filter_firBlock_left_firStep[30] );
xor U2503 ( my_IIR_filter_firBlock_right_N61, n2781, n2780 );
xor U2504 ( n2780, my_IIR_filter_firBlock_right_multProducts[90], my_IIR_filter_firBlock_right_firStep[90] );
xor U2505 ( my_IIR_filter_firBlock_right_N122, n345, n3318 );
xor U2506 ( n345, my_IIR_filter_firBlock_right_firStep[56], my_IIR_filter_firBlock_right_multProducts[56] );
xor U2507 ( n3509, my_IIR_filter_firBlock_right_multProducts[26], my_IIR_filter_firBlock_right_firStep[26] );
xor U2508 ( my_IIR_filter_firBlock_left_N156, n346, n2032 );
xor U2509 ( n346, my_IIR_filter_firBlock_left_firStep[155], my_IIR_filter_firBlock_left_multProducts[27] );
xor U2510 ( my_IIR_filter_firBlock_left_N124, n347, n1896 );
xor U2511 ( n347, my_IIR_filter_firBlock_left_firStep[187], my_IIR_filter_firBlock_left_multProducts[27] );
xor U2512 ( my_IIR_filter_firBlock_left_N250, n348, n2436 );
xor U2513 ( n348, my_IIR_filter_firBlock_left_firStep[57], my_IIR_filter_firBlock_left_multProducts[86] );
xor U2514 ( my_IIR_filter_firBlock_left_N26, n349, n1182 );
xor U2515 ( n349, my_IIR_filter_firBlock_left_firStep[281], my_IIR_filter_firBlock_left_multProducts[86] );
xor U2516 ( my_IIR_filter_firBlock_left_N189, n2175, n2174 );
xor U2517 ( n2174, my_IIR_filter_firBlock_left_multProducts[58], my_IIR_filter_firBlock_left_firStep[124] );
xor U2518 ( my_IIR_filter_firBlock_left_N93, n1599, n1598 );
xor U2519 ( n1598, my_IIR_filter_firBlock_left_multProducts[58], my_IIR_filter_firBlock_left_firStep[220] );
xor U2520 ( my_IIR_filter_firBlock_left_N220, n350, n2308 );
xor U2521 ( n350, my_IIR_filter_firBlock_left_firStep[91], my_IIR_filter_firBlock_left_multProducts[58] );
xor U2522 ( my_IIR_filter_firBlock_left_N60, n351, n1457 );
xor U2523 ( n351, my_IIR_filter_firBlock_left_firStep[251], my_IIR_filter_firBlock_left_multProducts[58] );
xor U2524 ( my_IIR_filter_firBlock_left_N287, n2607, n2605 );
xnor U2525 ( n2605, n526, my_IIR_filter_firBlock_left_firStep[30] );
xor U2526 ( my_IIR_filter_firBlock_right_N186, n352, n3505 );
xor U2527 ( n352, my_IIR_filter_firBlock_right_firStep[25], my_IIR_filter_firBlock_right_multProducts[25] );
xor U2528 ( my_IIR_filter_firBlock_right_N60, n353, n2776 );
xor U2529 ( n353, my_IIR_filter_firBlock_right_firStep[89], my_IIR_filter_firBlock_right_multProducts[89] );
xor U2530 ( my_IIR_filter_firBlock_right_N120, n354, n3309 );
xor U2531 ( n354, my_IIR_filter_firBlock_right_firStep[54], my_IIR_filter_firBlock_right_multProducts[54] );
xor U2532 ( my_IIR_filter_firBlock_left_N249, n2432, n2431 );
xor U2533 ( my_IIR_filter_firBlock_left_N25, n1178, n1177 );
xor U2534 ( my_IIR_filter_firBlock_left_N155, n2028, n2027 );
xor U2535 ( n2027, my_IIR_filter_firBlock_left_multProducts[26], my_IIR_filter_firBlock_left_firStep[154] );
xor U2536 ( my_IIR_filter_firBlock_left_N123, n1892, n1891 );
xor U2537 ( n1891, my_IIR_filter_firBlock_left_multProducts[26], my_IIR_filter_firBlock_left_firStep[186] );
xor U2538 ( my_IIR_filter_firBlock_left_N219, n2304, n2303 );
xor U2539 ( n2303, my_IIR_filter_firBlock_left_multProducts[57], my_IIR_filter_firBlock_left_firStep[90] );
xor U2540 ( my_IIR_filter_firBlock_left_N59, n1453, n1452 );
xor U2541 ( n1452, my_IIR_filter_firBlock_left_multProducts[57], my_IIR_filter_firBlock_left_firStep[250] );
xor U2542 ( my_IIR_filter_firBlock_left_N188, n355, n2170 );
xor U2543 ( n355, my_IIR_filter_firBlock_left_firStep[123], my_IIR_filter_firBlock_left_multProducts[57] );
xor U2544 ( my_IIR_filter_firBlock_left_N92, n356, n1594 );
xor U2545 ( n356, my_IIR_filter_firBlock_left_firStep[219], my_IIR_filter_firBlock_left_multProducts[57] );
xor U2546 ( n3500, my_IIR_filter_firBlock_right_multProducts[24], my_IIR_filter_firBlock_right_firStep[24] );
xnor U2547 ( my_IIR_filter_firBlock_left_N286, n2598, n2601 );
xnor U2548 ( n2598, my_IIR_filter_firBlock_left_firStep[29], n549 );
xor U2549 ( my_IIR_filter_firBlock_right_N59, n2772, n2771 );
xor U2550 ( n2771, my_IIR_filter_firBlock_right_multProducts[88], my_IIR_filter_firBlock_right_firStep[88] );
xor U2551 ( my_IIR_filter_firBlock_left_N154, n357, n2023 );
xor U2552 ( n357, my_IIR_filter_firBlock_left_firStep[153], my_IIR_filter_firBlock_left_multProducts[25] );
xor U2553 ( my_IIR_filter_firBlock_left_N122, n358, n1887 );
xor U2554 ( n358, my_IIR_filter_firBlock_left_firStep[185], my_IIR_filter_firBlock_left_multProducts[25] );
xor U2555 ( my_IIR_filter_firBlock_left_N187, n2166, n2165 );
xor U2556 ( n2165, my_IIR_filter_firBlock_left_multProducts[56], my_IIR_filter_firBlock_left_firStep[122] );
xor U2557 ( my_IIR_filter_firBlock_left_N91, n1590, n1589 );
xor U2558 ( n1589, my_IIR_filter_firBlock_left_multProducts[56], my_IIR_filter_firBlock_left_firStep[218] );
xor U2559 ( my_IIR_filter_firBlock_left_N218, n359, n2299 );
xor U2560 ( n359, my_IIR_filter_firBlock_left_firStep[89], my_IIR_filter_firBlock_left_multProducts[56] );
xor U2561 ( my_IIR_filter_firBlock_left_N58, n360, n1448 );
xor U2562 ( n360, my_IIR_filter_firBlock_left_firStep[249], my_IIR_filter_firBlock_left_multProducts[56] );
xor U2563 ( my_IIR_filter_firBlock_left_N248, n361, n2427 );
xor U2564 ( n361, my_IIR_filter_firBlock_left_firStep[55], my_IIR_filter_firBlock_left_multProducts[84] );
xor U2565 ( my_IIR_filter_firBlock_left_N24, n362, n1173 );
xor U2566 ( n362, my_IIR_filter_firBlock_left_firStep[279], my_IIR_filter_firBlock_left_multProducts[84] );
xor U2567 ( my_IIR_filter_firBlock_right_N184, n363, n3496 );
xor U2568 ( n363, my_IIR_filter_firBlock_right_firStep[23], my_IIR_filter_firBlock_right_multProducts[23] );
xor U2569 ( my_IIR_filter_firBlock_left_N285, n2594, n2593 );
xnor U2570 ( n2593, n526, my_IIR_filter_firBlock_left_firStep[28] );
xor U2571 ( my_IIR_filter_firBlock_right_N58, n364, n2767 );
xor U2572 ( n364, my_IIR_filter_firBlock_right_firStep[87], my_IIR_filter_firBlock_right_multProducts[87] );
xor U2573 ( n2422, my_IIR_filter_firBlock_left_multProducts[83], my_IIR_filter_firBlock_left_firStep[54] );
xor U2574 ( n1168, my_IIR_filter_firBlock_left_multProducts[83], my_IIR_filter_firBlock_left_firStep[278] );
xor U2575 ( my_IIR_filter_firBlock_right_N118, n365, n3300 );
xor U2576 ( n365, my_IIR_filter_firBlock_right_firStep[52], my_IIR_filter_firBlock_right_multProducts[52] );
xor U2577 ( my_IIR_filter_firBlock_left_N153, n2019, n2018 );
xor U2578 ( n2018, my_IIR_filter_firBlock_left_multProducts[24], my_IIR_filter_firBlock_left_firStep[152] );
xor U2579 ( my_IIR_filter_firBlock_left_N121, n1883, n1882 );
xor U2580 ( n1882, my_IIR_filter_firBlock_left_multProducts[24], my_IIR_filter_firBlock_left_firStep[184] );
xor U2581 ( n3295, my_IIR_filter_firBlock_right_multProducts[51], my_IIR_filter_firBlock_right_firStep[51] );
xor U2582 ( n3491, my_IIR_filter_firBlock_right_multProducts[22], my_IIR_filter_firBlock_right_firStep[22] );
xor U2583 ( my_IIR_filter_firBlock_left_N217, n2295, n2294 );
xor U2584 ( n2294, my_IIR_filter_firBlock_left_multProducts[55], my_IIR_filter_firBlock_left_firStep[88] );
xor U2585 ( my_IIR_filter_firBlock_left_N57, n1444, n1443 );
xor U2586 ( n1443, my_IIR_filter_firBlock_left_multProducts[55], my_IIR_filter_firBlock_left_firStep[248] );
xor U2587 ( my_IIR_filter_firBlock_left_N186, n366, n2161 );
xor U2588 ( n366, my_IIR_filter_firBlock_left_firStep[121], my_IIR_filter_firBlock_left_multProducts[55] );
xor U2589 ( my_IIR_filter_firBlock_left_N90, n367, n1585 );
xor U2590 ( n367, my_IIR_filter_firBlock_left_firStep[217], my_IIR_filter_firBlock_left_multProducts[55] );
xnor U2591 ( my_IIR_filter_firBlock_left_N284, n2588, n2589 );
xnor U2592 ( n2588, my_IIR_filter_firBlock_left_firStep[27], n549 );
xor U2593 ( my_IIR_filter_firBlock_right_N57, n2763, n2762 );
xor U2594 ( n2762, my_IIR_filter_firBlock_right_multProducts[86], my_IIR_filter_firBlock_right_firStep[86] );
xor U2595 ( my_IIR_filter_firBlock_left_N246, n368, n2418 );
xor U2596 ( n368, my_IIR_filter_firBlock_left_firStep[53], my_IIR_filter_firBlock_left_multProducts[82] );
xor U2597 ( my_IIR_filter_firBlock_left_N22, n369, n1164 );
xor U2598 ( n369, my_IIR_filter_firBlock_left_firStep[277], my_IIR_filter_firBlock_left_multProducts[82] );
xor U2599 ( my_IIR_filter_firBlock_right_N182, n370, n3487 );
xor U2600 ( n370, my_IIR_filter_firBlock_right_firStep[21], my_IIR_filter_firBlock_right_multProducts[21] );
xor U2601 ( my_IIR_filter_firBlock_left_N152, n371, n2014 );
xor U2602 ( n371, my_IIR_filter_firBlock_left_firStep[151], my_IIR_filter_firBlock_left_multProducts[23] );
xor U2603 ( my_IIR_filter_firBlock_left_N120, n372, n1878 );
xor U2604 ( n372, my_IIR_filter_firBlock_left_firStep[183], my_IIR_filter_firBlock_left_multProducts[23] );
xor U2605 ( my_IIR_filter_firBlock_left_N185, n2157, n2156 );
xor U2606 ( n2156, my_IIR_filter_firBlock_left_multProducts[54], my_IIR_filter_firBlock_left_firStep[120] );
xor U2607 ( my_IIR_filter_firBlock_left_N89, n1581, n1580 );
xor U2608 ( n1580, my_IIR_filter_firBlock_left_multProducts[54], my_IIR_filter_firBlock_left_firStep[216] );
xor U2609 ( my_IIR_filter_firBlock_right_N116, n373, n3291 );
xor U2610 ( n373, my_IIR_filter_firBlock_right_firStep[50], my_IIR_filter_firBlock_right_multProducts[50] );
xor U2611 ( my_IIR_filter_firBlock_left_N216, n374, n2290 );
xor U2612 ( n374, my_IIR_filter_firBlock_left_firStep[87], my_IIR_filter_firBlock_left_multProducts[54] );
xor U2613 ( my_IIR_filter_firBlock_left_N56, n375, n1439 );
xor U2614 ( n375, my_IIR_filter_firBlock_left_firStep[247], my_IIR_filter_firBlock_left_multProducts[54] );
xor U2615 ( my_IIR_filter_firBlock_left_N283, n2584, n2583 );
xnor U2616 ( n2583, n526, my_IIR_filter_firBlock_left_firStep[26] );
xor U2617 ( my_IIR_filter_firBlock_left_N245, n2414, n2413 );
xor U2618 ( n2413, my_IIR_filter_firBlock_left_multProducts[81], my_IIR_filter_firBlock_left_firStep[52] );
xor U2619 ( my_IIR_filter_firBlock_left_N21, n1160, n1159 );
xor U2620 ( n1159, my_IIR_filter_firBlock_left_multProducts[81], my_IIR_filter_firBlock_left_firStep[276] );
xor U2621 ( n3482, my_IIR_filter_firBlock_right_multProducts[20], my_IIR_filter_firBlock_right_firStep[20] );
xor U2622 ( n3284, my_IIR_filter_firBlock_right_multProducts[49], my_IIR_filter_firBlock_right_firStep[49] );
xor U2623 ( my_IIR_filter_firBlock_right_N56, n376, n2758 );
xor U2624 ( n376, my_IIR_filter_firBlock_right_firStep[85], my_IIR_filter_firBlock_right_multProducts[85] );
xor U2625 ( my_IIR_filter_firBlock_left_N151, n2010, n2009 );
xor U2626 ( n2009, my_IIR_filter_firBlock_left_multProducts[22], my_IIR_filter_firBlock_left_firStep[150] );
xor U2627 ( my_IIR_filter_firBlock_left_N119, n1874, n1873 );
xor U2628 ( n1873, my_IIR_filter_firBlock_left_multProducts[22], my_IIR_filter_firBlock_left_firStep[182] );
xor U2629 ( my_IIR_filter_firBlock_left_N215, n2286, n2285 );
xor U2630 ( n2285, my_IIR_filter_firBlock_left_multProducts[53], my_IIR_filter_firBlock_left_firStep[86] );
xor U2631 ( my_IIR_filter_firBlock_left_N55, n1435, n1434 );
xor U2632 ( n1434, my_IIR_filter_firBlock_left_multProducts[53], my_IIR_filter_firBlock_left_firStep[246] );
xor U2633 ( my_IIR_filter_firBlock_left_N184, n377, n2152 );
xor U2634 ( n377, my_IIR_filter_firBlock_left_firStep[119], my_IIR_filter_firBlock_left_multProducts[53] );
xor U2635 ( my_IIR_filter_firBlock_left_N88, n378, n1576 );
xor U2636 ( n378, my_IIR_filter_firBlock_left_firStep[215], my_IIR_filter_firBlock_left_multProducts[53] );
xor U2637 ( my_IIR_filter_firBlock_right_N180, n379, n3478 );
xor U2638 ( n379, my_IIR_filter_firBlock_right_firStep[19], my_IIR_filter_firBlock_right_multProducts[19] );
xnor U2639 ( my_IIR_filter_firBlock_left_N282, n2578, n2579 );
xnor U2640 ( n2578, my_IIR_filter_firBlock_left_firStep[25], n549 );
xor U2641 ( my_IIR_filter_firBlock_left_N244, n380, n2409 );
xor U2642 ( n380, my_IIR_filter_firBlock_left_firStep[51], my_IIR_filter_firBlock_left_multProducts[80] );
xor U2643 ( my_IIR_filter_firBlock_left_N20, n381, n1155 );
xor U2644 ( n381, my_IIR_filter_firBlock_left_firStep[275], my_IIR_filter_firBlock_left_multProducts[80] );
xor U2645 ( my_IIR_filter_firBlock_right_N55, n2754, n2753 );
xor U2646 ( n2753, my_IIR_filter_firBlock_right_multProducts[84], my_IIR_filter_firBlock_right_firStep[84] );
xor U2647 ( my_IIR_filter_firBlock_right_N114, n382, n3280 );
xor U2648 ( n382, my_IIR_filter_firBlock_right_firStep[48], my_IIR_filter_firBlock_right_multProducts[48] );
xor U2649 ( my_IIR_filter_firBlock_left_N150, n383, n2005 );
xor U2650 ( n383, my_IIR_filter_firBlock_left_firStep[149], my_IIR_filter_firBlock_left_multProducts[21] );
xor U2651 ( my_IIR_filter_firBlock_left_N118, n384, n1869 );
xor U2652 ( n384, my_IIR_filter_firBlock_left_firStep[181], my_IIR_filter_firBlock_left_multProducts[21] );
xor U2653 ( my_IIR_filter_firBlock_left_N183, n2148, n2147 );
xor U2654 ( n2147, my_IIR_filter_firBlock_left_multProducts[52], my_IIR_filter_firBlock_left_firStep[118] );
xor U2655 ( my_IIR_filter_firBlock_left_N87, n1572, n1571 );
xor U2656 ( n1571, my_IIR_filter_firBlock_left_multProducts[52], my_IIR_filter_firBlock_left_firStep[214] );
xor U2657 ( my_IIR_filter_firBlock_left_N214, n385, n2281 );
xor U2658 ( n385, my_IIR_filter_firBlock_left_firStep[85], my_IIR_filter_firBlock_left_multProducts[52] );
xor U2659 ( my_IIR_filter_firBlock_left_N54, n386, n1430 );
xor U2660 ( n386, my_IIR_filter_firBlock_left_firStep[245], my_IIR_filter_firBlock_left_multProducts[52] );
xor U2661 ( my_IIR_filter_firBlock_left_N243, n2403, n2402 );
xor U2662 ( n2402, my_IIR_filter_firBlock_left_multProducts[79], my_IIR_filter_firBlock_left_firStep[50] );
xor U2663 ( my_IIR_filter_firBlock_left_N19, n1149, n1148 );
xor U2664 ( n1148, my_IIR_filter_firBlock_left_multProducts[79], my_IIR_filter_firBlock_left_firStep[274] );
xor U2665 ( n3471, my_IIR_filter_firBlock_right_multProducts[18], my_IIR_filter_firBlock_right_firStep[18] );
xor U2666 ( my_IIR_filter_firBlock_left_N281, n2574, n2573 );
xor U2667 ( n2573, my_IIR_filter_firBlock_left_multProducts[114], my_IIR_filter_firBlock_left_firStep[24] );
xor U2668 ( my_IIR_filter_firBlock_right_N54, n387, n2749 );
xor U2669 ( n387, my_IIR_filter_firBlock_right_firStep[83], my_IIR_filter_firBlock_right_multProducts[83] );
xor U2670 ( my_IIR_filter_firBlock_left_N149, n2001, n2000 );
xor U2671 ( n2000, my_IIR_filter_firBlock_left_multProducts[20], my_IIR_filter_firBlock_left_firStep[148] );
xor U2672 ( my_IIR_filter_firBlock_left_N117, n1865, n1864 );
xor U2673 ( n1864, my_IIR_filter_firBlock_left_multProducts[20], my_IIR_filter_firBlock_left_firStep[180] );
xor U2674 ( my_IIR_filter_firBlock_left_N213, n2277, n2276 );
xor U2675 ( n2276, my_IIR_filter_firBlock_left_multProducts[51], my_IIR_filter_firBlock_left_firStep[84] );
xor U2676 ( my_IIR_filter_firBlock_left_N53, n1426, n1425 );
xor U2677 ( n1425, my_IIR_filter_firBlock_left_multProducts[51], my_IIR_filter_firBlock_left_firStep[244] );
xor U2678 ( my_IIR_filter_firBlock_left_N182, n388, n2143 );
xor U2679 ( n388, my_IIR_filter_firBlock_left_firStep[117], my_IIR_filter_firBlock_left_multProducts[51] );
xor U2680 ( my_IIR_filter_firBlock_left_N86, n389, n1567 );
xor U2681 ( n389, my_IIR_filter_firBlock_left_firStep[213], my_IIR_filter_firBlock_left_multProducts[51] );
xor U2682 ( my_IIR_filter_firBlock_right_N178, n390, n3467 );
xor U2683 ( n390, my_IIR_filter_firBlock_right_firStep[17], my_IIR_filter_firBlock_right_multProducts[17] );
xor U2684 ( my_IIR_filter_firBlock_right_N112, n391, n3271 );
xor U2685 ( n391, my_IIR_filter_firBlock_right_firStep[46], my_IIR_filter_firBlock_right_multProducts[46] );
xor U2686 ( my_IIR_filter_firBlock_left_N242, n392, n2398 );
xor U2687 ( n392, my_IIR_filter_firBlock_left_firStep[49], my_IIR_filter_firBlock_left_multProducts[78] );
xor U2688 ( my_IIR_filter_firBlock_left_N18, n393, n1144 );
xor U2689 ( n393, my_IIR_filter_firBlock_left_firStep[273], my_IIR_filter_firBlock_left_multProducts[78] );
xnor U2690 ( my_IIR_filter_firBlock_left_N280, n2568, n2569 );
xnor U2691 ( n2568, my_IIR_filter_firBlock_left_firStep[23], my_IIR_filter_firBlock_left_multProducts[113] );
xor U2692 ( my_IIR_filter_firBlock_right_N53, n2745, n2744 );
xor U2693 ( n2744, my_IIR_filter_firBlock_right_multProducts[82], my_IIR_filter_firBlock_right_firStep[82] );
xor U2694 ( n3462, my_IIR_filter_firBlock_right_multProducts[16], my_IIR_filter_firBlock_right_firStep[16] );
xor U2695 ( n3266, my_IIR_filter_firBlock_right_multProducts[45], my_IIR_filter_firBlock_right_firStep[45] );
xor U2696 ( my_IIR_filter_firBlock_left_N148, n394, n1996 );
xor U2697 ( n394, my_IIR_filter_firBlock_left_firStep[147], my_IIR_filter_firBlock_left_multProducts[19] );
xor U2698 ( my_IIR_filter_firBlock_left_N116, n395, n1860 );
xor U2699 ( n395, my_IIR_filter_firBlock_left_firStep[179], my_IIR_filter_firBlock_left_multProducts[19] );
xor U2700 ( my_IIR_filter_firBlock_left_N181, n2139, n2138 );
xor U2701 ( n2138, my_IIR_filter_firBlock_left_multProducts[50], my_IIR_filter_firBlock_left_firStep[116] );
xor U2702 ( my_IIR_filter_firBlock_left_N85, n1563, n1562 );
xor U2703 ( n1562, my_IIR_filter_firBlock_left_multProducts[50], my_IIR_filter_firBlock_left_firStep[212] );
xor U2704 ( my_IIR_filter_firBlock_left_N212, n396, n2272 );
xor U2705 ( n396, my_IIR_filter_firBlock_left_firStep[83], my_IIR_filter_firBlock_left_multProducts[50] );
xor U2706 ( my_IIR_filter_firBlock_left_N52, n397, n1421 );
xor U2707 ( n397, my_IIR_filter_firBlock_left_firStep[243], my_IIR_filter_firBlock_left_multProducts[50] );
xor U2708 ( my_IIR_filter_firBlock_left_N241, n2394, n2393 );
xor U2709 ( n2393, my_IIR_filter_firBlock_left_multProducts[77], my_IIR_filter_firBlock_left_firStep[48] );
xor U2710 ( my_IIR_filter_firBlock_left_N17, n1140, n1139 );
xor U2711 ( n1139, my_IIR_filter_firBlock_left_multProducts[77], my_IIR_filter_firBlock_left_firStep[272] );
xor U2712 ( my_IIR_filter_firBlock_left_N279, n2564, n2563 );
xor U2713 ( n2563, my_IIR_filter_firBlock_left_multProducts[112], my_IIR_filter_firBlock_left_firStep[22] );
xor U2714 ( my_IIR_filter_firBlock_right_N52, n398, n2740 );
xor U2715 ( n398, my_IIR_filter_firBlock_right_firStep[81], my_IIR_filter_firBlock_right_multProducts[81] );
xor U2716 ( my_IIR_filter_firBlock_left_N147, n1990, n1989 );
xor U2717 ( n1989, my_IIR_filter_firBlock_left_multProducts[18], my_IIR_filter_firBlock_left_firStep[146] );
xor U2718 ( my_IIR_filter_firBlock_left_N115, n1854, n1853 );
xor U2719 ( n1853, my_IIR_filter_firBlock_left_multProducts[18], my_IIR_filter_firBlock_left_firStep[178] );
xor U2720 ( my_IIR_filter_firBlock_right_N176, n399, n3458 );
xor U2721 ( n399, my_IIR_filter_firBlock_right_firStep[15], my_IIR_filter_firBlock_right_multProducts[15] );
xor U2722 ( my_IIR_filter_firBlock_left_N211, n2266, n2265 );
xor U2723 ( n2265, my_IIR_filter_firBlock_left_multProducts[49], my_IIR_filter_firBlock_left_firStep[82] );
xor U2724 ( my_IIR_filter_firBlock_left_N51, n1415, n1414 );
xor U2725 ( n1414, my_IIR_filter_firBlock_left_multProducts[49], my_IIR_filter_firBlock_left_firStep[242] );
xor U2726 ( my_IIR_filter_firBlock_right_N110, n400, n3262 );
xor U2727 ( n400, my_IIR_filter_firBlock_right_firStep[44], my_IIR_filter_firBlock_right_multProducts[44] );
xor U2728 ( my_IIR_filter_firBlock_left_N180, n401, n2134 );
xor U2729 ( n401, my_IIR_filter_firBlock_left_firStep[115], my_IIR_filter_firBlock_left_multProducts[49] );
xor U2730 ( my_IIR_filter_firBlock_left_N84, n402, n1558 );
xor U2731 ( n402, my_IIR_filter_firBlock_left_firStep[211], my_IIR_filter_firBlock_left_multProducts[49] );
xor U2732 ( my_IIR_filter_firBlock_left_N240, n403, n2389 );
xor U2733 ( n403, my_IIR_filter_firBlock_left_firStep[47], my_IIR_filter_firBlock_left_multProducts[76] );
xor U2734 ( my_IIR_filter_firBlock_left_N16, n404, n1135 );
xor U2735 ( n404, my_IIR_filter_firBlock_left_firStep[271], my_IIR_filter_firBlock_left_multProducts[76] );
xnor U2736 ( my_IIR_filter_firBlock_left_N278, n2558, n2559 );
xnor U2737 ( n2558, my_IIR_filter_firBlock_left_firStep[21], my_IIR_filter_firBlock_left_multProducts[111] );
xor U2738 ( my_IIR_filter_firBlock_right_N51, n2734, n2733 );
xor U2739 ( n2733, my_IIR_filter_firBlock_right_multProducts[80], my_IIR_filter_firBlock_right_firStep[80] );
xor U2740 ( n3453, my_IIR_filter_firBlock_right_multProducts[14], my_IIR_filter_firBlock_right_firStep[14] );
xor U2741 ( my_IIR_filter_firBlock_left_N239, n2385, n2384 );
xor U2742 ( n2384, my_IIR_filter_firBlock_left_multProducts[75], my_IIR_filter_firBlock_left_firStep[46] );
xor U2743 ( my_IIR_filter_firBlock_left_N15, n1131, n1130 );
xor U2744 ( n1130, my_IIR_filter_firBlock_left_multProducts[75], my_IIR_filter_firBlock_left_firStep[270] );
xor U2745 ( my_IIR_filter_firBlock_left_N146, n405, n1985 );
xor U2746 ( n405, my_IIR_filter_firBlock_left_firStep[145], my_IIR_filter_firBlock_left_multProducts[17] );
xor U2747 ( my_IIR_filter_firBlock_left_N114, n406, n1849 );
xor U2748 ( n406, my_IIR_filter_firBlock_left_firStep[177], my_IIR_filter_firBlock_left_multProducts[17] );
xor U2749 ( my_IIR_filter_firBlock_left_N179, n2128, n2127 );
xor U2750 ( n2127, my_IIR_filter_firBlock_left_multProducts[48], my_IIR_filter_firBlock_left_firStep[114] );
xor U2751 ( my_IIR_filter_firBlock_left_N83, n1552, n1551 );
xor U2752 ( n1551, my_IIR_filter_firBlock_left_multProducts[48], my_IIR_filter_firBlock_left_firStep[210] );
xor U2753 ( my_IIR_filter_firBlock_left_N210, n407, n2261 );
xor U2754 ( n407, my_IIR_filter_firBlock_left_firStep[81], my_IIR_filter_firBlock_left_multProducts[48] );
xor U2755 ( my_IIR_filter_firBlock_left_N50, n408, n1410 );
xor U2756 ( n408, my_IIR_filter_firBlock_left_firStep[241], my_IIR_filter_firBlock_left_multProducts[48] );
xor U2757 ( my_IIR_filter_firBlock_left_N277, n2554, n2553 );
xor U2758 ( n2553, my_IIR_filter_firBlock_left_multProducts[110], my_IIR_filter_firBlock_left_firStep[20] );
xor U2759 ( my_IIR_filter_firBlock_right_N108, n409, n3253 );
xor U2760 ( n409, my_IIR_filter_firBlock_right_firStep[42], my_IIR_filter_firBlock_right_multProducts[42] );
xor U2761 ( my_IIR_filter_firBlock_right_N174, n410, n3449 );
xor U2762 ( n410, my_IIR_filter_firBlock_right_firStep[13], my_IIR_filter_firBlock_right_multProducts[13] );
xor U2763 ( my_IIR_filter_firBlock_right_N50, n411, n2729 );
xor U2764 ( n411, my_IIR_filter_firBlock_right_firStep[79], my_IIR_filter_firBlock_right_multProducts[79] );
xor U2765 ( my_IIR_filter_firBlock_left_N145, n1981, n1980 );
xor U2766 ( n1980, my_IIR_filter_firBlock_left_multProducts[16], my_IIR_filter_firBlock_left_firStep[144] );
xor U2767 ( my_IIR_filter_firBlock_left_N113, n1845, n1844 );
xor U2768 ( n1844, my_IIR_filter_firBlock_left_multProducts[16], my_IIR_filter_firBlock_left_firStep[176] );
xor U2769 ( my_IIR_filter_firBlock_left_N209, n2257, n2256 );
xor U2770 ( n2256, my_IIR_filter_firBlock_left_multProducts[47], my_IIR_filter_firBlock_left_firStep[80] );
xor U2771 ( my_IIR_filter_firBlock_left_N49, n1406, n1405 );
xor U2772 ( n1405, my_IIR_filter_firBlock_left_multProducts[47], my_IIR_filter_firBlock_left_firStep[240] );
xor U2773 ( n3444, my_IIR_filter_firBlock_right_multProducts[12], my_IIR_filter_firBlock_right_firStep[12] );
xor U2774 ( my_IIR_filter_firBlock_left_N178, n412, n2123 );
xor U2775 ( n412, my_IIR_filter_firBlock_left_firStep[113], my_IIR_filter_firBlock_left_multProducts[47] );
xor U2776 ( my_IIR_filter_firBlock_left_N82, n413, n1547 );
xor U2777 ( n413, my_IIR_filter_firBlock_left_firStep[209], my_IIR_filter_firBlock_left_multProducts[47] );
xor U2778 ( my_IIR_filter_firBlock_left_N238, n414, n2380 );
xor U2779 ( n414, my_IIR_filter_firBlock_left_firStep[45], my_IIR_filter_firBlock_left_multProducts[74] );
xor U2780 ( my_IIR_filter_firBlock_left_N14, n415, n1126 );
xor U2781 ( n415, my_IIR_filter_firBlock_left_firStep[269], my_IIR_filter_firBlock_left_multProducts[74] );
xnor U2782 ( my_IIR_filter_firBlock_left_N276, n2546, n2549 );
xnor U2783 ( n2546, my_IIR_filter_firBlock_left_firStep[19], my_IIR_filter_firBlock_left_multProducts[109] );
xor U2784 ( my_IIR_filter_firBlock_right_N49, n2725, n2724 );
xor U2785 ( n2724, my_IIR_filter_firBlock_right_multProducts[78], my_IIR_filter_firBlock_right_firStep[78] );
xor U2786 ( my_IIR_filter_firBlock_left_N144, n416, n1976 );
xor U2787 ( n416, my_IIR_filter_firBlock_left_firStep[143], my_IIR_filter_firBlock_left_multProducts[15] );
xor U2788 ( my_IIR_filter_firBlock_left_N112, n417, n1840 );
xor U2789 ( n417, my_IIR_filter_firBlock_left_firStep[175], my_IIR_filter_firBlock_left_multProducts[15] );
xor U2790 ( my_IIR_filter_firBlock_left_N177, n2119, n2118 );
xor U2791 ( n2118, my_IIR_filter_firBlock_left_multProducts[46], my_IIR_filter_firBlock_left_firStep[112] );
xor U2792 ( my_IIR_filter_firBlock_left_N81, n1543, n1542 );
xor U2793 ( n1542, my_IIR_filter_firBlock_left_multProducts[46], my_IIR_filter_firBlock_left_firStep[208] );
xor U2794 ( my_IIR_filter_firBlock_left_N208, n418, n2252 );
xor U2795 ( n418, my_IIR_filter_firBlock_left_firStep[79], my_IIR_filter_firBlock_left_multProducts[46] );
xor U2796 ( my_IIR_filter_firBlock_left_N48, n419, n1401 );
xor U2797 ( n419, my_IIR_filter_firBlock_left_firStep[239], my_IIR_filter_firBlock_left_multProducts[46] );
xor U2798 ( my_IIR_filter_firBlock_right_N106, n420, n3355 );
xor U2799 ( n420, my_IIR_filter_firBlock_right_firStep[40], my_IIR_filter_firBlock_right_multProducts[40] );
xor U2800 ( my_IIR_filter_firBlock_right_N172, n421, n3440 );
xor U2801 ( n421, my_IIR_filter_firBlock_right_firStep[11], my_IIR_filter_firBlock_right_multProducts[11] );
xor U2802 ( my_IIR_filter_firBlock_left_N275, n2542, n2541 );
xor U2803 ( n2541, my_IIR_filter_firBlock_left_multProducts[108], my_IIR_filter_firBlock_left_firStep[18] );
xor U2804 ( my_IIR_filter_firBlock_left_N143, n1972, n1971 );
xor U2805 ( n1971, my_IIR_filter_firBlock_left_multProducts[14], my_IIR_filter_firBlock_left_firStep[142] );
xor U2806 ( my_IIR_filter_firBlock_left_N111, n1836, n1835 );
xor U2807 ( n1835, my_IIR_filter_firBlock_left_multProducts[14], my_IIR_filter_firBlock_left_firStep[174] );
xor U2808 ( my_IIR_filter_firBlock_right_N48, n422, n2720 );
xor U2809 ( n422, my_IIR_filter_firBlock_right_firStep[77], my_IIR_filter_firBlock_right_multProducts[77] );
xor U2810 ( n3353, my_IIR_filter_firBlock_right_multProducts[39], my_IIR_filter_firBlock_right_firStep[39] );
xor U2811 ( my_IIR_filter_firBlock_left_N236, n423, n2371 );
xor U2812 ( n423, my_IIR_filter_firBlock_left_firStep[43], my_IIR_filter_firBlock_left_multProducts[72] );
xor U2813 ( my_IIR_filter_firBlock_left_N12, n424, n1117 );
xor U2814 ( n424, my_IIR_filter_firBlock_left_firStep[267], my_IIR_filter_firBlock_left_multProducts[72] );
xor U2815 ( n3435, my_IIR_filter_firBlock_right_multProducts[10], my_IIR_filter_firBlock_right_firStep[10] );
xor U2816 ( my_IIR_filter_firBlock_left_N207, n2248, n2247 );
xor U2817 ( n2247, my_IIR_filter_firBlock_left_multProducts[45], my_IIR_filter_firBlock_left_firStep[78] );
xor U2818 ( my_IIR_filter_firBlock_left_N47, n1397, n1396 );
xor U2819 ( n1396, my_IIR_filter_firBlock_left_multProducts[45], my_IIR_filter_firBlock_left_firStep[238] );
xor U2820 ( my_IIR_filter_firBlock_left_N176, n425, n2114 );
xor U2821 ( n425, my_IIR_filter_firBlock_left_firStep[111], my_IIR_filter_firBlock_left_multProducts[45] );
xor U2822 ( my_IIR_filter_firBlock_left_N80, n426, n1538 );
xor U2823 ( n426, my_IIR_filter_firBlock_left_firStep[207], my_IIR_filter_firBlock_left_multProducts[45] );
xnor U2824 ( my_IIR_filter_firBlock_left_N274, n2536, n2537 );
xnor U2825 ( n2536, my_IIR_filter_firBlock_left_firStep[17], my_IIR_filter_firBlock_left_multProducts[107] );
xor U2826 ( my_IIR_filter_firBlock_right_N47, n2716, n2715 );
xor U2827 ( n2715, my_IIR_filter_firBlock_right_multProducts[76], my_IIR_filter_firBlock_right_firStep[76] );
xor U2828 ( my_IIR_filter_firBlock_left_N235, n2367, n2366 );
xor U2829 ( n2366, my_IIR_filter_firBlock_left_multProducts[71], my_IIR_filter_firBlock_left_firStep[42] );
xor U2830 ( my_IIR_filter_firBlock_left_N11, n1113, n1112 );
xor U2831 ( n1112, my_IIR_filter_firBlock_left_multProducts[71], my_IIR_filter_firBlock_left_firStep[266] );
xor U2832 ( my_IIR_filter_firBlock_left_N142, n427, n1967 );
xor U2833 ( n427, my_IIR_filter_firBlock_left_firStep[141], my_IIR_filter_firBlock_left_multProducts[13] );
xor U2834 ( my_IIR_filter_firBlock_left_N110, n428, n1831 );
xor U2835 ( n428, my_IIR_filter_firBlock_left_firStep[173], my_IIR_filter_firBlock_left_multProducts[13] );
xor U2836 ( my_IIR_filter_firBlock_right_N170, n429, n3542 );
xor U2837 ( n429, my_IIR_filter_firBlock_right_firStep[9], my_IIR_filter_firBlock_right_multProducts[9] );
xor U2838 ( my_IIR_filter_firBlock_right_N104, n430, n3352 );
xor U2839 ( n430, my_IIR_filter_firBlock_right_firStep[38], my_IIR_filter_firBlock_right_multProducts[38] );
xor U2840 ( my_IIR_filter_firBlock_left_N175, n2110, n2109 );
xor U2841 ( n2109, my_IIR_filter_firBlock_left_multProducts[44], my_IIR_filter_firBlock_left_firStep[110] );
xor U2842 ( my_IIR_filter_firBlock_left_N79, n1534, n1533 );
xor U2843 ( n1533, my_IIR_filter_firBlock_left_multProducts[44], my_IIR_filter_firBlock_left_firStep[206] );
xor U2844 ( my_IIR_filter_firBlock_left_N206, n431, n2243 );
xor U2845 ( n431, my_IIR_filter_firBlock_left_firStep[77], my_IIR_filter_firBlock_left_multProducts[44] );
xor U2846 ( my_IIR_filter_firBlock_left_N46, n432, n1392 );
xor U2847 ( n432, my_IIR_filter_firBlock_left_firStep[237], my_IIR_filter_firBlock_left_multProducts[44] );
xor U2848 ( n3350, my_IIR_filter_firBlock_right_multProducts[37], my_IIR_filter_firBlock_right_firStep[37] );
xor U2849 ( my_IIR_filter_firBlock_left_N273, n2532, n2531 );
xor U2850 ( n2531, my_IIR_filter_firBlock_left_multProducts[106], my_IIR_filter_firBlock_left_firStep[16] );
xor U2851 ( my_IIR_filter_firBlock_left_N141, n1963, n1962 );
xor U2852 ( n1962, my_IIR_filter_firBlock_left_multProducts[12], my_IIR_filter_firBlock_left_firStep[140] );
xor U2853 ( my_IIR_filter_firBlock_left_N109, n1827, n1826 );
xor U2854 ( n1826, my_IIR_filter_firBlock_left_multProducts[12], my_IIR_filter_firBlock_left_firStep[172] );
xor U2855 ( n3540, my_IIR_filter_firBlock_right_multProducts[8], my_IIR_filter_firBlock_right_firStep[8] );
xor U2856 ( my_IIR_filter_firBlock_right_N46, n433, n2711 );
xor U2857 ( n433, my_IIR_filter_firBlock_right_firStep[75], my_IIR_filter_firBlock_right_multProducts[75] );
xor U2858 ( my_IIR_filter_firBlock_left_N234, n434, n2475 );
xor U2859 ( n434, my_IIR_filter_firBlock_left_firStep[41], my_IIR_filter_firBlock_left_multProducts[70] );
xor U2860 ( my_IIR_filter_firBlock_left_N10, n435, n1221 );
xor U2861 ( n435, my_IIR_filter_firBlock_left_firStep[265], my_IIR_filter_firBlock_left_multProducts[70] );
xor U2862 ( my_IIR_filter_firBlock_left_N205, n2239, n2238 );
xor U2863 ( n2238, my_IIR_filter_firBlock_left_multProducts[43], my_IIR_filter_firBlock_left_firStep[76] );
xor U2864 ( my_IIR_filter_firBlock_left_N45, n1388, n1387 );
xor U2865 ( n1387, my_IIR_filter_firBlock_left_multProducts[43], my_IIR_filter_firBlock_left_firStep[236] );
xor U2866 ( my_IIR_filter_firBlock_left_N174, n436, n2105 );
xor U2867 ( n436, my_IIR_filter_firBlock_left_firStep[109], my_IIR_filter_firBlock_left_multProducts[43] );
xor U2868 ( my_IIR_filter_firBlock_left_N78, n437, n1529 );
xor U2869 ( n437, my_IIR_filter_firBlock_left_firStep[205], my_IIR_filter_firBlock_left_multProducts[43] );
xor U2870 ( my_IIR_filter_firBlock_right_N168, n438, n3539 );
xor U2871 ( n438, my_IIR_filter_firBlock_right_firStep[7], my_IIR_filter_firBlock_right_multProducts[7] );
xor U2872 ( my_IIR_filter_firBlock_right_N45, n2707, n2706 );
xor U2873 ( n2706, my_IIR_filter_firBlock_right_multProducts[74], my_IIR_filter_firBlock_right_firStep[74] );
xnor U2874 ( my_IIR_filter_firBlock_left_N272, n2526, n2527 );
xnor U2875 ( n2526, my_IIR_filter_firBlock_left_firStep[15], my_IIR_filter_firBlock_left_multProducts[105] );
xor U2876 ( my_IIR_filter_firBlock_right_N102, n439, n3349 );
xor U2877 ( n439, my_IIR_filter_firBlock_right_firStep[36], my_IIR_filter_firBlock_right_multProducts[36] );
xor U2878 ( my_IIR_filter_firBlock_left_N140, n440, n1958 );
xor U2879 ( n440, my_IIR_filter_firBlock_left_firStep[139], my_IIR_filter_firBlock_left_multProducts[11] );
xor U2880 ( my_IIR_filter_firBlock_left_N108, n441, n1822 );
xor U2881 ( n441, my_IIR_filter_firBlock_left_firStep[171], my_IIR_filter_firBlock_left_multProducts[11] );
xor U2882 ( my_IIR_filter_firBlock_left_N233, n2474, n2473 );
xor U2883 ( my_IIR_filter_firBlock_left_N9, n1220, n1219 );
xor U2884 ( my_IIR_filter_firBlock_left_N173, n2101, n2100 );
xor U2885 ( n2100, my_IIR_filter_firBlock_left_multProducts[42], my_IIR_filter_firBlock_left_firStep[108] );
xor U2886 ( my_IIR_filter_firBlock_left_N77, n1525, n1524 );
xor U2887 ( n1524, my_IIR_filter_firBlock_left_multProducts[42], my_IIR_filter_firBlock_left_firStep[204] );
xor U2888 ( n3347, my_IIR_filter_firBlock_right_multProducts[35], my_IIR_filter_firBlock_right_firStep[35] );
xor U2889 ( my_IIR_filter_firBlock_left_N204, n442, n2234 );
xor U2890 ( n442, my_IIR_filter_firBlock_left_firStep[75], my_IIR_filter_firBlock_left_multProducts[42] );
xor U2891 ( my_IIR_filter_firBlock_left_N44, n443, n1383 );
xor U2892 ( n443, my_IIR_filter_firBlock_left_firStep[235], my_IIR_filter_firBlock_left_multProducts[42] );
xor U2893 ( n3537, my_IIR_filter_firBlock_right_multProducts[6], my_IIR_filter_firBlock_right_firStep[6] );
xor U2894 ( my_IIR_filter_firBlock_left_N139, n1954, n1953 );
xor U2895 ( n1953, my_IIR_filter_firBlock_left_multProducts[10], my_IIR_filter_firBlock_left_firStep[138] );
xor U2896 ( my_IIR_filter_firBlock_left_N107, n1818, n1817 );
xor U2897 ( n1817, my_IIR_filter_firBlock_left_multProducts[10], my_IIR_filter_firBlock_left_firStep[170] );
xor U2898 ( my_IIR_filter_firBlock_left_N271, n2522, n2521 );
xor U2899 ( n2521, my_IIR_filter_firBlock_left_multProducts[104], my_IIR_filter_firBlock_left_firStep[14] );
xor U2900 ( my_IIR_filter_firBlock_left_N232, n444, n2472 );
xor U2901 ( n444, my_IIR_filter_firBlock_left_firStep[39], my_IIR_filter_firBlock_left_multProducts[68] );
xor U2902 ( my_IIR_filter_firBlock_left_N8, n445, n1218 );
xor U2903 ( n445, my_IIR_filter_firBlock_left_firStep[263], my_IIR_filter_firBlock_left_multProducts[68] );
xor U2904 ( my_IIR_filter_firBlock_right_N44, n446, n2702 );
xor U2905 ( n446, my_IIR_filter_firBlock_right_firStep[73], my_IIR_filter_firBlock_right_multProducts[73] );
xor U2906 ( my_IIR_filter_firBlock_right_N166, n447, n3536 );
xor U2907 ( n447, my_IIR_filter_firBlock_right_firStep[5], my_IIR_filter_firBlock_right_multProducts[5] );
xor U2908 ( my_IIR_filter_firBlock_left_N203, n2230, n2229 );
xor U2909 ( n2229, my_IIR_filter_firBlock_left_multProducts[41], my_IIR_filter_firBlock_left_firStep[74] );
xor U2910 ( my_IIR_filter_firBlock_left_N43, n1379, n1378 );
xor U2911 ( n1378, my_IIR_filter_firBlock_left_multProducts[41], my_IIR_filter_firBlock_left_firStep[234] );
xor U2912 ( my_IIR_filter_firBlock_left_N172, n448, n2096 );
xor U2913 ( n448, my_IIR_filter_firBlock_left_firStep[107], my_IIR_filter_firBlock_left_multProducts[41] );
xor U2914 ( my_IIR_filter_firBlock_left_N76, n449, n1520 );
xor U2915 ( n449, my_IIR_filter_firBlock_left_firStep[203], my_IIR_filter_firBlock_left_multProducts[41] );
xor U2916 ( my_IIR_filter_firBlock_right_N100, n450, n3346 );
xor U2917 ( n450, my_IIR_filter_firBlock_right_firStep[34], my_IIR_filter_firBlock_right_multProducts[34] );
xor U2918 ( my_IIR_filter_firBlock_left_N231, n2471, n2470 );
xor U2919 ( n2470, my_IIR_filter_firBlock_left_multProducts[67], my_IIR_filter_firBlock_left_firStep[38] );
xor U2920 ( my_IIR_filter_firBlock_left_N7, n1217, n1216 );
xor U2921 ( n1216, my_IIR_filter_firBlock_left_multProducts[67], my_IIR_filter_firBlock_left_firStep[262] );
xor U2922 ( my_IIR_filter_firBlock_left_N138, n451, n2063 );
xor U2923 ( n451, my_IIR_filter_firBlock_left_firStep[137], my_IIR_filter_firBlock_left_multProducts[9] );
xor U2924 ( my_IIR_filter_firBlock_left_N106, n452, n1925 );
xor U2925 ( n452, my_IIR_filter_firBlock_left_firStep[169], my_IIR_filter_firBlock_left_multProducts[9] );
xor U2926 ( my_IIR_filter_firBlock_right_N43, n2698, n2697 );
xor U2927 ( n2697, my_IIR_filter_firBlock_right_multProducts[72], my_IIR_filter_firBlock_right_firStep[72] );
xnor U2928 ( my_IIR_filter_firBlock_left_N270, n2516, n2517 );
xnor U2929 ( n2516, my_IIR_filter_firBlock_left_firStep[13], my_IIR_filter_firBlock_left_multProducts[103] );
xor U2930 ( n3534, my_IIR_filter_firBlock_right_multProducts[4], my_IIR_filter_firBlock_right_firStep[4] );
xor U2931 ( my_IIR_filter_firBlock_right_N99, n3336, n3335 );
xor U2932 ( n3335, my_IIR_filter_firBlock_right_multProducts[33], my_IIR_filter_firBlock_right_firStep[33] );
xor U2933 ( my_IIR_filter_firBlock_left_N171, n2092, n2091 );
xor U2934 ( n2091, my_IIR_filter_firBlock_left_multProducts[40], my_IIR_filter_firBlock_left_firStep[106] );
xor U2935 ( my_IIR_filter_firBlock_left_N75, n1516, n1515 );
xor U2936 ( n1515, my_IIR_filter_firBlock_left_multProducts[40], my_IIR_filter_firBlock_left_firStep[202] );
xor U2937 ( my_IIR_filter_firBlock_left_N137, n2062, n2061 );
xor U2938 ( n2061, my_IIR_filter_firBlock_left_multProducts[8], my_IIR_filter_firBlock_left_firStep[136] );
xor U2939 ( my_IIR_filter_firBlock_left_N105, n1924, n1923 );
xor U2940 ( n1923, my_IIR_filter_firBlock_left_multProducts[8], my_IIR_filter_firBlock_left_firStep[168] );
xor U2941 ( my_IIR_filter_firBlock_left_N202, n453, n2338 );
xor U2942 ( n453, my_IIR_filter_firBlock_left_firStep[73], my_IIR_filter_firBlock_left_multProducts[40] );
xor U2943 ( my_IIR_filter_firBlock_left_N42, n454, n1487 );
xor U2944 ( n454, my_IIR_filter_firBlock_left_firStep[233], my_IIR_filter_firBlock_left_multProducts[40] );
xor U2945 ( my_IIR_filter_firBlock_left_N269, n2512, n2511 );
xor U2946 ( n2511, my_IIR_filter_firBlock_left_multProducts[102], my_IIR_filter_firBlock_left_firStep[12] );
xor U2947 ( my_IIR_filter_firBlock_left_N230, n455, n2469 );
xor U2948 ( n455, my_IIR_filter_firBlock_left_firStep[37], my_IIR_filter_firBlock_left_multProducts[66] );
xor U2949 ( my_IIR_filter_firBlock_right_N42, n456, n2807 );
xor U2950 ( n456, my_IIR_filter_firBlock_right_firStep[71], my_IIR_filter_firBlock_right_multProducts[71] );
xor U2951 ( my_IIR_filter_firBlock_left_N6, n457, n1215 );
xor U2952 ( n457, my_IIR_filter_firBlock_left_firStep[261], my_IIR_filter_firBlock_left_multProducts[66] );
xor U2953 ( my_IIR_filter_firBlock_right_N164, n458, n3533 );
xor U2954 ( n458, my_IIR_filter_firBlock_right_firStep[3], my_IIR_filter_firBlock_right_multProducts[3] );
xor U2955 ( my_IIR_filter_firBlock_right_N98, n3290, n3289 );
xor U2956 ( my_IIR_filter_firBlock_left_N201, n2337, n2336 );
xor U2957 ( n2336, my_IIR_filter_firBlock_left_multProducts[39], my_IIR_filter_firBlock_left_firStep[72] );
xor U2958 ( my_IIR_filter_firBlock_left_N41, n1486, n1485 );
xor U2959 ( n1485, my_IIR_filter_firBlock_left_multProducts[39], my_IIR_filter_firBlock_left_firStep[232] );
xor U2960 ( my_IIR_filter_firBlock_left_N170, n459, n2201 );
xor U2961 ( n459, my_IIR_filter_firBlock_left_firStep[105], my_IIR_filter_firBlock_left_multProducts[39] );
xor U2962 ( my_IIR_filter_firBlock_left_N74, n460, n1625 );
xor U2963 ( n460, my_IIR_filter_firBlock_left_firStep[201], my_IIR_filter_firBlock_left_multProducts[39] );
xor U2964 ( my_IIR_filter_firBlock_left_N136, n461, n2060 );
xor U2965 ( n461, my_IIR_filter_firBlock_left_firStep[135], my_IIR_filter_firBlock_left_multProducts[7] );
xor U2966 ( my_IIR_filter_firBlock_left_N104, n462, n1922 );
xor U2967 ( n462, my_IIR_filter_firBlock_left_firStep[167], my_IIR_filter_firBlock_left_multProducts[7] );
xor U2968 ( my_IIR_filter_firBlock_left_N229, n2468, n2467 );
xor U2969 ( my_IIR_filter_firBlock_right_N41, n2806, n2805 );
xor U2970 ( n2805, my_IIR_filter_firBlock_right_multProducts[70], my_IIR_filter_firBlock_right_firStep[70] );
xnor U2971 ( my_IIR_filter_firBlock_left_N268, n2506, n2507 );
xnor U2972 ( n2506, my_IIR_filter_firBlock_left_firStep[11], my_IIR_filter_firBlock_left_multProducts[101] );
xor U2973 ( n3522, my_IIR_filter_firBlock_right_multProducts[2], my_IIR_filter_firBlock_right_firStep[2] );
xor U2974 ( my_IIR_filter_firBlock_left_N135, n2059, n2058 );
xor U2975 ( n2058, my_IIR_filter_firBlock_left_multProducts[6], my_IIR_filter_firBlock_left_firStep[134] );
xor U2976 ( my_IIR_filter_firBlock_left_N103, n1921, n1920 );
xor U2977 ( n1920, my_IIR_filter_firBlock_left_multProducts[6], my_IIR_filter_firBlock_left_firStep[166] );
xor U2978 ( my_IIR_filter_firBlock_left_N169, n2200, n2199 );
xor U2979 ( n2199, my_IIR_filter_firBlock_left_multProducts[38], my_IIR_filter_firBlock_left_firStep[104] );
xor U2980 ( my_IIR_filter_firBlock_left_N73, n1624, n1623 );
xor U2981 ( n1623, my_IIR_filter_firBlock_left_multProducts[38], my_IIR_filter_firBlock_left_firStep[200] );
xor U2982 ( my_IIR_filter_firBlock_left_N200, n463, n2335 );
xor U2983 ( n463, my_IIR_filter_firBlock_left_firStep[71], my_IIR_filter_firBlock_left_multProducts[38] );
xor U2984 ( my_IIR_filter_firBlock_left_N40, n464, n1484 );
xor U2985 ( n464, my_IIR_filter_firBlock_left_firStep[231], my_IIR_filter_firBlock_left_multProducts[38] );
xor U2986 ( my_IIR_filter_firBlock_right_N162, n3477, n3476 );
xor U2987 ( n3476, my_IIR_filter_firBlock_right_multProducts[1], my_IIR_filter_firBlock_right_firStep[1] );
xor U2988 ( my_IIR_filter_firBlock_right_N97, my_IIR_filter_firBlock_right_multProducts[31], my_IIR_filter_firBlock_right_firStep[31] );
xor U2989 ( my_IIR_filter_firBlock_left_N228, n465, n2466 );
xor U2990 ( n465, my_IIR_filter_firBlock_left_firStep[35], my_IIR_filter_firBlock_left_multProducts[64] );
xor U2991 ( my_IIR_filter_firBlock_left_N4, n466, n1212 );
xor U2992 ( n466, my_IIR_filter_firBlock_left_firStep[259], my_IIR_filter_firBlock_left_multProducts[64] );
xor U2993 ( my_IIR_filter_firBlock_left_N267, n2502, n2501 );
xor U2994 ( n2501, my_IIR_filter_firBlock_left_multProducts[100], my_IIR_filter_firBlock_left_firStep[10] );
xor U2995 ( my_IIR_filter_firBlock_right_N40, n467, n2804 );
xor U2996 ( n467, my_IIR_filter_firBlock_right_firStep[69], my_IIR_filter_firBlock_right_multProducts[69] );
xor U2997 ( my_IIR_filter_firBlock_left_N227, n2455, n2454 );
xor U2998 ( n2454, my_IIR_filter_firBlock_left_multProducts[63], my_IIR_filter_firBlock_left_firStep[34] );
xor U2999 ( my_IIR_filter_firBlock_left_N3, n1201, n1200 );
xor U3000 ( n1200, my_IIR_filter_firBlock_left_multProducts[63], my_IIR_filter_firBlock_left_firStep[258] );
xor U3001 ( my_IIR_filter_firBlock_left_N199, n2334, n2333 );
xor U3002 ( n2333, my_IIR_filter_firBlock_left_multProducts[37], my_IIR_filter_firBlock_left_firStep[70] );
xor U3003 ( my_IIR_filter_firBlock_left_N39, n1483, n1482 );
xor U3004 ( n1482, my_IIR_filter_firBlock_left_multProducts[37], my_IIR_filter_firBlock_left_firStep[230] );
xor U3005 ( my_IIR_filter_firBlock_left_N168, n468, n2198 );
xor U3006 ( n468, my_IIR_filter_firBlock_left_firStep[103], my_IIR_filter_firBlock_left_multProducts[37] );
xor U3007 ( my_IIR_filter_firBlock_left_N72, n469, n1622 );
xor U3008 ( n469, my_IIR_filter_firBlock_left_firStep[199], my_IIR_filter_firBlock_left_multProducts[37] );
xor U3009 ( my_IIR_filter_firBlock_left_N134, n470, n2057 );
xor U3010 ( n470, my_IIR_filter_firBlock_left_firStep[133], my_IIR_filter_firBlock_left_multProducts[5] );
xor U3011 ( my_IIR_filter_firBlock_left_N102, n471, n1919 );
xor U3012 ( n471, my_IIR_filter_firBlock_left_firStep[165], my_IIR_filter_firBlock_left_multProducts[5] );
xor U3013 ( my_IIR_filter_firBlock_right_N39, n2803, n2802 );
xor U3014 ( n2802, my_IIR_filter_firBlock_right_multProducts[68], my_IIR_filter_firBlock_right_firStep[68] );
xnor U3015 ( my_IIR_filter_firBlock_left_N266, n2624, n2623 );
xnor U3016 ( n2624, my_IIR_filter_firBlock_left_firStep[9], my_IIR_filter_firBlock_left_multProducts[99] );
xor U3017 ( my_IIR_filter_firBlock_left_N133, n2056, n2055 );
xor U3018 ( n2055, my_IIR_filter_firBlock_left_multProducts[4], my_IIR_filter_firBlock_left_firStep[132] );
xor U3019 ( my_IIR_filter_firBlock_left_N101, n1918, n1917 );
xor U3020 ( n1917, my_IIR_filter_firBlock_left_multProducts[4], my_IIR_filter_firBlock_left_firStep[164] );
xor U3021 ( my_IIR_filter_firBlock_left_N167, n2197, n2196 );
xor U3022 ( n2196, my_IIR_filter_firBlock_left_multProducts[36], my_IIR_filter_firBlock_left_firStep[102] );
xor U3023 ( my_IIR_filter_firBlock_left_N71, n1621, n1620 );
xor U3024 ( n1620, my_IIR_filter_firBlock_left_multProducts[36], my_IIR_filter_firBlock_left_firStep[198] );
xor U3025 ( my_IIR_filter_firBlock_left_N2, n1154, n1153 );
xor U3026 ( my_IIR_filter_firBlock_left_N226, n2408, n2407 );
xor U3027 ( my_IIR_filter_firBlock_left_N198, n472, n2332 );
xor U3028 ( n472, my_IIR_filter_firBlock_left_firStep[69], my_IIR_filter_firBlock_left_multProducts[36] );
xor U3029 ( my_IIR_filter_firBlock_left_N38, n473, n1481 );
xor U3030 ( n473, my_IIR_filter_firBlock_left_firStep[229], my_IIR_filter_firBlock_left_multProducts[36] );
xor U3031 ( my_IIR_filter_firBlock_left_N265, n2622, n2621 );
xor U3032 ( n2621, my_IIR_filter_firBlock_left_multProducts[98], my_IIR_filter_firBlock_left_firStep[8] );
xor U3033 ( my_IIR_filter_firBlock_right_N38, n474, n2801 );
xor U3034 ( n474, my_IIR_filter_firBlock_right_firStep[67], my_IIR_filter_firBlock_right_multProducts[67] );
xor U3035 ( my_IIR_filter_firBlock_left_N197, n2331, n2330 );
xor U3036 ( n2330, my_IIR_filter_firBlock_left_multProducts[35], my_IIR_filter_firBlock_left_firStep[68] );
xor U3037 ( my_IIR_filter_firBlock_left_N37, n1480, n1479 );
xor U3038 ( n1479, my_IIR_filter_firBlock_left_multProducts[35], my_IIR_filter_firBlock_left_firStep[228] );
xor U3039 ( my_IIR_filter_firBlock_left_N166, n475, n2195 );
xor U3040 ( n475, my_IIR_filter_firBlock_left_firStep[101], my_IIR_filter_firBlock_left_multProducts[35] );
xor U3041 ( my_IIR_filter_firBlock_left_N70, n476, n1619 );
xor U3042 ( n476, my_IIR_filter_firBlock_left_firStep[197], my_IIR_filter_firBlock_left_multProducts[35] );
xor U3043 ( my_IIR_filter_firBlock_right_N37, n2800, n2799 );
xor U3044 ( n2799, my_IIR_filter_firBlock_right_multProducts[66], my_IIR_filter_firBlock_right_firStep[66] );
xor U3045 ( my_IIR_filter_firBlock_left_N132, n477, n2054 );
xor U3046 ( n477, my_IIR_filter_firBlock_left_firStep[131], my_IIR_filter_firBlock_left_multProducts[3] );
xor U3047 ( my_IIR_filter_firBlock_left_N100, n478, n1916 );
xor U3048 ( n478, my_IIR_filter_firBlock_left_firStep[163], my_IIR_filter_firBlock_left_multProducts[3] );
xnor U3049 ( my_IIR_filter_firBlock_left_N264, n2620, n2619 );
xnor U3050 ( n2620, my_IIR_filter_firBlock_left_firStep[7], my_IIR_filter_firBlock_left_multProducts[97] );
xor U3051 ( my_IIR_filter_firBlock_left_N131, n2042, n2041 );
xor U3052 ( n2041, my_IIR_filter_firBlock_left_multProducts[2], my_IIR_filter_firBlock_left_firStep[130] );
xor U3053 ( my_IIR_filter_firBlock_left_N99, n1906, n1905 );
xor U3054 ( n1905, my_IIR_filter_firBlock_left_multProducts[2], my_IIR_filter_firBlock_left_firStep[162] );
xor U3055 ( my_IIR_filter_firBlock_left_N165, n2194, n2193 );
xor U3056 ( n2193, my_IIR_filter_firBlock_left_multProducts[34], my_IIR_filter_firBlock_left_firStep[100] );
xor U3057 ( my_IIR_filter_firBlock_left_N69, n1618, n1617 );
xor U3058 ( n1617, my_IIR_filter_firBlock_left_multProducts[34], my_IIR_filter_firBlock_left_firStep[196] );
xor U3059 ( my_IIR_filter_firBlock_left_N196, n479, n2329 );
xor U3060 ( n479, my_IIR_filter_firBlock_left_firStep[67], my_IIR_filter_firBlock_left_multProducts[34] );
xor U3061 ( my_IIR_filter_firBlock_left_N36, n480, n1478 );
xor U3062 ( n480, my_IIR_filter_firBlock_left_firStep[227], my_IIR_filter_firBlock_left_multProducts[34] );
xor U3063 ( my_IIR_filter_firBlock_right_N36, n481, n2798 );
xor U3064 ( n481, my_IIR_filter_firBlock_right_firStep[65], my_IIR_filter_firBlock_right_multProducts[65] );
xor U3065 ( my_IIR_filter_firBlock_left_N263, n2618, n2617 );
xor U3066 ( n2617, my_IIR_filter_firBlock_left_multProducts[96], my_IIR_filter_firBlock_left_firStep[6] );
xor U3067 ( my_IIR_filter_firBlock_right_N35, n2786, n2785 );
xor U3068 ( n2785, my_IIR_filter_firBlock_right_multProducts[64], my_IIR_filter_firBlock_right_firStep[64] );
xor U3069 ( my_IIR_filter_firBlock_left_N195, n2318, n2317 );
xor U3070 ( n2317, my_IIR_filter_firBlock_left_multProducts[33], my_IIR_filter_firBlock_left_firStep[66] );
xor U3071 ( my_IIR_filter_firBlock_left_N35, n1467, n1466 );
xor U3072 ( n1466, my_IIR_filter_firBlock_left_multProducts[33], my_IIR_filter_firBlock_left_firStep[226] );
xor U3073 ( my_IIR_filter_firBlock_left_N130, n1995, n1994 );
xor U3074 ( n1994, my_IIR_filter_firBlock_left_multProducts[1], my_IIR_filter_firBlock_left_firStep[129] );
xor U3075 ( my_IIR_filter_firBlock_left_N98, n1859, n1858 );
xor U3076 ( n1858, my_IIR_filter_firBlock_left_multProducts[1], my_IIR_filter_firBlock_left_firStep[161] );
xor U3077 ( my_IIR_filter_firBlock_left_N164, n482, n2192 );
xor U3078 ( n482, my_IIR_filter_firBlock_left_firStep[99], my_IIR_filter_firBlock_left_multProducts[33] );
xor U3079 ( my_IIR_filter_firBlock_left_N68, n483, n1616 );
xor U3080 ( n483, my_IIR_filter_firBlock_left_firStep[195], my_IIR_filter_firBlock_left_multProducts[33] );
xnor U3081 ( my_IIR_filter_firBlock_left_N262, n2616, n2615 );
xnor U3082 ( n2616, my_IIR_filter_firBlock_left_firStep[5], my_IIR_filter_firBlock_left_multProducts[95] );
xor U3083 ( my_IIR_filter_firBlock_right_N34, n2739, n2738 );
xor U3084 ( n2738, my_IIR_filter_firBlock_right_multProducts[63], my_IIR_filter_firBlock_right_firStep[63] );
xor U3085 ( my_IIR_filter_firBlock_left_N194, n2271, n2270 );
xor U3086 ( n2270, my_IIR_filter_firBlock_left_multProducts[32], my_IIR_filter_firBlock_left_firStep[65] );
xor U3087 ( my_IIR_filter_firBlock_left_N163, n2180, n2179 );
xor U3088 ( n2179, my_IIR_filter_firBlock_left_multProducts[32], my_IIR_filter_firBlock_left_firStep[98] );
xor U3089 ( my_IIR_filter_firBlock_left_N67, n1604, n1603 );
xor U3090 ( n1603, my_IIR_filter_firBlock_left_multProducts[32], my_IIR_filter_firBlock_left_firStep[194] );
xor U3091 ( my_IIR_filter_firBlock_left_N34, n1420, n1419 );
xor U3092 ( n1419, my_IIR_filter_firBlock_left_multProducts[32], my_IIR_filter_firBlock_left_firStep[225] );
xor U3093 ( my_IIR_filter_firBlock_left_N261, n2614, n2613 );
xor U3094 ( n2613, my_IIR_filter_firBlock_left_multProducts[94], my_IIR_filter_firBlock_left_firStep[4] );
xor U3095 ( my_IIR_filter_firBlock_left_N129, my_IIR_filter_firBlock_left_multProducts[0], my_IIR_filter_firBlock_left_firStep[128] );
xor U3096 ( my_IIR_filter_firBlock_left_N97, my_IIR_filter_firBlock_left_multProducts[0], my_IIR_filter_firBlock_left_firStep[160] );
xor U3097 ( my_IIR_filter_firBlock_left_N162, n2133, n2132 );
xor U3098 ( n2132, my_IIR_filter_firBlock_left_multProducts[31], my_IIR_filter_firBlock_left_firStep[97] );
xor U3099 ( my_IIR_filter_firBlock_left_N66, n1557, n1556 );
xor U3100 ( n1556, my_IIR_filter_firBlock_left_multProducts[31], my_IIR_filter_firBlock_left_firStep[193] );
xor U3101 ( my_IIR_filter_firBlock_right_N33, my_IIR_filter_firBlock_right_multProducts[62], my_IIR_filter_firBlock_right_firStep[62] );
xor U3102 ( my_IIR_filter_firBlock_left_N260, n484, n2612 );
xor U3103 ( n484, my_IIR_filter_firBlock_left_firStep[3], my_IIR_filter_firBlock_left_multProducts[93] );
xor U3104 ( my_IIR_filter_firBlock_left_N193, my_IIR_filter_firBlock_left_multProducts[31], my_IIR_filter_firBlock_left_firStep[64] );
xor U3105 ( my_IIR_filter_firBlock_left_N33, my_IIR_filter_firBlock_left_multProducts[31], my_IIR_filter_firBlock_left_firStep[224] );
xor U3106 ( my_IIR_filter_firBlock_left_N259, n2600, n2599 );
xor U3107 ( n2599, my_IIR_filter_firBlock_left_multProducts[92], my_IIR_filter_firBlock_left_firStep[2] );
xor U3108 ( my_IIR_filter_firBlock_left_N161, my_IIR_filter_firBlock_left_multProducts[30], my_IIR_filter_firBlock_left_firStep[96] );
xor U3109 ( my_IIR_filter_firBlock_left_N65, my_IIR_filter_firBlock_left_multProducts[30], my_IIR_filter_firBlock_left_firStep[192] );
xor U3110 ( my_IIR_filter_firBlock_left_N258, n2548, n2547 );
xor U3111 ( n2547, my_IIR_filter_firBlock_left_multProducts[91], my_IIR_filter_firBlock_left_firStep[1] );
xor U3112 ( my_IIR_filter_firBlock_left_N257, my_IIR_filter_firBlock_left_multProducts[90], my_IIR_filter_firBlock_left_firStep[0] );
buf U3113 ( n629, reset );
nand U3114 ( n2860, n496, n2857 );
or U3115 ( n2858, n2857, n495 );
nand U3116 ( n2857, n2856, n2855 );
nand U3117 ( n3642, n3640, n3639 );
nand U3118 ( n1016, my_IIR_filter_firBlock_left_multProducts[101], n1015 );
or U3119 ( n1015, n1014, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[26] );
nand U3120 ( n3002, n3000, n2999 );
nand U3121 ( n2999, n2998, n689 );
nand U3122 ( n936, n815, n814 );
nand U3123 ( n3618, n3617, n147 );
xnor U3124 ( my_IIR_filter_firBlock_right_multProducts[22], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[29], n3393 );
xor U3125 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[29], n3166, n3164 );
xor U3126 ( n3701, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[30], n647 );
xor U3127 ( n1055, my_IIR_filter_firBlock_left_multProducts[110], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[35] );
or U3128 ( n3596, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[5], n3595 );
not U3129 ( n669, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[35] );
nand U3130 ( n3048, n3047, n3046 );
xor U3131 ( n1064, my_IIR_filter_firBlock_left_multProducts[112], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[37] );
xor U3132 ( n1779, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[37], n526 );
nand U3133 ( n1783, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[37], n1780 );
or U3134 ( n1781, n1780, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[37] );
xor U3135 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[37], n927, n926 );
nand U3136 ( n727, leftOut[9], n810 );
xor U3137 ( n1028, my_IIR_filter_firBlock_left_multProducts[104], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[29] );
xor U3138 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[11], n3082, n3081 );
xor U3139 ( n1045, my_IIR_filter_firBlock_left_multProducts[108], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[33] );
xor U3140 ( n1759, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[33], n526 );
nand U3141 ( n1763, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[33], n1760 );
or U3142 ( n1761, n1760, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[33] );
nand U3143 ( n3208, n3207, n3206 );
xor U3144 ( n1121, my_IIR_filter_firBlock_left_multProducts[73], my_IIR_filter_firBlock_left_firStep[268] );
nand U3145 ( n1124, my_IIR_filter_firBlock_left_multProducts[73], n1123 );
xor U3146 ( n2375, my_IIR_filter_firBlock_left_multProducts[73], my_IIR_filter_firBlock_left_firStep[44] );
xor U3147 ( n1004, my_IIR_filter_firBlock_left_multProducts[99], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[24] );
xor U3148 ( n1714, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[24], n54 );
nand U3149 ( n1718, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[24], n1715 );
or U3150 ( n1716, n1715, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[24] );
buf U3151 ( n510, outData_in[12] );
buf U3152 ( n511, outData_in[12] );
nand U3153 ( n2819, n517, n2931 );
or U3154 ( n2817, n2931, n517 );
xor U3155 ( n3055, n706, n517 );
xor U3156 ( my_IIR_filter_firBlock_right_N123, n3323, n3322 );
nand U3157 ( n3326, my_IIR_filter_firBlock_right_firStep[57], n3323 );
xor U3158 ( n995, my_IIR_filter_firBlock_left_multProducts[97], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[22] );
xor U3159 ( n1704, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[22], n53 );
nand U3160 ( n1708, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[22], n1705 );
or U3161 ( n1706, n1705, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[22] );
xor U3162 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[22], n855, n854 );
xor U3163 ( n1037, my_IIR_filter_firBlock_left_multProducts[106], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[31] );
xor U3164 ( n1749, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[31], n526 );
nand U3165 ( n1753, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[31], n1750 );
or U3166 ( n1751, n1750, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[31] );
nand U3167 ( n905, n903, n902 );
xor U3168 ( n1040, my_IIR_filter_firBlock_left_multProducts[107], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[32] );
nand U3169 ( n1107, my_IIR_filter_firBlock_left_multProducts[69], n1106 );
xor U3170 ( n1219, my_IIR_filter_firBlock_left_multProducts[69], my_IIR_filter_firBlock_left_firStep[264] );
nand U3171 ( n2361, my_IIR_filter_firBlock_left_multProducts[69], n2360 );
xor U3172 ( n2473, my_IIR_filter_firBlock_left_multProducts[69], my_IIR_filter_firBlock_left_firStep[40] );
nand U3173 ( n1095, my_IIR_filter_firBlock_left_multProducts[65], n1094 );
xor U3174 ( n1213, my_IIR_filter_firBlock_left_multProducts[65], my_IIR_filter_firBlock_left_firStep[260] );
nand U3175 ( n2349, my_IIR_filter_firBlock_left_multProducts[65], n2348 );
xor U3176 ( n2467, my_IIR_filter_firBlock_left_multProducts[65], my_IIR_filter_firBlock_left_firStep[36] );
xor U3177 ( my_IIR_filter_firBlock_left_multProducts[65], n974, n973 );
xor U3178 ( n3687, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[27], n645 );
xor U3179 ( n1050, my_IIR_filter_firBlock_left_multProducts[109], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[34] );
nand U3180 ( n1054, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[34], n1051 );
or U3181 ( n1052, n1051, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[34] );
xor U3182 ( n1764, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[34], n526 );
nand U3183 ( n1768, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[34], n1765 );
or U3184 ( n1766, n1765, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[34] );
xor U3185 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[34], n910, n909 );
xor U3186 ( n3615, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[11], n147 );
xnor U3187 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[9], n3220, n3219 );
buf U3188 ( n485, outData_in[14] );
buf U3189 ( n486, outData_in[14] );
xor U3190 ( outData_in[14], n744, n743 );
xor U3191 ( n3682, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[26], n644 );
not U3192 ( n651, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[35] );
xor U3193 ( my_IIR_filter_firBlock_right_multProducts[28], n3402, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[35] );
nor U3194 ( n3401, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[35], n3402 );
or U3195 ( n3403, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[36], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[35] );
xor U3196 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[35], n3194, n3193 );
xor U3197 ( n1784, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[38], n526 );
or U3198 ( n1786, n1785, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[38] );
xor U3199 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[38], n932, n931 );
nand U3200 ( n1160, n1158, n1157 );
nand U3201 ( n1157, my_IIR_filter_firBlock_left_multProducts[80], n1156 );
nand U3202 ( n3442, my_IIR_filter_firBlock_right_multProducts[11], n3441 );
buf U3203 ( n487, n528 );
buf U3204 ( n488, n528 );
buf U3205 ( n528, outData_in[11] );
buf U3206 ( n489, outData_in[22] );
buf U3207 ( n490, outData_in[22] );
xor U3208 ( outData_in[22], n771, n770 );
xor U3209 ( n1177, my_IIR_filter_firBlock_left_multProducts[85], my_IIR_filter_firBlock_left_firStep[280] );
nand U3210 ( n1180, my_IIR_filter_firBlock_left_multProducts[85], n1179 );
xor U3211 ( n2431, my_IIR_filter_firBlock_left_multProducts[85], my_IIR_filter_firBlock_left_firStep[56] );
xor U3212 ( my_IIR_filter_firBlock_right_multProducts[24], n3396, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[31] );
nor U3213 ( n3395, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[31], n3396 );
xor U3214 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[31], n3174, n3173 );
nand U3215 ( n3469, my_IIR_filter_firBlock_right_multProducts[17], n3468 );
buf U3216 ( n493, outData_in[19] );
xnor U3217 ( my_IIR_filter_firBlock_right_multProducts[5], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[12], n3365 );
xnor U3218 ( my_IIR_filter_firBlock_right_multProducts[26], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[33], n3399 );
nor U3219 ( n3400, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[34], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[33] );
nand U3220 ( n3228, my_IIR_filter_firBlock_right_multProducts[34], n3227 );
nor U3221 ( n3358, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[4], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[3] );
or U3222 ( n3588, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[3], n3587 );
xor U3223 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[3], n3213, n167 );
nand U3224 ( n1036, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[30], n1033 );
or U3225 ( n1034, n1033, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[30] );
xor U3226 ( n1744, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[30], n61 );
nand U3227 ( n1748, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[30], n1745 );
or U3228 ( n1746, n1745, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[30] );
xor U3229 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[30], n891, n890 );
buf U3230 ( n495, outData_in[15] );
nand U3231 ( n1142, my_IIR_filter_firBlock_left_multProducts[77], n1141 );
or U3232 ( n1141, n1140, my_IIR_filter_firBlock_left_firStep[272] );
nand U3233 ( n3507, my_IIR_filter_firBlock_right_multProducts[25], n3506 );
xor U3234 ( my_IIR_filter_firBlock_left_N1, my_IIR_filter_firBlock_left_multProducts[61], my_IIR_filter_firBlock_left_firStep[256] );
xor U3235 ( my_IIR_filter_firBlock_left_N225, my_IIR_filter_firBlock_left_multProducts[61], my_IIR_filter_firBlock_left_firStep[32] );
and U3236 ( n2408, my_IIR_filter_firBlock_left_multProducts[61], my_IIR_filter_firBlock_left_firStep[32] );
nand U3237 ( n834, n832, n831 );
or U3238 ( n3356, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[2], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[1] );
nand U3239 ( n865, n863, n862 );
xor U3240 ( n1013, my_IIR_filter_firBlock_left_multProducts[101], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[26] );
xor U3241 ( n1023, my_IIR_filter_firBlock_left_multProducts[103], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[28] );
nand U3242 ( n1027, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[28], n1024 );
or U3243 ( n1025, n1024, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[28] );
xor U3244 ( n1734, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[28], n59 );
nand U3245 ( n1738, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[28], n1735 );
or U3246 ( n1736, n1735, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[28] );
xor U3247 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[28], n881, n880 );
xor U3248 ( n1018, my_IIR_filter_firBlock_left_multProducts[102], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[27] );
xor U3249 ( n1729, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[27], n57 );
nand U3250 ( n1733, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[27], n1730 );
or U3251 ( n1731, n1730, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[27] );
buf U3252 ( n497, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[1] );
xor U3253 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[1], rightOut[0], leftOut[0] );
nand U3254 ( n806, n720, n719 );
nand U3255 ( n1003, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[23], n1000 );
or U3256 ( n1001, n1000, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[23] );
xor U3257 ( n1709, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[23], n308 );
nand U3258 ( n1713, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[23], n1710 );
or U3259 ( n1711, n1710, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[23] );
xor U3260 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[23], n860, n859 );
nand U3261 ( n1110, my_IIR_filter_firBlock_left_multProducts[70], n1109 );
nand U3262 ( n876, n874, n873 );
xnor U3263 ( outData_in[13], n739, n740 );
xor U3264 ( n1694, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[20], n51 );
nand U3265 ( n1698, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[20], n1695 );
or U3266 ( n1696, n1695, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[20] );
buf U3267 ( n500, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[2] );
xor U3268 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[2], n760, n759 );
nand U3269 ( n1092, my_IIR_filter_firBlock_left_multProducts[64], n1091 );
nand U3270 ( n2346, my_IIR_filter_firBlock_left_multProducts[64], n2345 );
buf U3271 ( n502, outData_in[3] );
nand U3272 ( n847, n845, n844 );
nand U3273 ( n3075, n167, n3220 );
or U3274 ( n3073, n3220, n167 );
or U3275 ( n3065, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[10], n167 );
nor U3276 ( n3214, n167, n3213 );
buf U3277 ( n504, outData_in[25] );
nand U3278 ( n1128, my_IIR_filter_firBlock_left_multProducts[74], n1127 );
nand U3279 ( n2382, my_IIR_filter_firBlock_left_multProducts[74], n2381 );
xor U3280 ( my_IIR_filter_firBlock_left_multProducts[74], n1014, n1013 );
xor U3281 ( my_IIR_filter_firBlock_left_N29, n1196, n1195 );
nand U3282 ( n1199, my_IIR_filter_firBlock_left_firStep[284], n1196 );
or U3283 ( n1197, n1196, my_IIR_filter_firBlock_left_firStep[284] );
nand U3284 ( n1196, n1194, n1193 );
buf U3285 ( n506, outData_in[8] );
buf U3286 ( n507, outData_in[8] );
xor U3287 ( outData_in[8], n809, n808 );
buf U3288 ( n508, outData_in[10] );
xor U3289 ( outData_in[10], n729, n728 );
xnor U3290 ( my_IIR_filter_firBlock_right_multProducts[101], outData_in[16], n3558 );
or U3291 ( n3560, outData_in[16], n496 );
nor U3292 ( n2644, outData_in[16], n496 );
xor U3293 ( my_IIR_filter_firBlock_right_multProducts[75], n2642, outData_in[16] );
nand U3294 ( n2864, outData_in[16], n2861 );
or U3295 ( n2862, n2861, outData_in[16] );
nand U3296 ( n2855, outData_in[16], n2854 );
not U3297 ( n685, outData_in[16] );
buf U3298 ( n513, outData_in[17] );
xor U3299 ( n982, my_IIR_filter_firBlock_left_multProducts[94], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[19] );
nand U3300 ( n986, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[19], n983 );
or U3301 ( n984, n983, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[19] );
xor U3302 ( n1689, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[19], n304 );
nand U3303 ( n1693, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[19], n1690 );
or U3304 ( n1691, n1690, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[19] );
buf U3305 ( n514, outData_in[29] );
xor U3306 ( n973, my_IIR_filter_firBlock_left_multProducts[92], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[17] );
nand U3307 ( n977, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[17], n974 );
or U3308 ( n975, n974, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[17] );
xor U3309 ( n1679, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[17], n300 );
nand U3310 ( n1683, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[17], n1680 );
or U3311 ( n1681, n1680, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[17] );
xor U3312 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[17], n834, n833 );
buf U3313 ( n516, outData_in[4] );
buf U3314 ( n517, outData_in[4] );
xor U3315 ( outData_in[4], n803, n802 );
xnor U3316 ( outData_in[9], n811, n810 );
buf U3317 ( n520, outData_in[6] );
buf U3318 ( n521, outData_in[6] );
xor U3319 ( outData_in[6], n806, n805 );
xnor U3320 ( outData_in[11], n732, n733 );
not U3321 ( n529, n692 );
not U3322 ( n692, outData_in[23] );
nand U3323 ( n3398, n3399, n128 );
or U3324 ( n3102, n3099, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[21] );
nand U3325 ( n3100, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[21], n3099 );
nand U3326 ( n3080, n3077, n657 );
or U3327 ( n3078, n657, n3077 );
xnor U3328 ( my_IIR_filter_firBlock_right_multProducts[105], outData_in[20], n3564 );
xor U3329 ( n3257, my_IIR_filter_firBlock_right_multProducts[43], my_IIR_filter_firBlock_right_firStep[43] );
xor U3330 ( my_IIR_filter_firBlock_right_multProducts[79], n2648, outData_in[20] );
nand U3331 ( n2881, outData_in[20], n2878 );
or U3332 ( n2879, n2878, outData_in[20] );
or U3333 ( n3379, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[20], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[19] );
xnor U3334 ( my_IIR_filter_firBlock_right_multProducts[13], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[20], n3377 );
not U3335 ( n638, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[20] );
nand U3336 ( n2872, outData_in[20], n2871 );
not U3337 ( n689, outData_in[20] );
not U3338 ( n641, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[23] );
nand U3339 ( n3204, n3202, n3201 );
xnor U3340 ( my_IIR_filter_firBlock_right_multProducts[113], n209, n3576 );
xor U3341 ( my_IIR_filter_firBlock_right_multProducts[87], n2660, n209 );
nand U3342 ( n2916, n209, n2913 );
or U3343 ( n2914, n2913, n209 );
nand U3344 ( n2906, n209, n2905 );
not U3345 ( n697, outData_in[28] );
xor U3346 ( n3033, n695, outData_in[28] );
xnor U3347 ( n3127, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[27], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[21] );
xor U3348 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[21], n3128, n3127 );
nand U3349 ( n3662, n3661, n639 );
nand U3350 ( n3697, n3696, n3695 );
nand U3351 ( n3231, my_IIR_filter_firBlock_right_multProducts[35], n3230 );
nand U3352 ( n3246, my_IIR_filter_firBlock_right_multProducts[40], n3245 );
nand U3353 ( n3260, my_IIR_filter_firBlock_right_multProducts[43], n3259 );
nand U3354 ( n3008, n3007, n691 );
nand U3355 ( n3046, n3045, n699 );
nand U3356 ( n2989, n2988, n2987 );
not U3357 ( n699, outData_in[30] );
xnor U3358 ( my_IIR_filter_firBlock_right_multProducts[89], outData_in[30], n2663 );
nand U3359 ( n2915, outData_in[30], n2914 );
nand U3360 ( n2925, outData_in[30], n2922 );
or U3361 ( n2923, n2922, outData_in[30] );
xor U3362 ( my_IIR_filter_firBlock_right_multProducts[115], n3579, outData_in[30] );
or U3363 ( n2665, outData_in[30], n514 );
nor U3364 ( n3581, outData_in[30], n514 );
nand U3365 ( n3695, n3694, n646 );
nand U3366 ( n3678, n3676, n3675 );
nand U3367 ( n3273, n3272, my_IIR_filter_firBlock_right_multProducts[46] );
xnor U3368 ( my_IIR_filter_firBlock_right_multProducts[14], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[21], n3381 );
not U3369 ( n639, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[21] );
nand U3370 ( n942, n823, n822 );
xor U3371 ( my_IIR_filter_firBlock_left_N256, n2465, n2464 );
nor U3372 ( n2464, n2463, n2462 );
nand U3373 ( n940, n821, n820 );
nand U3374 ( n820, n819, n45 );
nand U3375 ( n2403, n2401, n2400 );
nand U3376 ( n2400, my_IIR_filter_firBlock_left_multProducts[78], n2399 );
nand U3377 ( n2441, n2439, n2438 );
nand U3378 ( n2438, my_IIR_filter_firBlock_left_multProducts[86], n2437 );
nand U3379 ( n2367, n2365, n2364 );
nand U3380 ( n2364, my_IIR_filter_firBlock_left_multProducts[70], n2363 );
nand U3381 ( n2474, n2359, n2358 );
nand U3382 ( n2358, my_IIR_filter_firBlock_left_multProducts[68], n2357 );
nand U3383 ( n2425, my_IIR_filter_firBlock_left_multProducts[83], n2424 );
nand U3384 ( n2434, my_IIR_filter_firBlock_left_multProducts[85], n2433 );
or U3385 ( n2433, n2432, my_IIR_filter_firBlock_left_firStep[56] );
nand U3386 ( n2416, my_IIR_filter_firBlock_left_multProducts[81], n2415 );
or U3387 ( n2415, n2414, my_IIR_filter_firBlock_left_firStep[52] );
nand U3388 ( n2396, my_IIR_filter_firBlock_left_multProducts[77], n2395 );
or U3389 ( n2395, n2394, my_IIR_filter_firBlock_left_firStep[48] );
nand U3390 ( n2378, my_IIR_filter_firBlock_left_multProducts[73], n2377 );
nand U3391 ( n2411, my_IIR_filter_firBlock_left_multProducts[80], n2410 );
nand U3392 ( n2373, my_IIR_filter_firBlock_left_multProducts[72], n2372 );
or U3393 ( n2357, n2472, my_IIR_filter_firBlock_left_firStep[39] );
nor U3394 ( n2460, my_IIR_filter_firBlock_left_firStep[62], n2461 );
xor U3395 ( my_IIR_filter_firBlock_left_multProducts[63], n1084, n1083 );
xor U3396 ( n1083, my_IIR_filter_firBlock_left_multProducts[90], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[15] );
xor U3397 ( my_IIR_filter_firBlock_right_multProducts[112], n3577, n492 );
nor U3398 ( n3576, n491, n3577 );
or U3399 ( n3578, n209, n492 );
nor U3400 ( n2662, n209, n491 );
nand U3401 ( n2912, n492, n2909 );
xnor U3402 ( n2908, n491, n515 );
or U3403 ( n2910, n2909, n492 );
nand U3404 ( n2902, n491, n2901 );
not U3405 ( n696, n491 );
nand U3406 ( n3526, my_IIR_filter_firBlock_right_multProducts[29], n3525 );
nand U3407 ( n3494, my_IIR_filter_firBlock_right_multProducts[22], n3493 );
nand U3408 ( n3524, n3521, n3520 );
nand U3409 ( n3478, n3475, n3474 );
nand U3410 ( n3472, n3470, n3469 );
nand U3411 ( n3467, n3466, n3465 );
xnor U3412 ( my_IIR_filter_firBlock_right_multProducts[109], n157, n3570 );
xor U3413 ( n3275, my_IIR_filter_firBlock_right_multProducts[47], my_IIR_filter_firBlock_right_firStep[47] );
or U3414 ( n3572, n157, n529 );
nor U3415 ( n2656, n157, n529 );
xor U3416 ( my_IIR_filter_firBlock_right_multProducts[83], n2654, n157 );
nand U3417 ( n2898, n157, n2895 );
or U3418 ( n2896, n2895, n157 );
or U3419 ( n3385, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[24], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[23] );
xnor U3420 ( my_IIR_filter_firBlock_right_multProducts[17], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[24], n3383 );
not U3421 ( n642, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[24] );
nand U3422 ( n2888, n157, n2887 );
not U3423 ( n693, outData_in[24] );
xor U3424 ( n3015, n691, outData_in[24] );
nand U3425 ( n3264, my_IIR_filter_firBlock_right_multProducts[44], n3263 );
nand U3426 ( n3114, n3112, n3111 );
nand U3427 ( n3111, n3110, n661 );
xor U3428 ( n3715, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[33], n128 );
xnor U3429 ( my_IIR_filter_firBlock_right_multProducts[110], n505, n3574 );
nor U3430 ( n2657, n504, n2658 );
xor U3431 ( my_IIR_filter_firBlock_right_multProducts[84], n2658, n505 );
nor U3432 ( n3388, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[26], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[25] );
xnor U3433 ( n2899, n505, n491 );
nand U3434 ( n2903, n504, n2900 );
or U3435 ( n2901, n2900, n504 );
xnor U3436 ( my_IIR_filter_firBlock_right_multProducts[18], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[25], n3387 );
xnor U3437 ( n2890, n529, n504 );
nand U3438 ( n2893, n505, n2892 );
nand U3439 ( n3699, n3698, n140 );
nand U3440 ( n3666, n3665, n640 );
xor U3441 ( n3637, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[16], n635 );
xnor U3442 ( my_IIR_filter_firBlock_right_multProducts[9], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[16], n3371 );
not U3443 ( n635, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[16] );
nand U3444 ( n3520, my_IIR_filter_firBlock_right_multProducts[28], n3519 );
nand U3445 ( n3465, my_IIR_filter_firBlock_right_multProducts[16], n3464 );
xor U3446 ( my_IIR_filter_firBlock_right_multProducts[16], n3384, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[23] );
nand U3447 ( n3685, n3684, n644 );
nand U3448 ( n3207, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[37], n3204 );
xor U3449 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[37], n3204, n3203 );
or U3450 ( n3205, n3204, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[37] );
nand U3451 ( n3123, n3121, n3120 );
not U3452 ( n658, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[18] );
xor U3453 ( n3692, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[28], n646 );
xnor U3454 ( n3160, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[28], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[34] );
xor U3455 ( my_IIR_filter_firBlock_right_multProducts[111], n3573, n158 );
nor U3456 ( n3575, n158, n504 );
xnor U3457 ( n3178, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[32], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[38] );
or U3458 ( n2659, n158, n505 );
xnor U3459 ( my_IIR_filter_firBlock_right_multProducts[85], n158, n2657 );
nand U3460 ( n2907, n158, n2904 );
or U3461 ( n2905, n2904, n158 );
nand U3462 ( n2897, n158, n2896 );
not U3463 ( n667, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[32] );
xnor U3464 ( n3150, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[26], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[32] );
not U3465 ( n695, outData_in[26] );
xor U3466 ( n3024, n693, outData_in[26] );
nand U3467 ( n2987, n2986, n686 );
not U3468 ( n686, n512 );
nand U3469 ( n2985, n2983, n2982 );
nand U3470 ( n3022, n3021, n694 );
not U3471 ( n694, n505 );
nand U3472 ( n3044, n3042, n3041 );
nand U3473 ( n3041, n3040, n698 );
xor U3474 ( n3711, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[32], n649 );
nand U3475 ( n3027, n3026, n695 );
nand U3476 ( n3053, n3051, n3050 );
xor U3477 ( n3010, n690, outData_in[23] );
nor U3478 ( n531, n790, leftOut[28] );
nand U3479 ( n532, n3315, n534 );
and U3480 ( n3321, n532, n533 );
or U3481 ( n533, n537, n3317 );
and U3482 ( n534, my_IIR_filter_firBlock_right_multProducts[55], my_IIR_filter_firBlock_right_firStep[56] );
nand U3483 ( n3709, n3708, n648 );
nand U3484 ( n3712, n3710, n3709 );
nand U3485 ( n3741, n3740, n654 );
nand U3486 ( n3211, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[38], n3208 );
or U3487 ( n3209, n3208, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[38] );
nand U3488 ( n3133, n3131, n3130 );
nand U3489 ( n3130, n664, n3129 );
nand U3490 ( n3120, n3119, n662 );
xor U3491 ( my_IIR_filter_firBlock_right_multProducts[99], n3555, n486 );
xnor U3492 ( n3122, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[26], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[20] );
xnor U3493 ( my_IIR_filter_firBlock_right_multProducts[73], n486, n2639 );
nand U3494 ( n2856, n485, n2853 );
or U3495 ( n2854, n2853, n486 );
not U3496 ( n659, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[20] );
nand U3497 ( n2847, n486, n2846 );
not U3498 ( n683, n485 );
nand U3499 ( n535, n3315, my_IIR_filter_firBlock_right_multProducts[55] );
nand U3500 ( n3319, n535, n536 );
and U3501 ( n536, n537, n3317 );
nand U3502 ( n3436, n3434, n3433 );
nand U3503 ( n3447, my_IIR_filter_firBlock_right_multProducts[12], n3446 );
nand U3504 ( n3516, my_IIR_filter_firBlock_right_multProducts[27], n3515 );
nand U3505 ( n3480, my_IIR_filter_firBlock_right_multProducts[19], n3479 );
nand U3506 ( n3498, my_IIR_filter_firBlock_right_multProducts[23], n3497 );
nand U3507 ( n3460, my_IIR_filter_firBlock_right_multProducts[15], n3459 );
nand U3508 ( n3424, my_IIR_filter_firBlock_right_multProducts[6], n3423 );
nand U3509 ( n3485, my_IIR_filter_firBlock_right_multProducts[20], n3484 );
nand U3510 ( n3430, my_IIR_filter_firBlock_right_multProducts[8], n3429 );
nand U3511 ( n3318, n3317, n3316 );
xor U3512 ( outData_in[2], n792, n791 );
xor U3513 ( my_IIR_filter_firBlock_left_N27, n1187, n1186 );
nor U3514 ( n1209, n1206, n631 );
nand U3515 ( n1778, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[36], n1775 );
or U3516 ( n1776, n1775, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[36] );
xor U3517 ( n1774, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[36], n527 );
nand U3518 ( n1190, my_IIR_filter_firBlock_left_firStep[282], n1187 );
or U3519 ( n1188, n1187, my_IIR_filter_firBlock_left_firStep[282] );
nand U3520 ( n1187, n1185, n1184 );
nand U3521 ( n2429, my_IIR_filter_firBlock_left_multProducts[84], n2428 );
nand U3522 ( n1175, my_IIR_filter_firBlock_left_multProducts[84], n1174 );
nand U3523 ( n1063, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[36], n1060 );
or U3524 ( n1061, n1060, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[36] );
nand U3525 ( n913, my_IIR_filter_firBlock_left_multProducts[110], n910 );
or U3526 ( n911, n910, my_IIR_filter_firBlock_left_multProducts[110] );
nand U3527 ( n908, my_IIR_filter_firBlock_left_multProducts[109], n905 );
xor U3528 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[33], n905, n904 );
or U3529 ( n906, n905, my_IIR_filter_firBlock_left_multProducts[109] );
nand U3530 ( n900, n899, n898 );
xor U3531 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[31], n896, n895 );
nand U3532 ( n899, my_IIR_filter_firBlock_left_multProducts[107], n896 );
or U3533 ( n897, n896, my_IIR_filter_firBlock_left_multProducts[107] );
nand U3534 ( n884, my_IIR_filter_firBlock_left_multProducts[104], n881 );
or U3535 ( n882, n881, my_IIR_filter_firBlock_left_multProducts[104] );
nand U3536 ( n879, my_IIR_filter_firBlock_left_multProducts[103], n876 );
xor U3537 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[27], n876, n875 );
or U3538 ( n877, n876, my_IIR_filter_firBlock_left_multProducts[103] );
xor U3539 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[24], n865, n864 );
or U3540 ( n866, n865, my_IIR_filter_firBlock_left_multProducts[100] );
nand U3541 ( n863, my_IIR_filter_firBlock_left_multProducts[99], n860 );
or U3542 ( n861, n860, my_IIR_filter_firBlock_left_multProducts[99] );
xor U3543 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[20], n847, n846 );
or U3544 ( n848, n847, my_IIR_filter_firBlock_left_multProducts[96] );
nand U3545 ( n845, my_IIR_filter_firBlock_left_multProducts[95], n842 );
or U3546 ( n843, n842, my_IIR_filter_firBlock_left_multProducts[95] );
nand U3547 ( n838, n836, n835 );
nand U3548 ( n836, n834, n49 );
xor U3549 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[14], n944, n943 );
or U3550 ( n827, n944, my_IIR_filter_firBlock_left_multProducts[90] );
xor U3551 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[9], n934, n933 );
xor U3552 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[10], n936, n935 );
nand U3553 ( n818, inData_in[2], n936 );
or U3554 ( n816, n936, inData_in[2] );
or U3555 ( n815, n40, n934 );
nand U3556 ( n813, n934, n40 );
nand U3557 ( n709, rightOut[1], n708 );
or U3558 ( n708, leftOut[1], n760 );
nand U3559 ( n792, n709, n710 );
nand U3560 ( n780, leftOut[24], n778 );
xor U3561 ( my_IIR_filter_firBlock_right_N101, n3348, n3347 );
nand U3562 ( n3296, n3294, n3293 );
nand U3563 ( n3262, n3260, n3261 );
nand U3564 ( n3258, n3256, n3255 );
nand U3565 ( n3249, n3247, n3246 );
nand U3566 ( n3355, n3244, n3243 );
nand U3567 ( n3232, my_IIR_filter_firBlock_right_firStep[35], n3348 );
or U3568 ( n3230, n3348, my_IIR_filter_firBlock_right_firStep[35] );
nand U3569 ( n3229, my_IIR_filter_firBlock_right_firStep[34], n3346 );
or U3570 ( n3227, n3346, my_IIR_filter_firBlock_right_firStep[34] );
nand U3571 ( n778, n777, n776 );
xor U3572 ( n1186, my_IIR_filter_firBlock_left_multProducts[87], my_IIR_filter_firBlock_left_firStep[282] );
xor U3573 ( n2440, my_IIR_filter_firBlock_left_multProducts[87], my_IIR_filter_firBlock_left_firStep[58] );
nor U3574 ( n2463, n2460, n631 );
nand U3575 ( n1189, my_IIR_filter_firBlock_left_multProducts[87], n1188 );
nand U3576 ( n2443, my_IIR_filter_firBlock_left_multProducts[87], n2442 );
nand U3577 ( n1070, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[38], n1067 );
or U3578 ( n1068, n1067, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[38] );
xor U3579 ( my_IIR_filter_firBlock_left_multProducts[85], n1065, n1064 );
or U3580 ( n1066, n1065, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[37] );
xor U3581 ( my_IIR_filter_firBlock_left_multProducts[83], n1056, n1055 );
nand U3582 ( n1059, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[35], n1056 );
or U3583 ( n1057, n1056, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[35] );
xor U3584 ( my_IIR_filter_firBlock_left_multProducts[81], n1046, n1045 );
nand U3585 ( n1049, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[33], n1046 );
or U3586 ( n1047, n1046, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[33] );
xor U3587 ( my_IIR_filter_firBlock_left_multProducts[80], n1041, n1040 );
nand U3588 ( n1044, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[32], n1041 );
or U3589 ( n1042, n1041, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[32] );
xor U3590 ( my_IIR_filter_firBlock_left_multProducts[79], n1038, n1037 );
or U3591 ( n1039, n1038, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[31] );
xor U3592 ( my_IIR_filter_firBlock_left_multProducts[77], n1029, n1028 );
nand U3593 ( n1032, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[29], n1029 );
or U3594 ( n1030, n1029, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[29] );
xor U3595 ( my_IIR_filter_firBlock_left_multProducts[75], n1019, n1018 );
nand U3596 ( n1022, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[27], n1019 );
or U3597 ( n1020, n1019, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[27] );
nand U3598 ( n1012, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[25], n1009 );
or U3599 ( n1010, n1009, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[25] );
xor U3600 ( my_IIR_filter_firBlock_left_multProducts[72], n1005, n1004 );
nand U3601 ( n1008, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[24], n1005 );
or U3602 ( n1006, n1005, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[24] );
xor U3603 ( my_IIR_filter_firBlock_left_multProducts[70], n996, n995 );
nand U3604 ( n999, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[22], n996 );
or U3605 ( n997, n996, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[22] );
nand U3606 ( n994, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[21], n991 );
or U3607 ( n992, n991, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[21] );
nand U3608 ( n990, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[20], n987 );
or U3609 ( n988, n987, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[20] );
xor U3610 ( my_IIR_filter_firBlock_left_multProducts[64], n969, n968 );
nand U3611 ( n972, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[16], n969 );
or U3612 ( n970, n969, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[16] );
nand U3613 ( n969, n967, n966 );
nand U3614 ( n1648, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[10], n1645 );
or U3615 ( n1646, n1645, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[10] );
xor U3616 ( my_IIR_filter_firBlock_left_multProducts[61], n1080, n1079 );
xor U3617 ( n1644, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[10], n48 );
nand U3618 ( n961, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[13], n1080 );
or U3619 ( n959, n1080, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[13] );
nand U3620 ( n955, n954, n953 );
nand U3621 ( n3030, n3028, n3027 );
nand U3622 ( n3063, n2951, n2950 );
nand U3623 ( n2950, n2949, n701 );
not U3624 ( n704, n516 );
nand U3625 ( n3004, n3003, n690 );
nand U3626 ( n803, n715, n714 );
or U3627 ( n716, n539, n540 );
nand U3628 ( n3739, n3738, n3737 );
nand U3629 ( n3730, n3728, n3727 );
nand U3630 ( n3716, n3714, n3713 );
nand U3631 ( n3683, n3681, n3680 );
nand U3632 ( n3674, n3672, n3671 );
nand U3633 ( n3656, n3654, n3653 );
nand U3634 ( n3638, n3636, n3635 );
nand U3635 ( n3626, n3625, n115 );
nand U3636 ( n3616, n3614, n3613 );
xnor U3637 ( my_IIR_filter_firBlock_right_multProducts[31], n3745, n3744 );
nand U3638 ( n3607, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[8], n3745 );
nand U3639 ( n3597, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[5], n3594 );
nor U3640 ( n3595, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[5], n3594 );
nand U3641 ( n3593, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[4], n3590 );
nor U3642 ( n3591, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[4], n3590 );
nor U3643 ( n3585, n501, n656 );
nand U3644 ( n2810, n501, n2926 );
nor U3645 ( n3165, n498, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[7] );
or U3646 ( n2808, n501, n2926 );
not U3647 ( n678, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[7] );
not U3648 ( n707, n500 );
xor U3649 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[7], n500, n497 );
nand U3650 ( n3327, n3325, n3326 );
nand U3651 ( n3325, my_IIR_filter_firBlock_right_multProducts[57], n3324 );
nand U3652 ( n3334, my_IIR_filter_firBlock_right_firStep[59], n3331 );
xor U3653 ( my_IIR_filter_firBlock_right_N163, n3523, n3522 );
xor U3654 ( my_IIR_filter_firBlock_right_N161, my_IIR_filter_firBlock_right_multProducts[0], my_IIR_filter_firBlock_right_firStep[0] );
nor U3655 ( n3532, n3531, n3530 );
nand U3656 ( n3501, n3499, n3498 );
nand U3657 ( n3487, n3486, n3485 );
nand U3658 ( n3483, n3481, n3480 );
nand U3659 ( n3463, n3461, n3460 );
nand U3660 ( n3542, n3431, n3430 );
nand U3661 ( n3539, n3425, n3424 );
nand U3662 ( n3413, my_IIR_filter_firBlock_right_firStep[2], n3523 );
or U3663 ( n3411, n3523, my_IIR_filter_firBlock_right_firStep[2] );
nand U3664 ( n3331, n3330, n3329 );
xor U3665 ( n3668, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[23], n641 );
xnor U3666 ( n3136, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[23], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[29] );
xor U3667 ( my_IIR_filter_firBlock_right_multProducts[104], n3565, n494 );
nor U3668 ( n3564, n493, n3565 );
or U3669 ( n3566, outData_in[20], n494 );
xor U3670 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[36], n3044, n3043 );
nand U3671 ( n3047, n209, n3044 );
or U3672 ( n3045, n3044, n209 );
nand U3673 ( n3034, n3032, n3031 );
nor U3674 ( n2650, outData_in[20], n493 );
nand U3675 ( n2648, n2649, n688 );
xor U3676 ( my_IIR_filter_firBlock_right_multProducts[78], n688, n2649 );
nand U3677 ( n2877, n493, n2874 );
or U3678 ( n2875, n2874, n494 );
xnor U3679 ( n2865, n513, n493 );
nand U3680 ( n2868, n493, n2867 );
nand U3681 ( n2995, n2994, n688 );
not U3682 ( n688, n494 );
nand U3683 ( n738, leftOut[12], n736 );
nand U3684 ( n3141, n3139, n3138 );
nand U3685 ( n3179, n3177, n3176 );
nand U3686 ( n3176, n3175, n670 );
nand U3687 ( n3161, n3159, n3158 );
nand U3688 ( n3158, n3157, n668 );
nand U3689 ( n3174, n3172, n3171 );
not U3690 ( n681, outData_in[12] );
xor U3691 ( n3720, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[34], n650 );
nand U3692 ( n3189, n3187, n3186 );
nand U3693 ( n736, n735, n734 );
xor U3694 ( my_IIR_filter_firBlock_right_multProducts[107], n3567, n490 );
nand U3695 ( n3737, n3736, n653 );
nor U3696 ( n3569, n489, n154 );
nand U3697 ( n3727, n3726, n651 );
nand U3698 ( n3680, n3679, n643 );
or U3699 ( n2653, n490, n154 );
xnor U3700 ( my_IIR_filter_firBlock_right_multProducts[81], n489, n2651 );
nand U3701 ( n3671, n3670, n641 );
nand U3702 ( n2889, n489, n2886 );
or U3703 ( n2887, n2886, n490 );
nor U3704 ( n3382, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[22], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[21] );
xor U3705 ( my_IIR_filter_firBlock_right_multProducts[15], n3380, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[22] );
nand U3706 ( n2880, n490, n2879 );
not U3707 ( n691, n489 );
or U3708 ( n741, n541, n542 );
nor U3709 ( n542, n740, leftOut[13] );
or U3710 ( n782, n543, n544 );
nor U3711 ( n544, n781, leftOut[25] );
or U3712 ( n785, n545, n546 );
nor U3713 ( n546, n784, leftOut[26] );
nand U3714 ( n797, n795, n794 );
xnor U3715 ( n3164, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[29], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[35] );
and U3716 ( n798, n797, leftOut[30] );
nand U3717 ( n801, n711, n712 );
xor U3718 ( my_IIR_filter_firBlock_left_N5, n1214, n1213 );
xor U3719 ( my_IIR_filter_firBlock_left_N13, n1122, n1121 );
xor U3720 ( my_IIR_filter_firBlock_left_N23, n1169, n1168 );
xor U3721 ( n1153, my_IIR_filter_firBlock_left_multProducts[62], my_IIR_filter_firBlock_left_firStep[257] );
xor U3722 ( n2407, my_IIR_filter_firBlock_left_multProducts[62], my_IIR_filter_firBlock_left_firStep[33] );
and U3723 ( n1208, n1207, my_IIR_filter_firBlock_left_firStep[286] );
nand U3724 ( n1205, my_IIR_filter_firBlock_left_firStep[285], n1202 );
or U3725 ( n1203, n1202, my_IIR_filter_firBlock_left_firStep[285] );
nand U3726 ( n1194, my_IIR_filter_firBlock_left_firStep[283], n1191 );
or U3727 ( n1192, n1191, my_IIR_filter_firBlock_left_firStep[283] );
nand U3728 ( n1185, my_IIR_filter_firBlock_left_firStep[281], n1182 );
or U3729 ( n1183, n1182, my_IIR_filter_firBlock_left_firStep[281] );
nand U3730 ( n1176, my_IIR_filter_firBlock_left_firStep[279], n1173 );
or U3731 ( n1174, n1173, my_IIR_filter_firBlock_left_firStep[279] );
nand U3732 ( n1172, my_IIR_filter_firBlock_left_firStep[278], n1169 );
or U3733 ( n1170, n1169, my_IIR_filter_firBlock_left_firStep[278] );
nand U3734 ( n1167, my_IIR_filter_firBlock_left_firStep[277], n1164 );
or U3735 ( n1165, n1164, my_IIR_filter_firBlock_left_firStep[277] );
nand U3736 ( n1158, my_IIR_filter_firBlock_left_firStep[275], n1155 );
or U3737 ( n1156, n1155, my_IIR_filter_firBlock_left_firStep[275] );
nand U3738 ( n1147, my_IIR_filter_firBlock_left_firStep[273], n1144 );
or U3739 ( n1145, n1144, my_IIR_filter_firBlock_left_firStep[273] );
nand U3740 ( n1138, my_IIR_filter_firBlock_left_firStep[271], n1135 );
or U3741 ( n1136, n1135, my_IIR_filter_firBlock_left_firStep[271] );
nand U3742 ( n1129, my_IIR_filter_firBlock_left_firStep[269], n1126 );
or U3743 ( n1127, n1126, my_IIR_filter_firBlock_left_firStep[269] );
nand U3744 ( n1125, my_IIR_filter_firBlock_left_firStep[268], n1122 );
or U3745 ( n1123, n1122, my_IIR_filter_firBlock_left_firStep[268] );
nand U3746 ( n1120, my_IIR_filter_firBlock_left_firStep[267], n1117 );
or U3747 ( n1118, n1117, my_IIR_filter_firBlock_left_firStep[267] );
nand U3748 ( n1111, my_IIR_filter_firBlock_left_firStep[265], n1221 );
or U3749 ( n1109, n1221, my_IIR_filter_firBlock_left_firStep[265] );
nand U3750 ( n1105, my_IIR_filter_firBlock_left_firStep[263], n1218 );
or U3751 ( n1103, n1218, my_IIR_filter_firBlock_left_firStep[263] );
nand U3752 ( n1668, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[14], n1665 );
or U3753 ( n1666, n1665, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[14] );
nand U3754 ( n1099, my_IIR_filter_firBlock_left_firStep[261], n1215 );
xor U3755 ( n1664, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[14], n294 );
or U3756 ( n1097, n1215, my_IIR_filter_firBlock_left_firStep[261] );
nand U3757 ( n1096, my_IIR_filter_firBlock_left_firStep[260], n1214 );
or U3758 ( n1094, n1214, my_IIR_filter_firBlock_left_firStep[260] );
nand U3759 ( n1093, my_IIR_filter_firBlock_left_firStep[259], n1212 );
or U3760 ( n1091, n1212, my_IIR_filter_firBlock_left_firStep[259] );
nand U3761 ( n2340, my_IIR_filter_firBlock_left_multProducts[62], n2339 );
nand U3762 ( n1086, my_IIR_filter_firBlock_left_multProducts[62], n1085 );
nand U3763 ( n964, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[14], n1082 );
or U3764 ( n962, n1082, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[14] );
xor U3765 ( n1081, inData_in[5], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[14] );
xor U3766 ( n1343, inData_in[5], inData_in[1] );
xor U3767 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[8], n916, n915 );
nand U3768 ( n1224, inData_in[1], n1344 );
or U3769 ( n1222, inData_in[1], n1344 );
nand U3770 ( n950, inData_in[1], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[10] );
or U3771 ( n947, inData_in[1], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[10] );
xor U3772 ( n933, inData_in[3], inData_in[1] );
nand U3773 ( n714, rightOut[3], n713 );
or U3774 ( n3157, n3156, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[27] );
or U3775 ( n3152, n3151, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[26] );
not U3776 ( n664, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[27] );
xor U3777 ( n3001, n688, outData_in[21] );
nand U3778 ( n3298, n3297, my_IIR_filter_firBlock_right_multProducts[51] );
nand U3779 ( n3278, n3277, my_IIR_filter_firBlock_right_multProducts[47] );
nand U3780 ( n3042, n492, n3039 );
or U3781 ( n3040, n3039, n492 );
nand U3782 ( n3039, n3037, n3036 );
nand U3783 ( n3016, n3014, n3013 );
nand U3784 ( n3006, n3005, n3004 );
nand U3785 ( n2993, n2992, n2991 );
nand U3786 ( n2981, n2980, n2979 );
nand U3787 ( n2958, n2955, n679 );
nor U3788 ( n2627, outData_in[5], n2628 );
or U3789 ( n2956, n679, n2955 );
xor U3790 ( my_IIR_filter_firBlock_right_multProducts[64], n2628, outData_in[5] );
nand U3791 ( n2822, outData_in[5], n2932 );
nand U3792 ( n3062, n2948, n2947 );
or U3793 ( n2820, n2932, outData_in[5] );
nand U3794 ( n2945, n3059, n518 );
nand U3795 ( n2815, outData_in[5], n2814 );
nand U3796 ( n2942, n2941, n133 );
nand U3797 ( n758, leftOut[18], n756 );
nand U3798 ( n720, leftOut[5], n804 );
xor U3799 ( my_IIR_filter_firBlock_left_N237, n2376, n2375 );
xor U3800 ( my_IIR_filter_firBlock_left_N247, n2423, n2422 );
and U3801 ( n2462, n2461, my_IIR_filter_firBlock_left_firStep[62] );
nand U3802 ( n2459, my_IIR_filter_firBlock_left_firStep[61], n2456 );
or U3803 ( n2457, n2456, my_IIR_filter_firBlock_left_firStep[61] );
nand U3804 ( n2448, my_IIR_filter_firBlock_left_firStep[59], n2445 );
or U3805 ( n2446, n2445, my_IIR_filter_firBlock_left_firStep[59] );
nand U3806 ( n2439, my_IIR_filter_firBlock_left_firStep[57], n2436 );
or U3807 ( n2437, n2436, my_IIR_filter_firBlock_left_firStep[57] );
nand U3808 ( n2430, my_IIR_filter_firBlock_left_firStep[55], n2427 );
or U3809 ( n2428, n2427, my_IIR_filter_firBlock_left_firStep[55] );
nand U3810 ( n2426, my_IIR_filter_firBlock_left_firStep[54], n2423 );
or U3811 ( n2424, n2423, my_IIR_filter_firBlock_left_firStep[54] );
nand U3812 ( n2421, my_IIR_filter_firBlock_left_firStep[53], n2418 );
or U3813 ( n2419, n2418, my_IIR_filter_firBlock_left_firStep[53] );
nand U3814 ( n2412, my_IIR_filter_firBlock_left_firStep[51], n2409 );
or U3815 ( n2410, n2409, my_IIR_filter_firBlock_left_firStep[51] );
nand U3816 ( n2401, my_IIR_filter_firBlock_left_firStep[49], n2398 );
or U3817 ( n2399, n2398, my_IIR_filter_firBlock_left_firStep[49] );
nand U3818 ( n2392, my_IIR_filter_firBlock_left_firStep[47], n2389 );
or U3819 ( n2390, n2389, my_IIR_filter_firBlock_left_firStep[47] );
nand U3820 ( n2383, my_IIR_filter_firBlock_left_firStep[45], n2380 );
or U3821 ( n2381, n2380, my_IIR_filter_firBlock_left_firStep[45] );
nand U3822 ( n2379, my_IIR_filter_firBlock_left_firStep[44], n2376 );
or U3823 ( n2377, n2376, my_IIR_filter_firBlock_left_firStep[44] );
nand U3824 ( n2374, my_IIR_filter_firBlock_left_firStep[43], n2371 );
or U3825 ( n2372, n2371, my_IIR_filter_firBlock_left_firStep[43] );
nand U3826 ( n1688, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[18], n1685 );
or U3827 ( n1686, n1685, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[18] );
nand U3828 ( n2365, my_IIR_filter_firBlock_left_firStep[41], n2475 );
xor U3829 ( n1684, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[18], n296 );
or U3830 ( n2363, n2475, my_IIR_filter_firBlock_left_firStep[41] );
nand U3831 ( n1098, my_IIR_filter_firBlock_left_multProducts[66], n1097 );
nand U3832 ( n2352, my_IIR_filter_firBlock_left_multProducts[66], n2351 );
nand U3833 ( n981, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[18], n978 );
or U3834 ( n979, n978, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[18] );
nand U3835 ( n841, my_IIR_filter_firBlock_left_multProducts[94], n838 );
xor U3836 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[18], n838, n837 );
or U3837 ( n839, n838, my_IIR_filter_firBlock_left_multProducts[94] );
or U3838 ( n828, n946, my_IIR_filter_firBlock_left_multProducts[91] );
nand U3839 ( n826, inData_in[5], n942 );
or U3840 ( n824, n942, inData_in[5] );
xor U3841 ( n915, inData_in[2], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[6] );
xor U3842 ( my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[7], inData_in[1], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nor U3843 ( n1632, my_IIR_filter_firBlock_left_multProducts[90], n41 );
and U3844 ( n1344, inData_in[4], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nor U3845 ( n1629, inData_in[1], my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nand U3846 ( n1628, my_IIR_filter_firBlock_left_multProducts[90], n41 );
nand U3847 ( n949, n948, my_IIR_filter_firBlock_left_my_IIR_filter_firBlock_left_MultiplyBlock_w192[6] );
nand U3848 ( n812, n41, n916 );
nand U3849 ( n916, n41, n40 );
xor U3850 ( my_IIR_filter_firBlock_right_N109, n3258, n3257 );
nand U3851 ( n3300, n3299, n3298 );
nand U3852 ( n3261, my_IIR_filter_firBlock_right_firStep[43], n3258 );
or U3853 ( n3259, n3258, my_IIR_filter_firBlock_right_firStep[43] );
nand U3854 ( n3256, my_IIR_filter_firBlock_right_firStep[42], n3253 );
or U3855 ( n3254, n3253, my_IIR_filter_firBlock_right_firStep[42] );
nand U3856 ( n3240, n3239, my_IIR_filter_firBlock_right_multProducts[38] );
or U3857 ( n3373, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[16], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[15] );
nor U3858 ( n3371, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[15], n3372 );
xor U3859 ( my_IIR_filter_firBlock_right_multProducts[8], n3372, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[15] );
not U3860 ( n634, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[15] );
nand U3861 ( n804, n716, n717 );
nand U3862 ( n790, n789, n788 );
nand U3863 ( n774, leftOut[22], n771 );
nand U3864 ( n756, n755, n754 );
nand U3865 ( n752, leftOut[16], n750 );
xor U3866 ( n3304, my_IIR_filter_firBlock_right_multProducts[53], my_IIR_filter_firBlock_right_firStep[53] );
nand U3867 ( n3202, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[36], n3199 );
or U3868 ( n3200, n3199, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[36] );
nor U3869 ( n3394, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[30], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[29] );
xor U3870 ( my_IIR_filter_firBlock_right_multProducts[23], n3392, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[30] );
not U3871 ( n647, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[30] );
xor U3872 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[33], n3030, n3029 );
nand U3873 ( n3032, n505, n3030 );
nand U3874 ( n3028, n157, n3025 );
or U3875 ( n3026, n3025, n157 );
nand U3876 ( n3013, n3012, n692 );
nand U3877 ( n2642, n2643, n684 );
xor U3878 ( my_IIR_filter_firBlock_right_multProducts[74], n684, n2643 );
nand U3879 ( n2988, n495, n2985 );
xor U3880 ( n2984, n684, outData_in[17] );
or U3881 ( n2986, n2985, n496 );
nand U3882 ( n2979, n2978, n684 );
nand U3883 ( n3742, n525, n3739 );
or U3884 ( n3740, n3739, n525 );
or U3885 ( n3543, n523, n501 );
nand U3886 ( n3702, n3700, n3699 );
nand U3887 ( n3700, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[29], n3697 );
or U3888 ( n3698, n3697, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[29] );
xor U3889 ( my_IIR_filter_firBlock_right_multProducts[48], n3678, n3677 );
nand U3890 ( n3681, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[25], n3678 );
or U3891 ( n3679, n3678, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[25] );
nand U3892 ( n3653, n3652, n637 );
nand U3893 ( n3644, n3643, n125 );
nand U3894 ( n3635, n3634, n634 );
nand U3895 ( n3636, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[15], n3633 );
or U3896 ( n3634, n3633, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[15] );
nand U3897 ( n3610, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[9], n3746 );
or U3898 ( n3608, n3746, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[9] );
nand U3899 ( n3072, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[8], n3218 );
nand U3900 ( n3605, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[7], n3602 );
nor U3901 ( n3603, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[7], n3602 );
or U3902 ( n3070, n3218, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[8] );
or U3903 ( n2625, n523, n501 );
xor U3904 ( n2927, n518, n523 );
nand U3905 ( n2813, n523, n2928 );
or U3906 ( n2811, n2928, n522 );
xor U3907 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[3], n522, n498 );
nand U3908 ( n2940, n522, n3056 );
nor U3909 ( n3064, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[8], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[7] );
xnor U3910 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[2], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[8], n3165 );
and U3911 ( n2926, n522, n498 );
not U3912 ( n706, n523 );
nand U3913 ( n3210, n3209, n547 );
nand U3914 ( n3206, n3205, n547 );
nand U3915 ( n3201, n3200, n547 );
nand U3916 ( n3186, n3185, n547 );
nand U3917 ( n786, leftOut[26], n784 );
nand U3918 ( n771, n769, n768 );
nand U3919 ( n750, n749, n748 );
xor U3920 ( my_IIR_filter_firBlock_right_N115, n3285, n3284 );
xor U3921 ( my_IIR_filter_firBlock_right_multProducts[103], n3561, outData_in[18] );
xor U3922 ( n3248, my_IIR_filter_firBlock_right_multProducts[41], my_IIR_filter_firBlock_right_firStep[41] );
nand U3923 ( n3339, my_IIR_filter_firBlock_right_multProducts[60], n3338 );
nor U3924 ( n3563, outData_in[18], n512 );
nand U3925 ( n3291, n3288, n3287 );
nand U3926 ( n3288, my_IIR_filter_firBlock_right_firStep[49], n3285 );
nand U3927 ( n3280, n3279, n3278 );
nand U3928 ( n3276, n3274, n3273 );
xnor U3929 ( n3140, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[24], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[30] );
or U3930 ( n2647, outData_in[18], n513 );
xnor U3931 ( my_IIR_filter_firBlock_right_multProducts[77], outData_in[18], n2645 );
nand U3932 ( n2873, outData_in[18], n2870 );
nor U3933 ( n3376, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[18], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[17] );
xor U3934 ( my_IIR_filter_firBlock_right_multProducts[11], n3374, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[18] );
or U3935 ( n2871, n2870, outData_in[18] );
not U3936 ( n636, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[18] );
nand U3937 ( n2863, outData_in[18], n2862 );
xnor U3938 ( n3113, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[24], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[18] );
not U3939 ( n687, outData_in[18] );
nand U3940 ( n725, leftOut[8], n809 );
xor U3941 ( my_IIR_filter_firBlock_right_N187, n3510, n3509 );
xor U3942 ( my_IIR_filter_firBlock_right_N177, n3463, n3462 );
xor U3943 ( my_IIR_filter_firBlock_right_N169, n3541, n3540 );
xor U3944 ( my_IIR_filter_firBlock_right_N181, n3483, n3482 );
xor U3945 ( my_IIR_filter_firBlock_right_N167, n3538, n3537 );
xor U3946 ( my_IIR_filter_firBlock_right_N171, n3436, n3435 );
xor U3947 ( my_IIR_filter_firBlock_right_N175, n3454, n3453 );
xor U3948 ( my_IIR_filter_firBlock_right_N179, n3472, n3471 );
xor U3949 ( my_IIR_filter_firBlock_right_N183, n3492, n3491 );
nor U3950 ( n3531, n3528, n215 );
nand U3951 ( n3521, my_IIR_filter_firBlock_right_firStep[28], n3518 );
or U3952 ( n3519, n3518, my_IIR_filter_firBlock_right_firStep[28] );
nand U3953 ( n3513, my_IIR_filter_firBlock_right_firStep[26], n3510 );
or U3954 ( n3511, n3510, my_IIR_filter_firBlock_right_firStep[26] );
nand U3955 ( n3510, n3508, n3507 );
nand U3956 ( n3495, my_IIR_filter_firBlock_right_firStep[22], n3492 );
or U3957 ( n3493, n3492, my_IIR_filter_firBlock_right_firStep[22] );
nand U3958 ( n3486, my_IIR_filter_firBlock_right_firStep[20], n3483 );
or U3959 ( n3484, n3483, my_IIR_filter_firBlock_right_firStep[20] );
nand U3960 ( n3475, my_IIR_filter_firBlock_right_firStep[18], n3472 );
or U3961 ( n3473, n3472, my_IIR_filter_firBlock_right_firStep[18] );
nand U3962 ( n3466, my_IIR_filter_firBlock_right_firStep[16], n3463 );
or U3963 ( n3464, n3463, my_IIR_filter_firBlock_right_firStep[16] );
nand U3964 ( n3457, my_IIR_filter_firBlock_right_firStep[14], n3454 );
or U3965 ( n3455, n3454, my_IIR_filter_firBlock_right_firStep[14] );
nand U3966 ( n3445, n3443, n3442 );
nand U3967 ( n3439, my_IIR_filter_firBlock_right_firStep[10], n3436 );
or U3968 ( n3437, n3436, my_IIR_filter_firBlock_right_firStep[10] );
nand U3969 ( n3431, my_IIR_filter_firBlock_right_firStep[8], n3541 );
or U3970 ( n3429, n3541, my_IIR_filter_firBlock_right_firStep[8] );
nand U3971 ( n3425, my_IIR_filter_firBlock_right_firStep[6], n3538 );
or U3972 ( n3423, n3538, my_IIR_filter_firBlock_right_firStep[6] );
nand U3973 ( n3092, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[13], n3091 );
nand U3974 ( n3536, n3419, n3418 );
or U3975 ( n3361, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[8], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[7] );
or U3976 ( n3604, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[7], n3603 );
nor U3977 ( n3407, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[7], n3406 );
xor U3978 ( my_IIR_filter_firBlock_right_multProducts[0], n3406, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[7] );
not U3979 ( n674, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[13] );
nand U3980 ( n3337, n3334, n3333 );
nand U3981 ( n3305, n3302, n3303 );
nand U3982 ( n3302, my_IIR_filter_firBlock_right_multProducts[52], n3301 );
nand U3983 ( n784, n783, n782 );
nand U3984 ( n729, n727, n726 );
nand U3985 ( n809, n723, n722 );
xor U3986 ( my_IIR_filter_firBlock_right_multProducts[92], n3583, outData_in[7] );
nor U3987 ( n3584, outData_in[7], n3583 );
nand U3988 ( n3342, n3340, n3339 );
nand U3989 ( n3187, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[33], n3184 );
nand U3990 ( n3309, n3308, n3307 );
or U3991 ( n3185, n3184, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[33] );
xnor U3992 ( n3183, n525, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[33] );
or U3993 ( n3391, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[28], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[27] );
nor U3994 ( n3389, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[27], n3390 );
nand U3995 ( n3293, my_IIR_filter_firBlock_right_multProducts[50], n3292 );
xor U3996 ( my_IIR_filter_firBlock_right_multProducts[20], n3390, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[27] );
not U3997 ( n645, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[27] );
not U3998 ( n668, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[33] );
xnor U3999 ( n3155, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[27], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[33] );
nand U4000 ( n3014, n154, n3011 );
or U4001 ( n3012, n3011, n154 );
nand U4002 ( n3009, outData_in[20], n3006 );
or U4003 ( n3007, n3006, outData_in[20] );
nand U4004 ( n2997, n2996, n2995 );
nand U4005 ( n2996, n513, n2993 );
or U4006 ( n2994, n2993, n512 );
nand U4007 ( n2983, n485, n2981 );
xor U4008 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[20], n2972, n2971 );
nand U4009 ( n2630, n2631, n702 );
xor U4010 ( my_IIR_filter_firBlock_right_multProducts[66], n702, n2631 );
nand U4011 ( n2962, n2959, n680 );
nand U4012 ( n2827, outData_in[7], n2826 );
nand U4013 ( n2954, outData_in[7], n3063 );
nand U4014 ( n2821, outData_in[7], n2820 );
nand U4015 ( n2947, n2946, n702 );
not U4016 ( n702, outData_in[7] );
nand U4017 ( n810, n725, n724 );
nand U4018 ( n3109, n3107, n3106 );
nand U4019 ( n3106, n3105, n660 );
nand U4020 ( n3118, n3116, n3115 );
nand U4021 ( n3166, n3163, n3162 );
nand U4022 ( n3194, n3192, n3191 );
nand U4023 ( n3191, n3190, n547 );
nand U4024 ( n3128, n3126, n3125 );
nand U4025 ( n3125, n3124, n663 );
nand U4026 ( n3146, n3144, n3143 );
nand U4027 ( n3143, n3142, n665 );
nand U4028 ( n3156, n3154, n3153 );
nand U4029 ( n3153, n3152, n667 );
nand U4030 ( n3170, n3169, n3168 );
nand U4031 ( n3168, n3167, n669 );
nand U4032 ( n3184, n3182, n3181 );
nand U4033 ( n3181, n3180, n671 );
nand U4034 ( n3151, n3149, n3148 );
nand U4035 ( n3148, n3147, n666 );
nand U4036 ( n3137, n3135, n3134 );
nand U4037 ( n3199, n3197, n3196 );
nand U4038 ( n3196, n3195, n547 );
nand U4039 ( n2972, n2970, n2969 );
nand U4040 ( n787, n786, n785 );
nor U4041 ( n800, n799, n798 );
xor U4042 ( n3706, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[31], n648 );
xnor U4043 ( my_IIR_filter_firBlock_right_multProducts[93], n507, n3584 );
xor U4044 ( my_IIR_filter_firBlock_right_multProducts[60], n3735, n3734 );
nand U4045 ( n3738, n525, n3735 );
or U4046 ( n3736, n3735, n525 );
nand U4047 ( n3725, n3723, n3722 );
or U4048 ( n3548, n506, outData_in[7] );
xor U4049 ( my_IIR_filter_firBlock_right_multProducts[54], n3707, n3706 );
nand U4050 ( n3710, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[31], n3707 );
or U4051 ( n3708, n3707, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[31] );
xor U4052 ( my_IIR_filter_firBlock_right_multProducts[51], n3693, n3692 );
nand U4053 ( n3696, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[28], n3693 );
or U4054 ( n3694, n3693, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[28] );
xor U4055 ( my_IIR_filter_firBlock_right_multProducts[50], n3688, n3687 );
nand U4056 ( n3691, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[27], n3688 );
or U4057 ( n3689, n3688, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[27] );
xor U4058 ( my_IIR_filter_firBlock_right_multProducts[47], n3674, n3673 );
nand U4059 ( n3676, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[24], n3674 );
nand U4060 ( n3669, n3667, n3666 );
nand U4061 ( n3663, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[21], n3660 );
or U4062 ( n3661, n3660, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[21] );
xor U4063 ( my_IIR_filter_firBlock_right_multProducts[42], n3651, n3650 );
nand U4064 ( n3654, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[19], n3651 );
or U4065 ( n3652, n3651, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[19] );
xor U4066 ( my_IIR_filter_firBlock_right_multProducts[40], n3642, n3641 );
nand U4067 ( n3645, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[17], n3642 );
or U4068 ( n3643, n3642, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[17] );
nand U4069 ( n3627, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[13], n3624 );
nand U4070 ( n3097, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[14], n3096 );
or U4071 ( n3625, n3624, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[13] );
xnor U4072 ( n3094, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[14], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[20] );
xor U4073 ( my_IIR_filter_firBlock_right_multProducts[34], n3616, n3615 );
nand U4074 ( n3623, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[12], n3620 );
or U4075 ( n3621, n3620, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[12] );
xor U4076 ( my_IIR_filter_firBlock_right_multProducts[33], n3612, n3611 );
nor U4077 ( n2632, n507, outData_in[7] );
nand U4078 ( n3619, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[11], n3616 );
xor U4079 ( my_IIR_filter_firBlock_right_multProducts[67], n2630, n506 );
or U4080 ( n3617, n3616, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[11] );
nand U4081 ( n3614, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[10], n3612 );
nand U4082 ( n2832, n506, n2829 );
or U4083 ( n2830, n2829, n507 );
nand U4084 ( n2957, n506, n2956 );
nand U4085 ( n2825, n506, n2934 );
not U4086 ( n673, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[14] );
or U4087 ( n2823, n2934, n507 );
not U4088 ( n701, n506 );
nand U4089 ( n3307, my_IIR_filter_firBlock_right_multProducts[53], n3306 );
nand U4090 ( n3287, n3286, my_IIR_filter_firBlock_right_multProducts[49] );
or U4091 ( n3286, n3285, my_IIR_filter_firBlock_right_firStep[49] );
nand U4092 ( n3243, n3242, my_IIR_filter_firBlock_right_multProducts[39] );
nand U4093 ( n3329, my_IIR_filter_firBlock_right_multProducts[58], n3328 );
nand U4094 ( n3323, n3321, n3320 );
nand U4095 ( n3320, n3319, my_IIR_filter_firBlock_right_multProducts[56] );
nand U4096 ( n3285, n3283, n3282 );
nand U4097 ( n3282, my_IIR_filter_firBlock_right_multProducts[48], n3281 );
nand U4098 ( n3269, n3268, my_IIR_filter_firBlock_right_multProducts[45] );
nand U4099 ( n3253, n3252, n3251 );
nand U4100 ( n3251, n3250, my_IIR_filter_firBlock_right_multProducts[41] );
nand U4101 ( n747, n746, n745 );
nand U4102 ( n3721, n3719, n3718 );
nand U4103 ( n3718, n3717, n128 );
nand U4104 ( n767, n766, n765 );
nand U4105 ( n733, n731, n730 );
nand U4106 ( n753, n752, n751 );
nand U4107 ( n764, n763, n762 );
nand U4108 ( n744, n741, n742 );
nand U4109 ( n3693, n3691, n3690 );
nand U4110 ( n3690, n3689, n645 );
nand U4111 ( n3735, n3733, n3732 );
nand U4112 ( n3732, n3731, n652 );
nand U4113 ( n3707, n3705, n3704 );
nand U4114 ( n3704, n3703, n647 );
nand U4115 ( n3743, n3742, n3741 );
nand U4116 ( n773, rightOut[22], n772 );
xnor U4117 ( n3145, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[25], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[31] );
nand U4118 ( n781, n780, n779 );
xor U4119 ( n3313, my_IIR_filter_firBlock_right_multProducts[55], my_IIR_filter_firBlock_right_firStep[55] );
nand U4120 ( n3316, my_IIR_filter_firBlock_right_multProducts[55], n3315 );
or U4121 ( n3397, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[32], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[31] );
xnor U4122 ( my_IIR_filter_firBlock_right_multProducts[25], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[32], n3395 );
not U4123 ( n649, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[32] );
nor U4124 ( n3545, n518, n503 );
nand U4125 ( n3050, n3049, n548 );
nand U4126 ( n3051, n514, n3048 );
or U4127 ( n3049, n3048, n514 );
nand U4128 ( n3036, n3035, n697 );
nand U4129 ( n3037, n158, n3034 );
or U4130 ( n3035, n3034, n158 );
nand U4131 ( n3023, outData_in[23], n3020 );
or U4132 ( n3021, n3020, outData_in[23] );
nand U4133 ( n3018, n489, n3016 );
nand U4134 ( n3005, n494, n3002 );
or U4135 ( n3003, n3002, n494 );
nand U4136 ( n3000, outData_in[18], n2997 );
or U4137 ( n2998, n2997, outData_in[18] );
nand U4138 ( n2991, n2990, n687 );
nand U4139 ( n2992, outData_in[16], n2989 );
or U4140 ( n2990, n2989, outData_in[16] );
nand U4141 ( n2975, n510, n2972 );
or U4142 ( n2973, n2972, n510 );
nand U4143 ( n2963, n2962, n2961 );
nand U4144 ( n2959, n2957, n2958 );
nor U4145 ( n2626, n518, n503 );
nand U4146 ( n2669, n2668, n705 );
xor U4147 ( my_IIR_filter_firBlock_right_multProducts[62], n705, n2668 );
xor U4148 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[13], n3061, n3060 );
nand U4149 ( n2948, outData_in[5], n3061 );
nand U4150 ( n2816, n503, n2929 );
or U4151 ( n2814, n2929, n503 );
nand U4152 ( n2943, n503, n3058 );
nand U4153 ( n2809, n503, n2808 );
or U4154 ( n2941, n3058, n503 );
nand U4155 ( n2937, n2936, n705 );
not U4156 ( n705, n502 );
xor U4157 ( my_IIR_filter_firBlock_right_N173, n3445, n3444 );
xor U4158 ( my_IIR_filter_firBlock_right_N165, n3535, n3534 );
xor U4159 ( my_IIR_filter_firBlock_right_N185, n3501, n3500 );
and U4160 ( n3530, n3529, my_IIR_filter_firBlock_right_firStep[30] );
nand U4161 ( n3527, my_IIR_filter_firBlock_right_firStep[29], n3524 );
or U4162 ( n3525, n3524, my_IIR_filter_firBlock_right_firStep[29] );
nand U4163 ( n3517, my_IIR_filter_firBlock_right_firStep[27], n3514 );
or U4164 ( n3515, n3514, my_IIR_filter_firBlock_right_firStep[27] );
nand U4165 ( n3508, my_IIR_filter_firBlock_right_firStep[25], n3505 );
or U4166 ( n3506, n3505, my_IIR_filter_firBlock_right_firStep[25] );
nand U4167 ( n3504, my_IIR_filter_firBlock_right_firStep[24], n3501 );
or U4168 ( n3502, n3501, my_IIR_filter_firBlock_right_firStep[24] );
nor U4169 ( n3544, n521, outData_in[5] );
nand U4170 ( n3499, my_IIR_filter_firBlock_right_firStep[23], n3496 );
or U4171 ( n3497, n3496, my_IIR_filter_firBlock_right_firStep[23] );
nand U4172 ( n3490, my_IIR_filter_firBlock_right_firStep[21], n3487 );
or U4173 ( n3488, n3487, my_IIR_filter_firBlock_right_firStep[21] );
nand U4174 ( n3481, my_IIR_filter_firBlock_right_firStep[19], n3478 );
or U4175 ( n3479, n3478, my_IIR_filter_firBlock_right_firStep[19] );
nand U4176 ( n3470, my_IIR_filter_firBlock_right_firStep[17], n3467 );
or U4177 ( n3468, n3467, my_IIR_filter_firBlock_right_firStep[17] );
nand U4178 ( n3461, my_IIR_filter_firBlock_right_firStep[15], n3458 );
or U4179 ( n3459, n3458, my_IIR_filter_firBlock_right_firStep[15] );
nand U4180 ( n3452, my_IIR_filter_firBlock_right_firStep[13], n3449 );
or U4181 ( n3450, n3449, my_IIR_filter_firBlock_right_firStep[13] );
nand U4182 ( n3448, my_IIR_filter_firBlock_right_firStep[12], n3445 );
or U4183 ( n3446, n3445, my_IIR_filter_firBlock_right_firStep[12] );
nand U4184 ( n3443, my_IIR_filter_firBlock_right_firStep[11], n3440 );
or U4185 ( n3441, n3440, my_IIR_filter_firBlock_right_firStep[11] );
nand U4186 ( n3434, my_IIR_filter_firBlock_right_firStep[9], n3542 );
or U4187 ( n3432, n3542, my_IIR_filter_firBlock_right_firStep[9] );
nand U4188 ( n3428, my_IIR_filter_firBlock_right_firStep[7], n3539 );
or U4189 ( n3426, n3539, my_IIR_filter_firBlock_right_firStep[7] );
nand U4190 ( n3422, my_IIR_filter_firBlock_right_firStep[5], n3536 );
or U4191 ( n3420, n3536, my_IIR_filter_firBlock_right_firStep[5] );
nand U4192 ( n3088, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[12], n3087 );
nand U4193 ( n3419, my_IIR_filter_firBlock_right_firStep[4], n3535 );
or U4194 ( n3417, n3535, my_IIR_filter_firBlock_right_firStep[4] );
nand U4195 ( n3416, my_IIR_filter_firBlock_right_firStep[3], n3533 );
or U4196 ( n3414, n3533, my_IIR_filter_firBlock_right_firStep[3] );
or U4197 ( n2629, n520, outData_in[5] );
xnor U4198 ( my_IIR_filter_firBlock_right_multProducts[65], n521, n2627 );
xor U4199 ( n2933, n520, n507 );
nand U4200 ( n2824, n520, n2823 );
or U4201 ( n3600, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[6], n3599 );
xor U4202 ( n2930, n521, n517 );
nor U4203 ( n3357, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[6], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[5] );
nand U4204 ( n2951, n521, n3062 );
nand U4205 ( n2818, n521, n2817 );
or U4206 ( n2949, n3062, n520 );
not U4207 ( n675, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[12] );
not U4208 ( n703, n520 );
xor U4209 ( my_IIR_filter_firBlock_right_N113, n3276, n3275 );
xor U4210 ( my_IIR_filter_firBlock_right_N103, n3351, n3350 );
xor U4211 ( my_IIR_filter_firBlock_right_N105, n3354, n3353 );
xor U4212 ( my_IIR_filter_firBlock_right_N119, n3305, n3304 );
xor U4213 ( my_IIR_filter_firBlock_right_N121, n3314, n3313 );
xor U4214 ( my_IIR_filter_firBlock_right_N111, n3267, n3266 );
xnor U4215 ( my_IIR_filter_firBlock_right_multProducts[94], n519, n3550 );
and U4216 ( n3343, n3342, my_IIR_filter_firBlock_right_firStep[61] );
xor U4217 ( n3289, my_IIR_filter_firBlock_right_multProducts[32], my_IIR_filter_firBlock_right_firStep[32] );
nand U4218 ( n3340, my_IIR_filter_firBlock_right_firStep[60], n3337 );
nand U4219 ( n3317, my_IIR_filter_firBlock_right_firStep[55], n3314 );
nand U4220 ( n3308, my_IIR_filter_firBlock_right_firStep[53], n3305 );
or U4221 ( n3306, n3305, my_IIR_filter_firBlock_right_firStep[53] );
nand U4222 ( n3303, my_IIR_filter_firBlock_right_firStep[52], n3300 );
or U4223 ( n3301, n3300, my_IIR_filter_firBlock_right_firStep[52] );
nand U4224 ( n3279, my_IIR_filter_firBlock_right_firStep[47], n3276 );
or U4225 ( n3277, n3276, my_IIR_filter_firBlock_right_firStep[47] );
nand U4226 ( n3274, my_IIR_filter_firBlock_right_firStep[46], n3271 );
or U4227 ( n3272, n3271, my_IIR_filter_firBlock_right_firStep[46] );
nand U4228 ( n3271, n3270, n3269 );
nand U4229 ( n3270, my_IIR_filter_firBlock_right_firStep[45], n3267 );
nand U4230 ( n3244, my_IIR_filter_firBlock_right_firStep[39], n3354 );
or U4231 ( n3242, n3354, my_IIR_filter_firBlock_right_firStep[39] );
nand U4232 ( n3241, my_IIR_filter_firBlock_right_firStep[38], n3352 );
nand U4233 ( n3238, my_IIR_filter_firBlock_right_firStep[37], n3351 );
or U4234 ( n3236, n3351, my_IIR_filter_firBlock_right_firStep[37] );
nand U4235 ( n3101, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[15], n3100 );
nand U4236 ( n3235, my_IIR_filter_firBlock_right_firStep[36], n3349 );
nor U4237 ( n2633, n519, n2634 );
or U4238 ( n3233, n3349, my_IIR_filter_firBlock_right_firStep[36] );
xor U4239 ( my_IIR_filter_firBlock_right_multProducts[68], n2634, n519 );
nand U4240 ( n2836, n519, n2833 );
nor U4241 ( n3364, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[10], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[9] );
nand U4242 ( n3222, my_IIR_filter_firBlock_right_multProducts[32], n3221 );
or U4243 ( n2834, n2833, n519 );
xnor U4244 ( my_IIR_filter_firBlock_right_multProducts[2], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[9], n3363 );
nand U4245 ( n2961, n519, n2960 );
nand U4246 ( n2828, n519, n2935 );
not U4247 ( n655, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[9] );
or U4248 ( n2826, n2935, n519 );
nand U4249 ( n719, rightOut[5], n718 );
xor U4250 ( my_IIR_filter_firBlock_right_multProducts[95], n3549, n509 );
xor U4251 ( my_IIR_filter_firBlock_right_multProducts[30], n3405, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[38] );
not U4252 ( n654, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[38] );
nand U4253 ( n3197, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[35], n3194 );
or U4254 ( n3195, n3194, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[35] );
nor U4255 ( n3551, n509, n519 );
nand U4256 ( n3192, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[34], n3189 );
or U4257 ( n3190, n3189, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[34] );
xor U4258 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[32], n3179, n3178 );
nand U4259 ( n3182, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[32], n3179 );
or U4260 ( n3180, n3179, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[32] );
nand U4261 ( n3177, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[31], n3174 );
or U4262 ( n3175, n3174, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[31] );
nand U4263 ( n3169, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[29], n3166 );
or U4264 ( n3167, n3166, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[29] );
nand U4265 ( n3163, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[28], n3161 );
nand U4266 ( n3149, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[25], n3146 );
or U4267 ( n3147, n3146, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[25] );
xor U4268 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[24], n3141, n3140 );
nand U4269 ( n3144, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[24], n3141 );
or U4270 ( n3142, n3141, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[24] );
xor U4271 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[22], n3133, n3132 );
nand U4272 ( n3135, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[22], n3133 );
nand U4273 ( n3131, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[21], n3128 );
or U4274 ( n3129, n3128, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[21] );
xor U4275 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[20], n3123, n3122 );
nand U4276 ( n3126, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[20], n3123 );
or U4277 ( n3124, n3123, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[20] );
xor U4278 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[18], n3114, n3113 );
nand U4279 ( n3116, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[18], n3114 );
xor U4280 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[16], n3104, n3103 );
nand U4281 ( n3107, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[16], n3104 );
xnor U4282 ( n3103, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[22], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[16] );
or U4283 ( n3105, n3104, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[16] );
or U4284 ( n2635, n509, n519 );
xnor U4285 ( my_IIR_filter_firBlock_right_multProducts[69], n509, n2633 );
xor U4286 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[14], n3095, n3094 );
nand U4287 ( n3098, n3095, n659 );
or U4288 ( n3096, n659, n3095 );
nand U4289 ( n2840, n509, n2837 );
or U4290 ( n2838, n2837, n509 );
nand U4291 ( n3089, n3086, n658 );
or U4292 ( n3087, n658, n3086 );
nand U4293 ( n3084, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[11], n3083 );
nand U4294 ( n2966, n509, n2963 );
nand U4295 ( n2831, n509, n2830 );
xnor U4296 ( n3076, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[10], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[16] );
not U4297 ( n657, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[16] );
not U4298 ( n679, n508 );
nand U4299 ( n710, leftOut[1], n760 );
xor U4300 ( my_IIR_filter_firBlock_right_multProducts[96], n3553, n488 );
nor U4301 ( n3552, n487, n3553 );
xor U4302 ( my_IIR_filter_firBlock_right_multProducts[58], n3725, n3724 );
nand U4303 ( n3728, n525, n3725 );
or U4304 ( n3726, n3725, n525 );
xor U4305 ( my_IIR_filter_firBlock_right_multProducts[56], n3716, n3715 );
or U4306 ( n3554, n510, n488 );
nand U4307 ( n3719, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[33], n3716 );
or U4308 ( n3717, n3716, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[33] );
xor U4309 ( my_IIR_filter_firBlock_right_multProducts[55], n3712, n3711 );
nand U4310 ( n3714, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[32], n3712 );
xor U4311 ( my_IIR_filter_firBlock_right_multProducts[53], n3702, n3701 );
nand U4312 ( n3705, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[30], n3702 );
or U4313 ( n3703, n3702, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[30] );
xor U4314 ( my_IIR_filter_firBlock_right_multProducts[49], n3683, n3682 );
nand U4315 ( n3688, n3686, n3685 );
nand U4316 ( n3686, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[26], n3683 );
or U4317 ( n3684, n3683, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[26] );
xor U4318 ( my_IIR_filter_firBlock_right_multProducts[46], n3669, n3668 );
nand U4319 ( n3672, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[23], n3669 );
or U4320 ( n3670, n3669, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[23] );
nand U4321 ( n3667, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[22], n3664 );
or U4322 ( n3665, n3664, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[22] );
xor U4323 ( my_IIR_filter_firBlock_right_multProducts[43], n3656, n3655 );
nand U4324 ( n3659, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[20], n3656 );
or U4325 ( n3657, n3656, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[20] );
nand U4326 ( n3649, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[18], n3646 );
or U4327 ( n3647, n3646, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[18] );
xor U4328 ( my_IIR_filter_firBlock_right_multProducts[39], n3638, n3637 );
nor U4329 ( n2638, n510, n488 );
nand U4330 ( n3640, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[16], n3638 );
nand U4331 ( n3112, n163, n3109 );
or U4332 ( n3110, n3109, n163 );
xnor U4333 ( n3108, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[23], n163 );
xor U4334 ( my_IIR_filter_firBlock_right_multProducts[37], n3629, n3628 );
nand U4335 ( n3632, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[14], n3629 );
or U4336 ( n3630, n3629, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[14] );
nand U4337 ( n2844, n488, n2841 );
or U4338 ( n3367, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[12], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[11] );
nor U4339 ( n3365, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[11], n3366 );
or U4340 ( n2842, n2841, n487 );
xor U4341 ( my_IIR_filter_firBlock_right_multProducts[4], n3366, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[11] );
nand U4342 ( n2970, n487, n2967 );
nand U4343 ( n2835, n487, n2834 );
or U4344 ( n2968, n2967, n487 );
or U4345 ( n3085, n3082, n163 );
nand U4346 ( n3083, n163, n3082 );
xnor U4347 ( n3081, n676, n163 );
not U4348 ( n680, n528 );
nor U4349 ( my_IIR_filter_firBlock_right_multProducts[117], n3582, n525 );
xor U4350 ( n3734, n653, n524 );
xor U4351 ( my_IIR_filter_firBlock_right_multProducts[59], n3730, n3729 );
xor U4352 ( n3729, n652, n524 );
nand U4353 ( n3733, n525, n3730 );
or U4354 ( n3731, n3730, n525 );
xnor U4355 ( n3203, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[37], n524 );
nor U4356 ( my_IIR_filter_firBlock_right_multProducts[91], n2666, n525 );
xor U4357 ( n3724, n651, n524 );
xor U4358 ( my_IIR_filter_firBlock_right_multProducts[57], n3721, n3720 );
xnor U4359 ( n3198, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[36], n524 );
nand U4360 ( n3723, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10[34], n3721 );
xnor U4361 ( n3193, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[35], n524 );
xnor U4362 ( n3188, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[34], n524 );
xnor U4363 ( n2917, n514, n524 );
not U4364 ( n548, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w10_39 );
nor U4365 ( n799, n796, n58 );
nand U4366 ( n789, leftOut[27], n787 );
nand U4367 ( n783, leftOut[25], n781 );
nand U4368 ( n777, leftOut[23], n775 );
nand U4369 ( n769, leftOut[21], n767 );
nand U4370 ( n755, leftOut[17], n753 );
nand U4371 ( n749, leftOut[15], n747 );
nand U4372 ( n742, leftOut[13], n740 );
nand U4373 ( n735, leftOut[11], n733 );
nand U4374 ( n712, leftOut[2], n792 );
xor U4375 ( my_IIR_filter_firBlock_right_N107, n3249, n3248 );
xor U4376 ( my_IIR_filter_firBlock_right_N117, n3296, n3295 );
xnor U4377 ( my_IIR_filter_firBlock_right_multProducts[98], n499, n3556 );
nand U4378 ( n3330, my_IIR_filter_firBlock_right_firStep[58], n3327 );
nor U4379 ( n3557, n485, n499 );
nand U4380 ( n3314, n3312, n3311 );
nand U4381 ( n3312, my_IIR_filter_firBlock_right_firStep[54], n3309 );
or U4382 ( n3310, n3309, my_IIR_filter_firBlock_right_firStep[54] );
nand U4383 ( n3299, my_IIR_filter_firBlock_right_firStep[51], n3296 );
nand U4384 ( n3294, my_IIR_filter_firBlock_right_firStep[50], n3291 );
or U4385 ( n3292, n3291, my_IIR_filter_firBlock_right_firStep[50] );
nand U4386 ( n3283, my_IIR_filter_firBlock_right_firStep[48], n3280 );
or U4387 ( n3281, n3280, my_IIR_filter_firBlock_right_firStep[48] );
nand U4388 ( n3267, n3265, n3264 );
nand U4389 ( n3265, my_IIR_filter_firBlock_right_firStep[44], n3262 );
or U4390 ( n3263, n3262, my_IIR_filter_firBlock_right_firStep[44] );
nand U4391 ( n3252, my_IIR_filter_firBlock_right_firStep[41], n3249 );
or U4392 ( n2641, n485, n499 );
nor U4393 ( n2639, n499, n2640 );
nand U4394 ( n3121, n160, n3118 );
nand U4395 ( n3247, my_IIR_filter_firBlock_right_firStep[40], n3355 );
or U4396 ( n3119, n3118, n160 );
or U4397 ( n3245, n3355, my_IIR_filter_firBlock_right_firStep[40] );
xor U4398 ( my_IIR_filter_firBlock_right_multProducts[72], n2640, n499 );
xnor U4399 ( n3117, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[25], n160 );
nor U4400 ( n3370, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[14], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[13] );
nand U4401 ( n2852, n499, n2849 );
or U4402 ( n2850, n2849, n499 );
nand U4403 ( n3234, my_IIR_filter_firBlock_right_multProducts[36], n3233 );
xnor U4404 ( my_IIR_filter_firBlock_right_multProducts[6], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w189[13], n3369 );
nand U4405 ( n2980, n499, n2977 );
nand U4406 ( n2843, n499, n2842 );
or U4407 ( n2978, n2977, n499 );
or U4408 ( n3093, n3090, n160 );
nand U4409 ( n3091, n160, n3090 );
not U4410 ( n682, outData_in[13] );
nand U4411 ( n731, leftOut[10], n729 );
nand U4412 ( n723, leftOut[7], n807 );
nand U4413 ( n717, leftOut[4], n803 );
nand U4414 ( n715, leftOut[3], n801 );
or U4415 ( n3315, n3314, my_IIR_filter_firBlock_right_firStep[55] );
nor U4416 ( n796, leftOut[30], n797 );
nand U4417 ( n3311, n3310, my_IIR_filter_firBlock_right_multProducts[54] );
nor U4418 ( n3345, n3344, n3343 );
nand U4419 ( n775, n774, n773 );
nand U4420 ( n740, n738, n737 );
or U4421 ( n772, n771, leftOut[22] );
or U4422 ( n721, n806, leftOut[6] );
or U4423 ( n3332, n3331, my_IIR_filter_firBlock_right_firStep[59] );
nor U4424 ( n3344, n3341, n210 );
or U4425 ( n3338, n3337, my_IIR_filter_firBlock_right_firStep[60] );
or U4426 ( n3328, n3327, my_IIR_filter_firBlock_right_firStep[58] );
xnor U4427 ( n3173, my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[31], my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[37] );
xor U4428 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[21], n2977, n2976 );
xor U4429 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[27], n3002, n3001 );
xor U4430 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[30], n3016, n3015 );
xor U4431 ( my_IIR_filter_firBlock_right_my_IIR_filter_firBlock_right_MultiplyBlock_w192[38], n3053, n3052 );
endmodule

