module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule

module s38417_ori ( clk, reset, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214,
g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224,
g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234,
g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437,
g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657,
g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442,
g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837,
g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229,
g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956,
g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106,
g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263,
g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273,
g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420,
g25435, g25442, g25489, g26104, g26135, g26149, g27380 );
input clk, reset, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216,
g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226,
g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234;
output g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437,
g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657,
g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442,
g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837,
g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229,
g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956,
g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106,
g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263,
g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273,
g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420,
g25435, g25442, g25489, g26104, g26135, g26149, g27380;
wire g165, g305, g401, g309, g550, g499, g629, g630, g853, g992, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, ex_wire25, ex_wire26, ex_wire27, ex_wire28, ex_wire29, ex_wire30, ex_wire31, ex_wire32, ex_wire33, ex_wire34, ex_wire35, ex_wire36, ex_wire37, ex_wire38, ex_wire39, ex_wire40, ex_wire41, ex_wire42, ex_wire43, ex_wire44, ex_wire45, ex_wire46, ex_wire47, ex_wire48, ex_wire49, ex_wire50, ex_wire51, g1088,
g996, g1236, g1186, g1315, g1316, g1547, g1686, g1782, g1690, g1930,
g1880, g2009, g2010, g2241, g2380, g2476, g2384, g2624, g2574, g2703,
g2704, g2879, g2950, g2987, g3080, g150, g155, g157, g171, g176, g178,
g408, g455, g699, g726, g835, g840, g842, g856, g861, g863, g1526,
g1531, g1533, g1552, g1554, g2217, g2222, g2224, g2245, g3064, g3073,
g3204, g153, g158, g160, g174, g179, g411, g417, g427, g700, g702,
g727, g838, g843, g845, g859, g864, g866, g1095, g1142, g1385, g1412,
g1529, g1534, g1536, g1550, g1555, g1557, g2220, g2225, g2227, g2246,
g2248, g3074, g3207, g130, g156, g161, g163, g177, g414, g420, g428,
g698, g703, g705, g725, g841, g846, g848, g862, g867, g1098, g1104,
g1114, g1386, g1388, g1413, g1532, g1537, g1539, g1553, g1558, g1560,
g1789, g1836, g2079, g2106, g2223, g2228, g2230, g2244, g2249, g2251,
g3188, g131, g133, g159, g164, g354, g423, g426, g429, g701, g706,
g708, g818, g844, g849, g851, g865, g1101, g1107, g1115, g1384, g1389,
g1391, g1411, g1535, g1540, g1542, g1556, g1561, g1792, g1798, g1808,
g2080, g2082, g2107, g2226, g2231, g2233, g2247, g2252, g2254, g2483,
g2530, g2773, g2800, g181, g129, g134, g162, g101, g105, g343, g369,
g432, g438, g704, g709, g711, g729, g819, g821, g847, g852, g1041,
g1110, g1113, g1116, g1387, g1392, g1394, g1512, g1538, g1543, g1545,
g1559, g1795, g1801, g1809, g2078, g2083, g2085, g2105, g2229, g2234,
g2236, g2250, g2255, g2486, g2492, g2502, g2774, g2776, g2801, g132,
g346, g358, g384, g435, g441, g576, g587, g707, g712, g714, g730,
g732, g869, g817, g822, g850, g789, g793, g1030, g1056, g1119, g1125,
g1390, g1395, g1397, g1415, g1513, g1515, g1541, g1546, g1735, g1804,
g1807, g1810, g2081, g2086, g2088, g2206, g2232, g2237, g2239, g2253,
g2489, g2495, g2503, g2772, g2777, g2779, g2799, g361, g373, g398,
g444, g577, g579, g590, g596, g710, g715, g717, g728, g733, g735,
g820, g1033, g1045, g1071, g1122, g1128, g1262, g1273, g1393, g1398,
g1400, g1416, g1418, g1563, g1511, g1516, g1544, g1476, g1481, g1724,
g1750, g1813, g1819, g2084, g2089, g2091, g2109, g2207, g2209, g2235,
g2240, g2429, g2498, g2501, g2504, g2775, g2780, g2782, g121, g125,
g376, g388, g575, g580, g582, g593, g599, g713, g718, g720, g731,
g736, g1048, g1060, g1085, g1131, g1263, g1265, g1276, g1282, g1396,
g1401, g1403, g1414, g1419, g1421, g1514, g1727, g1739, g1765, g1816,
g1822, g1956, g1967, g2087, g2092, g2094, g2110, g2112, g2257, g2205,
g2210, g2238, g2170, g2175, g2418, g2444, g2507, g2513, g2778, g2783,
g2785, g2803, g391, g448, g578, g583, g585, g602, g605, g716, g721,
g723, g734, g809, g813, g1063, g1075, g1261, g1266, g1268, g1279,
g1285, g1399, g1404, g1406, g1417, g1422, g1742, g1754, g1779, g1825,
g1957, g1959, g1970, g1976, g2090, g2095, g2097, g2108, g2113, g2115,
g2208, g2421, g2433, g2459, g2510, g2516, g2650, g2661, g2781, g2786,
g2788, g2804, g2806, g449, g581, g586, g608, g614, g719, g724, g1078,
g1135, g1264, g1269, g1271, g1288, g1291, g1402, g1407, g1409, g1420,
g1501, g1506, g1757, g1769, g1955, g1960, g1962, g1973, g1979, g2093,
g2098, g2100, g2111, g2116, g2436, g2448, g2473, g2519, g2651, g2653,
g2664, g2670, g2784, g2789, g2791, g2802, g2807, g2809, g109, g447,
g584, g611, g617, g722, g1136, g1267, g1272, g1294, g1300, g1405,
g1410, g1772, g1829, g1958, g1963, g1965, g1982, g1985, g2096, g2101,
g2103, g2114, g2195, g2200, g2451, g2463, g2649, g2654, g2656, g2667,
g2673, g2787, g2792, g2794, g2805, g2810, g620, g797, g1134, g1270,
g1297, g1303, g1408, g1830, g1961, g1966, g1988, g1994, g2099, g2104,
g2466, g2523, g2652, g2657, g2659, g2676, g2679, g2790, g2795, g2797,
g2808, g2857, g738, g1306, g1486, g1828, g1964, g1991, g1997, g2102,
g2524, g2655, g2660, g2682, g2688, g2793, g2798, g2873, g739, g1424,
g2000, g2180, g2522, g2658, g2685, g2691, g2796, g3106, g2877, g737,
g1425, g2118, g2694, g3107, g2878, g1423, g2119, g2812, g2933, g3108,
g2117, g2813, g2811, g3054, g3079, g3210, g3211, g3084, g3085, g3086,
g3155, g3087, g3164, g3091, g3158, g3173, g3092, g3167, g3182, g79,
g3093, g3161, g3176, g70, g767, g3170, g3185, g61, g213, g758, g1453,
g3179, g65, g216, g222, g299, g749, g900, g1444, g2147, g3088, g56,
g219, g225, g231, g113, g507, g541, g753, g903, g909, g986, g1192,
g1435, g1594, g2138, g92, g52, g228, g234, g240, g744, g906, g912,
g918, g801, g1227, g1439, g1597, g1603, g1680, g1886, g2129, g2288,
g83, g117, g237, g243, g249, g780, g740, g915, g921, g927, g1430,
g1600, g1606, g1612, g1491, g1921, g2133, g2291, g2297, g74, g246,
g252, g258, g97, g538, g771, g805, g924, g930, g936, g1466, g1426,
g1609, g1615, g1621, g2124, g2294, g2300, g2306, g2185, g2581, g2615,
g88, g186, g255, g261, g267, g762, g933, g939, g945, g785, g1224,
g1457, g1496, g1618, g1624, g1630, g2160, g2120, g2303, g2309, g2315,
g189, g195, g264, g270, g776, g873, g942, g948, g954, g1448, g1627,
g1633, g1639, g1471, g1918, g2151, g2190, g2312, g2318, g2324, g192,
g198, g204, g273, g876, g882, g951, g957, g1462, g1567, g1636, g1642,
g1648, g2142, g2321, g2327, g2333, g2165, g2612, g201, g207, g879,
g885, g891, g960, g1570, g1576, g1645, g1651, g2156, g2261, g2330,
g2336, g2342, g210, g888, g894, g1573, g1579, g1585, g1654, g2264,
g2270, g2339, g2345, g471, g897, g1582, g1588, g2267, g2273, g2279,
g2348, g1158, g1591, g2276, g2282, g1852, g2285, g3142, g2546, g458,
g461, g1145, g465, g1148, g1839, g468, g1152, g1842, g2533, g1155,
g1846, g2536, g1849, g2540, g2543, g672, g524, g554, g679, g1358,
g3097, g3147, g686, g1210, g1240, g1365, g2052, g3098, g557, g633,
g692, g1372, g1904, g1934, g2059, g2746, g3099, g542, g646, g1243,
g1319, g1378, g2066, g2598, g2628, g2753, g3100, g510, g640, g1228,
g1332, g1937, g2013, g2072, g2760, g3101, g653, g1196, g1326, g1922,
g2026, g2631, g2707, g2766, g3102, g544, g660, g1339, g1890, g2020,
g2616, g2720, g3103, g464, g559, g666, g1230, g1346, g2033, g2584,
g2714, g2993, g3006, g3104, g484, g1151, g1245, g1352, g1924, g2040,
g2727, g2998, g3013, g3105, g3136, g480, g1171, g1845, g1939, g2046,
g2618, g2734, g3002, g3139, g490, g1167, g1865, g2539, g2633, g2740,
g2912, g3010, g3036, g493, g1177, g1861, g2559, g2917, g3018, g496,
g1180, g1871, g2555, g2883, g2920, g2990, g3028, g3114, g1183, g1874,
g2565, g2888, g2896, g3032, g3120, g3128, g1877, g2568, g2892, g2903,
g2571, g2900, g2908, g3133, g2924, g312, g3123, g313, g999, g314,
g315, g403, g1000, g1693, g3094, g3125, g316, g318, g404, g1001,
g1002, g1090, g1694, g2387, g3095, g317, g319, g402, g1003, g1005,
g1091, g1695, g1696, g1784, g2388, g3096, g320, g1004, g1006, g1089,
g1697, g1699, g1785, g2389, g2390, g2478, g1007, g1698, g1700, g1783,
g2391, g2393, g2479, g322, g1701, g2392, g2394, g2477, g323, g659,
g1009, g2395, g321, g1010, g1345, g1703, g1008, g1704, g2039, g2397,
g1702, g2398, g2733, g479, g2396, g478, g1166, g2953, g3044, g477,
g1165, g1860, g2956, g2981, g3045, g3055, g1164, g1859, g2554, g2959,
g2874, g3046, g3056, g3065, g3201, g1858, g2553, g3047, g3057, g3066,
g3075, g3151, g488, g2552, g2935, g2963, g3048, g3058, g3067, g3076,
g142, g487, g1175, g2938, g2966, g3049, g3059, g3068, g3077, g3109,
g3191, g143, g145, g486, g485, g830, g1174, g1869, g2941, g2969,
g3050, g3060, g3069, g3078, g3083, g3194, g141, g146, g148, g169,
g831, g833, g1173, g1172, g1524, g1868, g2563, g2944, g2972, g3051,
g3061, g3070, g2997, g185, g3197, g144, g149, g151, g170, g172, g829,
g834, g836, g857, g1525, g1527, g1867, g1866, g2218, g2562, g2947,
g2975, g3043, g3052, g3062, g3071, g3198, g147, g152, g154, g168,
g173, g175, g832, g837, g839, g858, g860, g1523, g1528, g1530, g1551,
g2219, g2221, g2561, g2560, g2978, g3053, g3063, g3072, new_g13149_,
new_g13111_, new_g13155_, new_g13160_, new_g13124_, new_g13164_,
new_g12487_, new_g13171_, new_g13135_, new_g13175_, new_g12507_,
new_g13182_, new_g13143_, new_g12524_, new_g13194_, new_g12457_,
new_g12539_, new_g12467_, new_g12482_, new_g12499_, new_g13110_,
new_g12433_, new_g16132_, new_g16181_, new_g18669_, new_g18678_,
new_g18707_, new_g18719_, new_g18726_, new_g18743_, new_g18755_,
new_g18763_, new_g18780_, new_g18782_, new_g18794_, new_g18821_,
new_g18804_, new_g18820_, new_g18835_, new_g18852_, new_g18836_,
new_g18975_, new_g18837_, new_g18866_, new_g18968_, new_g18883_,
new_g18867_, new_g18868_, new_g18885_, new_g18754_, new_g18906_,
new_g18907_, new_g18781_, new_g18542_, new_g18803_, new_g18942_,
new_g18957_, new_g16654_, new_g16671_, new_g16692_, new_g16718_,
new_g16860_, new_g16866_, new_g16803_, new_g16566_, new_g16824_,
new_g16835_, new_g16844_, new_g16845_, new_g16851_, new_g16853_,
new_g16854_, new_g16857_, new_g16861_, new_g16880_, new_g16802_,
new_g16823_, new_g17222_, new_g17224_, new_g17225_, new_g17226_,
new_g17228_, new_g17229_, new_g17234_, new_g17235_, new_g17236_,
new_g17246_, new_g17247_, new_g17248_, new_g17269_, new_g17270_,
new_g17271_, new_g17302_, new_g17303_, new_g17340_, new_g17341_,
new_g17383_, new_g17429_, new_g20310_, new_g20314_, new_g20333_,
new_g20343_, new_g20353_, new_g20375_, new_g20376_, new_g20417_,
new_g19144_, new_g19149_, new_g19153_, new_g19154_, new_g19157_,
new_g19162_, new_g19163_, new_g19167_, new_g19172_, new_g19173_,
new_g19178_, new_g19184_, new_g19152_, new_g20497_, new_g21842_,
new_g21843_, new_g21845_, new_g21847_, new_g21851_, new_g21878_,
new_g21880_, new_g21882_, new_g20874_, new_g20875_, new_g20876_,
new_g20879_, new_g20880_, new_g20881_, new_g20882_, new_g20883_,
new_g20682_, new_g20891_, new_g20892_, new_g20893_, new_g20894_,
new_g20896_, new_g20897_, new_g20898_, new_g20899_, new_g20900_,
new_g20901_, new_g20902_, new_g20903_, new_g20717_, new_g20910_,
new_g20911_, new_g20912_, new_g20913_, new_g20915_, new_g20916_,
new_g20917_, new_g20918_, new_g20919_, new_g20921_, new_g20922_,
new_g20923_, new_g20924_, new_g20925_, new_g20926_, new_g20927_,
new_g20752_, new_g20934_, new_g20935_, new_g20936_, new_g20937_,
new_g20939_, new_g20940_, new_g20941_, new_g20944_, new_g20945_,
new_g20946_, new_g20947_, new_g20948_, new_g20949_, new_g20950_,
new_g20951_, new_g20952_, new_g20953_, new_g20954_, new_g20955_,
new_g20789_, new_g20962_, new_g20963_, new_g20964_, new_g20965_,
new_g20966_, new_g20967_, new_g20968_, new_g20969_, new_g20970_,
new_g20972_, new_g20973_, new_g20974_, new_g20975_, new_g20976_,
new_g20977_, new_g20978_, new_g20979_, new_g20980_, new_g20981_,
new_g20982_, new_g20983_, new_g20989_, new_g20990_, new_g20991_,
new_g20992_, new_g20993_, new_g20994_, new_g20995_, new_g20996_,
new_g20997_, new_g20999_, new_g21000_, new_g21001_, new_g21002_,
new_g21003_, new_g21004_, new_g21005_, new_g21006_, new_g21007_,
new_g21009_, new_g21010_, new_g21011_, new_g21015_, new_g21016_,
new_g21017_, new_g21018_, new_g21019_, new_g21020_, new_g21021_,
new_g21022_, new_g21023_, new_g21025_, new_g21026_, new_g21027_,
new_g21028_, new_g21029_, new_g21031_, new_g21032_, new_g21033_,
new_g21034_, new_g21035_, new_g21039_, new_g21040_, new_g21041_,
new_g21042_, new_g21043_, new_g21044_, new_g21045_, new_g21046_,
new_g21047_, new_g21051_, new_g21052_, new_g21053_, new_g21054_,
new_g21055_, new_g21056_, new_g21060_, new_g21061_, new_g21062_,
new_g21063_, new_g20825_, new_g21070_, new_g21071_, new_g21072_,
new_g21073_, new_g21074_, new_g21075_, new_g21080_, new_g21081_,
new_g21082_, new_g21094_, new_g20877_, new_g20884_, new_g21346_,
new_g23000_, new_g23117_, new_g23014_, new_g23126_, new_g23022_,
new_g23030_, new_g23137_, new_g23039_, new_g23047_, new_g21970_,
new_g23058_, new_g23067_, new_g23076_, new_g23081_, new_g23092_,
new_g23093_, new_g23097_, new_g23110_, new_g23111_, new_g23114_,
new_g23123_, new_g23124_, new_g23132_, new_g23133_, new_g22025_,
new_g22027_, new_g22028_, new_g22029_, new_g22030_, new_g22031_,
new_g22032_, new_g22033_, new_g22034_, new_g22035_, new_g22037_,
new_g22038_, new_g22039_, new_g22040_, new_g22041_, new_g22042_,
new_g22043_, new_g22044_, new_g22045_, new_g22047_, new_g22048_,
new_g22049_, new_g23136_, new_g22054_, new_g22055_, new_g22056_,
new_g22057_, new_g22058_, new_g22059_, new_g22060_, new_g22061_,
new_g22063_, new_g22064_, new_g22065_, new_g22066_, new_g22067_,
new_g22068_, new_g21969_, new_g22073_, new_g22074_, new_g22075_,
new_g22076_, new_g22077_, new_g22078_, new_g22079_, new_g22080_,
new_g22081_, new_g22087_, new_g22088_, new_g22089_, new_g22090_,
new_g22091_, new_g22092_, new_g21972_, new_g22097_, new_g22098_,
new_g22099_, new_g22100_, new_g22101_, new_g22102_, new_g22103_,
new_g22104_, new_g22105_, new_g22106_, new_g22112_, new_g22113_,
new_g22114_, new_g22115_, new_g22116_, new_g22117_, new_g21974_,
new_g22122_, new_g22123_, new_g22124_, new_g22125_, new_g22126_,
new_g22127_, new_g22128_, new_g22129_, new_g22130_, new_g22131_,
new_g22132_, new_g22138_, new_g22139_, new_g22140_, new_g22141_,
new_g22142_, new_g22143_, new_g22145_, new_g22146_, new_g22147_,
new_g22148_, new_g22149_, new_g22150_, new_g22151_, new_g22152_,
new_g22153_, new_g22154_, new_g22155_, new_g22161_, new_g22162_,
new_g22163_, new_g22164_, new_g22166_, new_g22167_, new_g22168_,
new_g22169_, new_g22170_, new_g22171_, new_g22172_, new_g22173_,
new_g22177_, new_g22178_, new_g22179_, new_g22180_, new_g22182_,
new_g22183_, new_g22184_, new_g22185_, new_g22191_, new_g22192_,
new_g22193_, new_g22194_, new_g22200_, new_g21989_, new_g22578_,
new_g22002_, new_g22615_, new_g22651_, new_g22026_, new_g22218_,
new_g22687_, new_g22231_, new_g22234_, new_g22242_, new_g22247_,
new_g22249_, new_g22263_, new_g22267_, new_g22269_, new_g22280_,
new_g22284_, new_g22299_, new_g23399_, new_g23406_, new_g24174_,
new_g23413_, new_g24178_, new_g24179_, new_g23418_, new_g24181_,
new_g24182_, new_g24206_, new_g24207_, new_g24208_, new_g24209_,
new_g24212_, new_g24213_, new_g24214_, new_g24215_, new_g24216_,
new_g24218_, new_g24219_, new_g24222_, new_g24223_, new_g24225_,
new_g24226_, new_g24228_, new_g24230_, new_g24231_, new_g24235_,
new_g24237_, new_g24238_, new_g24243_, new_g24250_, new_g23385_,
new_g23392_, new_g23400_, new_g23324_, new_g23407_, new_g23329_,
new_g23330_, new_g23339_, new_g23348_, new_g23357_, new_g23358_,
new_g23359_, new_g24059_, new_g24072_, new_g24083_, new_g24092_,
new_g25027_, new_g25042_, new_g25056_, new_g25067_, new_g24426_,
new_g24430_, new_g24434_, new_g24438_, new_g24491_, new_g24498_,
new_g24499_, new_g24501_, new_g24507_, new_g24508_, new_g24510_,
new_g24511_, new_g24513_, new_g24445_, new_g24446_, new_g24519_,
new_g24521_, new_g24522_, new_g24524_, new_g24525_, new_g24527_,
new_g24532_, new_g24534_, new_g24535_, new_g24537_, new_g24538_,
new_g24545_, new_g24547_, new_g24548_, new_g24557_, new_g24473_,
new_g24476_, new_g25932_, new_g25935_, new_g25938_, new_g25940_,
new_g25204_, new_g25206_, new_g25207_, new_g25209_, new_g25211_,
new_g25212_, new_g25213_, new_g25214_, new_g25215_, new_g25217_,
new_g25218_, new_g25219_, new_g25220_, new_g25221_, new_g25222_,
new_g25223_, new_g25224_, new_g25225_, new_g25227_, new_g25228_,
new_g25229_, new_g25230_, new_g25231_, new_g25232_, new_g25233_,
new_g25234_, new_g25235_, new_g25236_, new_g25237_, new_g25239_,
new_g25240_, new_g25241_, new_g25242_, new_g25243_, new_g25244_,
new_g25245_, new_g25246_, new_g25247_, new_g25248_, new_g25249_,
new_g25250_, new_g25251_, new_g25252_, new_g25253_, new_g25185_,
new_g25255_, new_g25256_, new_g25257_, new_g25189_, new_g25259_,
new_g25265_, new_g25191_, new_g25260_, new_g25194_, new_g25262_,
new_g25263_, new_g25197_, new_g25266_, new_g25267_, new_g25268_,
new_g25270_, new_g25271_, new_g25272_, new_g25279_, new_g25280_,
new_g25199_, new_g25288_, new_g25201_, new_g25202_, new_g25450_,
new_g25451_, new_g25452_, new_g26541_, new_g26545_, new_g26547_,
new_g26553_, new_g26557_, new_g26559_, new_g26569_, new_g26573_,
new_g26575_, new_g26592_, new_g26596_, new_g26616_, new_g26529_,
new_g26530_, new_g26655_, new_g26531_, new_g26659_, new_g26661_,
new_g26532_, new_g26664_, new_g26665_, new_g26667_, new_g26669_,
new_g26670_, new_g26672_, new_g26675_, new_g26676_, new_g26025_,
new_g26660_, new_g26666_, new_g26671_, new_g26677_, new_g26048_,
new_g26031_, new_g26037_, new_g26106_, new_g26120_, new_g26130_,
new_g26144_, new_g27120_, new_g27123_, new_g27129_, new_g27131_,
new_g26803_, new_g26804_, new_g26805_, new_g26806_, new_g26807_,
new_g26808_, new_g26776_, new_g26809_, new_g26810_, new_g26811_,
new_g26812_, new_g26813_, new_g26814_, new_g26781_, new_g26815_,
new_g26816_, new_g26817_, new_g26786_, new_g26818_, new_g26820_,
new_g26821_, new_g26789_, new_g26822_, new_g26823_, new_g26824_,
new_g26825_, new_g26826_, new_g26795_, new_g26827_, new_g26798_,
new_g27594_, new_g27603_, new_g27612_, new_g27621_, new_g27672_,
new_g27678_, new_g27682_, new_g27243_, new_g27253_, new_g27255_,
new_g27256_, new_g27257_, new_g27258_, new_g27259_, new_g27260_,
new_g27261_, new_g27262_, new_g27263_, new_g27264_, new_g27265_,
new_g27266_, new_g27267_, new_g27268_, new_g27269_, new_g27270_,
new_g27271_, new_g27272_, new_g27273_, new_g27274_, new_g27275_,
new_g27276_, new_g27277_, new_g27278_, new_g27279_, new_g27280_,
new_g27281_, new_g27282_, new_g27283_, new_g27284_, new_g27285_,
new_g27286_, new_g27287_, new_g27288_, new_g27289_, new_g27290_,
new_g27291_, new_g27292_, new_g27293_, new_g27294_, new_g27295_,
new_g27296_, new_g27297_, new_g27298_, new_g27299_, new_g27300_,
new_g27301_, new_g27302_, new_g27303_, new_g27304_, new_g27305_,
new_g27306_, new_g27307_, new_g27308_, new_g27309_, new_g27310_,
new_g27311_, new_g27312_, new_g27313_, new_g27314_, new_g27315_,
new_g27316_, new_g27317_, new_g27318_, new_g27319_, new_g27320_,
new_g27321_, new_g27322_, new_g27323_, new_g27324_, new_g27325_,
new_g27326_, new_g27327_, new_g27328_, new_g27329_, new_g27330_,
new_g27331_, new_g27332_, new_g27333_, new_g27334_, new_g27335_,
new_g27336_, new_g27337_, new_g27338_, new_g27339_, new_g27340_,
new_g27341_, new_g27342_, new_g27343_, new_g27344_, new_g27345_,
new_g27346_, new_g27347_, new_g27348_, new_g27354_, new_g28145_,
new_g28146_, new_g28147_, new_g28148_, new_g28199_, new_g27718_,
new_g27722_, new_g27724_, new_g27759_, new_g27760_, new_g27761_,
new_g27762_, new_g27763_, new_g27764_, new_g27765_, new_g27766_,
new_g27767_, new_g27768_, new_g27769_, new_g27771_, new_g28634_,
new_g28635_, new_g28636_, new_g28637_, new_g28668_, new_g28321_,
new_g28325_, new_g28328_, new_g28342_, new_g28344_, new_g28345_,
new_g28346_, new_g28348_, new_g28349_, new_g28350_, new_g28351_,
new_g28352_, new_g28353_, new_g28354_, new_g28355_, new_g28356_,
new_g28357_, new_g28358_, new_g28360_, new_g28361_, new_g28362_,
new_g28363_, new_g28364_, new_g28366_, new_g28367_, new_g28368_,
new_g28371_, new_g28420_, new_g28421_, new_g28425_, new_g29109_,
new_g29110_, new_g29111_, new_g29112_, new_g28732_, new_g28735_,
new_g28736_, new_g28738_, new_g28744_, new_g28745_, new_g28746_,
new_g28747_, new_g28749_, new_g28754_, new_g28758_, new_g28759_,
new_g28760_, new_g28761_, new_g28990_, new_g28763_, new_g28767_,
new_g28771_, new_g28772_, new_g28773_, new_g28774_, new_g28778_,
new_g28782_, new_g28783_, new_g28788_, new_g28903_, new_g29353_,
new_g29354_, new_g29355_, new_g29357_, new_g29167_, new_g29169_,
new_g29170_, new_g29172_, new_g29173_, new_g29178_, new_g29179_,
new_g29181_, new_g29182_, new_g29184_, new_g29185_, new_g29187_,
new_g29194_, new_g29197_, new_g29198_, new_g29201_, new_g29204_,
new_g29205_, new_g29209_, new_g29212_, new_g29213_, new_g29218_,
new_g29221_, new_g29226_, new_g29579_, new_g29606_, new_g29608_,
new_g29580_, new_g29609_, new_g29611_, new_g29612_, new_g29581_,
new_g29613_, new_g29616_, new_g29617_, new_g29582_, new_g29618_,
new_g29620_, new_g29621_, new_g29623_, new_g29936_, new_g29939_,
new_g29941_, new_g30055_, new_g30061_, new_g30267_, new_g30268_,
new_g30269_, new_g30270_, new_g30271_, new_g30272_, new_g30273_,
new_g30274_, new_g30275_, new_g30276_, new_g30277_, new_g30278_,
new_g30279_, new_g30280_, new_g30281_, new_g30282_, new_g30283_,
new_g30284_, new_g30285_, new_g30286_, new_g30287_, new_g30288_,
new_g30289_, new_g30290_, new_g30291_, new_g30292_, new_g30293_,
new_g30294_, new_g30295_, new_g30296_, new_g30297_, new_g30298_,
new_g30299_, new_g30300_, new_g30301_, new_g30302_, new_g30303_,
new_g30304_, new_g30245_, new_g30246_, new_g30247_, new_g30248_,
new_g30249_, new_g30250_, new_g30251_, new_g30252_, new_g30253_,
new_g30254_, new_g30255_, new_g30256_, new_g30257_, new_g30258_,
new_g30259_, new_g30260_, new_g30261_, new_g30262_, new_g30263_,
new_g30264_, new_g30265_, new_g30266_, new_g30455_, new_g30468_,
new_g30470_, new_g30482_, new_g30485_, new_g30487_, new_g30500_,
new_g30503_, new_g30505_, new_g30338_, new_g30341_, new_g30356_,
new_g30668_, new_g30669_, new_g30670_, new_g30671_, new_g30672_,
new_g30673_, new_g30674_, new_g30675_, new_g30676_, new_g30677_,
new_g30678_, new_g30679_, new_g30680_, new_g30681_, new_g30682_,
new_g30683_, new_g30684_, new_g30686_, new_g30687_, new_g30688_,
new_g30689_, new_g30690_, new_g30691_, new_g30692_, new_g30693_,
new_g30694_, new_g30695_, new_g30699_, new_g30700_, new_g30701_,
new_g30702_, new_g30703_, new_g30704_, new_g30705_, new_g30706_,
new_g30707_, new_g30708_, new_g30709_, new_g30566_, new_g30635_,
new_g30636_, new_g30637_, new_g30638_, new_g30639_, new_g30640_,
new_g30641_, new_g30642_, new_g30643_, new_g30644_, new_g30645_,
new_g30646_, new_g30647_, new_g30648_, new_g30649_, new_g30650_,
new_g30651_, new_g30652_, new_g30653_, new_g30654_, new_g30655_,
new_g30656_, new_g30657_, new_g30658_, new_g30659_, new_g30660_,
new_g30661_, new_g30662_, new_g30663_, new_g30664_, new_g30665_,
new_g30666_, new_g30667_, new_g30796_, new_g30798_, new_g30801_, g349,
g351, g364, g1036, g337, g353, g366, g379, g1038, g1051, g1730, g368,
g381, g394, g1024, g1040, g1053, g1066, g1732, g1745, g2424, g383,
g396, g1055, g1068, g1081, g1718, g1734, g1747, g1760, g2426, g2439,
g324, g1070, g1083, g1749, g1762, g1775, g2412, g2428, g2441, g2454,
g1011, g1764, g1777, g2443, g2456, g2469, g1705, g2458, g2471, g2399,
g565, g567, g1251, g489, g1253, g1945, g1176, g1947, g2639, g1870,
g2641, g2564, g569, g571, g1255, g573, g1257, g1949, g1259, g1951,
g2643, g1953, g2645, g2647, g298, g985, g1679, g2373, g548, g1234,
g1928, g2622, g3124, g3111, g3110, g3126, g3112, g3113, g3135, g3127,
g3134, g3132, g2962, g2934, g2984, g2985, g537, g529, g530, g531,
g532, g533, g534, g536, g1223, g1215, g1216, g1217, g1218, g1219,
g1220, g1222, g1917, g1909, g1910, g1911, g1912, g1913, g1914, g1916,
g2611, g2603, g2604, g2605, g2606, g2607, g2608, g2610, n1058, n1062,
n1481, n1737, n1746, n1755, n1764, n1773, n1782, n1791, n1800, n1809,
n1883, n1892, n1901, n1910, n1919, n1928, n1937, n1946, n1955, n1964,
n1973, n1982, n2032, n2036, n2045, n2054, n2063, n2072, n2081, n2090,
n2187, n2191, n2200, n2214, n2223, n2759, n2763, n3182, n3438, n3447,
n3456, n3465, n3474, n3483, n3492, n3501, n3510, n3584, n3593, n3602,
n3611, n3620, n3629, n3638, n3647, n3656, n3665, n3674, n3683, n3733,
n3737, n3746, n3755, n3764, n3773, n3782, n3791, n3888, n3892, n3901,
n3915, n3924, n4460, n4464, n4883, n5139, n5148, n5157, n5166, n5175,
n5184, n5193, n5202, n5211, n5285, n5294, n5303, n5312, n5321, n5330,
n5339, n5348, n5357, n5366, n5375, n5384, n5434, n5438, n5447, n5456,
n5465, n5474, n5483, n5492, n5589, n5593, n5602, n5616, n5625, n6161,
n6165, n6584, n6840, n6849, n6858, n6867, n6876, n6885, n6894, n6903,
n6912, n6986, n6995, n7004, n7013, n7022, n7031, n7040, n7049, n7058,
n7067, n7076, n7085, n7135, n7139, n7148, n7157, n7166, n7175, n7184,
n7193, n7290, n7294, n7303, n7317, n7326, n1, n2, n5, n7, n10, n11,
n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n23, n24, n25, n26,
n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
n41, n42, n43, n48, n49, n52, n53, n54, n55, n56, n57, n58, n59, n60,
n62, n63, n65, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84, n85,
n87, n96, n97, n98, n99, n100, n101, n102, n103, n104, n106, n107,
n109, n118, n119, n120, n121, n122, n123, n124, n125, n126, n128,
n129, n131, n143, n145, n146, n147, n148, n149, n151, n155, n158,
n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
n171, n172, n173, n176, n178, n179, n180, n184, n185, n186, n187,
n188, n189, n190, n191, n192, n193, n195, n196, n197, n198, n199,
n200, n201, n202, n203, n204, n205, n216, n217, n218, n219, n220,
n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
n246, n247, n255, n256, n257, n259, n260, n261, n262, n263, n264,
n265, n267, n269, n281, n282, n283, n284, n285, n286, n287, n288,
n289, n290, n291, n292, n293, n294, n297, n299, n300, n301, n305,
n306, n307, n308, n309, n310, n311, n312, n313, n314, n316, n317,
n318, n319, n320, n321, n322, n323, n324, n325, n337, n338, n339,
n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
n354, n355, n364, n365, n366, n368, n369, n370, n371, n372, n373,
n374, n376, n378, n390, n391, n392, n393, n394, n395, n396, n397,
n398, n399, n400, n401, n402, n403, n406, n408, n409, n410, n414,
n415, n416, n417, n418, n419, n420, n421, n422, n423, n425, n426,
n427, n428, n429, n430, n431, n432, n433, n434, n446, n447, n448,
n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
n463, n464, n472, n473, n474, n476, n477, n478, n479, n480, n481,
n482, n484, n486, n498, n499, n500, n501, n502, n503, n504, n505,
n506, n507, n509, n510, n511, n512, n515, n518, n519, n520, n524,
n525, n527, n528, n529, n530, n531, n532, n533, n534, n537, n538,
n539, n540, n541, n542, n543, n545, n546, n547, n560, n561, n563,
n564, n565, n566, n567, n568, n569, n570, n572, n573, n574, n575,
n579, n581, n590, n591, n592, n594, n595, n596, n597, n599, n600,
n601, n603, n605, n619, n620, n621, n622, n624, n628, n637, n638,
n639, n640, n641, n642, n644, n645, n646, n647, n648, n649, n650,
n651, n653, n654, n655, n656, n657, n658, n659, n660, n662, n663,
n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
n708, n709, n710, n711, n712, n713, n714, n716, n717, n718, n720,
n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1059, n1060, n1061, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
n1478, n1479, n1480, n1482, n1483, n1484, n1486, n1487, n1488, n1489,
n1490, n1491, n1492, n1493, n1495, n1496, n1497, n1499, n1500, n1501,
n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
n1732, n1733, n1734, n1735, n1736, n1738, n1739, n1740, n1741, n1742,
n1743, n1744, n1745, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
n1754, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1765,
n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1774, n1775, n1778,
n1779, n1780, n1781, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
n1790, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1801,
n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1810, n1811, n1812,
n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1884, n1885,
n1886, n1887, n1888, n1889, n1890, n1891, n1893, n1894, n1895, n1896,
n1897, n1898, n1899, n1900, n1902, n1903, n1904, n1905, n1906, n1907,
n1908, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1920, n1921,
n1922, n1923, n1924, n1925, n1926, n1927, n1929, n1930, n1931, n1932,
n1933, n1934, n1935, n1936, n1938, n1939, n1940, n1941, n1942, n1943,
n1944, n1945, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1965, n1966,
n1967, n1968, n1969, n1970, n1971, n1972, n1974, n1977, n1978, n1979,
n1980, n1981, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
n1992, n1993, n1994, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
n2003, n2005, n2006, n2007, n2009, n2010, n2011, n2012, n2013, n2014,
n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2033, n2034, n2035,
n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2046, n2047,
n2048, n2049, n2050, n2051, n2052, n2053, n2055, n2056, n2057, n2058,
n2059, n2060, n2061, n2062, n2064, n2065, n2066, n2067, n2068, n2069,
n2070, n2071, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2091, n2092,
n2093, n2094, n2095, n2096, n2097, n2098, n2100, n2101, n2102, n2104,
n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
n2185, n2186, n2188, n2189, n2190, n2192, n2193, n2194, n2195, n2196,
n2197, n2198, n2199, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
n2208, n2209, n2210, n2211, n2212, n2213, n2215, n2216, n2217, n2218,
n2219, n2220, n2221, n2222, n2224, n2225, n2226, n2227, n2228, n2229,
n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2418, n2419, n2420,
n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
n2471, n2472, n2473, n2474, n2475, n2477, n2478, n2479, n2481, n2482,
n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2743,
n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
n2754, n2755, n2756, n2757, n2758, n2760, n2761, n2762, n2764, n2766,
n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2787,
n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
n2798, n2799, n2800, n2801, n2803, n2804, n2805, n2806, n2807, n2808,
n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
n3179, n3180, n3181, n3183, n3184, n3185, n3187, n3188, n3189, n3190,
n3191, n3192, n3193, n3194, n3196, n3197, n3198, n3200, n3201, n3202,
n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
n3433, n3434, n3435, n3436, n3437, n3439, n3440, n3441, n3442, n3443,
n3444, n3445, n3446, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
n3455, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3466,
n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3475, n3476, n3477,
n3478, n3479, n3480, n3481, n3482, n3484, n3485, n3486, n3487, n3488,
n3489, n3490, n3491, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
n3500, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3511,
n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3594, n3597,
n3598, n3599, n3600, n3601, n3603, n3604, n3605, n3606, n3607, n3608,
n3609, n3610, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3630, n3631,
n3632, n3633, n3634, n3635, n3636, n3637, n3639, n3640, n3641, n3642,
n3643, n3644, n3645, n3646, n3648, n3649, n3650, n3651, n3652, n3653,
n3654, n3655, n3657, n3658, n3659, n3660, n3661, n3662, n3666, n3667,
n3668, n3669, n3670, n3671, n3672, n3673, n3675, n3676, n3677, n3678,
n3679, n3680, n3681, n3682, n3684, n3685, n3686, n3687, n3688, n3689,
n3690, n3691, n3693, n3694, n3695, n3697, n3698, n3701, n3702, n3703,
n3704, n3706, n3707, n3708, n3710, n3711, n3712, n3713, n3714, n3715,
n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3734, n3735, n3736,
n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3747, n3748,
n3749, n3750, n3751, n3752, n3753, n3754, n3756, n3757, n3758, n3759,
n3760, n3761, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3783, n3784,
n3785, n3786, n3787, n3788, n3789, n3790, n3792, n3793, n3794, n3795,
n3796, n3799, n3801, n3802, n3803, n3805, n3806, n3807, n3808, n3809,
n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
n3880, n3881, n3882, n3885, n3886, n3887, n3889, n3890, n3891, n3893,
n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3902, n3903, n3904,
n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3925, n3926,
n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
n4117, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4178,
n4179, n4180, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
n4190, n4191, n4192, n4193, n4194, n4195, n4198, n4199, n4200, n4201,
n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
n4222, n4223, n4224, n4225, n4226, n4229, n4230, n4231, n4232, n4233,
n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
n4324, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
n4458, n4459, n4461, n4462, n4463, n4465, n4466, n4467, n4468, n4469,
n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
n4880, n4881, n4882, n4884, n4885, n4886, n4888, n4889, n4890, n4891,
n4892, n4893, n4894, n4895, n4897, n4898, n4899, n4901, n4902, n4903,
n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
n5134, n5135, n5136, n5137, n5138, n5140, n5141, n5142, n5143, n5144,
n5145, n5146, n5147, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
n5156, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5167,
n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5176, n5177, n5178,
n5179, n5180, n5181, n5182, n5183, n5185, n5186, n5187, n5188, n5189,
n5190, n5191, n5192, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
n5201, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5212,
n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
n5283, n5284, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5304, n5305,
n5306, n5307, n5308, n5309, n5310, n5311, n5313, n5314, n5315, n5316,
n5317, n5318, n5319, n5320, n5322, n5323, n5324, n5325, n5326, n5327,
n5328, n5329, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5349, n5350,
n5351, n5352, n5353, n5354, n5355, n5356, n5358, n5359, n5360, n5361,
n5362, n5363, n5364, n5365, n5367, n5368, n5369, n5370, n5371, n5372,
n5373, n5374, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5394, n5395,
n5396, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5407,
n5408, n5409, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
n5429, n5430, n5431, n5432, n5433, n5435, n5436, n5437, n5439, n5440,
n5441, n5442, n5443, n5444, n5445, n5446, n5448, n5449, n5450, n5451,
n5452, n5453, n5454, n5455, n5457, n5458, n5459, n5460, n5461, n5462,
n5463, n5464, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5484, n5485,
n5486, n5487, n5488, n5489, n5490, n5491, n5493, n5494, n5495, n5496,
n5497, n5498, n5499, n5500, n5502, n5503, n5504, n5506, n5507, n5508,
n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
n5590, n5591, n5592, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
n5601, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
n5612, n5613, n5614, n5615, n5617, n5618, n5619, n5620, n5621, n5622,
n5623, n5624, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
n5814, n5815, n5816, n5817, n5818, n5820, n5821, n5822, n5823, n5824,
n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
n5875, n5876, n5877, n5879, n5880, n5881, n5883, n5884, n5885, n5886,
n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
n6137, n6138, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
n6159, n6160, n6162, n6163, n6164, n6166, n6167, n6168, n6169, n6170,
n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6391, n6392,
n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
n6583, n6587, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
n6598, n6599, n6600, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6841,
n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6850, n6851, n6852,
n6853, n6854, n6855, n6856, n6857, n6859, n6860, n6861, n6862, n6863,
n6864, n6865, n6866, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
n6875, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6886,
n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6895, n6896, n6897,
n6898, n6899, n6900, n6901, n6902, n6904, n6905, n6906, n6907, n6908,
n6909, n6910, n6911, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6981,
n6982, n6983, n6984, n6985, n6987, n6988, n6989, n6990, n6991, n6992,
n6993, n6994, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7014, n7015,
n7016, n7017, n7018, n7019, n7020, n7021, n7023, n7024, n7025, n7026,
n7027, n7028, n7029, n7030, n7032, n7033, n7034, n7035, n7036, n7037,
n7038, n7039, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7059, n7060,
n7061, n7062, n7063, n7064, n7065, n7066, n7068, n7069, n7070, n7071,
n7072, n7073, n7074, n7075, n7077, n7078, n7079, n7080, n7081, n7082,
n7083, n7084, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
n7095, n7096, n7097, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
n7106, n7108, n7109, n7110, n7112, n7113, n7114, n7115, n7116, n7117,
n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7136, n7137, n7138,
n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7149, n7150,
n7151, n7152, n7153, n7154, n7155, n7156, n7158, n7159, n7160, n7161,
n7162, n7163, n7164, n7165, n7167, n7168, n7169, n7170, n7171, n7172,
n7173, n7174, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7194, n7195,
n7196, n7197, n7198, n7199, n7200, n7201, n7203, n7204, n7205, n7207,
n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
n7288, n7289, n7291, n7292, n7293, n7295, n7296, n7297, n7298, n7299,
n7300, n7301, n7302, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
n7311, n7312, n7313, n7314, n7315, n7316, n7318, n7319, n7320, n7321,
n7322, n7323, n7324, n7325, n7327, n7328, n7329, n7330, n7331, n7332,
n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
n7473, n7474, n7476, n7477, n7479, n7480, n7482, n7483, n7485, n7486,
n7488, n7489, n7491, n7492, n7494, n7495, n7497, n7498, n7499, n7500,
n7501;

dff g2814_reg ( clk, reset, ex_wire0, g51 );
not U_inv0 ( n7246, ex_wire0 );
dff g2817_reg ( clk, reset, ex_wire1, new_g16802_ );
not U_inv1 ( n7295, ex_wire1 );
dff g2933_reg ( clk, reset, g2933, new_g16823_ );
dff g2908_reg ( clk, reset, g2908, new_g26798_ );
dff g2883_reg ( clk, reset, g2883, new_g20825_ );
not U_inv2 ( n7105, g2883 );
dff g2888_reg ( clk, reset, g2888, new_g22026_ );
not U_inv3 ( n7381, g2888 );
dff g2896_reg ( clk, reset, g2896, new_g23358_ );
not U_inv4 ( n7106, g2896 );
dff g2892_reg ( clk, reset, g2892, new_g24473_ );
dff g2903_reg ( clk, reset, g2903, new_g25201_ );
not U_inv5 ( n7241, g2903 );
dff g2900_reg ( clk, reset, g2900, new_g26037_ );
not U_inv6 ( n7223, g2900 );
dff g2920_reg ( clk, reset, g2920, new_g25199_ );
dff g2912_reg ( clk, reset, g2912, new_g21989_ );
not U_inv7 ( n7238, g2912 );
dff g2917_reg ( clk, reset, g2917, new_g23357_ );
dff g2924_reg ( clk, reset, g2924, new_g24476_ );
not U_inv8 ( n7218, g2924 );
dff g2930_reg ( clk, reset, g8021, g51 );
dff g2929_reg ( clk, reset, ex_wire2, g8021 );
not U_inv9 ( n7293, ex_wire2 );
dff g2879_reg ( clk, reset, g2879, new_g12433_ );
not U_inv10 ( n7244, g2879 );
dff g2934_reg ( clk, reset, g2934, g3212 );
dff g2935_reg ( clk, reset, g2935, g3228 );
dff g2938_reg ( clk, reset, g2938, g3227 );
dff g2941_reg ( clk, reset, g2941, g3226 );
dff g2944_reg ( clk, reset, g2944, g3225 );
dff g2947_reg ( clk, reset, g2947, g3224 );
dff g2953_reg ( clk, reset, g2953, g3223 );
dff g2956_reg ( clk, reset, g2956, g3222 );
dff g2959_reg ( clk, reset, g2959, g3221 );
dff g2984_reg ( clk, reset, g2984, new_g16181_ );
dff g2962_reg ( clk, reset, g2962, g3232 );
dff g2963_reg ( clk, reset, g2963, g3220 );
dff g2966_reg ( clk, reset, g2966, g3219 );
dff g2969_reg ( clk, reset, g2969, g3218 );
dff g2972_reg ( clk, reset, g2972, g3217 );
dff g2975_reg ( clk, reset, g2975, g3216 );
dff g2978_reg ( clk, reset, g2978, g3215 );
dff g2981_reg ( clk, reset, g2981, g3214 );
dff g2874_reg ( clk, reset, g2874, g3213 );
dff g2985_reg ( clk, reset, g2985, new_g16132_ );
dff g1506_reg ( clk, reset, g1506, new_g18754_ );
not U_inv11 ( n7143, g1506 );
dff g1501_reg ( clk, reset, g1501, new_g18781_ );
not U_inv12 ( n7145, g1501 );
dff g1496_reg ( clk, reset, g1496, new_g18803_ );
not U_inv13 ( n7150, g1496 );
dff g1491_reg ( clk, reset, g1491, new_g18821_ );
not U_inv14 ( n7093, g1491 );
dff g1486_reg ( clk, reset, g1486, new_g18835_ );
not U_inv15 ( n7133, g1486 );
dff g1481_reg ( clk, reset, g1481, new_g18852_ );
not U_inv16 ( n7129, g1481 );
dff g1476_reg ( clk, reset, g1476, new_g18866_ );
not U_inv17 ( n7125, g1476 );
dff g1471_reg ( clk, reset, g1471, new_g18883_ );
not U_inv18 ( n7131, g1471 );
dff g2861_reg ( clk, reset, g8251, new_g19154_ );
dff g813_reg ( clk, reset, g813, g8251 );
not U_inv19 ( n7146, g813 );
dff g2864_reg ( clk, reset, g4090, new_g19163_ );
dff g809_reg ( clk, reset, g809, g4090 );
not U_inv20 ( n7151, g809 );
dff g2867_reg ( clk, reset, g4323, new_g19173_ );
dff g805_reg ( clk, reset, g805, g4323 );
not U_inv21 ( n7153, g805 );
dff g2870_reg ( clk, reset, g4590, new_g19184_ );
dff g801_reg ( clk, reset, g801, g4590 );
not U_inv22 ( n7095, g801 );
dff g2818_reg ( clk, reset, g6225, new_g20310_ );
dff g797_reg ( clk, reset, g797, g6225 );
not U_inv23 ( n7140, g797 );
dff g2821_reg ( clk, reset, g6442, new_g20343_ );
dff g793_reg ( clk, reset, g793, g6442 );
not U_inv24 ( n7134, g793 );
dff g2824_reg ( clk, reset, g6895, new_g20376_ );
dff g789_reg ( clk, reset, g789, g6895 );
not U_inv25 ( n7126, g789 );
dff g2827_reg ( clk, reset, g7334, new_g20417_ );
dff g785_reg ( clk, reset, g785, g7334 );
not U_inv26 ( n7137, g785 );
dff g2833_reg ( clk, reset, g8249, new_g19153_ );
dff g125_reg ( clk, reset, g125, g8249 );
not U_inv27 ( n7147, g125 );
dff g2836_reg ( clk, reset, g4088, new_g19162_ );
dff g121_reg ( clk, reset, g121, g4088 );
not U_inv28 ( n7152, g121 );
dff g2839_reg ( clk, reset, g4321, new_g19172_ );
dff g117_reg ( clk, reset, g117, g4321 );
not U_inv29 ( n7154, g117 );
dff g2842_reg ( clk, reset, g8023, new_g19144_ );
dff g113_reg ( clk, reset, g113, g8023 );
not U_inv30 ( n7096, g113 );
dff g2845_reg ( clk, reset, g8175, new_g19149_ );
dff g109_reg ( clk, reset, g109, g8175 );
not U_inv31 ( n7141, g109 );
dff g2848_reg ( clk, reset, g3993, new_g19157_ );
dff g105_reg ( clk, reset, g105, g3993 );
not U_inv32 ( n7136, g105 );
dff g2851_reg ( clk, reset, g4200, new_g19167_ );
dff g101_reg ( clk, reset, g101, g4200 );
not U_inv33 ( n7127, g101 );
dff g2854_reg ( clk, reset, g4450, new_g19178_ );
dff g97_reg ( clk, reset, g97, g4450 );
not U_inv34 ( n7138, g97 );
dff g2200_reg ( clk, reset, g2200, new_g18885_ );
not U_inv35 ( n7142, g2200 );
dff g2195_reg ( clk, reset, g2195, new_g18975_ );
not U_inv36 ( n7144, g2195 );
dff g2190_reg ( clk, reset, g2190, new_g18968_ );
not U_inv37 ( n7149, g2190 );
dff g2185_reg ( clk, reset, g2185, new_g18942_ );
not U_inv38 ( n7092, g2185 );
dff g2180_reg ( clk, reset, g2180, new_g18906_ );
not U_inv39 ( n7132, g2180 );
dff g2175_reg ( clk, reset, g2175, new_g18867_ );
not U_inv40 ( n7128, g2175 );
dff g2170_reg ( clk, reset, g2170, new_g18836_ );
not U_inv41 ( n7124, g2170 );
dff g2165_reg ( clk, reset, g2165, new_g18957_ );
not U_inv42 ( n7130, g2165 );
dff g138_reg ( clk, reset, n1058, g2950 );
not U_inv43 ( n7120, n1058 );
dff g135_reg ( clk, reset, n1062, g6231 );
not U_inv44 ( n7116, n1062 );
dff g165_reg ( clk, reset, g165, g6313 );
dff g169_reg ( clk, reset, g169, new_g25204_ );
dff g170_reg ( clk, reset, g170, new_g25206_ );
dff g168_reg ( clk, reset, g168, new_g25211_ );
dff g172_reg ( clk, reset, g172, new_g25207_ );
dff g173_reg ( clk, reset, g173, new_g25212_ );
dff g171_reg ( clk, reset, g171, new_g25218_ );
dff g175_reg ( clk, reset, g175, new_g25213_ );
dff g176_reg ( clk, reset, g176, new_g25219_ );
dff g174_reg ( clk, reset, g174, new_g25228_ );
dff g178_reg ( clk, reset, g178, new_g25220_ );
dff g179_reg ( clk, reset, g179, new_g25229_ );
dff g177_reg ( clk, reset, g177, new_g25239_ );
dff g180_reg ( clk, reset, n1481, new_g13110_ );
dff g182_reg ( clk, reset, g5549, n1481 );
dff g181_reg ( clk, reset, g181, g5549 );
not U_inv45 ( n7358, g181 );
dff g92_reg ( clk, reset, g92, new_g25027_ );
dff g88_reg ( clk, reset, g88, new_g25932_ );
dff g83_reg ( clk, reset, g83, new_g26529_ );
not U_inv46 ( n7192, g83 );
dff g79_reg ( clk, reset, g79, new_g27120_ );
dff g74_reg ( clk, reset, g74, new_g27594_ );
not U_inv47 ( n7213, g74 );
dff g70_reg ( clk, reset, g70, new_g28145_ );
dff g65_reg ( clk, reset, g65, new_g28634_ );
not U_inv48 ( n7233, g65 );
dff g61_reg ( clk, reset, g61, new_g29109_ );
dff g56_reg ( clk, reset, g56, new_g29353_ );
dff g52_reg ( clk, reset, g52, new_g29579_ );
dff g132_reg ( clk, reset, g132, new_g22161_ );
dff g162_reg ( clk, reset, g162, new_g22143_ );
dff g129_reg ( clk, reset, g129, new_g22141_ );
dff g159_reg ( clk, reset, g159, new_g22124_ );
dff g156_reg ( clk, reset, g156, new_g22101_ );
dff g153_reg ( clk, reset, g153, new_g22079_ );
dff g150_reg ( clk, reset, g150, new_g22063_ );
dff g147_reg ( clk, reset, g147, new_g22047_ );
dff g144_reg ( clk, reset, g144, new_g22037_ );
dff g141_reg ( clk, reset, g141, new_g22030_ );
dff g134_reg ( clk, reset, g134, new_g22142_ );
dff g164_reg ( clk, reset, g164, new_g22125_ );
dff g131_reg ( clk, reset, g131, new_g22122_ );
dff g161_reg ( clk, reset, g161, new_g22102_ );
dff g158_reg ( clk, reset, g158, new_g22080_ );
dff g155_reg ( clk, reset, g155, new_g22064_ );
dff g152_reg ( clk, reset, g152, new_g22048_ );
dff g149_reg ( clk, reset, g149, new_g22038_ );
dff g146_reg ( clk, reset, g146, new_g22031_ );
dff g143_reg ( clk, reset, g143, new_g22027_ );
dff g133_reg ( clk, reset, g133, new_g22123_ );
dff g163_reg ( clk, reset, g163, new_g22103_ );
dff g130_reg ( clk, reset, g130, new_g22100_ );
dff g160_reg ( clk, reset, g160, new_g22081_ );
dff g157_reg ( clk, reset, g157, new_g22065_ );
dff g154_reg ( clk, reset, g154, new_g22049_ );
dff g151_reg ( clk, reset, g151, new_g22039_ );
dff g148_reg ( clk, reset, g148, new_g22032_ );
dff g145_reg ( clk, reset, g145, new_g22028_ );
dff g142_reg ( clk, reset, g142, new_g22025_ );
dff g309_reg ( clk, reset, g309, g5549 );
not U_inv49 ( n7217, g309 );
dff g426_reg ( clk, reset, g426, new_g28754_ );
dff g414_reg ( clk, reset, g414, new_g28744_ );
dff g411_reg ( clk, reset, g411, new_g28735_ );
dff g408_reg ( clk, reset, g408, new_g28732_ );
dff g423_reg ( clk, reset, g423, new_g29201_ );
dff g420_reg ( clk, reset, g420, new_g29197_ );
dff g417_reg ( clk, reset, g417, new_g29194_ );
dff g428_reg ( clk, reset, g428, new_g28745_ );
dff g427_reg ( clk, reset, g427, new_g28736_ );
dff g435_reg ( clk, reset, g435, new_g26807_ );
dff g432_reg ( clk, reset, g432, new_g26804_ );
dff g429_reg ( clk, reset, g429, new_g26803_ );
dff g447_reg ( clk, reset, g447, new_g27762_ );
dff g444_reg ( clk, reset, g444, new_g26812_ );
dff g441_reg ( clk, reset, g441, new_g26808_ );
dff g438_reg ( clk, reset, g438, new_g26805_ );
dff g449_reg ( clk, reset, g449, new_g27760_ );
dff g448_reg ( clk, reset, g448, new_g27759_ );
dff g402_reg ( clk, reset, g402, new_g26664_ );
dff g219_reg ( clk, reset, g219, new_g30248_ );
dff g216_reg ( clk, reset, g216, new_g30246_ );
dff g213_reg ( clk, reset, g213, new_g30245_ );
dff g228_reg ( clk, reset, g228, new_g30639_ );
dff g225_reg ( clk, reset, g225, new_g30636_ );
dff g222_reg ( clk, reset, g222, new_g30635_ );
dff g273_reg ( clk, reset, g273, new_g30675_ );
dff g270_reg ( clk, reset, g270, new_g30669_ );
dff g267_reg ( clk, reset, g267, new_g30661_ );
dff g322_reg ( clk, reset, g322, new_g29167_ );
dff g317_reg ( clk, reset, g317, new_g30702_ );
dff g316_reg ( clk, reset, g316, new_g30700_ );
dff g315_reg ( clk, reset, g315, new_g30699_ );
dff g192_reg ( clk, reset, g192, new_g30275_ );
dff g189_reg ( clk, reset, g189, new_g30267_ );
dff g186_reg ( clk, reset, g186, new_g30261_ );
dff g320_reg ( clk, reset, g320, new_g30482_ );
dff g319_reg ( clk, reset, g319, new_g30468_ );
dff g318_reg ( clk, reset, g318, new_g30455_ );
dff g314_reg ( clk, reset, g314, new_g29611_ );
dff g313_reg ( clk, reset, g313, new_g29608_ );
dff g312_reg ( clk, reset, g312, new_g29606_ );
dff g237_reg ( clk, reset, g237, new_g30645_ );
dff g234_reg ( clk, reset, g234, new_g30640_ );
dff g231_reg ( clk, reset, g231, new_g30637_ );
dff g201_reg ( clk, reset, g201, new_g30680_ );
dff g198_reg ( clk, reset, g198, new_g30674_ );
dff g195_reg ( clk, reset, g195, new_g30668_ );
dff g246_reg ( clk, reset, g246, new_g30653_ );
dff g243_reg ( clk, reset, g243, new_g30646_ );
dff g240_reg ( clk, reset, g240, new_g30641_ );
dff g210_reg ( clk, reset, g210, new_g30292_ );
dff g207_reg ( clk, reset, g207, new_g30284_ );
dff g204_reg ( clk, reset, g204, new_g30276_ );
dff g255_reg ( clk, reset, g255, new_g30262_ );
dff g252_reg ( clk, reset, g252, new_g30257_ );
dff g249_reg ( clk, reset, g249, new_g30254_ );
dff g264_reg ( clk, reset, g264, new_g30268_ );
dff g261_reg ( clk, reset, g261, new_g30263_ );
dff g258_reg ( clk, reset, g258, new_g30258_ );
dff g321_reg ( clk, reset, g321, new_g29172_ );
dff g323_reg ( clk, reset, g323, new_g29169_ );
dff g354_reg ( clk, reset, g354, new_g27253_ );
dff g361_reg ( clk, reset, g361, new_g27265_ );
dff g358_reg ( clk, reset, g358, new_g27259_ );
dff g369_reg ( clk, reset, g369, new_g27256_ );
dff g376_reg ( clk, reset, g376, new_g27277_ );
dff g373_reg ( clk, reset, g373, new_g27266_ );
dff g384_reg ( clk, reset, g384, new_g27260_ );
dff g391_reg ( clk, reset, g391, new_g27293_ );
dff g388_reg ( clk, reset, g388, new_g27278_ );
dff g398_reg ( clk, reset, g398, new_g27267_ );
dff g346_reg ( clk, reset, g346, new_g27258_ );
dff g343_reg ( clk, reset, g343, new_g27255_ );
dff g404_reg ( clk, reset, g404, new_g26659_ );
dff g403_reg ( clk, reset, g403, new_g26655_ );
dff g450_reg ( clk, reset, n1737, n7147 );
dff g451_reg ( clk, reset, ex_wire3, n1737 );
not U_inv50 ( n7330, ex_wire3 );
dff g452_reg ( clk, reset, n1746, n7152 );
dff g453_reg ( clk, reset, ex_wire4, n1746 );
not U_inv51 ( n7329, ex_wire4 );
dff g454_reg ( clk, reset, n1755, n7154 );
dff g279_reg ( clk, reset, ex_wire5, n1755 );
not U_inv52 ( n7328, ex_wire5 );
dff g280_reg ( clk, reset, n1764, n7096 );
dff g281_reg ( clk, reset, ex_wire6, n1764 );
not U_inv53 ( n7327, ex_wire6 );
dff g282_reg ( clk, reset, n1773, n7141 );
dff g283_reg ( clk, reset, ex_wire7, n1773 );
not U_inv54 ( n7325, ex_wire7 );
dff g284_reg ( clk, reset, n1782, n7136 );
dff g285_reg ( clk, reset, ex_wire8, n1782 );
not U_inv55 ( n7324, ex_wire8 );
dff g286_reg ( clk, reset, n1791, n7127 );
dff g287_reg ( clk, reset, ex_wire9, n1791 );
not U_inv56 ( n7323, ex_wire9 );
dff g288_reg ( clk, reset, n1800, n7138 );
dff g289_reg ( clk, reset, ex_wire10, n1800 );
not U_inv57 ( n7322, ex_wire10 );
dff g299_reg ( clk, reset, g299, n7044 );
dff g298_reg ( clk, reset, g298, new_g26106_ );
dff g305_reg ( clk, reset, g305, new_g21346_ );
dff g342_reg ( clk, reset, n1883, g354 );
dff g349_reg ( clk, reset, g349, n1883 );
dff g350_reg ( clk, reset, n1892, g343 );
dff g351_reg ( clk, reset, g351, n1892 );
dff g352_reg ( clk, reset, n1901, g346 );
dff g353_reg ( clk, reset, g353, n1901 );
dff g357_reg ( clk, reset, n1910, g369 );
dff g364_reg ( clk, reset, g364, n1910 );
dff g365_reg ( clk, reset, n1919, g358 );
dff g366_reg ( clk, reset, g366, n1919 );
dff g367_reg ( clk, reset, n1928, g361 );
dff g368_reg ( clk, reset, g368, n1928 );
dff g372_reg ( clk, reset, n1937, g384 );
dff g379_reg ( clk, reset, g379, n1937 );
dff g380_reg ( clk, reset, n1946, g373 );
dff g381_reg ( clk, reset, g381, n1946 );
dff g382_reg ( clk, reset, n1955, g376 );
dff g383_reg ( clk, reset, g383, n1955 );
dff g387_reg ( clk, reset, n1964, g398 );
dff g394_reg ( clk, reset, g394, n1964 );
dff g395_reg ( clk, reset, n1973, g388 );
dff g396_reg ( clk, reset, g396, n1973 );
dff g397_reg ( clk, reset, n1982, g391 );
dff g324_reg ( clk, reset, g324, n1982 );
dff g474_reg ( clk, reset, g7909, g2950 );
not U_inv58 ( n7269, g7909 );
dff g481_reg ( clk, reset, g7956, g7909 );
not U_inv59 ( n7268, g7956 );
dff g485_reg ( clk, reset, g485, g7956 );
not U_inv60 ( n7273, g485 );
dff g486_reg ( clk, reset, g486, new_g23067_ );
dff g487_reg ( clk, reset, g487, new_g23093_ );
dff g488_reg ( clk, reset, g488, new_g23117_ );
dff g455_reg ( clk, reset, g455, new_g23385_ );
dff g564_reg ( clk, reset, n2045, g455 );
dff g569_reg ( clk, reset, g569, n2045 );
dff g458_reg ( clk, reset, g458, new_g23399_ );
dff g570_reg ( clk, reset, n2054, g458 );
dff g571_reg ( clk, reset, g571, n2054 );
dff g461_reg ( clk, reset, g461, new_g24174_ );
dff g572_reg ( clk, reset, n2063, g461 );
dff g573_reg ( clk, reset, g573, n2063 );
dff g477_reg ( clk, reset, g477, new_g24178_ );
dff g478_reg ( clk, reset, g478, new_g24207_ );
dff g479_reg ( clk, reset, g479, new_g24216_ );
dff g480_reg ( clk, reset, g480, new_g23092_ );
dff g484_reg ( clk, reset, g484, new_g23000_ );
dff g464_reg ( clk, reset, g464, new_g23022_ );
dff g465_reg ( clk, reset, g465, new_g24206_ );
dff g574_reg ( clk, reset, n2072, g465 );
dff g565_reg ( clk, reset, g565, n2072 );
dff g468_reg ( clk, reset, g468, new_g24215_ );
dff g566_reg ( clk, reset, n2081, g468 );
dff g567_reg ( clk, reset, g567, n2081 );
dff g471_reg ( clk, reset, g471, new_g24228_ );
dff g568_reg ( clk, reset, n2090, g471 );
dff g489_reg ( clk, reset, g489, n2090 );
dff g529_reg ( clk, reset, g529, n7330 );
dff g530_reg ( clk, reset, g530, n7329 );
dff g531_reg ( clk, reset, g531, n7328 );
dff g532_reg ( clk, reset, g532, n7327 );
dff g533_reg ( clk, reset, g533, n7325 );
dff g534_reg ( clk, reset, g534, n7324 );
dff g536_reg ( clk, reset, g536, n7323 );
dff g537_reg ( clk, reset, g537, n7322 );
dff g826_reg ( clk, reset, n2759, g2950 );
not U_inv61 ( n7119, n2759 );
dff g823_reg ( clk, reset, n2763, g6368 );
not U_inv62 ( n7115, n2763 );
dff g853_reg ( clk, reset, g853, g6518 );
dff g857_reg ( clk, reset, g857, new_g25209_ );
dff g858_reg ( clk, reset, g858, new_g25214_ );
dff g856_reg ( clk, reset, g856, new_g25221_ );
dff g860_reg ( clk, reset, g860, new_g25215_ );
dff g861_reg ( clk, reset, g861, new_g25222_ );
dff g859_reg ( clk, reset, g859, new_g25230_ );
dff g863_reg ( clk, reset, g863, new_g25223_ );
dff g864_reg ( clk, reset, g864, new_g25231_ );
dff g862_reg ( clk, reset, g862, new_g25240_ );
dff g866_reg ( clk, reset, g866, new_g25232_ );
dff g867_reg ( clk, reset, g867, new_g25241_ );
dff g865_reg ( clk, reset, g865, new_g25248_ );
dff g868_reg ( clk, reset, n3182, new_g13110_ );
dff g870_reg ( clk, reset, g5595, n3182 );
dff g869_reg ( clk, reset, g869, g5595 );
not U_inv63 ( n7357, g869 );
dff g780_reg ( clk, reset, g780, new_g25042_ );
dff g776_reg ( clk, reset, g776, new_g25935_ );
dff g771_reg ( clk, reset, g771, new_g26530_ );
not U_inv64 ( n7191, g771 );
dff g767_reg ( clk, reset, g767, new_g27123_ );
dff g762_reg ( clk, reset, g762, new_g27603_ );
not U_inv65 ( n7212, g762 );
dff g758_reg ( clk, reset, g758, new_g28146_ );
dff g753_reg ( clk, reset, g753, new_g28635_ );
not U_inv66 ( n7232, g753 );
dff g749_reg ( clk, reset, g749, new_g29110_ );
dff g744_reg ( clk, reset, g744, new_g29354_ );
dff g740_reg ( clk, reset, g740, new_g29580_ );
dff g820_reg ( clk, reset, g820, new_g22177_ );
dff g850_reg ( clk, reset, g850, new_g22164_ );
dff g817_reg ( clk, reset, g817, new_g22162_ );
dff g847_reg ( clk, reset, g847, new_g22147_ );
dff g844_reg ( clk, reset, g844, new_g22127_ );
dff g841_reg ( clk, reset, g841, new_g22104_ );
dff g838_reg ( clk, reset, g838, new_g22087_ );
dff g835_reg ( clk, reset, g835, new_g22066_ );
dff g832_reg ( clk, reset, g832, new_g22054_ );
dff g829_reg ( clk, reset, g829, new_g22040_ );
dff g822_reg ( clk, reset, g822, new_g22163_ );
dff g852_reg ( clk, reset, g852, new_g22148_ );
dff g819_reg ( clk, reset, g819, new_g22145_ );
dff g849_reg ( clk, reset, g849, new_g22128_ );
dff g846_reg ( clk, reset, g846, new_g22105_ );
dff g843_reg ( clk, reset, g843, new_g22088_ );
dff g840_reg ( clk, reset, g840, new_g22067_ );
dff g837_reg ( clk, reset, g837, new_g22055_ );
dff g834_reg ( clk, reset, g834, new_g22041_ );
dff g831_reg ( clk, reset, g831, new_g22033_ );
dff g821_reg ( clk, reset, g821, new_g22146_ );
dff g851_reg ( clk, reset, g851, new_g22129_ );
dff g818_reg ( clk, reset, g818, new_g22126_ );
dff g848_reg ( clk, reset, g848, new_g22106_ );
dff g845_reg ( clk, reset, g845, new_g22089_ );
dff g842_reg ( clk, reset, g842, new_g22068_ );
dff g839_reg ( clk, reset, g839, new_g22056_ );
dff g836_reg ( clk, reset, g836, new_g22042_ );
dff g833_reg ( clk, reset, g833, new_g22034_ );
dff g830_reg ( clk, reset, g830, new_g22029_ );
dff g996_reg ( clk, reset, g996, g5595 );
not U_inv67 ( n7214, g996 );
dff g1113_reg ( clk, reset, g1113, new_g28767_ );
dff g1101_reg ( clk, reset, g1101, new_g28758_ );
dff g1098_reg ( clk, reset, g1098, new_g28746_ );
dff g1095_reg ( clk, reset, g1095, new_g28738_ );
dff g1110_reg ( clk, reset, g1110, new_g29209_ );
dff g1107_reg ( clk, reset, g1107, new_g29204_ );
dff g1104_reg ( clk, reset, g1104, new_g29198_ );
dff g1115_reg ( clk, reset, g1115, new_g28759_ );
dff g1114_reg ( clk, reset, g1114, new_g28747_ );
dff g1122_reg ( clk, reset, g1122, new_g26813_ );
dff g1119_reg ( clk, reset, g1119, new_g26809_ );
dff g1116_reg ( clk, reset, g1116, new_g26806_ );
dff g1134_reg ( clk, reset, g1134, new_g27765_ );
dff g1131_reg ( clk, reset, g1131, new_g26818_ );
dff g1128_reg ( clk, reset, g1128, new_g26814_ );
dff g1125_reg ( clk, reset, g1125, new_g26810_ );
dff g1136_reg ( clk, reset, g1136, new_g27763_ );
dff g1135_reg ( clk, reset, g1135, new_g27761_ );
dff g1089_reg ( clk, reset, g1089, new_g26669_ );
dff g906_reg ( clk, reset, g906, new_g30251_ );
dff g903_reg ( clk, reset, g903, new_g30249_ );
dff g900_reg ( clk, reset, g900, new_g30247_ );
dff g915_reg ( clk, reset, g915, new_g30647_ );
dff g912_reg ( clk, reset, g912, new_g30642_ );
dff g909_reg ( clk, reset, g909, new_g30638_ );
dff g960_reg ( clk, reset, g960, new_g30682_ );
dff g957_reg ( clk, reset, g957, new_g30677_ );
dff g954_reg ( clk, reset, g954, new_g30670_ );
dff g1009_reg ( clk, reset, g1009, new_g29170_ );
dff g1004_reg ( clk, reset, g1004, new_g30705_ );
dff g1003_reg ( clk, reset, g1003, new_g30703_ );
dff g1002_reg ( clk, reset, g1002, new_g30701_ );
dff g879_reg ( clk, reset, g879, new_g30285_ );
dff g876_reg ( clk, reset, g876, new_g30277_ );
dff g873_reg ( clk, reset, g873, new_g30269_ );
dff g1007_reg ( clk, reset, g1007, new_g30500_ );
dff g1006_reg ( clk, reset, g1006, new_g30485_ );
dff g1005_reg ( clk, reset, g1005, new_g30470_ );
dff g1001_reg ( clk, reset, g1001, new_g29616_ );
dff g1000_reg ( clk, reset, g1000, new_g29612_ );
dff g999_reg ( clk, reset, g999, new_g29609_ );
dff g924_reg ( clk, reset, g924, new_g30654_ );
dff g921_reg ( clk, reset, g921, new_g30648_ );
dff g918_reg ( clk, reset, g918, new_g30643_ );
dff g888_reg ( clk, reset, g888, new_g30687_ );
dff g885_reg ( clk, reset, g885, new_g30681_ );
dff g882_reg ( clk, reset, g882, new_g30676_ );
dff g933_reg ( clk, reset, g933, new_g30662_ );
dff g930_reg ( clk, reset, g930, new_g30655_ );
dff g927_reg ( clk, reset, g927, new_g30649_ );
dff g897_reg ( clk, reset, g897, new_g30298_ );
dff g894_reg ( clk, reset, g894, new_g30293_ );
dff g891_reg ( clk, reset, g891, new_g30286_ );
dff g942_reg ( clk, reset, g942, new_g30270_ );
dff g939_reg ( clk, reset, g939, new_g30264_ );
dff g936_reg ( clk, reset, g936, new_g30259_ );
dff g951_reg ( clk, reset, g951, new_g30278_ );
dff g948_reg ( clk, reset, g948, new_g30271_ );
dff g945_reg ( clk, reset, g945, new_g30265_ );
dff g1008_reg ( clk, reset, g1008, new_g29179_ );
dff g1010_reg ( clk, reset, g1010, new_g29173_ );
dff g1041_reg ( clk, reset, g1041, new_g27257_ );
dff g1048_reg ( clk, reset, g1048, new_g27282_ );
dff g1045_reg ( clk, reset, g1045, new_g27271_ );
dff g1056_reg ( clk, reset, g1056, new_g27263_ );
dff g1063_reg ( clk, reset, g1063, new_g27297_ );
dff g1060_reg ( clk, reset, g1060, new_g27283_ );
dff g1071_reg ( clk, reset, g1071, new_g27272_ );
dff g1078_reg ( clk, reset, g1078, new_g27313_ );
dff g1075_reg ( clk, reset, g1075, new_g27298_ );
dff g1085_reg ( clk, reset, g1085, new_g27284_ );
dff g1033_reg ( clk, reset, g1033, new_g27270_ );
dff g1030_reg ( clk, reset, g1030, new_g27262_ );
dff g1091_reg ( clk, reset, g1091, new_g26665_ );
dff g1090_reg ( clk, reset, g1090, new_g26661_ );
dff g1137_reg ( clk, reset, n3438, n7146 );
dff g1138_reg ( clk, reset, ex_wire11, n3438 );
not U_inv68 ( n7321, ex_wire11 );
dff g1139_reg ( clk, reset, n3447, n7151 );
dff g1140_reg ( clk, reset, ex_wire12, n3447 );
not U_inv69 ( n7320, ex_wire12 );
dff g1141_reg ( clk, reset, n3456, n7153 );
dff g966_reg ( clk, reset, ex_wire13, n3456 );
not U_inv70 ( n7319, ex_wire13 );
dff g967_reg ( clk, reset, n3465, n7095 );
dff g968_reg ( clk, reset, ex_wire14, n3465 );
not U_inv71 ( n7318, ex_wire14 );
dff g969_reg ( clk, reset, n3474, n7140 );
dff g970_reg ( clk, reset, ex_wire15, n3474 );
not U_inv72 ( n7316, ex_wire15 );
dff g971_reg ( clk, reset, n3483, n7134 );
dff g972_reg ( clk, reset, ex_wire16, n3483 );
not U_inv73 ( n7315, ex_wire16 );
dff g973_reg ( clk, reset, n3492, n7126 );
dff g974_reg ( clk, reset, ex_wire17, n3492 );
not U_inv74 ( n7314, ex_wire17 );
dff g975_reg ( clk, reset, n3501, n7137 );
dff g976_reg ( clk, reset, ex_wire18, n3501 );
not U_inv75 ( n7313, ex_wire18 );
dff g986_reg ( clk, reset, g986, n7086 );
not U_inv76 ( n7228, g986 );
dff g985_reg ( clk, reset, g985, new_g26120_ );
dff g992_reg ( clk, reset, g992, n203 );
dff g1029_reg ( clk, reset, n3584, g1041 );
dff g1036_reg ( clk, reset, g1036, n3584 );
dff g1037_reg ( clk, reset, n3593, g1030 );
dff g1038_reg ( clk, reset, g1038, n3593 );
dff g1039_reg ( clk, reset, n3602, g1033 );
dff g1040_reg ( clk, reset, g1040, n3602 );
dff g1044_reg ( clk, reset, n3611, g1056 );
dff g1051_reg ( clk, reset, g1051, n3611 );
dff g1052_reg ( clk, reset, n3620, g1045 );
dff g1053_reg ( clk, reset, g1053, n3620 );
dff g1054_reg ( clk, reset, n3629, g1048 );
dff g1055_reg ( clk, reset, g1055, n3629 );
dff g1059_reg ( clk, reset, n3638, g1071 );
dff g1066_reg ( clk, reset, g1066, n3638 );
dff g1067_reg ( clk, reset, n3647, g1060 );
dff g1068_reg ( clk, reset, g1068, n3647 );
dff g1069_reg ( clk, reset, n3656, g1063 );
dff g1070_reg ( clk, reset, g1070, n3656 );
dff g1074_reg ( clk, reset, n3665, g1085 );
dff g1081_reg ( clk, reset, g1081, n3665 );
dff g1082_reg ( clk, reset, n3674, g1075 );
dff g1083_reg ( clk, reset, g1083, n3674 );
dff g1084_reg ( clk, reset, n3683, g1078 );
dff g1011_reg ( clk, reset, g1011, n3683 );
dff g1161_reg ( clk, reset, g7961, g2950 );
not U_inv77 ( n7265, g7961 );
dff g1168_reg ( clk, reset, g8007, g7961 );
not U_inv78 ( n7264, g8007 );
dff g1172_reg ( clk, reset, g1172, g8007 );
not U_inv79 ( n7270, g1172 );
dff g1173_reg ( clk, reset, g1173, new_g23081_ );
dff g1174_reg ( clk, reset, g1174, new_g23111_ );
dff g1175_reg ( clk, reset, g1175, new_g23126_ );
dff g1142_reg ( clk, reset, g1142, new_g23392_ );
dff g1250_reg ( clk, reset, n3746, g1142 );
dff g1255_reg ( clk, reset, g1255, n3746 );
dff g1145_reg ( clk, reset, g1145, new_g23406_ );
dff g1256_reg ( clk, reset, n3755, g1145 );
dff g1257_reg ( clk, reset, g1257, n3755 );
dff g1148_reg ( clk, reset, g1148, new_g24179_ );
dff g1258_reg ( clk, reset, n3764, g1148 );
dff g1259_reg ( clk, reset, g1259, n3764 );
dff g1164_reg ( clk, reset, g1164, new_g24181_ );
dff g1165_reg ( clk, reset, g1165, new_g24213_ );
dff g1166_reg ( clk, reset, g1166, new_g24223_ );
dff g1167_reg ( clk, reset, g1167, new_g23110_ );
dff g1171_reg ( clk, reset, g1171, new_g23014_ );
dff g1151_reg ( clk, reset, g1151, new_g23039_ );
dff g1152_reg ( clk, reset, g1152, new_g24212_ );
dff g1260_reg ( clk, reset, n3773, g1152 );
dff g1251_reg ( clk, reset, g1251, n3773 );
dff g1155_reg ( clk, reset, g1155, new_g24222_ );
dff g1252_reg ( clk, reset, n3782, g1155 );
dff g1253_reg ( clk, reset, g1253, n3782 );
dff g1158_reg ( clk, reset, g1158, new_g24235_ );
dff g1254_reg ( clk, reset, n3791, g1158 );
dff g1176_reg ( clk, reset, g1176, n3791 );
dff g1215_reg ( clk, reset, g1215, n7321 );
dff g1216_reg ( clk, reset, g1216, n7320 );
dff g1217_reg ( clk, reset, g1217, n7319 );
dff g1218_reg ( clk, reset, g1218, n7318 );
dff g1219_reg ( clk, reset, g1219, n7316 );
dff g1220_reg ( clk, reset, g1220, n7315 );
dff g1222_reg ( clk, reset, g1222, n7314 );
dff g1223_reg ( clk, reset, g1223, n7313 );
dff g1520_reg ( clk, reset, n4460, g2950 );
not U_inv80 ( n7118, n4460 );
dff g1517_reg ( clk, reset, n4464, g6573 );
not U_inv81 ( n7114, n4464 );
dff g1547_reg ( clk, reset, g1547, g6782 );
dff g1551_reg ( clk, reset, g1551, new_g25217_ );
dff g1552_reg ( clk, reset, g1552, new_g25224_ );
dff g1550_reg ( clk, reset, g1550, new_g25233_ );
dff g1554_reg ( clk, reset, g1554, new_g25225_ );
dff g1555_reg ( clk, reset, g1555, new_g25234_ );
dff g1553_reg ( clk, reset, g1553, new_g25242_ );
dff g1557_reg ( clk, reset, g1557, new_g25235_ );
dff g1558_reg ( clk, reset, g1558, new_g25243_ );
dff g1556_reg ( clk, reset, g1556, new_g25249_ );
dff g1560_reg ( clk, reset, g1560, new_g25244_ );
dff g1561_reg ( clk, reset, g1561, new_g25250_ );
dff g1559_reg ( clk, reset, g1559, new_g25255_ );
dff g1562_reg ( clk, reset, n4883, new_g13110_ );
dff g1564_reg ( clk, reset, g5612, n4883 );
dff g1563_reg ( clk, reset, g1563, g5612 );
not U_inv82 ( n7356, g1563 );
dff g1466_reg ( clk, reset, g1466, new_g25056_ );
dff g1462_reg ( clk, reset, g1462, new_g25938_ );
dff g1457_reg ( clk, reset, g1457, new_g26531_ );
not U_inv83 ( n7190, g1457 );
dff g1453_reg ( clk, reset, g1453, new_g27129_ );
dff g1448_reg ( clk, reset, g1448, new_g27612_ );
not U_inv84 ( n7211, g1448 );
dff g1444_reg ( clk, reset, g1444, new_g28147_ );
dff g1439_reg ( clk, reset, g1439, new_g28636_ );
not U_inv85 ( n7231, g1439 );
dff g1435_reg ( clk, reset, g1435, new_g29111_ );
dff g1430_reg ( clk, reset, g1430, new_g29355_ );
dff g1426_reg ( clk, reset, g1426, new_g29581_ );
dff g1514_reg ( clk, reset, g1514, new_g22191_ );
dff g1544_reg ( clk, reset, g1544, new_g22180_ );
dff g1511_reg ( clk, reset, g1511, new_g22178_ );
dff g1541_reg ( clk, reset, g1541, new_g22168_ );
dff g1538_reg ( clk, reset, g1538, new_g22150_ );
dff g1535_reg ( clk, reset, g1535, new_g22130_ );
dff g1532_reg ( clk, reset, g1532, new_g22112_ );
dff g1529_reg ( clk, reset, g1529, new_g22090_ );
dff g1526_reg ( clk, reset, g1526, new_g22073_ );
dff g1523_reg ( clk, reset, g1523, new_g22057_ );
dff g1516_reg ( clk, reset, g1516, new_g22179_ );
dff g1546_reg ( clk, reset, g1546, new_g22169_ );
dff g1513_reg ( clk, reset, g1513, new_g22166_ );
dff g1543_reg ( clk, reset, g1543, new_g22151_ );
dff g1540_reg ( clk, reset, g1540, new_g22131_ );
dff g1537_reg ( clk, reset, g1537, new_g22113_ );
dff g1534_reg ( clk, reset, g1534, new_g22091_ );
dff g1531_reg ( clk, reset, g1531, new_g22074_ );
dff g1528_reg ( clk, reset, g1528, new_g22058_ );
dff g1525_reg ( clk, reset, g1525, new_g22043_ );
dff g1515_reg ( clk, reset, g1515, new_g22167_ );
dff g1545_reg ( clk, reset, g1545, new_g22152_ );
dff g1512_reg ( clk, reset, g1512, new_g22149_ );
dff g1542_reg ( clk, reset, g1542, new_g22132_ );
dff g1539_reg ( clk, reset, g1539, new_g22114_ );
dff g1536_reg ( clk, reset, g1536, new_g22092_ );
dff g1533_reg ( clk, reset, g1533, new_g22075_ );
dff g1530_reg ( clk, reset, g1530, new_g22059_ );
dff g1527_reg ( clk, reset, g1527, new_g22044_ );
dff g1524_reg ( clk, reset, g1524, new_g22035_ );
dff g1690_reg ( clk, reset, g1690, g5612 );
not U_inv86 ( n7216, g1690 );
dff g1807_reg ( clk, reset, g1807, new_g28778_ );
dff g1795_reg ( clk, reset, g1795, new_g28771_ );
dff g1792_reg ( clk, reset, g1792, new_g28760_ );
dff g1789_reg ( clk, reset, g1789, new_g28749_ );
dff g1804_reg ( clk, reset, g1804, new_g29218_ );
dff g1801_reg ( clk, reset, g1801, new_g29212_ );
dff g1798_reg ( clk, reset, g1798, new_g29205_ );
dff g1809_reg ( clk, reset, g1809, new_g28772_ );
dff g1808_reg ( clk, reset, g1808, new_g28761_ );
dff g1816_reg ( clk, reset, g1816, new_g26820_ );
dff g1813_reg ( clk, reset, g1813, new_g26815_ );
dff g1810_reg ( clk, reset, g1810, new_g26811_ );
dff g1828_reg ( clk, reset, g1828, new_g27768_ );
dff g1825_reg ( clk, reset, g1825, new_g26824_ );
dff g1822_reg ( clk, reset, g1822, new_g26821_ );
dff g1819_reg ( clk, reset, g1819, new_g26816_ );
dff g1830_reg ( clk, reset, g1830, new_g27766_ );
dff g1829_reg ( clk, reset, g1829, new_g27764_ );
dff g1783_reg ( clk, reset, g1783, new_g26675_ );
dff g1600_reg ( clk, reset, g1600, new_g30255_ );
dff g1597_reg ( clk, reset, g1597, new_g30252_ );
dff g1594_reg ( clk, reset, g1594, new_g30250_ );
dff g1609_reg ( clk, reset, g1609, new_g30656_ );
dff g1606_reg ( clk, reset, g1606, new_g30650_ );
dff g1603_reg ( clk, reset, g1603, new_g30644_ );
dff g1654_reg ( clk, reset, g1654, new_g30689_ );
dff g1651_reg ( clk, reset, g1651, new_g30684_ );
dff g1648_reg ( clk, reset, g1648, new_g30678_ );
dff g1703_reg ( clk, reset, g1703, new_g29178_ );
dff g1698_reg ( clk, reset, g1698, new_g30708_ );
dff g1697_reg ( clk, reset, g1697, new_g30706_ );
dff g1696_reg ( clk, reset, g1696, new_g30704_ );
dff g1573_reg ( clk, reset, g1573, new_g30294_ );
dff g1570_reg ( clk, reset, g1570, new_g30287_ );
dff g1567_reg ( clk, reset, g1567, new_g30279_ );
dff g1700_reg ( clk, reset, g1700, new_g30503_ );
dff g1699_reg ( clk, reset, g1699, new_g30487_ );
dff g1701_reg ( clk, reset, g1701, new_g30338_ );
dff g1695_reg ( clk, reset, g1695, new_g29620_ );
dff g1694_reg ( clk, reset, g1694, new_g29617_ );
dff g1693_reg ( clk, reset, g1693, new_g29613_ );
dff g1618_reg ( clk, reset, g1618, new_g30663_ );
dff g1615_reg ( clk, reset, g1615, new_g30657_ );
dff g1612_reg ( clk, reset, g1612, new_g30651_ );
dff g1582_reg ( clk, reset, g1582, new_g30692_ );
dff g1579_reg ( clk, reset, g1579, new_g30688_ );
dff g1576_reg ( clk, reset, g1576, new_g30683_ );
dff g1627_reg ( clk, reset, g1627, new_g30671_ );
dff g1624_reg ( clk, reset, g1624, new_g30664_ );
dff g1621_reg ( clk, reset, g1621, new_g30658_ );
dff g1591_reg ( clk, reset, g1591, new_g30302_ );
dff g1588_reg ( clk, reset, g1588, new_g30299_ );
dff g1585_reg ( clk, reset, g1585, new_g30295_ );
dff g1636_reg ( clk, reset, g1636, new_g30280_ );
dff g1633_reg ( clk, reset, g1633, new_g30272_ );
dff g1630_reg ( clk, reset, g1630, new_g30266_ );
dff g1645_reg ( clk, reset, g1645, new_g30288_ );
dff g1642_reg ( clk, reset, g1642, new_g30281_ );
dff g1639_reg ( clk, reset, g1639, new_g30273_ );
dff g1702_reg ( clk, reset, g1702, new_g29184_ );
dff g1704_reg ( clk, reset, g1704, new_g29181_ );
dff g1735_reg ( clk, reset, g1735, new_g27264_ );
dff g1742_reg ( clk, reset, g1742, new_g27302_ );
dff g1739_reg ( clk, reset, g1739, new_g27288_ );
dff g1750_reg ( clk, reset, g1750, new_g27275_ );
dff g1757_reg ( clk, reset, g1757, new_g27317_ );
dff g1754_reg ( clk, reset, g1754, new_g27303_ );
dff g1765_reg ( clk, reset, g1765, new_g27289_ );
dff g1772_reg ( clk, reset, g1772, new_g27330_ );
dff g1769_reg ( clk, reset, g1769, new_g27318_ );
dff g1779_reg ( clk, reset, g1779, new_g27304_ );
dff g1727_reg ( clk, reset, g1727, new_g27287_ );
dff g1724_reg ( clk, reset, g1724, new_g27274_ );
dff g1785_reg ( clk, reset, g1785, new_g26670_ );
dff g1784_reg ( clk, reset, g1784, new_g26667_ );
dff g1831_reg ( clk, reset, n5139, n7143 );
dff g1832_reg ( clk, reset, ex_wire19, n5139 );
not U_inv87 ( n7312, ex_wire19 );
dff g1833_reg ( clk, reset, n5148, n7145 );
dff g1834_reg ( clk, reset, ex_wire20, n5148 );
not U_inv88 ( n7311, ex_wire20 );
dff g1835_reg ( clk, reset, n5157, n7150 );
dff g1660_reg ( clk, reset, ex_wire21, n5157 );
not U_inv89 ( n7310, ex_wire21 );
dff g1661_reg ( clk, reset, n5166, n7093 );
dff g1662_reg ( clk, reset, ex_wire22, n5166 );
not U_inv90 ( n7309, ex_wire22 );
dff g1663_reg ( clk, reset, n5175, n7133 );
dff g1664_reg ( clk, reset, ex_wire23, n5175 );
not U_inv91 ( n7308, ex_wire23 );
dff g1665_reg ( clk, reset, n5184, n7129 );
dff g1666_reg ( clk, reset, ex_wire24, n5184 );
not U_inv92 ( n7307, ex_wire24 );
dff g1667_reg ( clk, reset, n5193, n7125 );
dff g1668_reg ( clk, reset, ex_wire25, n5193 );
not U_inv93 ( n7306, ex_wire25 );
dff g1669_reg ( clk, reset, n5202, n7131 );
dff g1670_reg ( clk, reset, ex_wire26, n5202 );
not U_inv94 ( n7305, ex_wire26 );
dff g1680_reg ( clk, reset, g1680, n7087 );
not U_inv95 ( n7247, g1680 );
dff g1679_reg ( clk, reset, g1679, new_g26130_ );
dff g1686_reg ( clk, reset, g1686, new_g28903_ );
dff g1723_reg ( clk, reset, n5285, g1735 );
dff g1730_reg ( clk, reset, g1730, n5285 );
dff g1731_reg ( clk, reset, n5294, g1724 );
dff g1732_reg ( clk, reset, g1732, n5294 );
dff g1733_reg ( clk, reset, n5303, g1727 );
dff g1734_reg ( clk, reset, g1734, n5303 );
dff g1738_reg ( clk, reset, n5312, g1750 );
dff g1745_reg ( clk, reset, g1745, n5312 );
dff g1746_reg ( clk, reset, n5321, g1739 );
dff g1747_reg ( clk, reset, g1747, n5321 );
dff g1748_reg ( clk, reset, n5330, g1742 );
dff g1749_reg ( clk, reset, g1749, n5330 );
dff g1753_reg ( clk, reset, n5339, g1765 );
dff g1760_reg ( clk, reset, g1760, n5339 );
dff g1761_reg ( clk, reset, n5348, g1754 );
dff g1762_reg ( clk, reset, g1762, n5348 );
dff g1763_reg ( clk, reset, n5357, g1757 );
dff g1764_reg ( clk, reset, g1764, n5357 );
dff g1768_reg ( clk, reset, n5366, g1779 );
dff g1775_reg ( clk, reset, g1775, n5366 );
dff g1776_reg ( clk, reset, n5375, g1769 );
dff g1777_reg ( clk, reset, g1777, n5375 );
dff g1778_reg ( clk, reset, n5384, g1772 );
dff g1705_reg ( clk, reset, g1705, n5384 );
dff g1855_reg ( clk, reset, g8012, g2950 );
not U_inv96 ( n7267, g8012 );
dff g1862_reg ( clk, reset, g8082, g8012 );
not U_inv97 ( n7266, g8082 );
dff g1866_reg ( clk, reset, g1866, g8082 );
not U_inv98 ( n7272, g1866 );
dff g1867_reg ( clk, reset, g1867, new_g23097_ );
dff g1868_reg ( clk, reset, g1868, new_g23124_ );
dff g1869_reg ( clk, reset, g1869, new_g23137_ );
dff g1836_reg ( clk, reset, g1836, new_g23400_ );
dff g1944_reg ( clk, reset, n5447, g1836 );
dff g1949_reg ( clk, reset, g1949, n5447 );
dff g1839_reg ( clk, reset, g1839, new_g23413_ );
dff g1950_reg ( clk, reset, n5456, g1839 );
dff g1951_reg ( clk, reset, g1951, n5456 );
dff g1842_reg ( clk, reset, g1842, new_g24182_ );
dff g1952_reg ( clk, reset, n5465, g1842 );
dff g1953_reg ( clk, reset, g1953, n5465 );
dff g1858_reg ( clk, reset, g1858, new_g24208_ );
dff g1859_reg ( clk, reset, g1859, new_g24219_ );
dff g1860_reg ( clk, reset, g1860, new_g24231_ );
dff g1861_reg ( clk, reset, g1861, new_g23123_ );
dff g1865_reg ( clk, reset, g1865, new_g23030_ );
dff g1845_reg ( clk, reset, g1845, new_g23058_ );
dff g1846_reg ( clk, reset, g1846, new_g24218_ );
dff g1954_reg ( clk, reset, n5474, g1846 );
dff g1945_reg ( clk, reset, g1945, n5474 );
dff g1849_reg ( clk, reset, g1849, new_g24230_ );
dff g1946_reg ( clk, reset, n5483, g1849 );
dff g1947_reg ( clk, reset, g1947, n5483 );
dff g1852_reg ( clk, reset, g1852, new_g24243_ );
dff g1948_reg ( clk, reset, n5492, g1852 );
dff g1870_reg ( clk, reset, g1870, n5492 );
dff g1909_reg ( clk, reset, g1909, n7312 );
dff g1910_reg ( clk, reset, g1910, n7311 );
dff g1911_reg ( clk, reset, g1911, n7310 );
dff g1912_reg ( clk, reset, g1912, n7309 );
dff g1913_reg ( clk, reset, g1913, n7308 );
dff g1914_reg ( clk, reset, g1914, n7307 );
dff g1916_reg ( clk, reset, g1916, n7306 );
dff g1917_reg ( clk, reset, g1917, n7305 );
dff g2214_reg ( clk, reset, n6161, g2950 );
not U_inv99 ( n7117, n6161 );
dff g2211_reg ( clk, reset, n6165, g6837 );
not U_inv100 ( n7113, n6165 );
dff g2241_reg ( clk, reset, g2241, g7084 );
dff g2245_reg ( clk, reset, g2245, new_g25227_ );
dff g2246_reg ( clk, reset, g2246, new_g25236_ );
dff g2244_reg ( clk, reset, g2244, new_g25245_ );
dff g2248_reg ( clk, reset, g2248, new_g25237_ );
dff g2249_reg ( clk, reset, g2249, new_g25246_ );
dff g2247_reg ( clk, reset, g2247, new_g25251_ );
dff g2251_reg ( clk, reset, g2251, new_g25247_ );
dff g2252_reg ( clk, reset, g2252, new_g25252_ );
dff g2250_reg ( clk, reset, g2250, new_g25256_ );
dff g2254_reg ( clk, reset, g2254, new_g25253_ );
dff g2255_reg ( clk, reset, g2255, new_g25257_ );
dff g2253_reg ( clk, reset, g2253, new_g25259_ );
dff g2256_reg ( clk, reset, n6584, new_g13110_ );
dff g2258_reg ( clk, reset, g5637, n6584 );
dff g2257_reg ( clk, reset, g2257, g5637 );
not U_inv101 ( n7355, g2257 );
dff g2160_reg ( clk, reset, g2160, new_g25067_ );
dff g2156_reg ( clk, reset, g2156, new_g25940_ );
dff g2151_reg ( clk, reset, g2151, new_g26532_ );
not U_inv102 ( n7189, g2151 );
dff g2147_reg ( clk, reset, g2147, new_g27131_ );
dff g2142_reg ( clk, reset, g2142, new_g27621_ );
not U_inv103 ( n7210, g2142 );
dff g2138_reg ( clk, reset, g2138, new_g28148_ );
dff g2133_reg ( clk, reset, g2133, new_g28637_ );
not U_inv104 ( n7230, g2133 );
dff g2129_reg ( clk, reset, g2129, new_g29112_ );
dff g2124_reg ( clk, reset, g2124, new_g29357_ );
dff g2120_reg ( clk, reset, g2120, new_g29582_ );
dff g2208_reg ( clk, reset, g2208, new_g22200_ );
dff g2238_reg ( clk, reset, g2238, new_g22194_ );
dff g2205_reg ( clk, reset, g2205, new_g22192_ );
dff g2235_reg ( clk, reset, g2235, new_g22184_ );
dff g2232_reg ( clk, reset, g2232, new_g22171_ );
dff g2229_reg ( clk, reset, g2229, new_g22153_ );
dff g2226_reg ( clk, reset, g2226, new_g22138_ );
dff g2223_reg ( clk, reset, g2223, new_g22115_ );
dff g2220_reg ( clk, reset, g2220, new_g22097_ );
dff g2217_reg ( clk, reset, g2217, new_g22076_ );
dff g2210_reg ( clk, reset, g2210, new_g22193_ );
dff g2240_reg ( clk, reset, g2240, new_g22185_ );
dff g2207_reg ( clk, reset, g2207, new_g22182_ );
dff g2237_reg ( clk, reset, g2237, new_g22172_ );
dff g2234_reg ( clk, reset, g2234, new_g22154_ );
dff g2231_reg ( clk, reset, g2231, new_g22139_ );
dff g2228_reg ( clk, reset, g2228, new_g22116_ );
dff g2225_reg ( clk, reset, g2225, new_g22098_ );
dff g2222_reg ( clk, reset, g2222, new_g22077_ );
dff g2219_reg ( clk, reset, g2219, new_g22060_ );
dff g2209_reg ( clk, reset, g2209, new_g22183_ );
dff g2239_reg ( clk, reset, g2239, new_g22173_ );
dff g2206_reg ( clk, reset, g2206, new_g22170_ );
dff g2236_reg ( clk, reset, g2236, new_g22155_ );
dff g2233_reg ( clk, reset, g2233, new_g22140_ );
dff g2230_reg ( clk, reset, g2230, new_g22117_ );
dff g2227_reg ( clk, reset, g2227, new_g22099_ );
dff g2224_reg ( clk, reset, g2224, new_g22078_ );
dff g2221_reg ( clk, reset, g2221, new_g22061_ );
dff g2218_reg ( clk, reset, g2218, new_g22045_ );
dff g2384_reg ( clk, reset, g2384, g5637 );
not U_inv105 ( n7215, g2384 );
dff g2501_reg ( clk, reset, g2501, new_g28788_ );
dff g2489_reg ( clk, reset, g2489, new_g28782_ );
dff g2486_reg ( clk, reset, g2486, new_g28773_ );
dff g2483_reg ( clk, reset, g2483, new_g28763_ );
dff g2498_reg ( clk, reset, g2498, new_g29226_ );
dff g2495_reg ( clk, reset, g2495, new_g29221_ );
dff g2492_reg ( clk, reset, g2492, new_g29213_ );
dff g2503_reg ( clk, reset, g2503, new_g28783_ );
dff g2502_reg ( clk, reset, g2502, new_g28774_ );
dff g2510_reg ( clk, reset, g2510, new_g26825_ );
dff g2507_reg ( clk, reset, g2507, new_g26822_ );
dff g2504_reg ( clk, reset, g2504, new_g26817_ );
dff g2522_reg ( clk, reset, g2522, new_g27771_ );
dff g2519_reg ( clk, reset, g2519, new_g26827_ );
dff g2516_reg ( clk, reset, g2516, new_g26826_ );
dff g2513_reg ( clk, reset, g2513, new_g26823_ );
dff g2524_reg ( clk, reset, g2524, new_g27769_ );
dff g2523_reg ( clk, reset, g2523, new_g27767_ );
dff g2477_reg ( clk, reset, g2477, new_g26025_ );
dff g2294_reg ( clk, reset, g2294, new_g30260_ );
dff g2291_reg ( clk, reset, g2291, new_g30256_ );
dff g2288_reg ( clk, reset, g2288, new_g30253_ );
dff g2303_reg ( clk, reset, g2303, new_g30665_ );
dff g2300_reg ( clk, reset, g2300, new_g30659_ );
dff g2297_reg ( clk, reset, g2297, new_g30652_ );
dff g2348_reg ( clk, reset, g2348, new_g30694_ );
dff g2345_reg ( clk, reset, g2345, new_g30691_ );
dff g2342_reg ( clk, reset, g2342, new_g30686_ );
dff g2397_reg ( clk, reset, g2397, new_g29182_ );
dff g2391_reg ( clk, reset, g2391, new_g30709_ );
dff g2390_reg ( clk, reset, g2390, new_g30707_ );
dff g2392_reg ( clk, reset, g2392, new_g30566_ );
dff g2267_reg ( clk, reset, g2267, new_g30300_ );
dff g2264_reg ( clk, reset, g2264, new_g30296_ );
dff g2261_reg ( clk, reset, g2261, new_g30289_ );
dff g2393_reg ( clk, reset, g2393, new_g30505_ );
dff g2395_reg ( clk, reset, g2395, new_g30356_ );
dff g2394_reg ( clk, reset, g2394, new_g30341_ );
dff g2389_reg ( clk, reset, g2389, new_g29623_ );
dff g2388_reg ( clk, reset, g2388, new_g29621_ );
dff g2387_reg ( clk, reset, g2387, new_g29618_ );
dff g2312_reg ( clk, reset, g2312, new_g30672_ );
dff g2309_reg ( clk, reset, g2309, new_g30666_ );
dff g2306_reg ( clk, reset, g2306, new_g30660_ );
dff g2276_reg ( clk, reset, g2276, new_g30695_ );
dff g2273_reg ( clk, reset, g2273, new_g30693_ );
dff g2270_reg ( clk, reset, g2270, new_g30690_ );
dff g2321_reg ( clk, reset, g2321, new_g30679_ );
dff g2318_reg ( clk, reset, g2318, new_g30673_ );
dff g2315_reg ( clk, reset, g2315, new_g30667_ );
dff g2285_reg ( clk, reset, g2285, new_g30304_ );
dff g2282_reg ( clk, reset, g2282, new_g30303_ );
dff g2279_reg ( clk, reset, g2279, new_g30301_ );
dff g2330_reg ( clk, reset, g2330, new_g30290_ );
dff g2327_reg ( clk, reset, g2327, new_g30282_ );
dff g2324_reg ( clk, reset, g2324, new_g30274_ );
dff g2339_reg ( clk, reset, g2339, new_g30297_ );
dff g2336_reg ( clk, reset, g2336, new_g30291_ );
dff g2333_reg ( clk, reset, g2333, new_g30283_ );
dff g2396_reg ( clk, reset, g2396, new_g29187_ );
dff g2398_reg ( clk, reset, g2398, new_g29185_ );
dff g2429_reg ( clk, reset, g2429, new_g27276_ );
dff g2436_reg ( clk, reset, g2436, new_g27322_ );
dff g2433_reg ( clk, reset, g2433, new_g27308_ );
dff g2444_reg ( clk, reset, g2444, new_g27292_ );
dff g2451_reg ( clk, reset, g2451, new_g27334_ );
dff g2448_reg ( clk, reset, g2448, new_g27323_ );
dff g2459_reg ( clk, reset, g2459, new_g27309_ );
dff g2466_reg ( clk, reset, g2466, new_g27342_ );
dff g2463_reg ( clk, reset, g2463, new_g27335_ );
dff g2473_reg ( clk, reset, g2473, new_g27324_ );
dff g2421_reg ( clk, reset, g2421, new_g27307_ );
dff g2418_reg ( clk, reset, g2418, new_g27291_ );
dff g2479_reg ( clk, reset, g2479, new_g26676_ );
dff g2478_reg ( clk, reset, g2478, new_g26672_ );
dff g2525_reg ( clk, reset, n6840, n7142 );
dff g2526_reg ( clk, reset, ex_wire27, n6840 );
not U_inv106 ( n7304, ex_wire27 );
dff g2527_reg ( clk, reset, n6849, n7144 );
dff g2528_reg ( clk, reset, ex_wire28, n6849 );
not U_inv107 ( n7302, ex_wire28 );
dff g2529_reg ( clk, reset, n6858, n7149 );
dff g2354_reg ( clk, reset, ex_wire29, n6858 );
not U_inv108 ( n7301, ex_wire29 );
dff g2355_reg ( clk, reset, n6867, n7092 );
dff g2356_reg ( clk, reset, ex_wire30, n6867 );
not U_inv109 ( n7300, ex_wire30 );
dff g2357_reg ( clk, reset, n6876, n7132 );
dff g2358_reg ( clk, reset, ex_wire31, n6876 );
not U_inv110 ( n7299, ex_wire31 );
dff g2359_reg ( clk, reset, n6885, n7128 );
dff g2360_reg ( clk, reset, ex_wire32, n6885 );
not U_inv111 ( n7298, ex_wire32 );
dff g2361_reg ( clk, reset, n6894, n7124 );
dff g2362_reg ( clk, reset, ex_wire33, n6894 );
not U_inv112 ( n7297, ex_wire33 );
dff g2363_reg ( clk, reset, n6903, n7130 );
dff g2364_reg ( clk, reset, ex_wire34, n6903 );
not U_inv113 ( n7296, ex_wire34 );
dff g2374_reg ( clk, reset, ex_wire35, n7088 );
not U_inv114 ( n7287, ex_wire35 );
dff g2373_reg ( clk, reset, g2373, new_g26144_ );
dff g2380_reg ( clk, reset, g2380, new_g30055_ );
dff g2417_reg ( clk, reset, n6986, g2429 );
dff g2424_reg ( clk, reset, g2424, n6986 );
dff g2425_reg ( clk, reset, n6995, g2418 );
dff g2426_reg ( clk, reset, g2426, n6995 );
dff g2427_reg ( clk, reset, n7004, g2421 );
dff g2428_reg ( clk, reset, g2428, n7004 );
dff g2432_reg ( clk, reset, n7013, g2444 );
dff g2439_reg ( clk, reset, g2439, n7013 );
dff g2440_reg ( clk, reset, n7022, g2433 );
dff g2441_reg ( clk, reset, g2441, n7022 );
dff g2442_reg ( clk, reset, n7031, g2436 );
dff g2443_reg ( clk, reset, g2443, n7031 );
dff g2447_reg ( clk, reset, n7040, g2459 );
dff g2454_reg ( clk, reset, g2454, n7040 );
dff g2455_reg ( clk, reset, n7049, g2448 );
dff g2456_reg ( clk, reset, g2456, n7049 );
dff g2457_reg ( clk, reset, n7058, g2451 );
dff g2458_reg ( clk, reset, g2458, n7058 );
dff g2462_reg ( clk, reset, n7067, g2473 );
dff g2469_reg ( clk, reset, g2469, n7067 );
dff g2470_reg ( clk, reset, n7076, g2463 );
dff g2471_reg ( clk, reset, g2471, n7076 );
dff g2472_reg ( clk, reset, n7085, g2466 );
dff g2399_reg ( clk, reset, g2399, n7085 );
dff g2549_reg ( clk, reset, g8087, g2950 );
not U_inv115 ( n7263, g8087 );
dff g2556_reg ( clk, reset, g8167, g8087 );
not U_inv116 ( n7262, g8167 );
dff g2560_reg ( clk, reset, g2560, g8167 );
not U_inv117 ( n7271, g2560 );
dff g2561_reg ( clk, reset, g2561, new_g23114_ );
dff g2562_reg ( clk, reset, g2562, new_g23133_ );
dff g2563_reg ( clk, reset, g2563, new_g21970_ );
dff g2530_reg ( clk, reset, g2530, new_g23407_ );
dff g2638_reg ( clk, reset, n7148, g2530 );
dff g2643_reg ( clk, reset, g2643, n7148 );
dff g2533_reg ( clk, reset, g2533, new_g23418_ );
dff g2644_reg ( clk, reset, n7157, g2533 );
dff g2645_reg ( clk, reset, g2645, n7157 );
dff g2536_reg ( clk, reset, g2536, new_g24209_ );
dff g2646_reg ( clk, reset, n7166, g2536 );
dff g2647_reg ( clk, reset, g2647, n7166 );
dff g2552_reg ( clk, reset, g2552, new_g24214_ );
dff g2553_reg ( clk, reset, g2553, new_g24226_ );
dff g2554_reg ( clk, reset, g2554, new_g24238_ );
dff g2555_reg ( clk, reset, g2555, new_g23132_ );
dff g2559_reg ( clk, reset, g2559, new_g23047_ );
dff g2539_reg ( clk, reset, g2539, new_g23076_ );
dff g2540_reg ( clk, reset, g2540, new_g24225_ );
dff g2648_reg ( clk, reset, n7175, g2540 );
dff g2639_reg ( clk, reset, g2639, n7175 );
dff g2543_reg ( clk, reset, g2543, new_g24237_ );
dff g2640_reg ( clk, reset, n7184, g2543 );
dff g2641_reg ( clk, reset, g2641, n7184 );
dff g2546_reg ( clk, reset, g2546, new_g24250_ );
dff g2642_reg ( clk, reset, n7193, g2546 );
dff g2564_reg ( clk, reset, g2564, n7193 );
dff g2603_reg ( clk, reset, g2603, n7304 );
dff g2604_reg ( clk, reset, g2604, n7302 );
dff g2605_reg ( clk, reset, g2605, n7301 );
dff g2606_reg ( clk, reset, g2606, n7300 );
dff g2607_reg ( clk, reset, g2607, n7299 );
dff g2608_reg ( clk, reset, g2608, n7298 );
dff g2610_reg ( clk, reset, g2610, n7297 );
dff g2611_reg ( clk, reset, g2611, n7296 );
dff g325_reg ( clk, reset, g5629, g3080 );
dff g331_reg ( clk, reset, g5648, g5629 );
dff g337_reg ( clk, reset, g337, g5648 );
dff g1012_reg ( clk, reset, g5657, g3080 );
dff g1018_reg ( clk, reset, g5686, g5657 );
dff g1024_reg ( clk, reset, g1024, g5686 );
dff g1706_reg ( clk, reset, g5695, g3080 );
dff g1712_reg ( clk, reset, g5738, g5695 );
dff g1718_reg ( clk, reset, g1718, g5738 );
dff g2400_reg ( clk, reset, g5747, g3080 );
dff g2406_reg ( clk, reset, g5796, g5747 );
dff g2412_reg ( clk, reset, g2412, g5796 );
dff g558_reg ( clk, reset, n2223, new_g13160_ );
dff g559_reg ( clk, reset, g559, n2223 );
dff g543_reg ( clk, reset, n2200, new_g13149_ );
dff g544_reg ( clk, reset, g544, n2200 );
dff g549_reg ( clk, reset, n2214, new_g13111_ );
dff g506_reg ( clk, reset, ex_wire36, g499 );
not U_inv118 ( n7188, ex_wire36 );
dff g513_reg ( clk, reset, n2032, new_g12487_ );
dff g523_reg ( clk, reset, n2036, n2032 );
dff g524_reg ( clk, reset, g524, n2036 );
dff g528_reg ( clk, reset, n2187, new_g12457_ );
dff g535_reg ( clk, reset, n2191, n2187 );
dff g542_reg ( clk, reset, g542, n2191 );
dff g548_reg ( clk, reset, g548, new_g21851_ );
dff g623_reg ( clk, reset, g6677, g3080 );
not U_inv119 ( n7170, g6677 );
dff g626_reg ( clk, reset, g6911, g6677 );
not U_inv120 ( n7180, g6911 );
dff g629_reg ( clk, reset, g629, g6911 );
not U_inv121 ( n7181, g629 );
dff g1244_reg ( clk, reset, n3924, new_g13171_ );
dff g1245_reg ( clk, reset, g1245, n3924 );
dff g1229_reg ( clk, reset, n3901, new_g13155_ );
dff g1230_reg ( clk, reset, g1230, n3901 );
dff g1235_reg ( clk, reset, n3915, new_g13124_ );
dff g1186_reg ( clk, reset, g1186, n3915 );
not U_inv122 ( n7156, g1186 );
dff g1192_reg ( clk, reset, g1192, g1186 );
dff g1199_reg ( clk, reset, n3733, new_g12507_ );
dff g1209_reg ( clk, reset, n3737, n3733 );
dff g1210_reg ( clk, reset, g1210, n3737 );
dff g1214_reg ( clk, reset, n3888, new_g12467_ );
dff g1221_reg ( clk, reset, n3892, n3888 );
dff g1228_reg ( clk, reset, g1228, n3892 );
dff g1234_reg ( clk, reset, g1234, n241 );
dff g1309_reg ( clk, reset, g6979, g3080 );
not U_inv123 ( n7165, g6979 );
dff g1312_reg ( clk, reset, g7161, g6979 );
not U_inv124 ( n7174, g7161 );
dff g1315_reg ( clk, reset, g1315, g7161 );
not U_inv125 ( n7176, g1315 );
dff g1938_reg ( clk, reset, n5625, new_g13182_ );
dff g1939_reg ( clk, reset, g1939, n5625 );
dff g1923_reg ( clk, reset, n5602, new_g13164_ );
dff g1924_reg ( clk, reset, g1924, n5602 );
dff g1929_reg ( clk, reset, n5616, new_g13135_ );
dff g1880_reg ( clk, reset, g1880, n5616 );
not U_inv126 ( n7182, g1880 );
dff g1886_reg ( clk, reset, g1886, g1880 );
dff g1928_reg ( clk, reset, g1928, n238 );
dff g1893_reg ( clk, reset, n5434, new_g12524_ );
dff g1903_reg ( clk, reset, n5438, n5434 );
dff g1904_reg ( clk, reset, g1904, n5438 );
dff g1908_reg ( clk, reset, n5589, new_g12482_ );
dff g1915_reg ( clk, reset, n5593, n5589 );
dff g1922_reg ( clk, reset, g1922, n5593 );
dff g2003_reg ( clk, reset, g7229, g3080 );
not U_inv127 ( n7164, g7229 );
dff g2006_reg ( clk, reset, g7357, g7229 );
not U_inv128 ( n7173, g7357 );
dff g2009_reg ( clk, reset, g2009, g7357 );
not U_inv129 ( n7177, g2009 );
dff g2632_reg ( clk, reset, n7326, new_g13194_ );
dff g2633_reg ( clk, reset, g2633, n7326 );
dff g2617_reg ( clk, reset, n7303, new_g13175_ );
dff g2618_reg ( clk, reset, g2618, n7303 );
dff g2623_reg ( clk, reset, n7317, new_g13143_ );
dff g2574_reg ( clk, reset, g2574, n7317 );
not U_inv130 ( n7183, g2574 );
dff g2580_reg ( clk, reset, ex_wire37, g2574 );
not U_inv131 ( n7274, ex_wire37 );
dff g2622_reg ( clk, reset, g2622, n235 );
dff g2587_reg ( clk, reset, n7135, new_g12539_ );
dff g2597_reg ( clk, reset, n7139, n7135 );
dff g2598_reg ( clk, reset, g2598, n7139 );
dff g2602_reg ( clk, reset, n7290, new_g12499_ );
dff g2609_reg ( clk, reset, n7294, n7290 );
dff g2616_reg ( clk, reset, g2616, n7294 );
dff g2697_reg ( clk, reset, g7425, g3080 );
not U_inv132 ( n7163, g7425 );
dff g2700_reg ( clk, reset, g7487, g7425 );
not U_inv133 ( n7172, g7487 );
dff g2703_reg ( clk, reset, g2703, g7487 );
not U_inv134 ( n7178, g2703 );
dff g3108_reg ( clk, reset, g3108, new_g30801_ );
dff g3105_reg ( clk, reset, g3105, new_g29941_ );
dff g3102_reg ( clk, reset, g3102, new_g28425_ );
dff g3099_reg ( clk, reset, g3099, new_g25452_ );
dff g3084_reg ( clk, reset, g3084, new_g18782_ );
dff g3088_reg ( clk, reset, g3088, new_g17429_ );
dff g3179_reg ( clk, reset, g3179, new_g17383_ );
dff g3170_reg ( clk, reset, g3170, new_g17340_ );
dff g3161_reg ( clk, reset, g3161, new_g17302_ );
dff g3096_reg ( clk, reset, g3096, new_g17269_ );
dff g3093_reg ( clk, reset, g3093, new_g17246_ );
dff g3087_reg ( clk, reset, g3087, new_g17234_ );
dff g3107_reg ( clk, reset, g3107, new_g30798_ );
dff g3104_reg ( clk, reset, g3104, new_g29939_ );
dff g3101_reg ( clk, reset, g3101, new_g28421_ );
dff g3098_reg ( clk, reset, g3098, new_g25451_ );
dff g3211_reg ( clk, reset, g3211, new_g18719_ );
dff g3185_reg ( clk, reset, g3185, new_g17341_ );
dff g3176_reg ( clk, reset, g3176, new_g17303_ );
dff g3167_reg ( clk, reset, g3167, new_g17270_ );
dff g3158_reg ( clk, reset, g3158, new_g17247_ );
dff g3095_reg ( clk, reset, g3095, new_g17235_ );
dff g3092_reg ( clk, reset, g3092, new_g17228_ );
dff g3086_reg ( clk, reset, g3086, new_g17225_ );
dff g3106_reg ( clk, reset, g3106, new_g30796_ );
dff g3103_reg ( clk, reset, g3103, new_g29936_ );
dff g3100_reg ( clk, reset, g3100, new_g28420_ );
dff g3097_reg ( clk, reset, g3097, new_g25450_ );
not U_inv135 ( n7091, g3097 );
dff g3210_reg ( clk, reset, g3210, new_g18669_ );
dff g3182_reg ( clk, reset, g3182, new_g17271_ );
dff g3173_reg ( clk, reset, g3173, new_g17248_ );
dff g3164_reg ( clk, reset, g3164, new_g17236_ );
dff g3155_reg ( clk, reset, g3155, new_g17229_ );
dff g3094_reg ( clk, reset, g3094, new_g17226_ );
dff g3091_reg ( clk, reset, g3091, new_g17224_ );
dff g3085_reg ( clk, reset, g3085, new_g17222_ );
dff g3054_reg ( clk, reset, g3054, new_g20877_ );
dff g3079_reg ( clk, reset, g3079, new_g20884_ );
dff g3024_reg ( clk, reset, ex_wire38, new_g26786_ );
not U_inv136 ( n7100, ex_wire38 );
dff g2993_reg ( clk, reset, g2993, new_g25265_ );
not U_inv137 ( n7099, g2993 );
dff g2998_reg ( clk, reset, g2998, new_g26048_ );
dff g3006_reg ( clk, reset, g3006, new_g23330_ );
not U_inv138 ( n7097, g3006 );
dff g3002_reg ( clk, reset, g3002, new_g24445_ );
dff g3013_reg ( clk, reset, g3013, new_g25191_ );
not U_inv139 ( n7204, g3013 );
dff g3010_reg ( clk, reset, g3010, new_g26031_ );
not U_inv140 ( n7186, g3010 );
dff g2733_reg ( clk, reset, g2733, new_g20375_ );
dff g2039_reg ( clk, reset, g2039, new_g20353_ );
dff g1345_reg ( clk, reset, g1345, new_g20333_ );
dff g659_reg ( clk, reset, g659, new_g20314_ );
dff g3032_reg ( clk, reset, g3032, new_g25202_ );
dff g3018_reg ( clk, reset, g3018, new_g22002_ );
dff g3028_reg ( clk, reset, g3028, new_g23359_ );
not U_inv141 ( n7240, g3028 );
dff g3036_reg ( clk, reset, g3036, new_g24446_ );
dff g2628_reg ( clk, reset, g2628, new_g21847_ );
dff g2631_reg ( clk, reset, g2631, new_g18780_ );
not U_inv142 ( n7225, g2631 );
dff g2584_reg ( clk, reset, g2584, new_g18820_ );
not U_inv143 ( n7208, g2584 );
dff g2704_reg ( clk, reset, g2704, new_g16718_ );
dff g2714_reg ( clk, reset, g2714, new_g20789_ );
not U_inv144 ( n7254, g2714 );
dff g2707_reg ( clk, reset, g2707, new_g21974_ );
not U_inv145 ( n7199, g2707 );
dff g2727_reg ( clk, reset, g2727, new_g23348_ );
not U_inv146 ( n7194, g2727 );
dff g2720_reg ( clk, reset, g2720, new_g24438_ );
not U_inv147 ( n7279, g2720 );
dff g2734_reg ( clk, reset, g2734, new_g25197_ );
not U_inv148 ( n7219, g2734 );
dff g2746_reg ( clk, reset, g2746, new_g26677_ );
not U_inv149 ( n7280, g2746 );
dff g2740_reg ( clk, reset, g2740, new_g26795_ );
not U_inv150 ( n7234, g2740 );
dff g2753_reg ( clk, reset, g2753, new_g27243_ );
not U_inv151 ( n7275, g2753 );
dff g2760_reg ( clk, reset, g2760, new_g27724_ );
not U_inv152 ( n7249, g2760 );
dff g2766_reg ( clk, reset, g2766, new_g28328_ );
not U_inv153 ( n7258, g2766 );
dff g1934_reg ( clk, reset, g1934, new_g21845_ );
dff g1937_reg ( clk, reset, g1937, new_g18743_ );
not U_inv154 ( n7226, g1937 );
dff g1890_reg ( clk, reset, g1890, new_g18794_ );
not U_inv155 ( n7209, g1890 );
dff g2010_reg ( clk, reset, g2010, new_g16692_ );
dff g2020_reg ( clk, reset, g2020, new_g20752_ );
not U_inv156 ( n7255, g2020 );
dff g2013_reg ( clk, reset, g2013, new_g21972_ );
not U_inv157 ( n7200, g2013 );
dff g2033_reg ( clk, reset, g2033, new_g23339_ );
not U_inv158 ( n7195, g2033 );
dff g2026_reg ( clk, reset, g2026, new_g24434_ );
not U_inv159 ( n7281, g2026 );
dff g2040_reg ( clk, reset, g2040, new_g25194_ );
not U_inv160 ( n7220, g2040 );
dff g2052_reg ( clk, reset, g2052, new_g26671_ );
not U_inv161 ( n7282, g2052 );
dff g2046_reg ( clk, reset, g2046, new_g26789_ );
not U_inv162 ( n7235, g2046 );
dff g2059_reg ( clk, reset, g2059, new_g27682_ );
not U_inv163 ( n7276, g2059 );
dff g2066_reg ( clk, reset, g2066, new_g27722_ );
not U_inv164 ( n7250, g2066 );
dff g2072_reg ( clk, reset, g2072, new_g28325_ );
not U_inv165 ( n7259, g2072 );
dff g1240_reg ( clk, reset, g1240, new_g21843_ );
dff g1243_reg ( clk, reset, g1243, new_g18707_ );
not U_inv166 ( n7227, g1243 );
dff g1196_reg ( clk, reset, g1196, new_g18763_ );
not U_inv167 ( n7207, g1196 );
dff g1316_reg ( clk, reset, g1316, new_g16671_ );
dff g1326_reg ( clk, reset, g1326, new_g20717_ );
not U_inv168 ( n7256, g1326 );
dff g1319_reg ( clk, reset, g1319, new_g21969_ );
not U_inv169 ( n7201, g1319 );
dff g1339_reg ( clk, reset, g1339, new_g23329_ );
not U_inv170 ( n7196, g1339 );
dff g1332_reg ( clk, reset, g1332, new_g24430_ );
not U_inv171 ( n7283, g1332 );
dff g1346_reg ( clk, reset, g1346, new_g25189_ );
not U_inv172 ( n7221, g1346 );
dff g1358_reg ( clk, reset, g1358, new_g26666_ );
not U_inv173 ( n7284, g1358 );
dff g1352_reg ( clk, reset, g1352, new_g26781_ );
not U_inv174 ( n7236, g1352 );
dff g1365_reg ( clk, reset, g1365, new_g27678_ );
not U_inv175 ( n7277, g1365 );
dff g1372_reg ( clk, reset, g1372, new_g27718_ );
not U_inv176 ( n7251, g1372 );
dff g1378_reg ( clk, reset, g1378, new_g28321_ );
not U_inv177 ( n7260, g1378 );
dff g554_reg ( clk, reset, g554, new_g21842_ );
dff g557_reg ( clk, reset, g557, new_g18678_ );
not U_inv178 ( n7224, g557 );
dff g510_reg ( clk, reset, g510, new_g18726_ );
not U_inv179 ( n7205, g510 );
dff g630_reg ( clk, reset, g630, new_g16654_ );
dff g640_reg ( clk, reset, g640, new_g20682_ );
not U_inv180 ( n7257, g640 );
dff g633_reg ( clk, reset, g633, new_g23136_ );
not U_inv181 ( n7203, g633 );
dff g653_reg ( clk, reset, g653, new_g23324_ );
not U_inv182 ( n7197, g653 );
dff g646_reg ( clk, reset, g646, new_g24426_ );
not U_inv183 ( n7285, g646 );
dff g660_reg ( clk, reset, g660, new_g25185_ );
not U_inv184 ( n7222, g660 );
dff g672_reg ( clk, reset, g672, new_g26660_ );
not U_inv185 ( n7286, g672 );
dff g666_reg ( clk, reset, g666, new_g26776_ );
not U_inv186 ( n7237, g666 );
dff g679_reg ( clk, reset, g679, new_g27672_ );
not U_inv187 ( n7278, g679 );
dff g686_reg ( clk, reset, g686, new_g28199_ );
not U_inv188 ( n7252, g686 );
dff g692_reg ( clk, reset, g692, new_g28668_ );
not U_inv189 ( n7261, g692 );
dff g3040_reg ( clk, reset, g5388, g3234 );
dff g2986_reg ( clk, reset, ex_wire39, g5388 );
not U_inv190 ( n7123, ex_wire39 );
dff g2991_reg ( clk, reset, ex_wire40, n7090 );
not U_inv191 ( n7369, ex_wire40 );
dff g3134_reg ( clk, reset, g3134, g26135 );
dff g3147_reg ( clk, reset, g3147, g26135 );
dff g3114_reg ( clk, reset, g3114, g26135 );
dff g3204_reg ( clk, reset, g3204, g26135 );
not U_inv192 ( n7112, g3204 );
dff g3110_reg ( clk, reset, g3110, g25435 );
dff g3197_reg ( clk, reset, g3197, g25435 );
not U_inv193 ( n7108, g3197 );
dff g3111_reg ( clk, reset, g3111, g25442 );
dff g3124_reg ( clk, reset, g3124, g25442 );
dff g3194_reg ( clk, reset, g3194, g25442 );
dff g3112_reg ( clk, reset, g3112, g25420 );
dff g3126_reg ( clk, reset, g3126, g25420 );
dff g3198_reg ( clk, reset, g3198, g25420 );
dff g3123_reg ( clk, reset, g3123, n7043 );
dff g3191_reg ( clk, reset, g3191, g24734 );
dff g3136_reg ( clk, reset, g3136, g26104 );
dff g3142_reg ( clk, reset, g3142, g26104 );
dff g3120_reg ( clk, reset, g3120, g26104 );
dff g3132_reg ( clk, reset, g3132, g26104 );
dff g3207_reg ( clk, reset, g3207, g26104 );
not U_inv194 ( n7109, g3207 );
dff g3135_reg ( clk, reset, g3135, g26149 );
dff g3113_reg ( clk, reset, g3113, g26149 );
dff g3127_reg ( clk, reset, g3127, g26149 );
dff g3201_reg ( clk, reset, g3201, g26149 );
not U_inv195 ( n7110, g3201 );
dff g3139_reg ( clk, reset, g3139, g27380 );
dff g2878_reg ( clk, reset, g2878, new_g21882_ );
dff g2365_reg ( clk, reset, n6912, g2878 );
dff g2366_reg ( clk, reset, ex_wire41, n6912 );
not U_inv196 ( n7291, ex_wire41 );
dff g2615_reg ( clk, reset, g2615, n7291 );
dff g2612_reg ( clk, reset, g2612, new_g24092_ );
dff g2830_reg ( clk, reset, g7519, new_g21878_ );
dff g2873_reg ( clk, reset, g2873, g7519 );
dff g977_reg ( clk, reset, n3510, g2873 );
dff g978_reg ( clk, reset, ex_wire42, n3510 );
not U_inv197 ( n7292, ex_wire42 );
dff g1227_reg ( clk, reset, g1227, n7292 );
dff g1224_reg ( clk, reset, g1224, new_g24072_ );
dff g2877_reg ( clk, reset, g2877, new_g21880_ );
dff g1671_reg ( clk, reset, n5211, g2877 );
dff g1672_reg ( clk, reset, ex_wire43, n5211 );
not U_inv198 ( n7289, ex_wire43 );
dff g1921_reg ( clk, reset, g1921, n7289 );
dff g1918_reg ( clk, reset, g1918, new_g24083_ );
dff g2858_reg ( clk, reset, g8096, new_g20874_ );
dff g2857_reg ( clk, reset, g2857, g8096 );
dff g290_reg ( clk, reset, n1809, g2857 );
dff g291_reg ( clk, reset, ex_wire44, n1809 );
not U_inv199 ( n7288, ex_wire44 );
dff g541_reg ( clk, reset, g541, n7288 );
dff g538_reg ( clk, reset, g538, new_g24059_ );
dff g3151_reg ( clk, reset, g3151, g27380 );
not U_inv200 ( n7121, g3151 );
dff g3188_reg ( clk, reset, g3188, g27380 );
dff g185_reg ( clk, reset, g185, n48 );
not U_inv201 ( n7198, g185 );
dff g2676_reg ( clk, reset, g2676, new_g24557_ );
dff g2673_reg ( clk, reset, g2673, new_g24548_ );
dff g2670_reg ( clk, reset, g2670, new_g24538_ );
dff g2667_reg ( clk, reset, g2667, new_g24547_ );
dff g2664_reg ( clk, reset, g2664, new_g24537_ );
dff g2661_reg ( clk, reset, g2661, new_g24527_ );
dff g2685_reg ( clk, reset, g2685, new_g28367_ );
dff g2682_reg ( clk, reset, g2682, new_g28363_ );
dff g2679_reg ( clk, reset, g2679, new_g28358_ );
dff g2805_reg ( clk, reset, g2805, new_g21063_ );
dff g2807_reg ( clk, reset, g2807, new_g21047_ );
dff g2806_reg ( clk, reset, g2806, new_g21029_ );
dff g2581_reg ( clk, reset, g2581, new_g22687_ );
dff g2650_reg ( clk, reset, g2650, new_g27310_ );
dff g2652_reg ( clk, reset, g2652, new_g27343_ );
dff g2654_reg ( clk, reset, g2654, new_g27337_ );
dff g2653_reg ( clk, reset, g2653, new_g27326_ );
dff g2655_reg ( clk, reset, g2655, new_g27347_ );
dff g2657_reg ( clk, reset, g2657, new_g27344_ );
dff g2656_reg ( clk, reset, g2656, new_g27338_ );
dff g2658_reg ( clk, reset, g2658, new_g27354_ );
dff g2660_reg ( clk, reset, g2660, new_g27348_ );
dff g2659_reg ( clk, reset, g2659, new_g27345_ );
dff g2694_reg ( clk, reset, g2694, new_g28371_ );
dff g2691_reg ( clk, reset, g2691, new_g28368_ );
dff g2688_reg ( clk, reset, g2688, new_g28364_ );
dff g2571_reg ( clk, reset, g2571, new_g26616_ );
dff g2568_reg ( clk, reset, g2568, new_g26596_ );
dff g2565_reg ( clk, reset, g2565, new_g26575_ );
dff g2802_reg ( clk, reset, g2802, new_g21046_ );
dff g2804_reg ( clk, reset, g2804, new_g21028_ );
dff g2803_reg ( clk, reset, g2803, new_g21007_ );
dff g2649_reg ( clk, reset, g2649, new_g27336_ );
dff g2651_reg ( clk, reset, g2651, new_g27325_ );
dff g1982_reg ( clk, reset, g1982, new_g24545_ );
dff g1979_reg ( clk, reset, g1979, new_g24535_ );
dff g1976_reg ( clk, reset, g1976, new_g24525_ );
dff g1991_reg ( clk, reset, g1991, new_g28361_ );
dff g1988_reg ( clk, reset, g1988, new_g28356_ );
dff g1985_reg ( clk, reset, g1985, new_g28352_ );
dff g2111_reg ( clk, reset, g2111, new_g21042_ );
dff g2113_reg ( clk, reset, g2113, new_g21023_ );
dff g2112_reg ( clk, reset, g2112, new_g21003_ );
dff g1887_reg ( clk, reset, ex_wire45, new_g22651_ );
not U_inv202 ( n7248, ex_wire45 );
dff g1956_reg ( clk, reset, g1956, new_g27290_ );
dff g1958_reg ( clk, reset, g1958, new_g27331_ );
dff g1960_reg ( clk, reset, g1960, new_g27320_ );
dff g1959_reg ( clk, reset, g1959, new_g27306_ );
dff g1961_reg ( clk, reset, g1961, new_g27340_ );
dff g1963_reg ( clk, reset, g1963, new_g27332_ );
dff g1962_reg ( clk, reset, g1962, new_g27321_ );
dff g1964_reg ( clk, reset, g1964, new_g27346_ );
dff g1966_reg ( clk, reset, g1966, new_g27341_ );
dff g1965_reg ( clk, reset, g1965, new_g27333_ );
dff g2000_reg ( clk, reset, g2000, new_g28366_ );
dff g1997_reg ( clk, reset, g1997, new_g28362_ );
dff g1994_reg ( clk, reset, g1994, new_g28357_ );
dff g1877_reg ( clk, reset, g1877, new_g26592_ );
dff g1874_reg ( clk, reset, g1874, new_g26573_ );
dff g1871_reg ( clk, reset, g1871, new_g26559_ );
dff g2108_reg ( clk, reset, g2108, new_g21022_ );
dff g2110_reg ( clk, reset, g2110, new_g21002_ );
dff g2109_reg ( clk, reset, g2109, new_g20980_ );
dff g1955_reg ( clk, reset, g1955, new_g27319_ );
dff g1957_reg ( clk, reset, g1957, new_g27305_ );
dff g1973_reg ( clk, reset, g1973, new_g24534_ );
dff g1970_reg ( clk, reset, g1970, new_g24524_ );
dff g1967_reg ( clk, reset, g1967, new_g24513_ );
dff g1288_reg ( clk, reset, g1288, new_g24532_ );
dff g1285_reg ( clk, reset, g1285, new_g24522_ );
dff g1282_reg ( clk, reset, g1282, new_g24511_ );
dff g1297_reg ( clk, reset, g1297, new_g28354_ );
dff g1294_reg ( clk, reset, g1294, new_g28350_ );
dff g1291_reg ( clk, reset, g1291, new_g28346_ );
dff g1417_reg ( clk, reset, g1417, new_g21018_ );
dff g1419_reg ( clk, reset, g1419, new_g20997_ );
dff g1418_reg ( clk, reset, g1418, new_g20976_ );
dff g1193_reg ( clk, reset, ex_wire46, new_g22615_ );
not U_inv203 ( n7229, ex_wire46 );
dff g1262_reg ( clk, reset, g1262, new_g27273_ );
dff g1264_reg ( clk, reset, g1264, new_g27314_ );
dff g1266_reg ( clk, reset, g1266, new_g27300_ );
dff g1265_reg ( clk, reset, g1265, new_g27286_ );
dff g1267_reg ( clk, reset, g1267, new_g27328_ );
dff g1269_reg ( clk, reset, g1269, new_g27315_ );
dff g1268_reg ( clk, reset, g1268, new_g27301_ );
dff g1270_reg ( clk, reset, g1270, new_g27339_ );
dff g1272_reg ( clk, reset, g1272, new_g27329_ );
dff g1271_reg ( clk, reset, g1271, new_g27316_ );
dff g1306_reg ( clk, reset, g1306, new_g28360_ );
dff g1303_reg ( clk, reset, g1303, new_g28355_ );
dff g1300_reg ( clk, reset, g1300, new_g28351_ );
dff g1183_reg ( clk, reset, g1183, new_g26569_ );
dff g1180_reg ( clk, reset, g1180, new_g26557_ );
dff g1177_reg ( clk, reset, g1177, new_g26547_ );
dff g1414_reg ( clk, reset, g1414, new_g20996_ );
dff g1416_reg ( clk, reset, g1416, new_g20975_ );
dff g1415_reg ( clk, reset, g1415, new_g20952_ );
dff g1261_reg ( clk, reset, g1261, new_g27299_ );
dff g1263_reg ( clk, reset, g1263, new_g27285_ );
dff g1279_reg ( clk, reset, g1279, new_g24521_ );
dff g1276_reg ( clk, reset, g1276, new_g24510_ );
dff g1273_reg ( clk, reset, g1273, new_g24501_ );
dff g602_reg ( clk, reset, g602, new_g24519_ );
dff g599_reg ( clk, reset, g599, new_g24508_ );
dff g596_reg ( clk, reset, g596, new_g24499_ );
dff g611_reg ( clk, reset, g611, new_g28348_ );
dff g608_reg ( clk, reset, g608, new_g28344_ );
dff g605_reg ( clk, reset, g605, new_g28342_ );
dff g731_reg ( clk, reset, g731, new_g20992_ );
dff g733_reg ( clk, reset, g733, new_g20970_ );
dff g732_reg ( clk, reset, g732, new_g20948_ );
dff g507_reg ( clk, reset, g507, new_g22578_ );
dff g520_reg ( clk, reset, g16297, n242 );
dff g525_reg ( clk, reset, ex_wire47, g16297 );
not U_inv204 ( n7104, ex_wire47 );
dff g737_reg ( clk, reset, g737, new_g22242_ );
dff g722_reg ( clk, reset, g722, new_g21051_ );
dff g719_reg ( clk, reset, g719, new_g21031_ );
dff g716_reg ( clk, reset, g716, new_g21009_ );
dff g713_reg ( clk, reset, g713, new_g20989_ );
dff g710_reg ( clk, reset, g710, new_g20966_ );
dff g707_reg ( clk, reset, g707, new_g20944_ );
dff g704_reg ( clk, reset, g704, new_g20921_ );
dff g701_reg ( clk, reset, g701, new_g20901_ );
dff g725_reg ( clk, reset, g725, new_g20894_ );
dff g698_reg ( clk, reset, g698, new_g20891_ );
dff g739_reg ( clk, reset, g739, new_g22231_ );
dff g724_reg ( clk, reset, g724, new_g21032_ );
dff g721_reg ( clk, reset, g721, new_g21010_ );
dff g718_reg ( clk, reset, g718, new_g20990_ );
dff g715_reg ( clk, reset, g715, new_g20967_ );
dff g712_reg ( clk, reset, g712, new_g20945_ );
dff g709_reg ( clk, reset, g709, new_g20922_ );
dff g706_reg ( clk, reset, g706, new_g20902_ );
dff g703_reg ( clk, reset, g703, new_g20892_ );
dff g727_reg ( clk, reset, g727, new_g20881_ );
dff g700_reg ( clk, reset, g700, new_g20879_ );
dff g738_reg ( clk, reset, g738, new_g22218_ );
dff g723_reg ( clk, reset, g723, new_g21011_ );
dff g720_reg ( clk, reset, g720, new_g20991_ );
dff g717_reg ( clk, reset, g717, new_g20968_ );
dff g714_reg ( clk, reset, g714, new_g20946_ );
dff g711_reg ( clk, reset, g711, new_g20923_ );
dff g708_reg ( clk, reset, g708, new_g20903_ );
dff g705_reg ( clk, reset, g705, new_g20893_ );
dff g702_reg ( clk, reset, g702, new_g20880_ );
dff g726_reg ( clk, reset, g726, new_g20876_ );
dff g699_reg ( clk, reset, g699, new_g20875_ );
dff g1206_reg ( clk, reset, g16355, n243 );
dff g1211_reg ( clk, reset, ex_wire48, g16355 );
not U_inv205 ( n7103, ex_wire48 );
dff g1423_reg ( clk, reset, g1423, new_g22263_ );
dff g1408_reg ( clk, reset, g1408, new_g21070_ );
dff g1405_reg ( clk, reset, g1405, new_g21052_ );
dff g1402_reg ( clk, reset, g1402, new_g21033_ );
dff g1399_reg ( clk, reset, g1399, new_g21015_ );
dff g1396_reg ( clk, reset, g1396, new_g20993_ );
dff g1393_reg ( clk, reset, g1393, new_g20972_ );
dff g1390_reg ( clk, reset, g1390, new_g20949_ );
dff g1387_reg ( clk, reset, g1387, new_g20925_ );
dff g1411_reg ( clk, reset, g1411, new_g20913_ );
dff g1384_reg ( clk, reset, g1384, new_g20910_ );
dff g1425_reg ( clk, reset, g1425, new_g22247_ );
dff g1410_reg ( clk, reset, g1410, new_g21053_ );
dff g1407_reg ( clk, reset, g1407, new_g21034_ );
dff g1404_reg ( clk, reset, g1404, new_g21016_ );
dff g1401_reg ( clk, reset, g1401, new_g20994_ );
dff g1398_reg ( clk, reset, g1398, new_g20973_ );
dff g1395_reg ( clk, reset, g1395, new_g20950_ );
dff g1392_reg ( clk, reset, g1392, new_g20926_ );
dff g1389_reg ( clk, reset, g1389, new_g20911_ );
dff g1413_reg ( clk, reset, g1413, new_g20898_ );
dff g1386_reg ( clk, reset, g1386, new_g20896_ );
dff g1424_reg ( clk, reset, g1424, new_g22234_ );
dff g1409_reg ( clk, reset, g1409, new_g21035_ );
dff g1406_reg ( clk, reset, g1406, new_g21017_ );
dff g1403_reg ( clk, reset, g1403, new_g20995_ );
dff g1400_reg ( clk, reset, g1400, new_g20974_ );
dff g1397_reg ( clk, reset, g1397, new_g20951_ );
dff g1394_reg ( clk, reset, g1394, new_g20927_ );
dff g1391_reg ( clk, reset, g1391, new_g20912_ );
dff g1388_reg ( clk, reset, g1388, new_g20897_ );
dff g1412_reg ( clk, reset, g1412, new_g20883_ );
dff g1385_reg ( clk, reset, g1385, new_g20882_ );
dff g1420_reg ( clk, reset, g1420, new_g25270_ );
dff g1422_reg ( clk, reset, g1422, new_g25267_ );
dff g1421_reg ( clk, reset, g1421, new_g25263_ );
dff g3061_reg ( clk, reset, g3061, n7055 );
dff g3059_reg ( clk, reset, g3059, n7059 );
dff g3056_reg ( clk, reset, g3056, n7057 );
dff g3052_reg ( clk, reset, g3052, n7060 );
dff g3055_reg ( clk, reset, g3055, n7061 );
dff g3053_reg ( clk, reset, g3053, n7063 );
dff g3057_reg ( clk, reset, g3057, n7056 );
dff g3058_reg ( clk, reset, g3058, n7062 );
dff g3060_reg ( clk, reset, g3060, n7064 );
dff g1900_reg ( clk, reset, g16399, new_g28990_ );
dff g1905_reg ( clk, reset, ex_wire49, g16399 );
not U_inv206 ( n7102, ex_wire49 );
dff g2117_reg ( clk, reset, g2117, new_g22280_ );
dff g2102_reg ( clk, reset, g2102, new_g21080_ );
dff g2099_reg ( clk, reset, g2099, new_g21071_ );
dff g2096_reg ( clk, reset, g2096, new_g21054_ );
dff g2093_reg ( clk, reset, g2093, new_g21039_ );
dff g2090_reg ( clk, reset, g2090, new_g21019_ );
dff g2087_reg ( clk, reset, g2087, new_g20999_ );
dff g2084_reg ( clk, reset, g2084, new_g20977_ );
dff g2081_reg ( clk, reset, g2081, new_g20953_ );
dff g2105_reg ( clk, reset, g2105, new_g20937_ );
dff g2078_reg ( clk, reset, g2078, new_g20934_ );
dff g2119_reg ( clk, reset, g2119, new_g22267_ );
dff g2104_reg ( clk, reset, g2104, new_g21072_ );
dff g2101_reg ( clk, reset, g2101, new_g21055_ );
dff g2098_reg ( clk, reset, g2098, new_g21040_ );
dff g2095_reg ( clk, reset, g2095, new_g21020_ );
dff g2092_reg ( clk, reset, g2092, new_g21000_ );
dff g2089_reg ( clk, reset, g2089, new_g20978_ );
dff g2086_reg ( clk, reset, g2086, new_g20954_ );
dff g2083_reg ( clk, reset, g2083, new_g20935_ );
dff g2107_reg ( clk, reset, g2107, new_g20917_ );
dff g2080_reg ( clk, reset, g2080, new_g20915_ );
dff g2118_reg ( clk, reset, g2118, new_g22249_ );
dff g2103_reg ( clk, reset, g2103, new_g21056_ );
dff g2100_reg ( clk, reset, g2100, new_g21041_ );
dff g2097_reg ( clk, reset, g2097, new_g21021_ );
dff g2094_reg ( clk, reset, g2094, new_g21001_ );
dff g2091_reg ( clk, reset, g2091, new_g20979_ );
dff g2088_reg ( clk, reset, g2088, new_g20955_ );
dff g2085_reg ( clk, reset, g2085, new_g20936_ );
dff g2082_reg ( clk, reset, g2082, new_g20916_ );
dff g2106_reg ( clk, reset, g2106, new_g20900_ );
dff g2079_reg ( clk, reset, g2079, new_g20899_ );
dff g2114_reg ( clk, reset, g2114, new_g25279_ );
dff g2116_reg ( clk, reset, g2116, new_g25271_ );
dff g2115_reg ( clk, reset, g2115, new_g25268_ );
dff g3070_reg ( clk, reset, g3070, n7065 );
dff g3068_reg ( clk, reset, g3068, n7069 );
dff g3065_reg ( clk, reset, g3065, n7068 );
dff g3062_reg ( clk, reset, g3062, n7070 );
dff g3064_reg ( clk, reset, g3064, n7071 );
dff g3063_reg ( clk, reset, g3063, n7073 );
dff g3066_reg ( clk, reset, g3066, n7066 );
dff g3067_reg ( clk, reset, g3067, n7072 );
dff g3069_reg ( clk, reset, g3069, n7074 );
dff g2594_reg ( clk, reset, g16437, new_g30061_ );
dff g2599_reg ( clk, reset, ex_wire50, g16437 );
not U_inv207 ( n7101, ex_wire50 );
dff g2811_reg ( clk, reset, g2811, new_g22299_ );
dff g2796_reg ( clk, reset, g2796, new_g21094_ );
dff g2793_reg ( clk, reset, g2793, new_g21081_ );
dff g2790_reg ( clk, reset, g2790, new_g21073_ );
dff g2787_reg ( clk, reset, g2787, new_g21060_ );
dff g2784_reg ( clk, reset, g2784, new_g21043_ );
dff g2781_reg ( clk, reset, g2781, new_g21025_ );
dff g2778_reg ( clk, reset, g2778, new_g21004_ );
dff g2775_reg ( clk, reset, g2775, new_g20981_ );
dff g2799_reg ( clk, reset, g2799, new_g20965_ );
dff g2772_reg ( clk, reset, g2772, new_g20962_ );
dff g2813_reg ( clk, reset, g2813, new_g22284_ );
dff g2798_reg ( clk, reset, g2798, new_g21082_ );
dff g2795_reg ( clk, reset, g2795, new_g21074_ );
dff g2792_reg ( clk, reset, g2792, new_g21061_ );
dff g2789_reg ( clk, reset, g2789, new_g21044_ );
dff g2786_reg ( clk, reset, g2786, new_g21026_ );
dff g2783_reg ( clk, reset, g2783, new_g21005_ );
dff g2780_reg ( clk, reset, g2780, new_g20982_ );
dff g2777_reg ( clk, reset, g2777, new_g20963_ );
dff g2801_reg ( clk, reset, g2801, new_g20941_ );
dff g2774_reg ( clk, reset, g2774, new_g20939_ );
dff g2812_reg ( clk, reset, g2812, new_g22269_ );
dff g2797_reg ( clk, reset, g2797, new_g21075_ );
dff g2794_reg ( clk, reset, g2794, new_g21062_ );
dff g2791_reg ( clk, reset, g2791, new_g21045_ );
dff g2788_reg ( clk, reset, g2788, new_g21027_ );
dff g2785_reg ( clk, reset, g2785, new_g21006_ );
dff g2782_reg ( clk, reset, g2782, new_g20983_ );
dff g2779_reg ( clk, reset, g2779, new_g20964_ );
dff g2776_reg ( clk, reset, g2776, new_g20940_ );
dff g2800_reg ( clk, reset, g2800, new_g20919_ );
dff g2773_reg ( clk, reset, g2773, new_g20918_ );
dff g2808_reg ( clk, reset, g2808, new_g25288_ );
dff g2810_reg ( clk, reset, g2810, new_g25280_ );
dff g2809_reg ( clk, reset, g2809, new_g25272_ );
dff g2997_reg ( clk, reset, g2997, n7075 );
dff g2990_reg ( clk, reset, g2990, new_g18907_ );
dff g3077_reg ( clk, reset, g3077, n7079 );
dff g8_reg ( clk, reset, g8261, new_g18837_ );
dff g3074_reg ( clk, reset, g3074, n7078 );
dff g11_reg ( clk, reset, g8262, new_g16880_ );
dff g3071_reg ( clk, reset, g3071, n7080 );
dff g23_reg ( clk, reset, g8266, new_g16845_ );
dff g3073_reg ( clk, reset, g3073, n7081 );
dff g17_reg ( clk, reset, g8264, new_g16861_ );
dff g3072_reg ( clk, reset, g3072, n7083 );
dff g20_reg ( clk, reset, g8265, new_g16854_ );
dff g3075_reg ( clk, reset, g3075, n7077 );
dff g14_reg ( clk, reset, g8263, new_g18755_ );
dff g3076_reg ( clk, reset, g3076, n7082 );
dff g5_reg ( clk, reset, g8260, new_g18804_ );
dff g3078_reg ( clk, reset, g3078, n7084 );
dff g2_reg ( clk, reset, g8259, new_g18868_ );
dff g576_reg ( clk, reset, g576, new_g27261_ );
dff g578_reg ( clk, reset, g578, new_g27294_ );
dff g580_reg ( clk, reset, g580, new_g27280_ );
dff g579_reg ( clk, reset, g579, new_g27269_ );
dff g581_reg ( clk, reset, g581, new_g27311_ );
dff g583_reg ( clk, reset, g583, new_g27295_ );
dff g582_reg ( clk, reset, g582, new_g27281_ );
dff g584_reg ( clk, reset, g584, new_g27327_ );
dff g586_reg ( clk, reset, g586, new_g27312_ );
dff g585_reg ( clk, reset, g585, new_g27296_ );
dff g620_reg ( clk, reset, g620, new_g28353_ );
dff g617_reg ( clk, reset, g617, new_g28349_ );
dff g614_reg ( clk, reset, g614, new_g28345_ );
dff g496_reg ( clk, reset, g496, new_g26553_ );
dff g493_reg ( clk, reset, g493, new_g26545_ );
dff g490_reg ( clk, reset, g490, new_g26541_ );
dff g728_reg ( clk, reset, g728, new_g20969_ );
dff g730_reg ( clk, reset, g730, new_g20947_ );
dff g729_reg ( clk, reset, g729, new_g20924_ );
dff g734_reg ( clk, reset, g734, new_g25266_ );
dff g736_reg ( clk, reset, g736, new_g25262_ );
dff g735_reg ( clk, reset, g735, new_g25260_ );
dff g3046_reg ( clk, reset, g3046, n7048 );
dff g39_reg ( clk, reset, g8272, new_g16860_ );
dff g3050_reg ( clk, reset, g3050, n7046 );
dff g36_reg ( clk, reset, g8271, new_g16857_ );
dff g3048_reg ( clk, reset, g3048, n7047 );
dff g30_reg ( clk, reset, g8269, new_g16835_ );
dff g3044_reg ( clk, reset, g3044, n7050 );
dff g45_reg ( clk, reset, g8274, new_g16844_ );
dff g575_reg ( clk, reset, g575, new_g27279_ );
dff g577_reg ( clk, reset, g577, new_g27268_ );
dff g3045_reg ( clk, reset, g3045, n7053 );
dff g42_reg ( clk, reset, g8273, new_g16853_ );
dff g3043_reg ( clk, reset, g3043, n7054 );
dff g48_reg ( clk, reset, g8275, new_g16824_ );
dff g3049_reg ( clk, reset, g3049, n7051 );
dff g33_reg ( clk, reset, g8270, new_g16851_ );
dff g3051_reg ( clk, reset, g3051, n7045 );
dff g3083_reg ( clk, reset, g3083, new_g16866_ );
dff g3047_reg ( clk, reset, g3047, n7052 );
dff g27_reg ( clk, reset, g8268, new_g16803_ );
dff g26_reg ( clk, reset, g8267, new_g16566_ );
dff g2992_reg ( clk, reset, ex_wire51, n7089 );
not U_inv208 ( n7370, ex_wire51 );
dff g593_reg ( clk, reset, g593, new_g24507_ );
dff g590_reg ( clk, reset, g590, new_g24498_ );
dff g587_reg ( clk, reset, g587, new_g24491_ );
dff g3133_reg ( clk, reset, g3133, n48 );
dff g3125_reg ( clk, reset, g3125, n147 );
dff g3128_reg ( clk, reset, g3128, n143 );
dff g1_reg ( clk, reset, g8258, new_g18542_ );
dff g3109_reg ( clk, reset, g3109, g8030 );
not U_inv209 ( n7245, g3109 );
dff g2950_reg ( clk, reset, g2950, new_g19152_ );
not U_inv210 ( n7253, g2950 );
dff g3080_reg ( clk, reset, g3080, new_g20497_ );
not U_inv211 ( n7187, g3080 );
dff g3129_reg ( clk, reset, g8106, g3080 );
not U_inv212 ( n7242, g8106 );
dff g3117_reg ( clk, reset, g8030, g8106 );
not U_inv213 ( n7243, g8030 );
dff g2625_reg ( clk, reset, g7390, g7302 );
not U_inv214 ( n7161, g7390 );
dff g1237_reg ( clk, reset, g6944, g6750 );
not U_inv215 ( n7159, g6944 );
dff g1931_reg ( clk, reset, g7194, g7052 );
not U_inv216 ( n7158, g7194 );
dff g2619_reg ( clk, reset, g7302, g3080 );
not U_inv217 ( n7160, g7302 );
dff g1925_reg ( clk, reset, g7052, g3080 );
not U_inv218 ( n7155, g7052 );
dff g499_reg ( clk, reset, g499, n2214 );
not U_inv219 ( n7185, g499 );
dff g401_reg ( clk, reset, g401, g6447 );
dff g1088_reg ( clk, reset, g1088, g6712 );
dff g1782_reg ( clk, reset, g1782, g7014 );
dff g2476_reg ( clk, reset, g2476, g7264 );
dff g1786_reg ( clk, reset, g7014, g5511 );
dff g405_reg ( clk, reset, g6447, g5437 );
dff g276_reg ( clk, reset, g5437, g2950 );
dff g963_reg ( clk, reset, g5472, g2950 );
dff g1657_reg ( clk, reset, g5511, g2950 );
dff g2351_reg ( clk, reset, g5555, g2950 );
dff g2987_reg ( clk, reset, g2987, g16496 );
not U_inv220 ( n7239, g2987 );
dff g2624_reg ( clk, reset, g2624, g7390 );
not U_inv221 ( n7179, g2624 );
dff g551_reg ( clk, reset, g6642, g6485 );
not U_inv222 ( n7171, g6642 );
dff g550_reg ( clk, reset, g550, g6642 );
not U_inv223 ( n7169, g550 );
dff g1930_reg ( clk, reset, g1930, g7194 );
not U_inv224 ( n7168, g1930 );
dff g1236_reg ( clk, reset, g1236, g6944 );
not U_inv225 ( n7167, g1236 );
dff g545_reg ( clk, reset, g6485, g3080 );
not U_inv226 ( n7162, g6485 );
dff g1231_reg ( clk, reset, g6750, g3080 );
not U_inv227 ( n7122, g6750 );
dff g1092_reg ( clk, reset, g6712, g5472 );
dff g2480_reg ( clk, reset, g7264, g5555 );
buf U7973 ( n7477, n7476 );
buf U7974 ( n7483, n7482 );
buf U7975 ( n7489, n7488 );
buf U7976 ( n7495, n7494 );
buf U7977 ( n7474, n7473 );
buf U7978 ( n7480, n7479 );
buf U7979 ( n7486, n7485 );
buf U7980 ( n7492, n7491 );
buf U7981 ( n7500, n7497 );
buf U7982 ( n7499, n7497 );
nor U7983 ( n6238, n6315, n7185 );
not U7984 ( n7501, g3229 );
nand U7985 ( n2272, n5481, n5482 );
not U7986 ( n125, n971 );
not U7987 ( n59, n1012 );
not U7988 ( n81, n1048 );
not U7989 ( n103, n1073 );
not U7990 ( n529, n937 );
not U7991 ( n418, n981 );
not U7992 ( n309, n1022 );
not U7993 ( n188, n1059 );
not U7994 ( n126, n939 );
not U7995 ( n60, n983 );
not U7996 ( n82, n1024 );
not U7997 ( n104, n1061 );
nor U7998 ( n971, n126, n783 );
nor U7999 ( n1012, n60, n816 );
nor U8000 ( n1048, n82, n852 );
nor U8001 ( n1073, n104, n890 );
nor U8002 ( n806, n939, n531 );
nor U8003 ( n842, n983, n420 );
nor U8004 ( n880, n1024, n311 );
nor U8005 ( n926, n1061, n190 );
nor U8006 ( n786, n939, n972 );
nor U8007 ( n819, n983, n1013 );
nor U8008 ( n855, n1024, n1049 );
nor U8009 ( n893, n1061, n1074 );
nand U8010 ( n1821, n505, n499 );
nand U8011 ( n1885, n397, n391 );
nand U8012 ( n1956, n288, n282 );
nand U8013 ( n2021, n167, n161 );
not U8014 ( n531, n972 );
not U8015 ( n420, n1013 );
not U8016 ( n311, n1049 );
not U8017 ( n190, n1074 );
nand U8018 ( n937, n531, n530 );
nand U8019 ( n981, n420, n419 );
nand U8020 ( n1022, n311, n310 );
nand U8021 ( n1059, n190, n189 );
not U8022 ( n118, n2079 );
not U8023 ( n52, n2124 );
not U8024 ( n74, n2165 );
not U8025 ( n96, n2205 );
not U8026 ( n119, n1677 );
not U8027 ( n53, n1699 );
not U8028 ( n75, n1721 );
not U8029 ( n97, n1741 );
nand U8030 ( n935, n936, n937 );
nand U8031 ( n1020, n1021, n1022 );
nand U8032 ( n1056, n1057, n1059 );
nand U8033 ( n979, n980, n981 );
nor U8034 ( n6878, n579, n6797 );
nor U8035 ( n6682, n463, n6606 );
nor U8036 ( n6487, n354, n6411 );
not U8037 ( n528, n1437 );
not U8038 ( n308, n1529 );
not U8039 ( n187, n1570 );
not U8040 ( n417, n1482 );
not U8041 ( n527, n3141 );
not U8042 ( n307, n3298 );
not U8043 ( n416, n3230 );
not U8044 ( n186, n3330 );
not U8045 ( n27, n2033 );
not U8046 ( n25, n2039 );
not U8047 ( n23, n2044 );
not U8048 ( n29, n2027 );
nand U8049 ( n939, n1414, n1415 );
nor U8050 ( n1414, n529, n1416 );
and U8051 ( n1416, n1417, n1418 );
nand U8052 ( n983, n1458, n1459 );
nor U8053 ( n1458, n418, n1460 );
and U8054 ( n1460, n1461, n1462 );
nand U8055 ( n1024, n1506, n1507 );
nor U8056 ( n1506, n309, n1508 );
and U8057 ( n1508, n1509, n1510 );
nand U8058 ( n1061, n1547, n1548 );
nor U8059 ( n1547, n188, n1549 );
and U8060 ( n1549, n1550, n1551 );
nand U8061 ( n726, n1903, n84 );
and U8062 ( n1903, n725, n729 );
nand U8063 ( n759, n1968, n106 );
and U8064 ( n1968, n758, n762 );
nor U8065 ( n1936, n1938, n1939 );
nand U8066 ( n1939, n1940, n1941 );
nand U8067 ( n1941, n1934, n1942 );
nand U8068 ( n1940, n282, n1933 );
nor U8069 ( n2002, n2003, n2005 );
nand U8070 ( n2005, n2006, n2007 );
nand U8071 ( n2007, n2000, n2009 );
nand U8072 ( n2006, n161, n1999 );
nor U8073 ( n970, n510, n125 );
nor U8074 ( n1011, n401, n59 );
nor U8075 ( n1047, n292, n81 );
nor U8076 ( n1072, n171, n103 );
not U8077 ( n499, n1796 );
not U8078 ( n391, n1861 );
not U8079 ( n282, n1930 );
not U8080 ( n161, n1996 );
nor U8081 ( n1803, n1804, n1805 );
nand U8082 ( n1805, n1806, n1807 );
nand U8083 ( n1807, n1801, n1808 );
nand U8084 ( n1806, n499, n1799 );
nor U8085 ( n1867, n1868, n1869 );
nand U8086 ( n1869, n1870, n1871 );
nand U8087 ( n1871, n1865, n1872 );
nand U8088 ( n1870, n391, n1864 );
nand U8089 ( n1100, n1769, n128 );
and U8090 ( n1769, n1099, n1103 );
nand U8091 ( n688, n1837, n62 );
and U8092 ( n1837, n687, n691 );
nor U8093 ( n1802, n1801, n1810 );
nand U8094 ( n1810, n1811, n1812 );
nand U8095 ( n1812, n1799, n1804 );
nand U8096 ( n1811, n499, n1808 );
nor U8097 ( n1866, n1865, n1873 );
nand U8098 ( n1873, n1874, n1875 );
nand U8099 ( n1875, n1864, n1868 );
nand U8100 ( n1874, n391, n1872 );
nor U8101 ( n1935, n1934, n1943 );
nand U8102 ( n1943, n1944, n1945 );
nand U8103 ( n1945, n1933, n1938 );
nand U8104 ( n1944, n282, n1942 );
nor U8105 ( n2001, n2000, n2010 );
nand U8106 ( n2010, n2011, n2012 );
nand U8107 ( n2012, n1999, n2003 );
nand U8108 ( n2011, n161, n2009 );
and U8109 ( n783, n1415, n1420 );
nand U8110 ( n1420, n1421, n937 );
nand U8111 ( n1421, n1418, n1422 );
or U8112 ( n1422, n1417, n972 );
and U8113 ( n816, n1459, n1464 );
nand U8114 ( n1464, n1465, n981 );
nand U8115 ( n1465, n1462, n1466 );
or U8116 ( n1466, n1461, n1013 );
and U8117 ( n852, n1507, n1512 );
nand U8118 ( n1512, n1513, n1022 );
nand U8119 ( n1513, n1510, n1514 );
or U8120 ( n1514, n1509, n1049 );
and U8121 ( n890, n1548, n1553 );
nand U8122 ( n1553, n1554, n1059 );
nand U8123 ( n1554, n1551, n1555 );
or U8124 ( n1555, n1550, n1074 );
nor U8125 ( n1784, n1781, n1785 );
nand U8126 ( n1785, n1786, n1787 );
nand U8127 ( n1787, n1780, n1779 );
nand U8128 ( n1786, n505, n1778 );
nor U8129 ( n1850, n1848, n1851 );
nand U8130 ( n1851, n1852, n1853 );
nand U8131 ( n1853, n1847, n1846 );
nand U8132 ( n1852, n397, n1845 );
nor U8133 ( n1917, n1915, n1918 );
nand U8134 ( n1918, n1920, n1921 );
nand U8135 ( n1921, n1914, n1913 );
nand U8136 ( n1920, n288, n1912 );
nor U8137 ( n1983, n1980, n1984 );
nand U8138 ( n1984, n1985, n1986 );
nand U8139 ( n1986, n1979, n1978 );
nand U8140 ( n1985, n167, n1977 );
not U8141 ( n505, n1775 );
not U8142 ( n397, n1842 );
not U8143 ( n288, n1908 );
not U8144 ( n167, n1974 );
nor U8145 ( n1783, n1779, n1788 );
nand U8146 ( n1788, n1789, n1790 );
nand U8147 ( n1790, n1781, n1778 );
nand U8148 ( n1789, n505, n1780 );
nor U8149 ( n1849, n1846, n1854 );
nand U8150 ( n1854, n1855, n1856 );
nand U8151 ( n1856, n1848, n1845 );
nand U8152 ( n1855, n397, n1847 );
nor U8153 ( n1916, n1913, n1922 );
nand U8154 ( n1922, n1923, n1924 );
nand U8155 ( n1924, n1915, n1912 );
nand U8156 ( n1923, n288, n1914 );
nor U8157 ( n1981, n1978, n1987 );
nand U8158 ( n1987, n1988, n1989 );
nand U8159 ( n1989, n1980, n1977 );
nand U8160 ( n1988, n167, n1979 );
not U8161 ( n128, n1094 );
not U8162 ( n62, n682 );
not U8163 ( n84, n720 );
not U8164 ( n106, n753 );
nand U8165 ( n1095, n1098, n1099 );
or U8166 ( n1098, n1100, n541 );
nand U8167 ( n683, n686, n687 );
or U8168 ( n686, n688, n429 );
nand U8169 ( n721, n724, n725 );
or U8170 ( n724, n726, n320 );
nand U8171 ( n754, n757, n758 );
or U8172 ( n757, n759, n199 );
nand U8173 ( n711, n712, n313 );
nor U8174 ( n712, n713, n714 );
nor U8175 ( n714, n716, n717 );
nor U8176 ( n713, n721, n722 );
nand U8177 ( n746, n747, n192 );
nor U8178 ( n747, n748, n749 );
nor U8179 ( n749, n750, n751 );
nor U8180 ( n748, n754, n755 );
nand U8181 ( n1087, n1088, n533 );
nor U8182 ( n1088, n1089, n1090 );
nor U8183 ( n1090, n1091, n1092 );
nor U8184 ( n1089, n1095, n1096 );
nand U8185 ( n675, n676, n422 );
nor U8186 ( n676, n677, n678 );
nor U8187 ( n678, n679, n680 );
nor U8188 ( n677, n683, n684 );
nand U8189 ( n1096, n532, n1097 );
nand U8190 ( n684, n421, n685 );
nand U8191 ( n722, n312, n723 );
nand U8192 ( n755, n191, n756 );
nand U8193 ( n1179, n1816, n1817 );
nor U8194 ( n1817, n1818, n1819 );
nor U8195 ( n1816, n1820, n1821 );
nand U8196 ( n1819, n1778, n1801 );
nand U8197 ( n1197, n1879, n1880 );
nor U8198 ( n1880, n1881, n1882 );
nor U8199 ( n1879, n1884, n1885 );
nand U8200 ( n1882, n1845, n1865 );
nand U8201 ( n1139, n1950, n1951 );
nor U8202 ( n1951, n1952, n1953 );
nor U8203 ( n1950, n1954, n1956 );
nand U8204 ( n1953, n1912, n1934 );
nand U8205 ( n1159, n2016, n2017 );
nor U8206 ( n2017, n2018, n2019 );
nor U8207 ( n2016, n2020, n2021 );
nand U8208 ( n2019, n1977, n2000 );
nor U8209 ( n728, n730, n731 );
nand U8210 ( n731, n312, n725 );
nor U8211 ( n761, n763, n764 );
nand U8212 ( n764, n191, n758 );
nor U8213 ( n1102, n1104, n1105 );
nand U8214 ( n1105, n532, n1099 );
nor U8215 ( n690, n692, n693 );
nand U8216 ( n693, n421, n687 );
nand U8217 ( n1174, n1103, n1099 );
nand U8218 ( n1192, n691, n687 );
nand U8219 ( n1134, n729, n725 );
nand U8220 ( n1154, n762, n758 );
and U8221 ( n1108, n1164, n129 );
xor U8222 ( n1164, n1165, n532 );
nand U8223 ( n1165, n1166, n1167 );
nand U8224 ( n1166, n1168, n1169 );
and U8225 ( n1111, n1182, n63 );
xor U8226 ( n1182, n1183, n421 );
nand U8227 ( n1183, n1184, n1185 );
nand U8228 ( n1184, n1186, n1187 );
and U8229 ( n1114, n1124, n85 );
xor U8230 ( n1124, n1125, n312 );
nand U8231 ( n1125, n1126, n1127 );
nand U8232 ( n1126, n1128, n1129 );
and U8233 ( n1121, n1144, n107 );
xor U8234 ( n1144, n1145, n191 );
nand U8235 ( n1145, n1146, n1147 );
nand U8236 ( n1146, n1148, n1149 );
nor U8237 ( n1091, n541, n1094 );
nor U8238 ( n679, n429, n682 );
nor U8239 ( n716, n320, n720 );
nor U8240 ( n750, n199, n753 );
not U8241 ( n131, n1103 );
not U8242 ( n87, n729 );
not U8243 ( n230, n3105 );
not U8244 ( n349, n3017 );
not U8245 ( n458, n2930 );
not U8246 ( n574, n2875 );
not U8247 ( n65, n691 );
not U8248 ( n109, n762 );
nand U8249 ( n2908, n2627, n230 );
nand U8250 ( n2870, n2523, n349 );
nand U8251 ( n2848, n2411, n458 );
nand U8252 ( n2838, n2299, n574 );
nor U8253 ( n3243, g3229, n3189 );
nor U8254 ( n3154, g3229, n3086 );
nor U8255 ( n3053, g3229, n2998 );
nor U8256 ( n2965, g3229, n2911 );
nor U8257 ( n3122, g3229, n3043 );
nor U8258 ( n3211, g3229, n3144 );
nor U8259 ( n3279, g3229, n3233 );
nor U8260 ( n3311, g3229, n3301 );
and U8261 ( n1829, n1899, n1900 );
nand U8262 ( n1899, n308, n84 );
nand U8263 ( n1900, n1902, n312 );
nor U8264 ( n1902, n314, n726 );
and U8265 ( n1751, n1766, n1767 );
nand U8266 ( n1766, n528, n128 );
nand U8267 ( n1767, n1768, n532 );
nor U8268 ( n1768, n534, n1100 );
and U8269 ( n1760, n1834, n1835 );
nand U8270 ( n1834, n417, n62 );
nand U8271 ( n1835, n1836, n421 );
nor U8272 ( n1836, n423, n688 );
and U8273 ( n1894, n1965, n1966 );
nand U8274 ( n1965, n187, n106 );
nand U8275 ( n1966, n1967, n191 );
nor U8276 ( n1967, n193, n759 );
nor U8277 ( n972, n1167, n533 );
nor U8278 ( n1013, n1185, n422 );
nor U8279 ( n1049, n1127, n313 );
nor U8280 ( n1074, n1147, n192 );
nand U8281 ( n1167, n534, n532 );
nand U8282 ( n1185, n423, n421 );
nand U8283 ( n1127, n314, n312 );
nand U8284 ( n1147, n193, n191 );
nor U8285 ( n1212, n901, n1445 );
xor U8286 ( n1445, n503, n531 );
nor U8287 ( n803, n968, n969 );
xor U8288 ( n969, n504, n531 );
nor U8289 ( n1275, n1313, n1443 );
xor U8290 ( n1443, n507, n531 );
nor U8291 ( n1232, n948, n1491 );
xor U8292 ( n1491, n395, n420 );
nor U8293 ( n839, n1009, n1010 );
xor U8294 ( n1010, n396, n420 );
nor U8295 ( n1321, n1349, n1489 );
xor U8296 ( n1489, n399, n420 );
nor U8297 ( n1263, n992, n1537 );
xor U8298 ( n1537, n286, n311 );
nor U8299 ( n877, n1045, n1046 );
xor U8300 ( n1046, n287, n311 );
nor U8301 ( n1357, n1383, n1535 );
xor U8302 ( n1535, n290, n311 );
nor U8303 ( n1303, n1033, n1578 );
xor U8304 ( n1578, n165, n190 );
nor U8305 ( n923, n1070, n1071 );
xor U8306 ( n1071, n166, n190 );
nor U8307 ( n1391, n1408, n1576 );
xor U8308 ( n1576, n169, n190 );
and U8309 ( n785, n1447, n936 );
nor U8310 ( n1447, n529, n1448 );
xor U8311 ( n1448, n531, n502 );
and U8312 ( n818, n1493, n980 );
nor U8313 ( n1493, n418, n1495 );
xor U8314 ( n1495, n420, n394 );
and U8315 ( n854, n1539, n1021 );
nor U8316 ( n1539, n309, n1540 );
xor U8317 ( n1540, n311, n285 );
and U8318 ( n892, n1580, n1057 );
nor U8319 ( n1580, n188, n1581 );
xor U8320 ( n1581, n190, n164 );
nand U8321 ( n1677, n2117, n120 );
nor U8322 ( n2117, n510, n511 );
nand U8323 ( n1699, n2158, n54 );
nor U8324 ( n2158, n401, n402 );
nand U8325 ( n1721, n2197, n76 );
nor U8326 ( n2197, n292, n293 );
nand U8327 ( n1741, n2231, n98 );
nor U8328 ( n2231, n171, n172 );
nand U8329 ( n2079, n2082, n2083 );
nand U8330 ( n2124, n2126, n2127 );
nand U8331 ( n2165, n2167, n2168 );
nand U8332 ( n2205, n2207, n2208 );
nor U8333 ( n2107, n545, n119 );
nor U8334 ( n2148, n432, n53 );
nor U8335 ( n2185, n323, n75 );
nor U8336 ( n2220, n202, n97 );
and U8337 ( n1797, n1808, n1804 );
and U8338 ( n1862, n1872, n1868 );
and U8339 ( n1931, n1942, n1938 );
and U8340 ( n1997, n2009, n2003 );
nor U8341 ( n1795, n1797, n1798 );
and U8342 ( n1798, n1799, n1801 );
nor U8343 ( n1860, n1862, n1863 );
and U8344 ( n1863, n1864, n1865 );
nor U8345 ( n1929, n1931, n1932 );
and U8346 ( n1932, n1933, n1934 );
nor U8347 ( n1994, n1997, n1998 );
and U8348 ( n1998, n1999, n2000 );
and U8349 ( n1601, n1609, n129 );
nand U8350 ( n1609, n1611, n531 );
nand U8351 ( n1611, n1612, n1174 );
nor U8352 ( n1612, n534, n528 );
and U8353 ( n1606, n1620, n63 );
nand U8354 ( n1620, n1622, n420 );
nand U8355 ( n1622, n1623, n1192 );
nor U8356 ( n1623, n423, n417 );
and U8357 ( n1617, n1631, n85 );
nand U8358 ( n1631, n1633, n311 );
nand U8359 ( n1633, n1634, n1134 );
nor U8360 ( n1634, n314, n308 );
and U8361 ( n1628, n1639, n107 );
nand U8362 ( n1639, n1641, n190 );
nand U8363 ( n1641, n1642, n1154 );
nor U8364 ( n1642, n193, n187 );
and U8365 ( n1774, n7331, n7332 );
nand U8366 ( n7331, n1780, n1781 );
nand U8367 ( n7332, n1778, n1779 );
and U8368 ( n1841, n7333, n7334 );
nand U8369 ( n7333, n1847, n1848 );
nand U8370 ( n7334, n1845, n1846 );
and U8371 ( n1907, n7335, n7336 );
nand U8372 ( n7335, n1914, n1915 );
nand U8373 ( n7336, n1912, n1913 );
and U8374 ( n1972, n7337, n7338 );
nand U8375 ( n7337, n1979, n1980 );
nand U8376 ( n7338, n1977, n1978 );
not U8377 ( n530, n3887 );
not U8378 ( n419, n3963 );
not U8379 ( n310, n4033 );
not U8380 ( n189, n4103 );
or U8381 ( n1676, n1677, n1678 );
or U8382 ( n1698, n1699, n1700 );
or U8383 ( n1720, n1721, n1722 );
or U8384 ( n1740, n1741, n1742 );
nand U8385 ( n2064, n524, n2079 );
nand U8386 ( n2075, n414, n2124 );
nand U8387 ( n2095, n305, n2165 );
nand U8388 ( n2138, n184, n2205 );
nand U8389 ( n1681, n119, n545 );
nand U8390 ( n1703, n53, n432 );
nand U8391 ( n1725, n75, n323 );
nand U8392 ( n1745, n97, n202 );
not U8393 ( n129, n1435 );
not U8394 ( n63, n1479 );
not U8395 ( n85, n1527 );
not U8396 ( n107, n1568 );
xor U8397 ( n936, n972, n498 );
xor U8398 ( n980, n1013, n390 );
xor U8399 ( n1021, n1049, n281 );
xor U8400 ( n1057, n1074, n160 );
nand U8401 ( n1682, n512, n1683 );
nand U8402 ( n1704, n403, n1705 );
nand U8403 ( n1726, n294, n1727 );
nand U8404 ( n1747, n173, n1748 );
nand U8405 ( n1818, n1797, n1799 );
nand U8406 ( n1881, n1862, n1864 );
nand U8407 ( n1952, n1931, n1933 );
nand U8408 ( n2018, n1997, n1999 );
nand U8409 ( n1437, n4885, n533 );
nor U8410 ( n4885, n534, n532 );
nand U8411 ( n1482, n4895, n422 );
nor U8412 ( n4895, n423, n421 );
nand U8413 ( n1529, n4906, n313 );
nor U8414 ( n4906, n314, n312 );
nand U8415 ( n1570, n4911, n192 );
nor U8416 ( n4911, n193, n191 );
nand U8417 ( n1820, n1823, n1781 );
and U8418 ( n1823, n1779, n1780 );
nand U8419 ( n1884, n1887, n1848 );
and U8420 ( n1887, n1846, n1847 );
nand U8421 ( n1954, n1958, n1915 );
and U8422 ( n1958, n1913, n1914 );
nand U8423 ( n2020, n2023, n1980 );
and U8424 ( n2023, n1978, n1979 );
not U8425 ( n539, n2920 );
not U8426 ( n427, n3007 );
not U8427 ( n318, n3095 );
not U8428 ( n197, n3200 );
not U8429 ( n146, n4338 );
and U8430 ( n4305, n6150, n155 );
or U8431 ( n1427, n1428, n500 );
or U8432 ( n1471, n1472, n392 );
or U8433 ( n1519, n1520, n283 );
or U8434 ( n1560, n1561, n162 );
xor U8435 ( n6595, n6596, n6598 );
xor U8436 ( n6596, n6602, n6603 );
xor U8437 ( n6598, n6599, n6600 );
xor U8438 ( n6402, n6403, n6404 );
xor U8439 ( n6403, n6407, n6408 );
xor U8440 ( n6404, n6405, n6406 );
xor U8441 ( n6788, n6789, n6790 );
xor U8442 ( n6789, n6793, n6794 );
xor U8443 ( n6790, n6791, n6792 );
xor U8444 ( n6208, n6216, n6217 );
xor U8445 ( n6216, n6220, n6221 );
xor U8446 ( n6217, n6218, n6219 );
xor U8447 ( n6787, n6795, n6796 );
xor U8448 ( n6795, n6799, n6800 );
xor U8449 ( n6796, n6797, n6798 );
xor U8450 ( n6594, n6604, n6605 );
xor U8451 ( n6604, n6608, n6609 );
xor U8452 ( n6605, n6606, n6607 );
nand U8453 ( n6797, n6817, n6879 );
nand U8454 ( n6879, n6880, n6881 );
nand U8455 ( n6881, n601, n570 );
nor U8456 ( n6880, n6882, n6883 );
nand U8457 ( n6606, n6626, n6683 );
nand U8458 ( n6683, n6684, n6685 );
nand U8459 ( n6685, n482, n455 );
nor U8460 ( n6684, n6686, n6687 );
xor U8461 ( n6209, n6210, n6211 );
xnor U8462 ( n6210, n6214, n6215 );
xnor U8463 ( n6211, n6212, n6213 );
xor U8464 ( n6401, n6409, n6410 );
xnor U8465 ( n6409, n6413, n6414 );
xnor U8466 ( n6410, n6411, n6412 );
nand U8467 ( n6411, n6431, n6488 );
nand U8468 ( n6488, n6489, n6490 );
nand U8469 ( n6490, n374, n346 );
nor U8470 ( n6489, n6491, n6492 );
nand U8471 ( n3893, n501, n506 );
nand U8472 ( n3967, n393, n398 );
nand U8473 ( n4037, n284, n289 );
nand U8474 ( n4107, n163, n168 );
and U8475 ( n2995, n3140, n3141 );
nand U8476 ( n3140, n43, n530 );
and U8477 ( n3083, n3229, n3230 );
nand U8478 ( n3229, n43, n419 );
and U8479 ( n3185, n3297, n3298 );
nand U8480 ( n3297, n43, n310 );
and U8481 ( n3273, n3329, n3330 );
nand U8482 ( n3329, n43, n189 );
nor U8483 ( n6299, n246, n6218 );
nor U8484 ( n6307, n246, n6221 );
nor U8485 ( n6285, n246, n6219 );
nor U8486 ( n6273, n246, n6215 );
nor U8487 ( n6319, n246, n6220 );
nor U8488 ( n6237, n246, n6213 );
nor U8489 ( n6254, n246, n6212 );
nor U8490 ( n6264, n246, n6214 );
not U8491 ( n226, n6229 );
nor U8492 ( n6816, n579, n6792 );
nor U8493 ( n6625, n463, n6600 );
nor U8494 ( n6430, n354, n6406 );
nor U8495 ( n6475, n354, n6412 );
nor U8496 ( n6889, n579, n6800 );
nor U8497 ( n6864, n579, n6798 );
nor U8498 ( n6692, n463, n6609 );
nor U8499 ( n6670, n463, n6607 );
nor U8500 ( n6660, n463, n6602 );
nor U8501 ( n6637, n463, n6599 );
nor U8502 ( n6646, n463, n6603 );
nor U8503 ( n6513, n354, n6414 );
nor U8504 ( n6465, n354, n6407 );
nor U8505 ( n6442, n354, n6405 );
nor U8506 ( n6451, n354, n6408 );
nor U8507 ( n6907, n579, n6799 );
nor U8508 ( n6853, n579, n6793 );
nor U8509 ( n6828, n579, n6791 );
nor U8510 ( n6837, n579, n6794 );
nor U8511 ( n6708, n463, n6608 );
nor U8512 ( n6497, n354, n6413 );
not U8513 ( n233, n6808 );
not U8514 ( n236, n6617 );
not U8515 ( n239, n6422 );
nor U8516 ( n2645, n2646, n2647 );
nand U8517 ( n2647, n2648, n2649 );
nand U8518 ( n2649, n217, n2636 );
nand U8519 ( n2648, n2650, n229 );
and U8520 ( n2650, n2678, n228 );
nor U8521 ( n2678, n216, n218 );
nor U8522 ( n2541, n2542, n2543 );
nand U8523 ( n2543, n2544, n2545 );
nand U8524 ( n2545, n338, n2532 );
nand U8525 ( n2544, n2546, n348 );
nor U8526 ( n2430, n2431, n2432 );
nand U8527 ( n2432, n2433, n2434 );
nand U8528 ( n2434, n447, n2421 );
nand U8529 ( n2433, n2435, n457 );
and U8530 ( n2546, n2574, n347 );
nor U8531 ( n2574, n337, n339 );
and U8532 ( n2435, n2463, n456 );
nor U8533 ( n2463, n446, n448 );
nor U8534 ( n2289, n2269, n2292 );
nand U8535 ( n2292, n158, n2266 );
nor U8536 ( n2317, n2318, n2319 );
nand U8537 ( n2319, n2320, n2321 );
nand U8538 ( n2321, n561, n2308 );
nand U8539 ( n2320, n2322, n573 );
and U8540 ( n2322, n2350, n572 );
nor U8541 ( n2350, n560, n563 );
nand U8542 ( n3141, n4928, n534 );
nor U8543 ( n4928, n532, n533 );
nand U8544 ( n3298, n4962, n314 );
nor U8545 ( n4962, n312, n313 );
nand U8546 ( n3230, n4945, n423 );
nor U8547 ( n4945, n421, n422 );
nor U8548 ( n4264, n7435, n43 );
nor U8549 ( n4268, n7447, n43 );
nor U8550 ( n4272, n7459, n43 );
nor U8551 ( n4276, n7471, n43 );
nand U8552 ( n3330, n4977, n193 );
nor U8553 ( n4977, n191, n192 );
not U8554 ( n143, g26135 );
nor U8555 ( n6883, n601, n6884 );
nor U8556 ( n6687, n482, n6688 );
nor U8557 ( n6258, n265, n6249 );
nor U8558 ( n6492, n374, n6493 );
and U8559 ( n2419, n2420, n2421 );
not U8560 ( n48, g27380 );
and U8561 ( n2634, n2635, n2636 );
not U8562 ( n568, n6823 );
not U8563 ( n453, n6632 );
and U8564 ( n2530, n2531, n2532 );
not U8565 ( n569, n6884 );
not U8566 ( n454, n6688 );
not U8567 ( n345, n6493 );
not U8568 ( n225, n6291 );
not U8569 ( n344, n6437 );
and U8570 ( n2306, n2307, n2308 );
not U8571 ( n222, n6249 );
nor U8572 ( n2307, n561, n560 );
nor U8573 ( n2635, n217, n216 );
nor U8574 ( n2531, n338, n337 );
nor U8575 ( n2420, n447, n446 );
nand U8576 ( n2410, n2411, n448 );
nand U8577 ( n2626, n2627, n218 );
nand U8578 ( n2522, n2523, n339 );
nand U8579 ( n2298, n2299, n563 );
not U8580 ( n7498, n7499 );
not U8581 ( n260, n6259 );
not U8582 ( n595, n6848 );
not U8583 ( n477, n6656 );
not U8584 ( n369, n6461 );
not U8585 ( n10, n4541 );
not U8586 ( n11, n4544 );
not U8587 ( n13, n4552 );
not U8588 ( n12, n4549 );
not U8589 ( n14, n4565 );
not U8590 ( n16, n4580 );
not U8591 ( n15, n4570 );
not U8592 ( n17, n4593 );
not U8593 ( n19, n4612 );
not U8594 ( n18, n4598 );
not U8595 ( n20, n4625 );
not U8596 ( n21, n4645 );
buf U8597 ( n7382, n7500 );
buf U8598 ( n7384, n7500 );
buf U8599 ( n7383, n7500 );
nor U8600 ( n2796, n322, n306 );
nor U8601 ( n2752, n543, n525 );
nor U8602 ( n2775, n431, n415 );
nor U8603 ( n2812, n201, n185 );
nor U8604 ( n4717, n158, n624 );
not U8605 ( n591, n4367 );
not U8606 ( n592, n4364 );
not U8607 ( n473, n4410 );
not U8608 ( n474, n4371 );
not U8609 ( n365, n4453 );
not U8610 ( n366, n4414 );
not U8611 ( n256, n4502 );
not U8612 ( n257, n4457 );
not U8613 ( n590, n4407 );
not U8614 ( n472, n4450 );
not U8615 ( n364, n4499 );
not U8616 ( n255, n4538 );
nand U8617 ( n2033, n410, n43 );
nand U8618 ( n2039, n301, n43 );
nand U8619 ( n2044, n180, n43 );
nand U8620 ( n2027, n43, n520 );
not U8621 ( n247, n6227 );
not U8622 ( n581, n6806 );
not U8623 ( n464, n6615 );
not U8624 ( n355, n6420 );
nor U8625 ( n6243, n6327, n247 );
nor U8626 ( n6843, n6913, n581 );
nor U8627 ( n6651, n6713, n464 );
nor U8628 ( n6456, n6518, n355 );
not U8629 ( n622, n4696 );
not U8630 ( n7, n4826 );
not U8631 ( n246, n6327 );
not U8632 ( n579, n6913 );
not U8633 ( n463, n6713 );
not U8634 ( n354, n6518 );
not U8635 ( n5, n4688 );
xnor U8636 ( n1796, n808, n500 );
xnor U8637 ( n1861, n844, n392 );
xnor U8638 ( n1930, n882, n283 );
xnor U8639 ( n1996, n928, n162 );
nand U8640 ( n767, n780, n781 );
nand U8641 ( n781, n782, n783 );
nor U8642 ( n780, n786, n787 );
xor U8643 ( n782, n784, n785 );
nand U8644 ( n907, n965, n966 );
nand U8645 ( n966, n967, n783 );
nor U8646 ( n965, n786, n970 );
xor U8647 ( n967, n805, n803 );
nand U8648 ( n775, n813, n814 );
nand U8649 ( n814, n815, n816 );
nor U8650 ( n813, n819, n820 );
xor U8651 ( n815, n817, n818 );
nand U8652 ( n954, n1006, n1007 );
nand U8653 ( n1007, n1008, n816 );
nor U8654 ( n1006, n819, n1011 );
xor U8655 ( n1008, n841, n839 );
nand U8656 ( n795, n849, n850 );
nand U8657 ( n850, n851, n852 );
nor U8658 ( n849, n855, n856 );
xor U8659 ( n851, n853, n854 );
nand U8660 ( n998, n1042, n1043 );
nand U8661 ( n1043, n1044, n852 );
nor U8662 ( n1042, n855, n1047 );
xor U8663 ( n1044, n879, n877 );
nand U8664 ( n828, n887, n888 );
nand U8665 ( n888, n889, n890 );
nor U8666 ( n887, n893, n894 );
xor U8667 ( n889, n891, n892 );
nand U8668 ( n1039, n1067, n1068 );
nand U8669 ( n1068, n1069, n890 );
nor U8670 ( n1067, n893, n1072 );
xor U8671 ( n1069, n925, n923 );
nor U8672 ( n787, n7128, n125 );
nor U8673 ( n820, n7129, n59 );
nor U8674 ( n856, n7134, n81 );
nor U8675 ( n894, n7136, n103 );
nand U8676 ( n725, n1138, n1925 );
nand U8677 ( n1925, n1926, n1927 );
nand U8678 ( n1927, n1929, n1930 );
nor U8679 ( n1926, n1935, n1936 );
nand U8680 ( n758, n1158, n1990 );
nand U8681 ( n1990, n1992, n1993 );
nand U8682 ( n1993, n1994, n1996 );
nor U8683 ( n1992, n2001, n2002 );
nand U8684 ( n1431, n1093, n1432 );
nand U8685 ( n1432, n1433, n533 );
nor U8686 ( n1433, n541, n1100 );
nand U8687 ( n1475, n681, n1476 );
nand U8688 ( n1476, n1477, n422 );
nor U8689 ( n1477, n429, n688 );
nand U8690 ( n1523, n718, n1524 );
nand U8691 ( n1524, n1525, n313 );
nor U8692 ( n1525, n320, n726 );
nand U8693 ( n1564, n752, n1565 );
nand U8694 ( n1565, n1566, n192 );
nor U8695 ( n1566, n199, n759 );
nand U8696 ( n1099, n1178, n1792 );
nand U8697 ( n1792, n1793, n1794 );
nand U8698 ( n1794, n1795, n1796 );
nor U8699 ( n1793, n1802, n1803 );
nand U8700 ( n687, n1196, n1857 );
nand U8701 ( n1857, n1858, n1859 );
nand U8702 ( n1859, n1860, n1861 );
nor U8703 ( n1858, n1866, n1867 );
and U8704 ( n1415, n1429, n1430 );
nor U8705 ( n1429, n1435, n1436 );
nand U8706 ( n1430, n1431, n1082 );
nor U8707 ( n1436, n1437, n1438 );
and U8708 ( n1459, n1473, n1474 );
nor U8709 ( n1473, n1479, n1480 );
nand U8710 ( n1474, n1475, n670 );
nor U8711 ( n1480, n1482, n1483 );
and U8712 ( n1507, n1521, n1522 );
nor U8713 ( n1521, n1527, n1528 );
nand U8714 ( n1522, n1523, n706 );
nor U8715 ( n1528, n1529, n1530 );
and U8716 ( n1548, n1562, n1563 );
nor U8717 ( n1562, n1568, n1569 );
nand U8718 ( n1563, n1564, n741 );
nor U8719 ( n1569, n1570, n1571 );
nor U8720 ( n807, n808, n125 );
nor U8721 ( n843, n844, n59 );
nor U8722 ( n881, n882, n81 );
nor U8723 ( n927, n928, n103 );
and U8724 ( n831, n897, n898 );
nand U8725 ( n898, n783, n899 );
nor U8726 ( n897, n806, n902 );
xor U8727 ( n899, n900, n901 );
and U8728 ( n866, n931, n932 );
nand U8729 ( n932, n783, n933 );
nor U8730 ( n931, n806, n938 );
xor U8731 ( n933, n934, n935 );
and U8732 ( n770, n798, n799 );
nand U8733 ( n799, n783, n800 );
nor U8734 ( n798, n806, n807 );
xor U8735 ( n800, n801, n802 );
and U8736 ( n869, n944, n945 );
nand U8737 ( n945, n816, n946 );
nor U8738 ( n944, n842, n949 );
xor U8739 ( n946, n947, n948 );
and U8740 ( n912, n975, n976 );
nand U8741 ( n976, n816, n977 );
nor U8742 ( n975, n842, n982 );
xor U8743 ( n977, n978, n979 );
and U8744 ( n790, n834, n835 );
nand U8745 ( n835, n816, n836 );
nor U8746 ( n834, n842, n843 );
xor U8747 ( n836, n837, n838 );
and U8748 ( n915, n988, n989 );
nand U8749 ( n989, n852, n990 );
nor U8750 ( n988, n880, n993 );
xor U8751 ( n990, n991, n992 );
and U8752 ( n959, n1016, n1017 );
nand U8753 ( n1017, n852, n1018 );
nor U8754 ( n1016, n880, n1023 );
xor U8755 ( n1018, n1019, n1020 );
and U8756 ( n823, n872, n873 );
nand U8757 ( n873, n852, n874 );
nor U8758 ( n872, n880, n881 );
xor U8759 ( n874, n875, n876 );
and U8760 ( n962, n1029, n1030 );
nand U8761 ( n1030, n890, n1031 );
nor U8762 ( n1029, n926, n1034 );
xor U8763 ( n1031, n1032, n1033 );
and U8764 ( n1003, n1052, n1053 );
nand U8765 ( n1053, n890, n1054 );
nor U8766 ( n1052, n926, n1060 );
xor U8767 ( n1054, n1055, n1056 );
and U8768 ( n859, n918, n919 );
nand U8769 ( n919, n890, n920 );
nor U8770 ( n918, n926, n927 );
xor U8771 ( n920, n921, n922 );
xnor U8772 ( n1775, n1822, n506 );
xnor U8773 ( n1842, n1886, n398 );
xnor U8774 ( n1908, n1957, n289 );
xnor U8775 ( n1974, n2022, n168 );
nand U8776 ( n1103, n1178, n1770 );
nand U8777 ( n1770, n1771, n1772 );
nand U8778 ( n1772, n1774, n1775 );
nor U8779 ( n1771, n1783, n1784 );
nand U8780 ( n691, n1196, n1838 );
nand U8781 ( n1838, n1839, n1840 );
nand U8782 ( n1840, n1841, n1842 );
nor U8783 ( n1839, n1849, n1850 );
nand U8784 ( n729, n1138, n1904 );
nand U8785 ( n1904, n1905, n1906 );
nand U8786 ( n1906, n1907, n1908 );
nor U8787 ( n1905, n1916, n1917 );
nand U8788 ( n762, n1158, n1969 );
nand U8789 ( n1969, n1970, n1971 );
nand U8790 ( n1971, n1972, n1974 );
nor U8791 ( n1970, n1981, n1983 );
not U8792 ( n511, n808 );
not U8793 ( n402, n844 );
not U8794 ( n293, n882 );
not U8795 ( n172, n928 );
nand U8796 ( n4230, n4231, n4232 );
xor U8797 ( n4232, n4233, n510 );
xor U8798 ( n4231, n4238, n511 );
nand U8799 ( n4233, n4234, n4235 );
nand U8800 ( n3598, n3599, n3600 );
xor U8801 ( n3600, n3601, n401 );
xor U8802 ( n3599, n3607, n402 );
nand U8803 ( n3601, n3603, n3604 );
nand U8804 ( n3702, n3703, n3704 );
xor U8805 ( n3704, n3706, n292 );
xor U8806 ( n3703, n3712, n293 );
nand U8807 ( n3706, n3707, n3708 );
nand U8808 ( n3801, n3802, n3803 );
xor U8809 ( n3803, n3805, n171 );
xor U8810 ( n3802, n3810, n172 );
nand U8811 ( n3805, n3806, n3807 );
nand U8812 ( n1094, n4187, n4188 );
nor U8813 ( n4188, n4189, n4190 );
nor U8814 ( n4187, n4229, n4230 );
nand U8815 ( n4189, n4210, n4211 );
nand U8816 ( n682, n3553, n3554 );
nor U8817 ( n3554, n3555, n3556 );
nor U8818 ( n3553, n3597, n3598 );
nand U8819 ( n3555, n3576, n3577 );
nand U8820 ( n720, n3653, n3654 );
nor U8821 ( n3654, n3655, n3657 );
nor U8822 ( n3653, n3701, n3702 );
nand U8823 ( n3655, n3679, n3680 );
nand U8824 ( n753, n3752, n3753 );
nor U8825 ( n3753, n3754, n3756 );
nor U8826 ( n3752, n3799, n3801 );
nand U8827 ( n3754, n3778, n3779 );
not U8828 ( n510, n1822 );
not U8829 ( n401, n1886 );
not U8830 ( n292, n1957 );
not U8831 ( n171, n2022 );
nor U8832 ( n4210, n4217, n4218 );
xor U8833 ( n4217, n7130, n4224 );
xor U8834 ( n4218, n7128, n4219 );
nor U8835 ( n4224, n4225, n4226 );
nor U8836 ( n3576, n3583, n3585 );
xor U8837 ( n3583, n7131, n3591 );
xor U8838 ( n3585, n7129, n3586 );
nor U8839 ( n3591, n3592, n3594 );
nor U8840 ( n3679, n3687, n3688 );
xor U8841 ( n3687, n7137, n3695 );
xor U8842 ( n3688, n7134, n3689 );
nor U8843 ( n3695, n3697, n3698 );
nor U8844 ( n3778, n3786, n3787 );
xor U8845 ( n3786, n7138, n3794 );
xor U8846 ( n3787, n7136, n3788 );
nor U8847 ( n3794, n3795, n3796 );
nand U8848 ( n4229, n4243, n1178 );
nor U8849 ( n4243, n4248, n4249 );
xor U8850 ( n4248, n7142, n4255 );
xor U8851 ( n4249, n7149, n4250 );
nand U8852 ( n3597, n3613, n1196 );
nor U8853 ( n3613, n3618, n3619 );
xor U8854 ( n3618, n7143, n3626 );
xor U8855 ( n3619, n7150, n3621 );
nand U8856 ( n3701, n3717, n1138 );
nor U8857 ( n3717, n3722, n3723 );
xor U8858 ( n3722, n7146, n3729 );
xor U8859 ( n3723, n7153, n3724 );
nand U8860 ( n3799, n3815, n1158 );
nor U8861 ( n3815, n3820, n3821 );
xor U8862 ( n3820, n7147, n3827 );
xor U8863 ( n3821, n7154, n3822 );
nor U8864 ( n1079, n1085, n1086 );
nor U8865 ( n1085, n533, n1101 );
nand U8866 ( n1086, n1087, n1082 );
nor U8867 ( n1101, n1102, n131 );
nor U8868 ( n667, n673, n674 );
nor U8869 ( n673, n422, n689 );
nand U8870 ( n674, n675, n670 );
nor U8871 ( n689, n690, n65 );
nor U8872 ( n703, n709, n710 );
nor U8873 ( n709, n313, n727 );
nand U8874 ( n710, n711, n706 );
nor U8875 ( n727, n728, n87 );
nor U8876 ( n738, n744, n745 );
nor U8877 ( n744, n192, n760 );
nand U8878 ( n745, n746, n741 );
nor U8879 ( n760, n761, n109 );
and U8880 ( n662, n701, n85 );
xor U8881 ( n701, n313, n702 );
nor U8882 ( n702, n703, n704 );
nor U8883 ( n704, n705, n706 );
and U8884 ( n698, n736, n107 );
xor U8885 ( n736, n192, n737 );
nor U8886 ( n737, n738, n739 );
nor U8887 ( n739, n740, n741 );
and U8888 ( n650, n1077, n129 );
xor U8889 ( n1077, n533, n1078 );
nor U8890 ( n1078, n1079, n1080 );
nor U8891 ( n1080, n1081, n1082 );
and U8892 ( n654, n665, n63 );
xor U8893 ( n665, n422, n666 );
nor U8894 ( n666, n667, n668 );
nor U8895 ( n668, n669, n670 );
nand U8896 ( n1438, n128, n1434 );
nand U8897 ( n1483, n62, n1478 );
nand U8898 ( n1530, n84, n1526 );
nand U8899 ( n1571, n106, n1567 );
and U8900 ( n1245, n1309, n1310 );
nand U8901 ( n1310, n783, n1311 );
nor U8902 ( n1309, n126, n1314 );
xor U8903 ( n1311, n1312, n1313 );
and U8904 ( n1285, n1345, n1346 );
nand U8905 ( n1346, n816, n1347 );
nor U8906 ( n1345, n60, n1350 );
xor U8907 ( n1347, n1348, n1349 );
and U8908 ( n1331, n1379, n1380 );
nand U8909 ( n1380, n852, n1381 );
nor U8910 ( n1379, n82, n1384 );
xor U8911 ( n1381, n1382, n1383 );
and U8912 ( n1367, n1404, n1405 );
nand U8913 ( n1405, n890, n1406 );
nor U8914 ( n1404, n104, n1409 );
xor U8915 ( n1406, n1407, n1408 );
and U8916 ( n1223, n1271, n1272 );
nand U8917 ( n1272, n783, n1273 );
nor U8918 ( n1271, n126, n1278 );
xor U8919 ( n1273, n1274, n968 );
and U8920 ( n1254, n1317, n1318 );
nand U8921 ( n1318, n816, n1319 );
nor U8922 ( n1317, n60, n1324 );
xor U8923 ( n1319, n1320, n1009 );
and U8924 ( n1294, n1353, n1354 );
nand U8925 ( n1354, n852, n1355 );
nor U8926 ( n1353, n82, n1360 );
xor U8927 ( n1355, n1356, n1045 );
and U8928 ( n1340, n1387, n1388 );
nand U8929 ( n1388, n890, n1389 );
nor U8930 ( n1387, n104, n1394 );
xor U8931 ( n1389, n1390, n1070 );
nor U8932 ( n1435, n1094, n1610 );
nor U8933 ( n1479, n682, n1621 );
nor U8934 ( n1527, n720, n1632 );
nor U8935 ( n1568, n753, n1640 );
not U8936 ( n637, n4346 );
or U8937 ( g26149, n4277, n4278 );
nand U8938 ( n4277, n4298, n4299 );
nand U8939 ( n4278, n4279, n4280 );
nor U8940 ( n4298, n4309, n4310 );
and U8941 ( n1097, n1093, n1177 );
nand U8942 ( n1177, n124, n1178 );
not U8943 ( n124, n1179 );
and U8944 ( n685, n681, n1195 );
nand U8945 ( n1195, n58, n1196 );
not U8946 ( n58, n1197 );
and U8947 ( n723, n718, n1137 );
nand U8948 ( n1137, n80, n1138 );
not U8949 ( n80, n1139 );
and U8950 ( n756, n752, n1157 );
nand U8951 ( n1157, n102, n1158 );
not U8952 ( n102, n1159 );
nand U8953 ( g26135, n6141, n6142 );
nor U8954 ( n6142, n6143, n6144 );
nor U8955 ( n6141, n6174, n6175 );
nand U8956 ( n6143, n6156, n6157 );
nand U8957 ( g26104, n4319, n4320 );
nor U8958 ( n4320, n4321, n4322 );
nor U8959 ( n4319, n4339, n4340 );
nand U8960 ( n4322, n4323, n4324 );
nor U8961 ( n1186, n1189, n1190 );
nor U8962 ( n1189, n671, n1194 );
nor U8963 ( n1190, n1191, n672 );
nand U8964 ( n1194, n685, n672 );
nor U8965 ( n1128, n1131, n1132 );
nor U8966 ( n1131, n707, n1136 );
nor U8967 ( n1132, n1133, n708 );
nand U8968 ( n1136, n723, n708 );
nor U8969 ( n1148, n1151, n1152 );
nor U8970 ( n1151, n742, n1156 );
nor U8971 ( n1152, n1153, n743 );
nand U8972 ( n1156, n756, n743 );
nor U8973 ( n1168, n1171, n1172 );
nor U8974 ( n1171, n1083, n1176 );
nor U8975 ( n1172, n1173, n1084 );
nand U8976 ( n1176, n1097, n1084 );
xnor U8977 ( n3105, n2624, g3229 );
xnor U8978 ( n3017, n2520, g3229 );
xnor U8979 ( n2930, n2408, g3229 );
xnor U8980 ( n2875, n2296, g3229 );
and U8981 ( n2959, n3103, n3104 );
nand U8982 ( n3104, n2636, n3105 );
nand U8983 ( n3103, n230, n2632 );
and U8984 ( n2904, n3015, n3016 );
nand U8985 ( n3016, n2532, n3017 );
nand U8986 ( n3015, n349, n2528 );
and U8987 ( n2866, n2928, n2929 );
nand U8988 ( n2929, n2421, n2930 );
nand U8989 ( n2928, n458, n2416 );
and U8990 ( n2844, n2873, n2874 );
nand U8991 ( n2874, n2308, n2875 );
nand U8992 ( n2873, n574, n2304 );
not U8993 ( g24734, n7043 );
nand U8994 ( g27380, n6114, n6115 );
nor U8995 ( n6115, n6116, n6117 );
nor U8996 ( n6114, n4346, n6138 );
nand U8997 ( n6116, n6128, n6129 );
and U8998 ( n3036, n3189, n3190 );
nand U8999 ( n3190, n3105, n2639 );
and U9000 ( n2949, n3086, n3087 );
nand U9001 ( n3087, n3017, n2535 );
and U9002 ( n2894, n2998, n2999 );
nand U9003 ( n2999, n2930, n2424 );
and U9004 ( n2856, n2911, n2912 );
nand U9005 ( n2912, n2875, n2311 );
nand U9006 ( n1104, n1178, n1179 );
nand U9007 ( n730, n1138, n1139 );
nand U9008 ( n692, n1196, n1197 );
nand U9009 ( n763, n1158, n1159 );
and U9010 ( n3110, n3240, n3241 );
nand U9011 ( n3241, g3229, n2651 );
nor U9012 ( n3240, n3242, n3243 );
nor U9013 ( n3242, n2651, n3244 );
and U9014 ( n3022, n3151, n3152 );
nand U9015 ( n3152, g3229, n2547 );
nor U9016 ( n3151, n3153, n3154 );
nor U9017 ( n3153, n2547, n3155 );
and U9018 ( n2935, n3050, n3051 );
nand U9019 ( n3051, g3229, n2436 );
nor U9020 ( n3050, n3052, n3053 );
nor U9021 ( n3052, n2436, n3054 );
and U9022 ( n2880, n2962, n2963 );
nand U9023 ( n2963, g3229, n2323 );
nor U9024 ( n2962, n2964, n2965 );
nor U9025 ( n2964, n2323, n2966 );
and U9026 ( n2994, n3119, n3120 );
nand U9027 ( n3120, g3229, n2988 );
nor U9028 ( n3119, n3121, n3122 );
nor U9029 ( n3121, n2988, n3123 );
and U9030 ( n3082, n3208, n3209 );
nand U9031 ( n3209, g3229, n3076 );
nor U9032 ( n3208, n3210, n3211 );
nor U9033 ( n3210, n3076, n3212 );
and U9034 ( n3184, n3276, n3277 );
nand U9035 ( n3277, g3229, n3177 );
nor U9036 ( n3276, n3278, n3279 );
nor U9037 ( n3278, n3177, n3280 );
and U9038 ( n3272, n3308, n3309 );
nand U9039 ( n3309, g3229, n3266 );
nor U9040 ( n3308, n3310, n3311 );
nor U9041 ( n3310, n3266, n3312 );
nor U9042 ( n1169, n534, n1170 );
and U9043 ( n1170, n1083, n1104 );
nor U9044 ( n1129, n314, n1130 );
and U9045 ( n1130, n707, n730 );
nor U9046 ( n1187, n423, n1188 );
and U9047 ( n1188, n671, n692 );
nor U9048 ( n1149, n193, n1150 );
and U9049 ( n1150, n742, n763 );
xnor U9050 ( n1779, n7130, n498 );
xnor U9051 ( n1846, n7131, n390 );
xnor U9052 ( n1913, n7137, n281 );
xnor U9053 ( n1978, n7138, n160 );
not U9054 ( n498, n1251 );
not U9055 ( n390, n1291 );
not U9056 ( n281, n1337 );
not U9057 ( n160, n1373 );
not U9058 ( n500, n801 );
not U9059 ( n392, n837 );
not U9060 ( n283, n875 );
not U9061 ( n162, n921 );
xor U9062 ( n1801, n934, n7124 );
xor U9063 ( n1865, n978, n7125 );
xor U9064 ( n1934, n1019, n7126 );
xor U9065 ( n2000, n1055, n7127 );
not U9066 ( n532, n1083 );
not U9067 ( n421, n671 );
not U9068 ( n312, n707 );
not U9069 ( n191, n742 );
nand U9070 ( n968, n1275, n1276 );
xor U9071 ( n1276, n1277, n531 );
nand U9072 ( n1313, n1212, n1444 );
xor U9073 ( n1444, n1211, n531 );
nand U9074 ( n901, n785, n1446 );
xor U9075 ( n1446, n784, n531 );
nand U9076 ( n1009, n1321, n1322 );
xor U9077 ( n1322, n1323, n420 );
nand U9078 ( n1349, n1232, n1490 );
xor U9079 ( n1490, n1231, n420 );
nand U9080 ( n948, n818, n1492 );
xor U9081 ( n1492, n817, n420 );
nand U9082 ( n1045, n1357, n1358 );
xor U9083 ( n1358, n1359, n311 );
nand U9084 ( n1383, n1263, n1536 );
xor U9085 ( n1536, n1262, n311 );
nand U9086 ( n992, n854, n1538 );
xor U9087 ( n1538, n853, n311 );
nand U9088 ( n1070, n1391, n1392 );
xor U9089 ( n1392, n1393, n190 );
nand U9090 ( n1408, n1303, n1577 );
xor U9091 ( n1577, n1302, n190 );
nand U9092 ( n1033, n892, n1579 );
xor U9093 ( n1579, n891, n190 );
nand U9094 ( n802, n803, n804 );
xor U9095 ( n804, n805, n531 );
nand U9096 ( n838, n839, n840 );
xor U9097 ( n840, n841, n420 );
nand U9098 ( n876, n877, n878 );
xor U9099 ( n878, n879, n311 );
nand U9100 ( n922, n923, n924 );
xor U9101 ( n924, n925, n190 );
buf U9102 ( n7432, n7431 );
buf U9103 ( n7444, n7443 );
buf U9104 ( n7456, n7455 );
buf U9105 ( n7468, n7467 );
buf U9106 ( n7429, n7428 );
buf U9107 ( n7453, n7452 );
not U9108 ( n506, n805 );
not U9109 ( n398, n841 );
not U9110 ( n289, n879 );
not U9111 ( n168, n925 );
buf U9112 ( g6837, n7476 );
buf U9113 ( g6573, n7482 );
buf U9114 ( g6368, n7488 );
buf U9115 ( g6231, n7494 );
buf U9116 ( g7084, n7473 );
buf U9117 ( g6782, n7479 );
buf U9118 ( n7466, n7464 );
buf U9119 ( g6518, n7485 );
buf U9120 ( g6313, n7491 );
and U9121 ( n2082, n2104, n2105 );
nand U9122 ( n2105, n2106, n1678 );
nand U9123 ( n2104, n2107, n540 );
nor U9124 ( n2106, n7088, n1677 );
and U9125 ( n2126, n2145, n2146 );
nand U9126 ( n2146, n2147, n1700 );
nand U9127 ( n2145, n2148, n428 );
nor U9128 ( n2147, n7087, n1699 );
and U9129 ( n2167, n2182, n2183 );
nand U9130 ( n2183, n2184, n1722 );
nand U9131 ( n2182, n2185, n319 );
nor U9132 ( n2184, n7086, n1721 );
and U9133 ( n2207, n2217, n2218 );
nand U9134 ( n2218, n2219, n1742 );
nand U9135 ( n2217, n2220, n198 );
nor U9136 ( n2219, n7044, n1741 );
buf U9137 ( n7441, n7440 );
xor U9138 ( n1781, n7092, n1211 );
xor U9139 ( n1848, n7093, n1231 );
xor U9140 ( n1915, n7095, n1262 );
xor U9141 ( n1980, n7096, n1302 );
xor U9142 ( n1799, n900, n7132 );
xor U9143 ( n1864, n947, n7133 );
xor U9144 ( n1933, n991, n7140 );
xor U9145 ( n1999, n1032, n7141 );
xor U9146 ( n1778, n784, n7128 );
xor U9147 ( n1845, n817, n7129 );
xor U9148 ( n1912, n853, n7134 );
xor U9149 ( n1977, n891, n7136 );
xnor U9150 ( n1780, n7144, n509 );
xnor U9151 ( n1847, n7145, n400 );
xnor U9152 ( n1914, n7151, n291 );
xnor U9153 ( n1979, n7152, n170 );
not U9154 ( n534, n1082 );
not U9155 ( n423, n670 );
not U9156 ( n314, n706 );
buf U9157 ( n7442, n7440 );
not U9158 ( n193, n741 );
not U9159 ( n509, n1277 );
not U9160 ( n400, n1323 );
not U9161 ( n291, n1359 );
not U9162 ( n170, n1393 );
buf U9163 ( n7430, n7428 );
buf U9164 ( n7454, n7452 );
buf U9165 ( n7433, n7431 );
buf U9166 ( n7445, n7443 );
buf U9167 ( n7457, n7455 );
buf U9168 ( n7469, n7467 );
xnor U9169 ( n1804, n7149, n507 );
xnor U9170 ( n1868, n7150, n399 );
xnor U9171 ( n1938, n7153, n290 );
xnor U9172 ( n2003, n7154, n169 );
not U9173 ( n507, n1312 );
not U9174 ( n399, n1348 );
not U9175 ( n290, n1382 );
not U9176 ( n169, n1407 );
buf U9177 ( n7465, n7464 );
xnor U9178 ( n1808, n7142, n504 );
xnor U9179 ( n1872, n7143, n396 );
xnor U9180 ( n1942, n7146, n287 );
xnor U9181 ( n2009, n7147, n166 );
not U9182 ( n504, n1274 );
not U9183 ( n396, n1320 );
not U9184 ( n287, n1356 );
not U9185 ( n166, n1390 );
xor U9186 ( n2071, n2100, n2101 );
nand U9187 ( n2100, n2083, n2102 );
nand U9188 ( n2102, n2082, n524 );
xor U9189 ( n2092, n2142, n2143 );
nand U9190 ( n2142, n2127, n2144 );
nand U9191 ( n2144, n2126, n414 );
xor U9192 ( n2135, n2179, n2180 );
nand U9193 ( n2179, n2168, n2181 );
nand U9194 ( n2181, n2167, n305 );
xor U9195 ( n2176, n2213, n2215 );
nand U9196 ( n2213, n2208, n2216 );
nand U9197 ( n2216, n2207, n184 );
not U9198 ( n533, n1084 );
not U9199 ( n313, n708 );
nand U9200 ( n1092, n1093, n1083 );
nand U9201 ( n680, n681, n671 );
nand U9202 ( n717, n718, n707 );
nand U9203 ( n751, n752, n742 );
nor U9204 ( n3887, n1167, n1084 );
nor U9205 ( n3963, n1185, n672 );
nor U9206 ( n4033, n1127, n708 );
nor U9207 ( n4103, n1147, n743 );
not U9208 ( n422, n672 );
nand U9209 ( n2083, n1683, n2112 );
nand U9210 ( n2112, n2113, n2114 );
nand U9211 ( n2113, n1677, n7088 );
nand U9212 ( n2114, n2115, n119 );
nand U9213 ( n2127, n1705, n2153 );
nand U9214 ( n2153, n2154, n2155 );
nand U9215 ( n2154, n1699, n7087 );
nand U9216 ( n2155, n2156, n53 );
nand U9217 ( n2168, n1727, n2192 );
nand U9218 ( n2192, n2193, n2194 );
nand U9219 ( n2193, n1721, n7086 );
nand U9220 ( n2194, n2195, n75 );
nand U9221 ( n2208, n1748, n2226 );
nand U9222 ( n2226, n2227, n2228 );
nand U9223 ( n2227, n1741, n7044 );
nand U9224 ( n2228, n2229, n97 );
not U9225 ( n192, n743 );
xor U9226 ( n1661, n545, n1669 );
nor U9227 ( n1669, n1670, n1671 );
nor U9228 ( n1670, n1681, n1682 );
nor U9229 ( n1671, n1672, n1673 );
xor U9230 ( n1666, n432, n1691 );
nor U9231 ( n1691, n1692, n1693 );
nor U9232 ( n1692, n1703, n1704 );
nor U9233 ( n1693, n1694, n1695 );
xor U9234 ( n1688, n323, n1713 );
nor U9235 ( n1713, n1714, n1715 );
nor U9236 ( n1714, n1725, n1726 );
nor U9237 ( n1715, n1716, n1717 );
xor U9238 ( n1710, n202, n1732 );
nor U9239 ( n1732, n1733, n1734 );
nor U9240 ( n1733, n1745, n1747 );
nor U9241 ( n1734, n1735, n1736 );
nand U9242 ( n1673, n1674, n1675 );
nand U9243 ( n1674, n7088, n1679 );
nand U9244 ( n1675, n1676, n545 );
nand U9245 ( n1679, n1677, n1680 );
nand U9246 ( n1695, n1696, n1697 );
nand U9247 ( n1696, n7087, n1701 );
nand U9248 ( n1697, n1698, n432 );
nand U9249 ( n1701, n1699, n1702 );
nand U9250 ( n1717, n1718, n1719 );
nand U9251 ( n1718, n7086, n1723 );
nand U9252 ( n1719, n1720, n323 );
nand U9253 ( n1723, n1721, n1724 );
nand U9254 ( n1736, n1738, n1739 );
nand U9255 ( n1738, n7044, n1743 );
nand U9256 ( n1739, n1740, n202 );
nand U9257 ( n1743, n1741, n1744 );
not U9258 ( n512, n1093 );
not U9259 ( n403, n681 );
not U9260 ( n294, n718 );
not U9261 ( n173, n752 );
nor U9262 ( n1678, n1680, n512 );
nor U9263 ( n1700, n1702, n403 );
nor U9264 ( n1722, n1724, n294 );
nor U9265 ( n1742, n1744, n173 );
buf U9266 ( n7426, n7427 );
buf U9267 ( n7438, n7439 );
buf U9268 ( n7450, n7451 );
buf U9269 ( n7462, n7463 );
buf U9270 ( n7425, n7427 );
buf U9271 ( n7437, n7439 );
buf U9272 ( n7449, n7451 );
buf U9273 ( n7461, n7463 );
buf U9274 ( n7436, n7434 );
buf U9275 ( n7448, n7446 );
buf U9276 ( n7460, n7458 );
buf U9277 ( n7472, n7470 );
nand U9278 ( n1418, n1423, n1424 );
nor U9279 ( n1424, n1425, n1426 );
nor U9280 ( n1423, n531, n1427 );
nand U9281 ( n1425, n934, n900 );
nand U9282 ( n1462, n1467, n1468 );
nor U9283 ( n1468, n1469, n1470 );
nor U9284 ( n1467, n420, n1471 );
nand U9285 ( n1469, n978, n947 );
nand U9286 ( n1510, n1515, n1516 );
nor U9287 ( n1516, n1517, n1518 );
nor U9288 ( n1515, n311, n1519 );
nand U9289 ( n1517, n1019, n991 );
nand U9290 ( n1551, n1556, n1557 );
nor U9291 ( n1557, n1558, n1559 );
nor U9292 ( n1556, n190, n1560 );
nand U9293 ( n1558, n1055, n1032 );
nor U9294 ( n2115, n7088, n512 );
nor U9295 ( n2156, n7087, n403 );
nor U9296 ( n2195, n7086, n294 );
nor U9297 ( n2229, n7044, n173 );
nand U9298 ( n3526, n4182, n1610 );
nor U9299 ( n4182, n1094, n7215 );
nand U9300 ( n3530, n3548, n1621 );
nor U9301 ( n3548, n682, n7216 );
nand U9302 ( n3544, n3648, n1632 );
nor U9303 ( n3648, n720, n7214 );
nand U9304 ( n3643, n3747, n1640 );
nor U9305 ( n3747, n753, n7217 );
and U9306 ( n1753, n1814, n1815 );
nand U9307 ( n1814, n528, n7215 );
nand U9308 ( n1815, n1104, n1437 );
and U9309 ( n1762, n1877, n1878 );
nand U9310 ( n1877, n417, n7216 );
nand U9311 ( n1878, n692, n1482 );
and U9312 ( n1831, n1948, n1949 );
nand U9313 ( n1948, n308, n7214 );
nand U9314 ( n1949, n730, n1529 );
and U9315 ( n1896, n2014, n2015 );
nand U9316 ( n2014, n187, n7217 );
nand U9317 ( n2015, n763, n1570 );
buf U9318 ( n7435, n7434 );
buf U9319 ( n7447, n7446 );
buf U9320 ( n7459, n7458 );
buf U9321 ( n7471, n7470 );
xor U9322 ( n3354, n3365, n3366 );
nor U9323 ( n3366, n7215, n3367 );
nand U9324 ( n3367, n2744, n2743 );
xor U9325 ( n3362, n3402, n3403 );
nor U9326 ( n3403, n7216, n3404 );
nand U9327 ( n3404, n2767, n2766 );
xor U9328 ( n3385, n3440, n3441 );
nor U9329 ( n3441, n7214, n3442 );
nand U9330 ( n3442, n2788, n2787 );
xor U9331 ( n3422, n3478, n3479 );
nor U9332 ( n3479, n7217, n3480 );
nand U9333 ( n3480, n2804, n2803 );
nand U9334 ( n2744, n3372, n3373 );
nand U9335 ( n3372, n3375, n525 );
nand U9336 ( n3373, n3374, n543 );
and U9337 ( n3375, n3365, n2750 );
nand U9338 ( n2767, n3409, n3410 );
nand U9339 ( n3409, n3412, n415 );
nand U9340 ( n3410, n3411, n431 );
and U9341 ( n3412, n3402, n2773 );
nand U9342 ( n2788, n3448, n3449 );
nand U9343 ( n3448, n3451, n306 );
nand U9344 ( n3449, n3450, n322 );
and U9345 ( n3451, n3440, n2794 );
nand U9346 ( n2804, n3486, n3487 );
nand U9347 ( n3486, n3489, n185 );
nand U9348 ( n3487, n3488, n201 );
and U9349 ( n3489, n3478, n2810 );
nor U9350 ( n3374, n525, n2750 );
nor U9351 ( n3411, n415, n2773 );
nor U9352 ( n3450, n306, n2794 );
nor U9353 ( n3488, n185, n2810 );
nor U9354 ( n2749, n2750, n2751 );
nor U9355 ( n2772, n2773, n2774 );
nor U9356 ( n2793, n2794, n2795 );
nor U9357 ( n2809, n2810, n2811 );
xor U9358 ( n2920, n7501, n3045 );
xor U9359 ( n3007, n7501, n3146 );
xor U9360 ( n3095, n7501, n3235 );
xor U9361 ( n3200, n7501, n3303 );
and U9362 ( n2886, n2985, n2986 );
nand U9363 ( n2985, n539, n2989 );
nand U9364 ( n2986, n2987, n537 );
not U9365 ( n537, n2988 );
and U9366 ( n2941, n3073, n3074 );
nand U9367 ( n3073, n427, n3077 );
nand U9368 ( n3074, n3075, n425 );
not U9369 ( n425, n3076 );
and U9370 ( n3028, n3174, n3175 );
nand U9371 ( n3174, n318, n3178 );
nand U9372 ( n3175, n3176, n316 );
not U9373 ( n316, n3177 );
and U9374 ( n3116, n3263, n3264 );
nand U9375 ( n3263, n197, n3267 );
nand U9376 ( n3264, n3265, n195 );
not U9377 ( n195, n3266 );
nor U9378 ( n2987, n539, n2989 );
nor U9379 ( n3075, n427, n3077 );
nor U9380 ( n3176, n318, n3178 );
nor U9381 ( n3265, n197, n3267 );
nand U9382 ( n4338, n6150, n6155 );
and U9383 ( n6150, n6173, n7110 );
and U9384 ( n4314, n6154, n155 );
nand U9385 ( n2860, n2918, n538 );
nor U9386 ( n2918, n2919, n2920 );
nand U9387 ( n2898, n3005, n426 );
nor U9388 ( n3005, n3006, n3007 );
nand U9389 ( n2953, n3093, n317 );
nor U9390 ( n3093, n3094, n3095 );
nand U9391 ( n3040, n3197, n196 );
nor U9392 ( n3197, n3198, n3200 );
and U9393 ( n4289, n6154, n6149 );
and U9394 ( n4317, n6149, n6150 );
and U9395 ( n4304, n6150, n6172 );
nand U9396 ( n1428, n3894, n3895 );
nor U9397 ( n3894, n1277, n1211 );
nor U9398 ( n3895, n1251, n3896 );
nand U9399 ( n3896, n504, n507 );
nand U9400 ( n1472, n3968, n3969 );
nor U9401 ( n3968, n1323, n1231 );
nor U9402 ( n3969, n1291, n3970 );
nand U9403 ( n3970, n396, n399 );
nand U9404 ( n1520, n4038, n4039 );
nor U9405 ( n4038, n1359, n1262 );
nor U9406 ( n4039, n1337, n4040 );
nand U9407 ( n4040, n287, n290 );
nand U9408 ( n1561, n4108, n4109 );
nor U9409 ( n4108, n1393, n1302 );
nor U9410 ( n4109, n1373, n4110 );
nand U9411 ( n4110, n166, n169 );
and U9412 ( n4318, n6154, n6155 );
not U9413 ( n151, n4709 );
not U9414 ( n149, n6168 );
and U9415 ( n2925, n3043, n3044 );
nand U9416 ( n3044, n2920, n2919 );
and U9417 ( n3012, n3144, n3145 );
nand U9418 ( n3145, n3007, n3006 );
and U9419 ( n3100, n3233, n3234 );
nand U9420 ( n3234, n3095, n3094 );
and U9421 ( n3205, n3301, n3302 );
nand U9422 ( n3302, n3200, n3198 );
not U9423 ( n148, n6129 );
nand U9424 ( n6162, n148, n6137 );
nand U9425 ( n1417, n3889, n3890 );
nor U9426 ( n3890, n934, n3891 );
nor U9427 ( n3889, n1428, n3893 );
nand U9428 ( n3891, n500, n503 );
nand U9429 ( n1461, n3964, n3965 );
nor U9430 ( n3965, n978, n3966 );
nor U9431 ( n3964, n1472, n3967 );
nand U9432 ( n3966, n392, n395 );
nand U9433 ( n1509, n4034, n4035 );
nor U9434 ( n4035, n1019, n4036 );
nor U9435 ( n4034, n1520, n4037 );
nand U9436 ( n4036, n283, n286 );
nand U9437 ( n1550, n4104, n4105 );
nor U9438 ( n4105, n1055, n4106 );
nor U9439 ( n4104, n1561, n4107 );
nand U9440 ( n4106, n162, n165 );
not U9441 ( n502, n934 );
not U9442 ( n394, n978 );
not U9443 ( n285, n1019 );
not U9444 ( n164, n1055 );
not U9445 ( n145, n6125 );
and U9446 ( n4313, n6153, n6149 );
and U9447 ( n4296, n6153, n6172 );
and U9448 ( n4285, n6153, n155 );
nor U9449 ( n4297, n6198, n6132 );
nand U9450 ( n6198, n7110, n149 );
nor U9451 ( n6626, n6703, n7182 );
nor U9452 ( n6431, n6508, n7156 );
nor U9453 ( n6817, n6901, n7183 );
nand U9454 ( n6600, n6626, n6627 );
nand U9455 ( n6627, n6628, n6629 );
nand U9456 ( n6629, n4441, n452 );
nor U9457 ( n6628, n6630, n6631 );
nand U9458 ( n6406, n6431, n6432 );
nand U9459 ( n6432, n6433, n6434 );
nand U9460 ( n6434, n4490, n343 );
nor U9461 ( n6433, n6435, n6436 );
nand U9462 ( n6792, n6817, n6818 );
nand U9463 ( n6818, n6819, n6820 );
nand U9464 ( n6820, n4398, n567 );
nor U9465 ( n6819, n6821, n6822 );
nand U9466 ( n6219, n6238, n6286 );
nand U9467 ( n6286, n6287, n6288 );
nand U9468 ( n6288, n4535, n224 );
nor U9469 ( n6287, n6289, n6290 );
not U9470 ( n541, n1434 );
not U9471 ( n429, n1478 );
not U9472 ( n320, n1526 );
not U9473 ( n199, n1567 );
nand U9474 ( n6607, n6626, n6671 );
nand U9475 ( n6671, n6672, n6673 );
nand U9476 ( n6672, n479, n452 );
nand U9477 ( n6673, n453, n6674 );
nand U9478 ( n6603, n6626, n6647 );
nand U9479 ( n6647, n6648, n6649 );
nand U9480 ( n6649, n4447, n452 );
nor U9481 ( n6648, n6630, n6650 );
nand U9482 ( n6408, n6431, n6452 );
nand U9483 ( n6452, n6453, n6454 );
nand U9484 ( n6454, n4496, n343 );
nor U9485 ( n6453, n6435, n6455 );
nand U9486 ( n6798, n6817, n6865 );
nand U9487 ( n6865, n6866, n6868 );
nand U9488 ( n6866, n597, n567 );
nand U9489 ( n6868, n568, n6869 );
nand U9490 ( n6794, n6817, n6838 );
nand U9491 ( n6838, n6839, n6841 );
nand U9492 ( n6841, n4404, n567 );
nor U9493 ( n6839, n6821, n6842 );
nand U9494 ( n6791, n6817, n6829 );
nand U9495 ( n6829, n6830, n6831 );
nand U9496 ( n6830, n600, n570 );
nand U9497 ( n6831, n569, n6832 );
nand U9498 ( n6599, n6626, n6638 );
nand U9499 ( n6638, n6639, n6640 );
nand U9500 ( n6639, n481, n455 );
nand U9501 ( n6640, n454, n6641 );
nand U9502 ( n6405, n6431, n6443 );
nand U9503 ( n6443, n6444, n6445 );
nand U9504 ( n6444, n373, n346 );
nand U9505 ( n6445, n345, n6446 );
nand U9506 ( n6221, n6238, n6308 );
nand U9507 ( n6308, n6309, n6310 );
nand U9508 ( n6309, n262, n224 );
nand U9509 ( n6310, n225, n6311 );
nand U9510 ( n6218, n6238, n6300 );
nand U9511 ( n6300, n6301, n6302 );
nand U9512 ( n6302, n4529, n224 );
nor U9513 ( n6301, n6289, n6303 );
nand U9514 ( n6609, n6626, n6693 );
nand U9515 ( n6693, n6694, n6695 );
or U9516 ( n6694, n4436, n2385 );
nand U9517 ( n6695, n454, n4436 );
nand U9518 ( n6800, n6817, n6890 );
nand U9519 ( n6890, n6891, n6892 );
or U9520 ( n6891, n4393, n2273 );
nand U9521 ( n6892, n569, n4393 );
nand U9522 ( n6793, n6817, n6854 );
nand U9523 ( n6854, n6855, n6856 );
nand U9524 ( n6855, n596, n567 );
nand U9525 ( n6856, n568, n4392 );
nand U9526 ( n6602, n6626, n6661 );
nand U9527 ( n6661, n6662, n6663 );
nand U9528 ( n6662, n478, n452 );
nand U9529 ( n6663, n453, n4435 );
nand U9530 ( n6407, n6431, n6466 );
nand U9531 ( n6466, n6467, n6468 );
nand U9532 ( n6467, n370, n343 );
nand U9533 ( n6468, n344, n4484 );
and U9534 ( n4290, n6173, n6167 );
and U9535 ( n4335, n6166, n6167 );
nor U9536 ( n6166, n6168, n7112 );
nand U9537 ( n6213, n6238, n6239 );
nand U9538 ( n6239, n6240, n6241 );
nand U9539 ( n6240, n263, n223 );
nand U9540 ( n6241, n222, n6242 );
nand U9541 ( n6220, n6238, n6320 );
nand U9542 ( n6320, n6321, n6322 );
nand U9543 ( n6321, n261, n224 );
nand U9544 ( n6322, n225, n4523 );
nand U9545 ( n6799, n6817, n6908 );
nand U9546 ( n6908, n6909, n6910 );
nand U9547 ( n6909, n599, n570 );
nand U9548 ( n6910, n569, n6911 );
nand U9549 ( n6608, n6626, n6709 );
nand U9550 ( n6709, n6710, n6711 );
nand U9551 ( n6710, n480, n455 );
nand U9552 ( n6711, n454, n6712 );
nand U9553 ( n6212, n6238, n6255 );
nand U9554 ( n6255, n6256, n6257 );
nand U9555 ( n6257, n265, n223 );
nor U9556 ( n6256, n6247, n6258 );
nand U9557 ( n6215, n6238, n6274 );
nand U9558 ( n6274, n6275, n6276 );
or U9559 ( n6275, n4524, n2609 );
nand U9560 ( n6276, n222, n4524 );
nand U9561 ( n6412, n6431, n6476 );
nand U9562 ( n6476, n6477, n6478 );
nand U9563 ( n6477, n371, n343 );
nand U9564 ( n6478, n344, n6479 );
nand U9565 ( n6214, n6238, n6265 );
nand U9566 ( n6265, n6266, n6267 );
nand U9567 ( n6266, n264, n223 );
nand U9568 ( n6267, n222, n6268 );
nand U9569 ( n6414, n6431, n6514 );
nand U9570 ( n6514, n6515, n6516 );
nand U9571 ( n6515, n372, n346 );
nand U9572 ( n6516, n345, n6517 );
not U9573 ( n503, n900 );
not U9574 ( n395, n947 );
not U9575 ( n286, n991 );
not U9576 ( n165, n1032 );
nand U9577 ( n6413, n6431, n6498 );
nand U9578 ( n6498, n6499, n6500 );
or U9579 ( n6499, n4485, n2500 );
nand U9580 ( n6500, n345, n4485 );
not U9581 ( n501, n784 );
not U9582 ( n393, n817 );
not U9583 ( n284, n853 );
not U9584 ( n163, n891 );
not U9585 ( n155, n6126 );
nand U9586 ( n1426, n805, n784 );
nand U9587 ( n1470, n841, n817 );
nand U9588 ( n1518, n879, n853 );
nand U9589 ( n1559, n925, n891 );
nand U9590 ( n6226, n6238, n6292 );
nand U9591 ( n6292, n6293, n6294 );
nand U9592 ( n6294, n4518, n224 );
nor U9593 ( n6293, n6289, n6295 );
nor U9594 ( n6223, n6224, n7224 );
xnor U9595 ( n6224, n6225, n6226 );
nand U9596 ( n6805, n6817, n6914 );
nand U9597 ( n6914, n6915, n6916 );
nand U9598 ( n6916, n4386, n570 );
nor U9599 ( n6915, n6882, n6917 );
nand U9600 ( n6614, n6626, n6714 );
nand U9601 ( n6714, n6715, n6716 );
nand U9602 ( n6716, n4429, n455 );
nor U9603 ( n6715, n6686, n6717 );
nand U9604 ( n6419, n6431, n6519 );
nand U9605 ( n6519, n6520, n6521 );
nand U9606 ( n6521, n4478, n346 );
nor U9607 ( n6520, n6491, n6522 );
nor U9608 ( n6802, n6803, n7225 );
xnor U9609 ( n6803, n6804, n6805 );
nor U9610 ( n6611, n6612, n7226 );
xnor U9611 ( n6612, n6613, n6614 );
nor U9612 ( n6416, n6417, n7227 );
xnor U9613 ( n6417, n6418, n6419 );
not U9614 ( n41, n2883 );
not U9615 ( n35, n3025 );
not U9616 ( n40, n2917 );
not U9617 ( n38, n2938 );
not U9618 ( n37, n3004 );
not U9619 ( n34, n3092 );
not U9620 ( n32, n3113 );
not U9621 ( n31, n3196 );
not U9622 ( n42, n2859 );
not U9623 ( n39, n2897 );
not U9624 ( n36, n2952 );
not U9625 ( n33, n3039 );
nand U9626 ( n6225, n6238, n6244 );
nand U9627 ( n6244, n6245, n6246 );
nand U9628 ( n6246, n4517, n223 );
nor U9629 ( n6245, n6247, n6248 );
nand U9630 ( n6804, n6817, n6844 );
nand U9631 ( n6844, n6845, n6846 );
nand U9632 ( n6846, n4387, n567 );
nor U9633 ( n6845, n6821, n6847 );
nand U9634 ( n6613, n6626, n6652 );
nand U9635 ( n6652, n6653, n6654 );
nand U9636 ( n6654, n4430, n452 );
nor U9637 ( n6653, n6630, n6655 );
nand U9638 ( n6418, n6431, n6457 );
nand U9639 ( n6457, n6458, n6459 );
nand U9640 ( n6459, n4479, n343 );
nor U9641 ( n6458, n6435, n6460 );
nand U9642 ( n6128, n6130, n6131 );
nor U9643 ( n6130, n6125, n7110 );
nor U9644 ( n6131, n6132, n6133 );
nand U9645 ( n6133, n6134, n6135 );
nand U9646 ( n7051, n6281, n6282 );
nand U9647 ( n6281, n6243, n6226 );
nand U9648 ( n6282, n6283, n247 );
nor U9649 ( n6283, n6284, n6285 );
nand U9650 ( n7046, n6233, n6234 );
nand U9651 ( n6233, n6243, n6225 );
nand U9652 ( n6234, n6235, n247 );
nor U9653 ( n6235, n6236, n6237 );
nor U9654 ( n6229, n6327, n6315 );
nand U9655 ( n7064, n6509, n6510 );
nand U9656 ( n6509, n6456, n6419 );
nand U9657 ( n6510, n6511, n355 );
nor U9658 ( n6511, n6512, n6513 );
nand U9659 ( n7069, n6642, n6643 );
nand U9660 ( n6642, n6651, n6613 );
nand U9661 ( n6643, n6644, n464 );
nor U9662 ( n6644, n6645, n6646 );
nand U9663 ( n7059, n6447, n6448 );
nand U9664 ( n6447, n6456, n6418 );
nand U9665 ( n6448, n6449, n355 );
nor U9666 ( n6449, n6450, n6451 );
nand U9667 ( n7084, n6902, n6904 );
nand U9668 ( n6902, n6843, n6805 );
nand U9669 ( n6904, n6905, n581 );
nor U9670 ( n6905, n6906, n6907 );
nand U9671 ( n7079, n6833, n6834 );
nand U9672 ( n6833, n6843, n6804 );
nand U9673 ( n6834, n6835, n581 );
nor U9674 ( n6835, n6836, n6837 );
nand U9675 ( n7074, n6704, n6705 );
nand U9676 ( n6704, n6651, n6614 );
nand U9677 ( n6705, n6706, n464 );
nor U9678 ( n6706, n6707, n6708 );
nor U9679 ( n6808, n6913, n6901 );
nor U9680 ( n6617, n6713, n6703 );
nor U9681 ( n6422, n6518, n6508 );
not U9682 ( n49, n6136 );
not U9683 ( n228, n2639 );
nor U9684 ( n2646, n228, n2638 );
nand U9685 ( n2395, n2599, n2600 );
nand U9686 ( n2599, n2272, n2609 );
nand U9687 ( n2600, n2601, n2602 );
nor U9688 ( n2601, n2603, n2272 );
nor U9689 ( n2603, n2604, n2605 );
nor U9690 ( n2604, n2607, n2608 );
and U9691 ( n2605, n2606, n2607 );
nor U9692 ( n2676, n2677, n2650 );
nor U9693 ( n2677, n2646, n2656 );
nor U9694 ( n2670, n2628, n2671 );
nor U9695 ( n2671, n2672, n2673 );
nor U9696 ( n2673, n228, n2663 );
nor U9697 ( n2672, n229, n2676 );
nand U9698 ( n2606, n2657, n2658 );
nand U9699 ( n2658, n2628, n2659 );
nor U9700 ( n2657, n2669, n2670 );
nand U9701 ( n2659, n2660, n2661 );
nor U9702 ( n2617, n2606, n2620 );
or U9703 ( n2620, n2608, n2602 );
nor U9704 ( n2641, n2628, n2642 );
nor U9705 ( n2642, n2643, n2644 );
and U9706 ( n2643, n2651, n2635 );
nor U9707 ( n2644, n2645, n2624 );
and U9708 ( n2507, n2614, n2615 );
nand U9709 ( n2614, n224, n2272 );
nand U9710 ( n2615, n2616, n624 );
nor U9711 ( n2616, n2617, n2618 );
and U9712 ( n2602, n2621, n2622 );
nand U9713 ( n2622, n2623, n2624 );
nor U9714 ( n2621, n2640, n2641 );
nand U9715 ( n2623, n2625, n2626 );
not U9716 ( n347, n2535 );
not U9717 ( n456, n2424 );
nand U9718 ( n2497, n2553, n2554 );
nand U9719 ( n2554, n2524, n2555 );
nor U9720 ( n2553, n2565, n2566 );
nand U9721 ( n2555, n2556, n2557 );
nand U9722 ( n2382, n2442, n2443 );
nand U9723 ( n2443, n2412, n2444 );
nor U9724 ( n2442, n2454, n2455 );
nand U9725 ( n2444, n2445, n2446 );
nor U9726 ( n2542, n347, n2534 );
nor U9727 ( n2431, n456, n2423 );
nand U9728 ( n2283, n2490, n2491 );
nand U9729 ( n2490, n2272, n2500 );
nand U9730 ( n2491, n2492, n2493 );
nor U9731 ( n2492, n2494, n2272 );
nand U9732 ( n2259, n2375, n2376 );
nand U9733 ( n2375, n2272, n2385 );
nand U9734 ( n2376, n2377, n2378 );
nor U9735 ( n2377, n2379, n2272 );
nor U9736 ( n2494, n2495, n2496 );
nor U9737 ( n2495, n2498, n2499 );
and U9738 ( n2496, n2497, n2498 );
nor U9739 ( n2379, n2380, n2381 );
nor U9740 ( n2380, n2383, n2384 );
and U9741 ( n2381, n2382, n2383 );
nor U9742 ( n2566, n2524, n2567 );
nor U9743 ( n2567, n2568, n2569 );
nor U9744 ( n2569, n347, n2559 );
nor U9745 ( n2568, n348, n2572 );
nor U9746 ( n2572, n2573, n2546 );
nor U9747 ( n2573, n2542, n2552 );
nor U9748 ( n2461, n2462, n2435 );
nor U9749 ( n2462, n2431, n2441 );
nor U9750 ( n2455, n2412, n2456 );
nor U9751 ( n2456, n2457, n2458 );
nor U9752 ( n2458, n456, n2448 );
nor U9753 ( n2457, n457, n2461 );
not U9754 ( n572, n2311 );
nand U9755 ( n2269, n2329, n2330 );
nand U9756 ( n2330, n2300, n2331 );
nor U9757 ( n2329, n2341, n2342 );
nand U9758 ( n2331, n2332, n2333 );
nor U9759 ( n2318, n572, n2310 );
nor U9760 ( n2265, n2267, n2268 );
nor U9761 ( n2267, n2270, n2271 );
and U9762 ( n2268, n2269, n2270 );
nor U9763 ( n2348, n2349, n2322 );
nor U9764 ( n2349, n2318, n2328 );
nor U9765 ( n2342, n2300, n2343 );
nor U9766 ( n2343, n2344, n2345 );
nor U9767 ( n2345, n572, n2335 );
nor U9768 ( n2344, n573, n2348 );
nand U9769 ( n2251, n2262, n2263 );
nand U9770 ( n2262, n2272, n2273 );
nand U9771 ( n2263, n2264, n624 );
nor U9772 ( n2264, n2265, n2266 );
nor U9773 ( n2513, n2497, n2516 );
or U9774 ( n2516, n2499, n2493 );
nor U9775 ( n2401, n2382, n2404 );
or U9776 ( n2404, n2384, n2378 );
nor U9777 ( n2537, n2524, n2538 );
nor U9778 ( n2538, n2539, n2540 );
and U9779 ( n2539, n2547, n2531 );
nor U9780 ( n2540, n2541, n2520 );
nor U9781 ( n2426, n2412, n2427 );
nor U9782 ( n2427, n2428, n2429 );
and U9783 ( n2428, n2436, n2420 );
nor U9784 ( n2429, n2430, n2408 );
and U9785 ( n2392, n2510, n2511 );
nand U9786 ( n2510, n343, n2272 );
nand U9787 ( n2511, n2512, n624 );
nor U9788 ( n2512, n2513, n2514 );
and U9789 ( n2280, n2398, n2399 );
nand U9790 ( n2398, n452, n2272 );
nand U9791 ( n2399, n2400, n624 );
nor U9792 ( n2400, n2401, n2402 );
and U9793 ( n2493, n2517, n2518 );
nand U9794 ( n2518, n2519, n2520 );
nor U9795 ( n2517, n2536, n2537 );
nand U9796 ( n2519, n2521, n2522 );
and U9797 ( n2378, n2405, n2406 );
nand U9798 ( n2406, n2407, n2408 );
nor U9799 ( n2405, n2425, n2426 );
nand U9800 ( n2407, n2409, n2410 );
nand U9801 ( n2266, n2293, n2294 );
nand U9802 ( n2294, n2295, n2296 );
nor U9803 ( n2293, n2312, n2313 );
nand U9804 ( n2295, n2297, n2298 );
nor U9805 ( n2313, n2300, n2314 );
nor U9806 ( n2314, n2315, n2316 );
and U9807 ( n2315, n2323, n2307 );
nor U9808 ( n2316, n2317, n2296 );
and U9809 ( n2256, n2286, n2287 );
nand U9810 ( n2286, n567, n2272 );
nand U9811 ( n2287, n2288, n624 );
nor U9812 ( n2288, n2289, n2290 );
nor U9813 ( n2636, n2632, n2651 );
nor U9814 ( n2028, n7230, n2029 );
nor U9815 ( n2713, n7210, n2714 );
nor U9816 ( n2034, n7231, n2035 );
nor U9817 ( n2717, n7211, n2718 );
nor U9818 ( n2040, n7232, n2041 );
nor U9819 ( n2721, n7212, n2722 );
nor U9820 ( n2046, n7233, n2047 );
nor U9821 ( n2725, n7213, n2726 );
nor U9822 ( n3338, n7189, n3339 );
nor U9823 ( n3342, n7190, n3343 );
nor U9824 ( n3346, n7191, n3347 );
nor U9825 ( n3350, n7192, n3351 );
nor U9826 ( n2532, n2528, n2547 );
nor U9827 ( n2421, n2416, n2436 );
nor U9828 ( n2618, n2606, n2619 );
nand U9829 ( n2619, n2607, n2608 );
nor U9830 ( n2308, n2304, n2323 );
nor U9831 ( n2514, n2497, n2515 );
nand U9832 ( n2515, n2498, n2499 );
nor U9833 ( n2402, n2382, n2403 );
nand U9834 ( n2403, n2383, n2384 );
nor U9835 ( n2290, n2269, n2291 );
nand U9836 ( n2291, n2270, n2271 );
not U9837 ( n229, n2632 );
not U9838 ( n348, n2528 );
not U9839 ( n457, n2416 );
not U9840 ( n573, n2304 );
nand U9841 ( n6260, n6243, n6328 );
nand U9842 ( n6328, n6238, n6314 );
nand U9843 ( n6824, n6843, n6857 );
nand U9844 ( n6857, n6817, n6859 );
nand U9845 ( n6633, n6651, n6664 );
nand U9846 ( n6664, n6626, n6665 );
nand U9847 ( n6438, n6456, n6469 );
nand U9848 ( n6469, n6431, n6470 );
not U9849 ( n621, n4461 );
not U9850 ( n619, n4830 );
not U9851 ( n231, n2624 );
and U9852 ( n2663, n2674, n2675 );
nand U9853 ( n2674, n216, n2624 );
nand U9854 ( n2675, n2635, n231 );
not U9855 ( n350, n2520 );
not U9856 ( n459, n2408 );
and U9857 ( n2448, n2459, n2460 );
nand U9858 ( n2459, n446, n2408 );
nand U9859 ( n2460, n2420, n459 );
and U9860 ( n2559, n2570, n2571 );
nand U9861 ( n2570, n337, n2520 );
nand U9862 ( n2571, n2531, n350 );
not U9863 ( n575, n2296 );
and U9864 ( n2335, n2346, n2347 );
nand U9865 ( n2346, n560, n2296 );
nand U9866 ( n2347, n2307, n575 );
nand U9867 ( n4175, n621, n640 );
nand U9868 ( n6848, n6922, n6923 );
nor U9869 ( n6922, n6952, n6953 );
nor U9870 ( n6923, n6924, n6925 );
nand U9871 ( n6953, n6954, n600 );
nand U9872 ( n6656, n6722, n6723 );
nor U9873 ( n6722, n6752, n6753 );
nor U9874 ( n6723, n6724, n6725 );
nand U9875 ( n6753, n6754, n481 );
nand U9876 ( n6461, n6527, n6528 );
nor U9877 ( n6527, n6557, n6558 );
nor U9878 ( n6528, n6529, n6530 );
nand U9879 ( n6558, n6559, n373 );
nand U9880 ( n6823, n6848, n5070 );
nand U9881 ( n6632, n6656, n5079 );
nand U9882 ( n6437, n6461, n5088 );
nor U9883 ( n6822, n4398, n6823 );
nor U9884 ( n6631, n4441, n6632 );
nor U9885 ( n6436, n4490, n6437 );
nand U9886 ( n6925, n6926, n4406 );
nor U9887 ( n6926, n4404, n4398 );
nand U9888 ( n6725, n6726, n4449 );
nor U9889 ( n6726, n4447, n4441 );
nand U9890 ( n6530, n6531, n4498 );
nor U9891 ( n6531, n4496, n4490 );
nand U9892 ( n6924, n6939, n4403 );
nor U9893 ( n6939, n4386, n4387 );
nand U9894 ( n6724, n6739, n4446 );
nor U9895 ( n6739, n4429, n4430 );
nand U9896 ( n6529, n6544, n4495 );
nor U9897 ( n6544, n4478, n4479 );
nand U9898 ( n6259, n6332, n6333 );
nor U9899 ( n6332, n6362, n6363 );
nor U9900 ( n6333, n6334, n6335 );
nand U9901 ( n6363, n6364, n264 );
nand U9902 ( n3939, n3141, n3940 );
nand U9903 ( n4010, n3230, n3940 );
nand U9904 ( n4080, n3298, n3940 );
nand U9905 ( n3897, n3936, n3937 );
nor U9906 ( n3936, n3945, n3946 );
nor U9907 ( n3937, n3938, n3939 );
xor U9908 ( n3945, n7230, n509 );
nand U9909 ( n3971, n4007, n4008 );
nor U9910 ( n4007, n4015, n4016 );
nor U9911 ( n4008, n4009, n4010 );
xor U9912 ( n4015, n7231, n400 );
nand U9913 ( n4041, n4077, n4078 );
nor U9914 ( n4077, n4085, n4086 );
nor U9915 ( n4078, n4079, n4080 );
xor U9916 ( n4085, n7232, n291 );
nor U9917 ( new_g26144_, n3885, n3886 );
nor U9918 ( n3886, n1417, n530 );
nor U9919 ( n3885, n3897, n3898 );
nand U9920 ( n3898, n3899, n3900 );
nor U9921 ( new_g26130_, n3961, n3962 );
nor U9922 ( n3962, n1461, n419 );
nor U9923 ( n3961, n3971, n3972 );
nand U9924 ( n3972, n3973, n3974 );
nor U9925 ( new_g26120_, n4031, n4032 );
nor U9926 ( n4032, n1509, n310 );
nor U9927 ( n4031, n4041, n4042 );
nand U9928 ( n4042, n4043, n4044 );
nand U9929 ( n6291, n6259, n5097 );
nor U9930 ( n6290, n4535, n6291 );
nor U9931 ( n6842, n4404, n6823 );
nor U9932 ( n6650, n4447, n6632 );
nor U9933 ( n6455, n4496, n6437 );
nand U9934 ( n4151, n3330, n3940 );
nand U9935 ( n4111, n4148, n4149 );
nor U9936 ( n4148, n4156, n4157 );
nor U9937 ( n4149, n4150, n4151 );
xor U9938 ( n4156, n7233, n170 );
nand U9939 ( n6335, n6336, n4537 );
nor U9940 ( n6336, n4535, n4529 );
nor U9941 ( new_g26106_, n4101, n4102 );
nor U9942 ( n4102, n1550, n189 );
nor U9943 ( n4101, n4111, n4112 );
nand U9944 ( n4112, n4113, n4114 );
nand U9945 ( n6334, n6349, n4534 );
nor U9946 ( n6349, n4517, n4518 );
nor U9947 ( n6303, n4529, n6291 );
nand U9948 ( n6250, n6243, n6315 );
nand U9949 ( n6621, n6651, n6703 );
nand U9950 ( n6426, n6456, n6508 );
nand U9951 ( n6812, n6843, n6901 );
nand U9952 ( n6884, n6848, n2273 );
nand U9953 ( n6688, n6656, n2385 );
nor U9954 ( n6954, n6869, n6911 );
nor U9955 ( n6754, n6674, n6712 );
nor U9956 ( n6559, n6479, n6517 );
nor U9957 ( n6364, n6311, n6242 );
nand U9958 ( n3123, n3043, n3045 );
nand U9959 ( n3212, n3144, n3146 );
nand U9960 ( n3280, n3233, n3235 );
not U9961 ( n538, n2989 );
not U9962 ( n426, n3077 );
not U9963 ( n317, n3178 );
or U9964 ( n3043, n2919, n538 );
or U9965 ( n3144, n3006, n426 );
or U9966 ( n3233, n3094, n317 );
nand U9967 ( n6249, n6259, n2609 );
nand U9968 ( n3312, n3301, n3303 );
not U9969 ( n196, n3267 );
or U9970 ( n3301, n3198, n196 );
nand U9971 ( n6493, n6461, n2500 );
nor U9972 ( n2633, n218, n2637 );
nand U9973 ( n2637, n2638, n2639 );
nand U9974 ( n2625, n2628, n2629 );
nand U9975 ( n2629, n2630, n2631 );
nand U9976 ( n2631, n217, n2632 );
nor U9977 ( n2630, n2633, n2634 );
not U9978 ( n596, n4392 );
not U9979 ( n478, n4435 );
not U9980 ( n370, n4484 );
nand U9981 ( n2409, n2412, n2413 );
nand U9982 ( n2413, n2414, n2415 );
nand U9983 ( n2415, n447, n2416 );
nor U9984 ( n2414, n2418, n2419 );
not U9985 ( n600, n6832 );
not U9986 ( n481, n6641 );
not U9987 ( n373, n6446 );
nor U9988 ( n6821, n6848, n5070 );
nor U9989 ( n6630, n6656, n5079 );
nor U9990 ( n6435, n6461, n5088 );
nor U9991 ( n2529, n339, n2533 );
nand U9992 ( n2533, n2534, n2535 );
nor U9993 ( n2418, n448, n2422 );
nand U9994 ( n2422, n2423, n2424 );
nand U9995 ( n2521, n2524, n2525 );
nand U9996 ( n2525, n2526, n2527 );
nand U9997 ( n2527, n338, n2528 );
nor U9998 ( n2526, n2529, n2530 );
not U9999 ( n261, n4523 );
not U10000 ( n264, n6268 );
nor U10001 ( n6289, n6259, n5097 );
nor U10002 ( n1081, n1083, n1084 );
nor U10003 ( n705, n707, n708 );
xor U10004 ( n5463, n5470, n5471 );
not U10005 ( n43, n3940 );
nor U10006 ( n669, n671, n672 );
nand U10007 ( n2297, n2300, n2301 );
nand U10008 ( n2301, n2302, n2303 );
nand U10009 ( n2303, n561, n2304 );
nor U10010 ( n2302, n2305, n2306 );
nor U10011 ( n740, n742, n743 );
xor U10012 ( n5467, n5470, n5810 );
nor U10013 ( new_g26786_, n3515, n621 );
xor U10014 ( n3515, n7100, n3516 );
nor U10015 ( n3516, n3517, n7186 );
not U10016 ( n147, g25435 );
not U10017 ( n216, n2638 );
not U10018 ( n337, n2534 );
not U10019 ( n446, n2423 );
nor U10020 ( new_g25191_, n621, n4693 );
nand U10021 ( n4693, n4694, n3517 );
nand U10022 ( n4694, n4695, n7204 );
nor U10023 ( new_g23330_, n621, n4998 );
nand U10024 ( n4998, n4999, n622 );
nand U10025 ( n4999, n5000, n7097 );
nand U10026 ( n2661, n229, n2662 );
nand U10027 ( n2662, n2663, n2664 );
nand U10028 ( n2664, n2665, n217 );
nor U10029 ( n2665, n216, n2639 );
not U10030 ( n540, n1680 );
not U10031 ( n319, n1724 );
nor U10032 ( n2681, n2638, n2687 );
nand U10033 ( n2687, n2656, n2624 );
nor U10034 ( n2669, n2679, n2680 );
nor U10035 ( n2679, n2696, n2639 );
nor U10036 ( n2680, n2681, n2682 );
nor U10037 ( n2696, n2628, n2651 );
nor U10038 ( n6882, n6848, n2273 );
nor U10039 ( n6686, n6656, n2385 );
nor U10040 ( n2305, n563, n2309 );
nand U10041 ( n2309, n2310, n2311 );
nand U10042 ( n2557, n348, n2558 );
nand U10043 ( n2558, n2559, n2560 );
nand U10044 ( n2560, n2561, n338 );
nor U10045 ( n2561, n337, n2535 );
nand U10046 ( n2446, n457, n2447 );
nand U10047 ( n2447, n2448, n2449 );
nand U10048 ( n2449, n2450, n447 );
nor U10049 ( n2450, n446, n2424 );
not U10050 ( n428, n1702 );
not U10051 ( n198, n1744 );
nor U10052 ( n2353, n2310, n2359 );
nand U10053 ( n2359, n2328, n2296 );
nor U10054 ( n2341, n2351, n2352 );
nor U10055 ( n2351, n2368, n2311 );
nor U10056 ( n2352, n2353, n2354 );
nor U10057 ( n2368, n2300, n2323 );
nand U10058 ( n2333, n573, n2334 );
nand U10059 ( n2334, n2335, n2336 );
nand U10060 ( n2336, n2337, n561 );
nor U10061 ( n2337, n560, n2311 );
nor U10062 ( n2425, n2423, n2437 );
nand U10063 ( n2437, n2438, n2416 );
nand U10064 ( n2438, n2439, n2440 );
nand U10065 ( n2440, n459, n2441 );
nand U10066 ( n2439, n456, n2412 );
nor U10067 ( n2466, n2423, n2472 );
nand U10068 ( n2472, n2441, n2408 );
nor U10069 ( n2565, n2575, n2576 );
nor U10070 ( n2575, n2592, n2535 );
nor U10071 ( n2576, n2577, n2578 );
nor U10072 ( n2592, n2524, n2547 );
nor U10073 ( n2454, n2464, n2465 );
nor U10074 ( n2464, n2483, n2424 );
nor U10075 ( n2465, n2466, n2467 );
nor U10076 ( n2483, n2412, n2436 );
nor U10077 ( n2577, n2534, n2583 );
nand U10078 ( n2583, n2552, n2520 );
nor U10079 ( n2640, n2638, n2652 );
nand U10080 ( n2652, n2653, n2632 );
nand U10081 ( n2653, n2654, n2655 );
nand U10082 ( n2655, n231, n2656 );
nand U10083 ( n2654, n228, n2628 );
nor U10084 ( n6247, n6259, n2609 );
nor U10085 ( n2536, n2534, n2548 );
nand U10086 ( n2548, n2549, n2528 );
nand U10087 ( n2549, n2550, n2551 );
nand U10088 ( n2551, n350, n2552 );
nand U10089 ( n2550, n347, n2524 );
not U10090 ( n218, n2668 );
not U10091 ( n339, n2564 );
not U10092 ( n448, n2453 );
nor U10093 ( n6491, n6461, n2500 );
not U10094 ( n560, n2310 );
nor U10095 ( n2312, n2310, n2324 );
nand U10096 ( n2324, n2325, n2304 );
nand U10097 ( n2325, n2326, n2327 );
nand U10098 ( n2327, n575, n2328 );
nand U10099 ( n2326, n572, n2300 );
nor U10100 ( n2682, n2624, n2668 );
nor U10101 ( n6295, n4518, n6291 );
not U10102 ( n563, n2340 );
nor U10103 ( n2578, n2520, n2564 );
nor U10104 ( n2467, n2408, n2453 );
nor U10105 ( n2354, n2296, n2340 );
nor U10106 ( n6847, n4387, n6823 );
nor U10107 ( n6655, n4430, n6632 );
nor U10108 ( n6460, n4479, n6437 );
nor U10109 ( n6917, n4386, n6884 );
nor U10110 ( n6717, n4429, n6688 );
nor U10111 ( n6522, n4478, n6493 );
nor U10112 ( n6248, n4517, n6249 );
xor U10113 ( new_g18542_, n5933, n5934 );
xor U10114 ( new_g16566_, n5933, n6011 );
not U10115 ( n561, n2328 );
not U10116 ( n217, n2656 );
not U10117 ( n338, n2552 );
not U10118 ( n447, n2441 );
not U10119 ( n235, n1582 );
nand U10120 ( n2660, n2666, n2651 );
nand U10121 ( n2666, n2656, n2667 );
nand U10122 ( n2667, n2668, n2624 );
nand U10123 ( n2332, n2338, n2323 );
nand U10124 ( n2338, n2328, n2339 );
nand U10125 ( n2339, n2340, n2296 );
nand U10126 ( n2556, n2562, n2547 );
nand U10127 ( n2562, n2552, n2563 );
nand U10128 ( n2563, n2564, n2520 );
nand U10129 ( n2445, n2451, n2436 );
nand U10130 ( n2451, n2441, n2452 );
nand U10131 ( n2452, n2453, n2408 );
nor U10132 ( n2411, n2424, n2416 );
nor U10133 ( n2627, n2639, n2632 );
nor U10134 ( n2523, n2535, n2528 );
nor U10135 ( n2829, n7237, n2830 );
nor U10136 ( n3739, n7222, n3740 );
nor U10137 ( n2824, n7236, n2825 );
nor U10138 ( n3635, n7221, n3636 );
nor U10139 ( n2819, n7235, n2820 );
nor U10140 ( n3537, n7220, n3538 );
nor U10141 ( n3334, n7234, n3335 );
nor U10142 ( n3522, n7219, n3523 );
nor U10143 ( n4848, n7197, n4849 );
nor U10144 ( n4844, n7196, n4845 );
nor U10145 ( n4840, n7195, n4841 );
nor U10146 ( n4836, n7194, n4837 );
nor U10147 ( n2299, n2311, n2304 );
nor U10148 ( new_g28668_, n267, n2236 );
xor U10149 ( n2236, n7261, n2237 );
nor U10150 ( n2237, n2238, n7252 );
nor U10151 ( new_g28321_, n376, n2707 );
xor U10152 ( n2707, n7260, n2708 );
nor U10153 ( n2708, n2709, n7251 );
nor U10154 ( new_g28325_, n484, n2704 );
xor U10155 ( n2704, n7259, n2705 );
nor U10156 ( n2705, n2706, n7250 );
nor U10157 ( new_g28328_, n603, n2701 );
xor U10158 ( n2701, n7258, n2702 );
nor U10159 ( n2702, n2703, n7249 );
nand U10160 ( n3189, n228, n2632 );
nand U10161 ( n3244, n3189, n2624 );
not U10162 ( n601, n4403 );
not U10163 ( n482, n4446 );
nand U10164 ( n3086, n347, n2528 );
nand U10165 ( n2998, n456, n2416 );
nand U10166 ( n2911, n572, n2304 );
nand U10167 ( n3155, n3086, n2520 );
nand U10168 ( n3054, n2998, n2408 );
nand U10169 ( n2966, n2911, n2296 );
not U10170 ( n374, n4495 );
not U10171 ( n265, n4534 );
not U10172 ( n262, n6311 );
not U10173 ( n597, n6869 );
not U10174 ( n479, n6674 );
not U10175 ( n371, n6479 );
not U10176 ( n263, n6242 );
not U10177 ( n599, n6911 );
not U10178 ( n480, n6712 );
not U10179 ( n372, n6517 );
not U10180 ( n515, n5133 );
not U10181 ( n518, n5121 );
not U10182 ( n406, n5168 );
not U10183 ( n408, n5141 );
not U10184 ( n297, n5214 );
not U10185 ( n299, n5176 );
not U10186 ( n176, n5258 );
not U10187 ( n178, n5221 );
not U10188 ( n203, n2060 );
not U10189 ( n238, n2024 );
not U10190 ( n120, n3395 );
not U10191 ( n54, n3432 );
not U10192 ( n76, n3470 );
not U10193 ( n98, n3503 );
not U10194 ( n570, n2273 );
not U10195 ( n346, n2500 );
not U10196 ( n343, n5088 );
not U10197 ( n223, n2609 );
not U10198 ( n224, n5097 );
not U10199 ( n221, n2956 );
not U10200 ( n219, n3031 );
nor U10201 ( n5095, n223, n3868 );
not U10202 ( n455, n2385 );
not U10203 ( n220, n2907 );
not U10204 ( n567, n5070 );
not U10205 ( n452, n5079 );
not U10206 ( n340, n2944 );
nor U10207 ( n5086, n346, n3862 );
not U10208 ( n342, n2901 );
not U10209 ( n341, n2869 );
not U10210 ( n566, n2841 );
nor U10211 ( n5067, n570, n3844 );
not U10212 ( n565, n2837 );
not U10213 ( n564, n2851 );
nand U10214 ( n4541, new_g13110_, n7388 );
nand U10215 ( n4544, new_g13110_, n7474 );
nand U10216 ( n4552, new_g13110_, n7477 );
nand U10217 ( n4549, new_g13110_, n7398 );
nand U10218 ( n4565, new_g13110_, n7480 );
nand U10219 ( n4580, new_g13110_, n7483 );
nand U10220 ( n4570, new_g13110_, n7408 );
nand U10221 ( n4593, new_g13110_, n7486 );
nand U10222 ( n4612, new_g13110_, n7489 );
nand U10223 ( n4598, new_g13110_, n7418 );
nand U10224 ( n4625, new_g13110_, n7492 );
nand U10225 ( n4645, new_g13110_, n7495 );
not U10226 ( n158, n2271 );
not U10227 ( n450, n2847 );
not U10228 ( n451, n2863 );
not U10229 ( n449, n2889 );
nor U10230 ( n5077, n455, n3853 );
not U10231 ( n545, n7088 );
not U10232 ( n323, n7086 );
not U10233 ( n432, n7087 );
not U10234 ( n202, n7044 );
not U10235 ( n525, n2751 );
not U10236 ( n306, n2795 );
not U10237 ( n415, n2774 );
not U10238 ( n185, n2811 );
not U10239 ( n543, n3365 );
not U10240 ( n322, n3440 );
not U10241 ( n431, n3402 );
not U10242 ( n201, n3478 );
not U10243 ( n624, n2272 );
nand U10244 ( n5487, n7097, n7186 );
nor U10245 ( n1683, n2101, n7215 );
nor U10246 ( n1727, n2180, n7214 );
nor U10247 ( n4767, n2607, n624 );
nor U10248 ( n4739, n2498, n624 );
nor U10249 ( n4720, n2383, n624 );
nor U10250 ( n4712, n2270, n624 );
nor U10251 ( n1705, n2143, n7216 );
nor U10252 ( n1748, n2215, n7217 );
nor U10253 ( n4174, n7099, n7187 );
nor U10254 ( n4696, n7097, n5000 );
or U10255 ( n3517, n4695, n7204 );
nor U10256 ( n5426, n7187, n5431 );
nor U10257 ( n4367, n7172, n5691 );
nor U10258 ( n4364, n7178, n5691 );
nor U10259 ( n4410, n7173, n5731 );
nor U10260 ( n4371, n7177, n5731 );
nor U10261 ( n4453, n7174, n5765 );
nor U10262 ( n4414, n7176, n5765 );
nor U10263 ( n4502, n7180, n5791 );
nor U10264 ( n4457, n7181, n5791 );
not U10265 ( n524, n1672 );
not U10266 ( n305, n1716 );
nor U10267 ( n4407, n5691, n7163 );
nor U10268 ( n4450, n5731, n7164 );
nor U10269 ( n4499, n5765, n7165 );
nor U10270 ( n4538, n5791, n7170 );
not U10271 ( n414, n1694 );
not U10272 ( n184, n1735 );
not U10273 ( n241, n3869 );
not U10274 ( n410, n5126 );
not U10275 ( n301, n5146 );
not U10276 ( n180, n5181 );
not U10277 ( n520, n5116 );
nor U10278 ( n4688, n7106, n4993 );
or U10279 ( n3512, n4687, n7241 );
and U10280 ( n4792, n2608, n2272 );
and U10281 ( n4764, n2499, n2272 );
and U10282 ( n4736, n2384, n2272 );
nand U10283 ( n5435, n5813, n5814 );
nor U10284 ( n5814, n5815, n5816 );
nor U10285 ( n5813, n5817, n5818 );
nand U10286 ( n5815, n7106, n7223 );
nor U10287 ( n4826, n5435, n7238 );
nand U10288 ( n6227, n6396, n7224 );
nand U10289 ( n6396, n7104, n7205 );
nand U10290 ( n6806, n7002, n7225 );
nand U10291 ( n7002, n7101, n7208 );
nand U10292 ( n6615, n6782, n7226 );
nand U10293 ( n6782, n7102, n7209 );
nand U10294 ( n6420, n6589, n7227 );
nand U10295 ( n6589, n7103, n7207 );
nand U10296 ( n6327, n6397, n7205 );
nand U10297 ( n6397, n7224, n7104 );
nand U10298 ( n6913, n7003, n7208 );
nand U10299 ( n7003, n7225, n7101 );
nand U10300 ( n6713, n6783, n7209 );
nand U10301 ( n6783, n7226, n7102 );
nand U10302 ( n6518, n6590, n7207 );
nand U10303 ( n6590, n7227, n7103 );
nand U10304 ( n3509, n5435, n7246 );
not U10305 ( n2, n4824 );
and U10306 ( n3858, n3867, n223 );
nor U10307 ( n3867, n3868, n7205 );
and U10308 ( n3849, n3861, n346 );
nor U10309 ( n3861, n3862, n7207 );
and U10310 ( n3835, n3843, n570 );
nor U10311 ( n3843, n3844, n7208 );
nor U10312 ( new_g25201_, n3509, n4685 );
nand U10313 ( n4685, n4686, n3512 );
nand U10314 ( n4686, n4687, n7241 );
and U10315 ( n3840, n3852, n455 );
nor U10316 ( n3852, n3853, n7209 );
not U10317 ( n243, n2053 );
nand U10318 ( new_g21989_, n4824, n5432 );
nand U10319 ( n5432, n5433, n7 );
nand U10320 ( n5433, n7238, n5435 );
nor U10321 ( new_g23358_, n3509, n4991 );
nand U10322 ( n4991, n4992, n5 );
nand U10323 ( n4992, n4993, n7106 );
nand U10324 ( new_g20825_, n1, n5811 );
nand U10325 ( n5811, n5812, n4994 );
not U10326 ( n1, n3509 );
nand U10327 ( n5812, n7253, n7105 );
nor U10328 ( new_g20682_, n267, n5823 );
xor U10329 ( n5823, n5008, n7257 );
nor U10330 ( new_g20717_, n376, n5822 );
xor U10331 ( n5822, n5460, n7256 );
nor U10332 ( new_g20752_, n484, n5821 );
xor U10333 ( n5821, n5449, n7255 );
nor U10334 ( new_g20789_, n603, n5820 );
xor U10335 ( n5820, n5444, n7254 );
not U10336 ( n267, n2828 );
not U10337 ( n376, n2823 );
not U10338 ( n484, n2818 );
not U10339 ( n603, n3333 );
not U10340 ( n628, n5069 );
not U10341 ( n242, n3879 );
not U10342 ( n269, n5641 );
not U10343 ( n605, n5521 );
not U10344 ( n486, n5552 );
not U10345 ( n378, n5594 );
not U10346 ( n259, n5708 );
not U10347 ( n594, n5571 );
not U10348 ( n476, n5619 );
not U10349 ( n368, n5664 );
nand U10350 ( n808, n5150, n5151 );
or U10351 ( n5151, n7436, g2247 );
nor U10352 ( n5150, n5152, n5153 );
nor U10353 ( n5152, g2249, n7113 );
nand U10354 ( n844, n5196, n5197 );
or U10355 ( n5197, n7448, g1553 );
nor U10356 ( n5196, n5198, n5199 );
nor U10357 ( n5198, g1555, n7114 );
nand U10358 ( n882, n5242, n5243 );
or U10359 ( n5243, n7460, g859 );
nor U10360 ( n5242, n5244, n5245 );
nor U10361 ( n5244, g861, n7115 );
nand U10362 ( n928, n5286, n5287 );
or U10363 ( n5287, n7472, g171 );
nor U10364 ( n5286, n5288, n5289 );
nor U10365 ( n5288, g173, n7116 );
nor U10366 ( n5153, g2248, n7117 );
nor U10367 ( n5199, g1554, n7118 );
nor U10368 ( n5245, g860, n7119 );
nor U10369 ( n5289, g172, n7120 );
nand U10370 ( new_g30638_, n1040, n1041 );
nand U10371 ( n1040, g909, n7119 );
nand U10372 ( n1041, g6368, n998 );
nand U10373 ( new_g30647_, n996, n997 );
nand U10374 ( n996, g915, n7459 );
nand U10375 ( n997, n7412, n998 );
nand U10376 ( new_g30635_, n1065, n1066 );
nand U10377 ( n1065, g222, n7120 );
nand U10378 ( n1066, g6231, n1039 );
nand U10379 ( new_g30639_, n1037, n1038 );
nand U10380 ( n1037, g228, n7471 );
nand U10381 ( n1038, n7422, n1039 );
buf U10382 ( n7476, n6161 );
buf U10383 ( n7482, n4460 );
buf U10384 ( n7488, n2759 );
buf U10385 ( n7494, n1058 );
nand U10386 ( new_g30695_, n765, n766 );
nand U10387 ( n765, g2276, n7436 );
nand U10388 ( n766, n7394, n767 );
nand U10389 ( new_g30665_, n905, n906 );
nand U10390 ( n905, g2303, n7435 );
nand U10391 ( n906, n7392, n907 );
nand U10392 ( new_g30692_, n773, n774 );
nand U10393 ( n773, g1582, n7448 );
nand U10394 ( n774, n7404, n775 );
nand U10395 ( new_g30656_, n952, n953 );
nand U10396 ( n952, g1609, n7447 );
nand U10397 ( n953, n7402, n954 );
nand U10398 ( new_g30687_, n793, n794 );
nand U10399 ( n793, g888, n7460 );
nand U10400 ( n794, n7414, n795 );
nand U10401 ( new_g30680_, n826, n827 );
nand U10402 ( n826, g201, n7472 );
nand U10403 ( n827, n7424, n828 );
nand U10404 ( new_g30690_, n778, n779 );
nand U10405 ( n778, g2270, n7117 );
nand U10406 ( n779, g6837, n767 );
nand U10407 ( new_g30693_, n771, n772 );
nand U10408 ( n771, g2273, n7113 );
nand U10409 ( n772, g7084, n767 );
nand U10410 ( new_g30652_, n963, n964 );
nand U10411 ( n963, g2297, n7117 );
nand U10412 ( n964, g6837, n907 );
nand U10413 ( new_g30659_, n940, n941 );
nand U10414 ( n940, g2300, n7113 );
nand U10415 ( n941, g7084, n907 );
nand U10416 ( new_g30683_, n811, n812 );
nand U10417 ( n811, g1576, n7118 );
nand U10418 ( n812, g6573, n775 );
nand U10419 ( new_g30688_, n791, n792 );
nand U10420 ( n791, g1579, n7114 );
nand U10421 ( n792, g6782, n775 );
nand U10422 ( new_g30644_, n1004, n1005 );
nand U10423 ( n1004, g1603, n7118 );
nand U10424 ( n1005, g6573, n954 );
nand U10425 ( new_g30650_, n984, n985 );
nand U10426 ( n984, g1606, n7114 );
nand U10427 ( n985, g6782, n954 );
nand U10428 ( new_g30676_, n847, n848 );
nand U10429 ( n847, g882, n7119 );
nand U10430 ( n848, g6368, n795 );
nand U10431 ( new_g30681_, n824, n825 );
nand U10432 ( n824, g885, n7115 );
nand U10433 ( n825, g6518, n795 );
nand U10434 ( new_g30642_, n1025, n1026 );
nand U10435 ( n1025, g912, n7115 );
nand U10436 ( n1026, g6518, n998 );
nand U10437 ( new_g30668_, n885, n886 );
nand U10438 ( n885, g195, n7120 );
nand U10439 ( n886, g6231, n828 );
nand U10440 ( new_g30674_, n860, n861 );
nand U10441 ( n860, g198, n7116 );
nand U10442 ( n861, g6313, n828 );
nand U10443 ( new_g30636_, n1063, n1064 );
nand U10444 ( n1063, g225, n7116 );
nand U10445 ( n1064, g6313, n1039 );
buf U10446 ( n7473, n6165 );
buf U10447 ( n7479, n4464 );
buf U10448 ( n7485, n2763 );
buf U10449 ( n7491, n1062 );
nor U10450 ( n902, g2180, n125 );
nor U10451 ( n938, g2170, n125 );
nor U10452 ( n949, g1486, n59 );
nor U10453 ( n982, g1476, n59 );
nor U10454 ( n993, g797, n81 );
nor U10455 ( n1023, g789, n81 );
nor U10456 ( n1034, g109, n103 );
nor U10457 ( n1060, g101, n103 );
nand U10458 ( new_g30679_, n829, n830 );
nand U10459 ( n829, g2321, n7435 );
nand U10460 ( n830, n831, n7392 );
nand U10461 ( new_g30694_, n768, n769 );
nand U10462 ( n768, g2348, n7435 );
nand U10463 ( n769, n770, n7392 );
nand U10464 ( new_g30671_, n867, n868 );
nand U10465 ( n867, g1627, n7447 );
nand U10466 ( n868, n869, n7402 );
nand U10467 ( new_g30689_, n788, n789 );
nand U10468 ( n788, g1654, n7447 );
nand U10469 ( n789, n790, n7402 );
nand U10470 ( new_g30662_, n913, n914 );
nand U10471 ( n913, g933, n7459 );
nand U10472 ( n914, n915, n7412 );
nand U10473 ( new_g30682_, n821, n822 );
nand U10474 ( n821, g960, n7459 );
nand U10475 ( n822, n823, n7412 );
nand U10476 ( new_g30653_, n960, n961 );
nand U10477 ( n960, g246, n7471 );
nand U10478 ( n961, n962, n7422 );
nand U10479 ( new_g30675_, n857, n858 );
nand U10480 ( n857, g273, n7471 );
nand U10481 ( n858, n859, n7422 );
nand U10482 ( new_g30672_, n864, n865 );
nand U10483 ( n864, g2312, n7435 );
nand U10484 ( n865, n866, n7394 );
nand U10485 ( new_g30663_, n910, n911 );
nand U10486 ( n910, g1618, n7447 );
nand U10487 ( n911, n912, n7404 );
nand U10488 ( new_g30654_, n957, n958 );
nand U10489 ( n957, g924, n7459 );
nand U10490 ( n958, n959, n7414 );
nand U10491 ( new_g30645_, n1001, n1002 );
nand U10492 ( n1001, g237, n7471 );
nand U10493 ( n1002, n1003, n7424 );
nand U10494 ( new_g30667_, n895, n896 );
nand U10495 ( n895, g2315, n7117 );
nand U10496 ( n896, n831, n7477 );
nand U10497 ( new_g30673_, n862, n863 );
nand U10498 ( n862, g2318, n7113 );
nand U10499 ( n863, n831, n7474 );
nand U10500 ( new_g30660_, n929, n930 );
nand U10501 ( n929, g2306, n7117 );
nand U10502 ( n930, n866, n7477 );
nand U10503 ( new_g30666_, n903, n904 );
nand U10504 ( n903, g2309, n7113 );
nand U10505 ( n904, n866, n7474 );
nand U10506 ( new_g30686_, n796, n797 );
nand U10507 ( n796, g2342, n7117 );
nand U10508 ( n797, n770, n7477 );
nand U10509 ( new_g30691_, n776, n777 );
nand U10510 ( n776, g2345, n7113 );
nand U10511 ( n777, n770, n7474 );
nand U10512 ( new_g30658_, n942, n943 );
nand U10513 ( n942, g1621, n7118 );
nand U10514 ( n943, n869, n7483 );
nand U10515 ( new_g30664_, n908, n909 );
nand U10516 ( n908, g1624, n7114 );
nand U10517 ( n909, n869, n7480 );
nand U10518 ( new_g30651_, n973, n974 );
nand U10519 ( n973, g1612, n7118 );
nand U10520 ( n974, n912, n7483 );
nand U10521 ( new_g30657_, n950, n951 );
nand U10522 ( n950, g1615, n7114 );
nand U10523 ( n951, n912, n7480 );
nand U10524 ( new_g30678_, n832, n833 );
nand U10525 ( n832, g1648, n7118 );
nand U10526 ( n833, n790, n7483 );
nand U10527 ( new_g30684_, n809, n810 );
nand U10528 ( n809, g1651, n7114 );
nand U10529 ( n810, n790, n7480 );
nand U10530 ( new_g30649_, n986, n987 );
nand U10531 ( n986, g927, n7119 );
nand U10532 ( n987, n915, n7489 );
nand U10533 ( new_g30655_, n955, n956 );
nand U10534 ( n955, g930, n7115 );
nand U10535 ( n956, n915, n7486 );
nand U10536 ( new_g30643_, n1014, n1015 );
nand U10537 ( n1014, g918, n7119 );
nand U10538 ( n1015, n959, n7489 );
nand U10539 ( new_g30648_, n994, n995 );
nand U10540 ( n994, g921, n7115 );
nand U10541 ( n995, n959, n7486 );
nand U10542 ( new_g30670_, n870, n871 );
nand U10543 ( n870, g954, n7119 );
nand U10544 ( n871, n823, n7489 );
nand U10545 ( new_g30677_, n845, n846 );
nand U10546 ( n845, g957, n7115 );
nand U10547 ( n846, n823, n7486 );
nand U10548 ( new_g30641_, n1027, n1028 );
nand U10549 ( n1027, g240, n7120 );
nand U10550 ( n1028, n962, n7495 );
nand U10551 ( new_g30646_, n999, n1000 );
nand U10552 ( n999, g243, n7116 );
nand U10553 ( n1000, n962, n7492 );
nand U10554 ( new_g30637_, n1050, n1051 );
nand U10555 ( n1050, g231, n7120 );
nand U10556 ( n1051, n1003, n7495 );
nand U10557 ( new_g30640_, n1035, n1036 );
nand U10558 ( n1035, g234, n7116 );
nand U10559 ( n1036, n1003, n7492 );
nand U10560 ( new_g30661_, n916, n917 );
nand U10561 ( n916, g267, n7120 );
nand U10562 ( n917, n859, n7495 );
nand U10563 ( new_g30669_, n883, n884 );
nand U10564 ( n883, g270, n7116 );
nand U10565 ( n884, n859, n7492 );
nor U10566 ( n5188, g2251, n7117 );
nor U10567 ( n5235, g1557, n7118 );
nor U10568 ( n5278, g863, n7119 );
nor U10569 ( n5323, g175, n7120 );
nand U10570 ( n1822, n5185, n5186 );
or U10571 ( n5186, n7436, g2250 );
nor U10572 ( n5185, n5187, n5188 );
nor U10573 ( n5187, g2252, n7113 );
nand U10574 ( n1886, n5232, n5233 );
or U10575 ( n5233, n7448, g1556 );
nor U10576 ( n5232, n5234, n5235 );
nor U10577 ( n5234, g1558, n7114 );
nand U10578 ( n1957, n5275, n5276 );
or U10579 ( n5276, n7460, g862 );
nor U10580 ( n5275, n5277, n5278 );
nor U10581 ( n5277, g864, n7115 );
nand U10582 ( n2022, n5319, n5320 );
or U10583 ( n5320, n7472, g174 );
nor U10584 ( n5319, n5322, n5323 );
nor U10585 ( n5322, g176, n7116 );
xor U10586 ( n4199, n7132, n4200 );
nor U10587 ( n4200, n4201, n4202 );
nor U10588 ( n4201, g2220, n7435 );
nand U10589 ( n4202, n4203, n4204 );
xor U10590 ( n3565, n7133, n3566 );
nor U10591 ( n3566, n3567, n3568 );
nor U10592 ( n3567, g1526, n7447 );
nand U10593 ( n3568, n3569, n3570 );
xor U10594 ( n3667, n7140, n3668 );
nor U10595 ( n3668, n3669, n3670 );
nor U10596 ( n3669, g832, n7459 );
nand U10597 ( n3670, n3671, n3672 );
xor U10598 ( n3766, n7141, n3767 );
nor U10599 ( n3767, n3768, n3769 );
nor U10600 ( n3768, g144, n7471 );
nand U10601 ( n3769, n3770, n3771 );
nand U10602 ( n4190, n4191, n4192 );
xor U10603 ( n4192, g2195, n4193 );
nor U10604 ( n4191, n4198, n4199 );
nor U10605 ( n4193, n4194, n4195 );
nand U10606 ( n3556, n3557, n3558 );
xor U10607 ( n3558, g1501, n3559 );
nor U10608 ( n3557, n3564, n3565 );
nor U10609 ( n3559, n3560, n3561 );
nand U10610 ( n3657, n3658, n3659 );
xor U10611 ( n3659, g809, n3660 );
nor U10612 ( n3658, n3666, n3667 );
nor U10613 ( n3660, n3661, n3662 );
nand U10614 ( n3756, n3757, n3758 );
xor U10615 ( n3758, g121, n3759 );
nor U10616 ( n3757, n3765, n3766 );
nor U10617 ( n3759, n3760, n3761 );
or U10618 ( n4204, n7113, g2222 );
or U10619 ( n3570, n7114, g1528 );
or U10620 ( n3672, n7115, g834 );
or U10621 ( n3771, n7116, g146 );
or U10622 ( n4203, n7117, g2221 );
or U10623 ( n3569, n7118, g1527 );
or U10624 ( n3671, n7119, g833 );
or U10625 ( n3770, n7120, g145 );
xor U10626 ( n4198, n7124, n4205 );
nor U10627 ( n4205, n4206, n4207 );
nor U10628 ( n4206, g2208, n7435 );
nand U10629 ( n4207, n4208, n4209 );
xor U10630 ( n3564, n7125, n3571 );
nor U10631 ( n3571, n3572, n3573 );
nor U10632 ( n3572, g1514, n7447 );
nand U10633 ( n3573, n3574, n3575 );
xor U10634 ( n3666, n7126, n3673 );
nor U10635 ( n3673, n3675, n3676 );
nor U10636 ( n3675, g820, n7459 );
nand U10637 ( n3676, n3677, n3678 );
xor U10638 ( n3765, n7127, n3772 );
nor U10639 ( n3772, n3774, n3775 );
nor U10640 ( n3774, g132, n7471 );
nand U10641 ( n3775, n3776, n3777 );
or U10642 ( n4209, n7113, g2210 );
or U10643 ( n3575, n7114, g1516 );
or U10644 ( n3678, n7115, g822 );
or U10645 ( n3777, n7116, g134 );
nor U10646 ( n4219, n4220, n4221 );
nor U10647 ( n4220, g2217, n7435 );
nand U10648 ( n4221, n4222, n4223 );
or U10649 ( n4222, n7117, g2218 );
nor U10650 ( n3586, n3587, n3588 );
nor U10651 ( n3587, g1523, n7447 );
nand U10652 ( n3588, n3589, n3590 );
or U10653 ( n3589, n7118, g1524 );
or U10654 ( n4223, n7113, g2219 );
or U10655 ( n3590, n7114, g1525 );
nor U10656 ( n3689, n3690, n3691 );
nor U10657 ( n3690, g829, n7459 );
nand U10658 ( n3691, n3693, n3694 );
or U10659 ( n3693, n7119, g830 );
nor U10660 ( n3788, n3789, n3790 );
nor U10661 ( n3789, g141, n7471 );
nand U10662 ( n3790, n3792, n3793 );
or U10663 ( n3792, n7120, g142 );
or U10664 ( n3694, n7115, g831 );
or U10665 ( n3793, n7116, g143 );
or U10666 ( n4208, n7117, g2209 );
or U10667 ( n3574, n7118, g1515 );
or U10668 ( n3677, n7119, g821 );
or U10669 ( n3776, n7120, g133 );
nor U10670 ( n4250, n4251, n4252 );
nor U10671 ( n4251, g2226, n7435 );
nand U10672 ( n4252, n4253, n4254 );
or U10673 ( n4253, n7117, g2227 );
nor U10674 ( n3621, n3622, n3623 );
nor U10675 ( n3622, g1532, n7447 );
nand U10676 ( n3623, n3624, n3625 );
or U10677 ( n3624, n7118, g1533 );
nor U10678 ( n3724, n3725, n3726 );
nor U10679 ( n3725, g838, n7459 );
nand U10680 ( n3726, n3727, n3728 );
or U10681 ( n3727, n7119, g839 );
nor U10682 ( n3822, n3823, n3824 );
nor U10683 ( n3823, g150, n7471 );
nand U10684 ( n3824, n3825, n3826 );
or U10685 ( n3825, n7120, g151 );
or U10686 ( n4254, n7113, g2228 );
or U10687 ( n3625, n7114, g1534 );
or U10688 ( n3728, n7115, g840 );
or U10689 ( n3826, n7116, g152 );
nand U10690 ( new_g30703_, n694, n695 );
nand U10691 ( n694, g1003, n7454 );
nand U10692 ( n695, n662, g6712 );
nand U10693 ( new_g30701_, n699, n700 );
nand U10694 ( n699, g1002, n7457 );
nand U10695 ( n700, n662, g5472 );
nand U10696 ( new_g30699_, n734, n735 );
nand U10697 ( n734, g315, n7469 );
nand U10698 ( n735, n698, g5437 );
nand U10699 ( new_g30700_, n732, n733 );
nand U10700 ( n732, g316, n7466 );
nand U10701 ( n733, n698, g6447 );
or U10702 ( n4226, n7339, n7340 );
nor U10703 ( n7339, n7117, g2206 );
nor U10704 ( n7340, n7113, g2207 );
or U10705 ( n3594, n7341, n7342 );
nor U10706 ( n7341, n7118, g1512 );
nor U10707 ( n7342, n7114, g1513 );
nand U10708 ( new_g30709_, n648, n649 );
nand U10709 ( n648, g2391, n7430 );
nand U10710 ( n649, n650, g7264 );
nand U10711 ( new_g30707_, n655, n656 );
nand U10712 ( n655, g2390, n7433 );
nand U10713 ( n656, n650, g5555 );
nand U10714 ( new_g30704_, n663, n664 );
nand U10715 ( n663, g1696, n7445 );
nand U10716 ( n664, n654, g5511 );
nand U10717 ( new_g30706_, n657, n658 );
nand U10718 ( n657, g1697, n7442 );
nand U10719 ( n658, n654, g7014 );
nand U10720 ( new_g30566_, n1075, n1076 );
nand U10721 ( n1075, g2392, n7425 );
nand U10722 ( n1076, n650, g2476 );
nand U10723 ( new_g30708_, n651, n653 );
nand U10724 ( n651, g1698, n7437 );
nand U10725 ( n653, n654, g1782 );
nand U10726 ( new_g30705_, n659, n660 );
nand U10727 ( n659, g1004, n7449 );
nand U10728 ( n660, n662, g1088 );
nand U10729 ( new_g30702_, n696, n697 );
nand U10730 ( n696, g317, n7461 );
nand U10731 ( n697, n698, g401 );
or U10732 ( n3698, n7343, n7344 );
nor U10733 ( n7343, n7119, g818 );
nor U10734 ( n7344, n7115, g819 );
or U10735 ( n3796, n7345, n7346 );
nor U10736 ( n7345, n7120, g130 );
nor U10737 ( n7346, n7116, g131 );
nor U10738 ( n4255, n4256, n4257 );
nor U10739 ( n4256, g2232, n7435 );
nand U10740 ( n4257, n4258, n4259 );
or U10741 ( n4258, n7117, g2233 );
nor U10742 ( n3626, n3627, n3628 );
nor U10743 ( n3627, g1538, n7447 );
nand U10744 ( n3628, n3630, n3631 );
or U10745 ( n3630, n7118, g1539 );
nor U10746 ( n3729, n3730, n3731 );
nor U10747 ( n3730, g844, n7459 );
nand U10748 ( n3731, n3732, n3734 );
or U10749 ( n3732, n7119, g845 );
nor U10750 ( n3827, n3828, n3829 );
nor U10751 ( n3828, g156, n7471 );
nand U10752 ( n3829, n3830, n3831 );
or U10753 ( n3830, n7120, g157 );
or U10754 ( n4259, n7113, g2234 );
or U10755 ( n3631, n7114, g1540 );
or U10756 ( n3734, n7115, g846 );
or U10757 ( n3831, n7116, g158 );
nor U10758 ( n1314, g2190, n783 );
nor U10759 ( n1350, g1496, n816 );
nand U10760 ( new_g30290_, n1243, n1244 );
nand U10761 ( n1243, g2330, n7436 );
nand U10762 ( n1244, n1245, n7393 );
nand U10763 ( new_g30280_, n1283, n1284 );
nand U10764 ( n1283, g1636, n7448 );
nand U10765 ( n1284, n1285, n7403 );
nand U10766 ( new_g30274_, n1307, n1308 );
nand U10767 ( n1307, g2324, n7117 );
nand U10768 ( n1308, n1245, n7477 );
nand U10769 ( new_g30282_, n1279, n1280 );
nand U10770 ( n1279, g2327, n7113 );
nand U10771 ( n1280, n1245, n7474 );
nand U10772 ( new_g30266_, n1343, n1344 );
nand U10773 ( n1343, g1630, n7118 );
nand U10774 ( n1344, n1285, n7483 );
nand U10775 ( new_g30272_, n1325, n1326 );
nand U10776 ( n1325, g1633, n7114 );
nand U10777 ( n1326, n1285, n7480 );
nor U10778 ( n1384, g805, n852 );
nor U10779 ( n1409, g117, n890 );
nor U10780 ( n4234, n4236, n4237 );
nor U10781 ( n4236, g2237, n7113 );
nor U10782 ( n4237, g2236, n7117 );
nor U10783 ( n3603, n3605, n3606 );
nor U10784 ( n3605, g1543, n7114 );
nor U10785 ( n3606, g1542, n7118 );
nor U10786 ( n3707, n3710, n3711 );
nor U10787 ( n3710, g849, n7115 );
nor U10788 ( n3711, g848, n7119 );
nor U10789 ( n3806, n3808, n3809 );
nor U10790 ( n3808, g161, n7116 );
nor U10791 ( n3809, g160, n7120 );
nand U10792 ( new_g30270_, n1329, n1330 );
nand U10793 ( n1329, g942, n7460 );
nand U10794 ( n1330, n1331, n7413 );
nand U10795 ( new_g30262_, n1365, n1366 );
nand U10796 ( n1365, g255, n7472 );
nand U10797 ( n1366, n1367, n7423 );
nand U10798 ( new_g30259_, n1377, n1378 );
nand U10799 ( n1377, g936, n7119 );
nand U10800 ( n1378, n1331, n7489 );
nand U10801 ( new_g30264_, n1361, n1362 );
nand U10802 ( n1361, g939, n7115 );
nand U10803 ( n1362, n1331, n7486 );
nand U10804 ( new_g30254_, n1402, n1403 );
nand U10805 ( n1402, g249, n7120 );
nand U10806 ( n1403, n1367, n7495 );
nand U10807 ( new_g30257_, n1395, n1396 );
nand U10808 ( n1395, g252, n7116 );
nand U10809 ( n1396, n1367, n7492 );
nor U10810 ( n1278, g2200, n783 );
nor U10811 ( n1324, g1506, n816 );
nor U10812 ( n1360, g813, n852 );
nor U10813 ( n1394, g125, n890 );
nand U10814 ( new_g30297_, n1221, n1222 );
nand U10815 ( n1221, g2339, n7436 );
nand U10816 ( n1222, n1223, n7390 );
nand U10817 ( new_g30288_, n1252, n1253 );
nand U10818 ( n1252, g1645, n7448 );
nand U10819 ( n1253, n1254, n7400 );
nand U10820 ( new_g30278_, n1292, n1293 );
nand U10821 ( n1292, g951, n7460 );
nand U10822 ( n1293, n1294, n7410 );
nand U10823 ( new_g30268_, n1338, n1339 );
nand U10824 ( n1338, g264, n7472 );
nand U10825 ( n1339, n1340, n7420 );
nand U10826 ( new_g30283_, n1269, n1270 );
nand U10827 ( n1269, g2333, n7117 );
nand U10828 ( n1270, n1223, n7477 );
nand U10829 ( new_g30291_, n1241, n1242 );
nand U10830 ( n1241, g2336, n7113 );
nand U10831 ( n1242, n1223, n7474 );
nand U10832 ( new_g30273_, n1315, n1316 );
nand U10833 ( n1315, g1639, n7118 );
nand U10834 ( n1316, n1254, n7483 );
nand U10835 ( new_g30281_, n1281, n1282 );
nand U10836 ( n1281, g1642, n7114 );
nand U10837 ( n1282, n1254, n7480 );
nand U10838 ( new_g30265_, n1351, n1352 );
nand U10839 ( n1351, g945, n7119 );
nand U10840 ( n1352, n1294, n7489 );
nand U10841 ( new_g30271_, n1327, n1328 );
nand U10842 ( n1327, g948, n7115 );
nand U10843 ( n1328, n1294, n7486 );
nand U10844 ( new_g30258_, n1385, n1386 );
nand U10845 ( n1385, g258, n7120 );
nand U10846 ( n1386, n1340, n7495 );
nand U10847 ( new_g30263_, n1363, n1364 );
nand U10848 ( n1363, g261, n7116 );
nand U10849 ( n1364, n1340, n7492 );
nand U10850 ( n1376, n1412, n1413 );
nand U10851 ( n1412, n1419, n783 );
nand U10852 ( n1413, n971, g2195 );
xor U10853 ( n1419, n1277, n1275 );
nand U10854 ( n1401, n1456, n1457 );
nand U10855 ( n1456, n1463, n816 );
nand U10856 ( n1457, n1012, g1501 );
xor U10857 ( n1463, n1323, n1321 );
nand U10858 ( n1453, n1504, n1505 );
nand U10859 ( n1504, n1511, n852 );
nand U10860 ( n1505, n1048, g809 );
xor U10861 ( n1511, n1359, n1357 );
nand U10862 ( n1501, n1545, n1546 );
nand U10863 ( n1545, n1552, n890 );
nand U10864 ( n1546, n1073, g121 );
xor U10865 ( n1552, n1393, n1391 );
nand U10866 ( new_g30260_, n1374, n1375 );
nand U10867 ( n1374, g2294, n7436 );
nand U10868 ( n1375, n7390, n1376 );
nand U10869 ( new_g30255_, n1399, n1400 );
nand U10870 ( n1399, g1600, n7448 );
nand U10871 ( n1400, n7400, n1401 );
nand U10872 ( new_g30250_, n1454, n1455 );
nand U10873 ( n1454, g1594, n7118 );
nand U10874 ( n1455, g6573, n1401 );
nand U10875 ( new_g30252_, n1449, n1450 );
nand U10876 ( n1449, g1597, n7114 );
nand U10877 ( n1450, g6782, n1401 );
nand U10878 ( n1200, n1208, n1209 );
nand U10879 ( n1208, n1210, n783 );
nand U10880 ( n1209, n971, g2185 );
xor U10881 ( n1210, n1211, n1212 );
nand U10882 ( n1205, n1228, n1229 );
nand U10883 ( n1228, n1230, n816 );
nand U10884 ( n1229, n1012, g1491 );
xor U10885 ( n1230, n1231, n1232 );
nand U10886 ( new_g30251_, n1451, n1452 );
nand U10887 ( n1451, g906, n7460 );
nand U10888 ( n1452, n7410, n1453 );
nand U10889 ( new_g30248_, n1499, n1500 );
nand U10890 ( n1499, g219, n7472 );
nand U10891 ( n1500, n7420, n1501 );
nand U10892 ( new_g30253_, n1410, n1411 );
nand U10893 ( n1410, g2288, n7117 );
nand U10894 ( n1411, g6837, n1376 );
nand U10895 ( new_g30256_, n1397, n1398 );
nand U10896 ( n1397, g2291, n7113 );
nand U10897 ( n1398, g7084, n1376 );
nand U10898 ( new_g30247_, n1502, n1503 );
nand U10899 ( n1502, g900, n7119 );
nand U10900 ( n1503, g6368, n1453 );
nand U10901 ( new_g30249_, n1496, n1497 );
nand U10902 ( n1496, g903, n7115 );
nand U10903 ( n1497, g6518, n1453 );
nand U10904 ( n1220, n1259, n1260 );
nand U10905 ( n1259, n1261, n852 );
nand U10906 ( n1260, n1048, g801 );
xor U10907 ( n1261, n1262, n1263 );
nand U10908 ( n1240, n1299, n1300 );
nand U10909 ( n1299, n1301, n890 );
nand U10910 ( n1300, n1073, g113 );
xor U10911 ( n1301, n1302, n1303 );
nand U10912 ( n1215, n1248, n1249 );
nand U10913 ( n1248, n783, n1250 );
nand U10914 ( n1249, n971, g2165 );
xor U10915 ( n1250, n1251, n937 );
nand U10916 ( n1235, n1288, n1289 );
nand U10917 ( n1288, n816, n1290 );
nand U10918 ( n1289, n1012, g1471 );
xor U10919 ( n1290, n1291, n981 );
nor U10920 ( n4242, g2239, n7117 );
nor U10921 ( n3612, g1545, n7118 );
nand U10922 ( new_g30289_, n1246, n1247 );
nand U10923 ( n1246, g2261, n7117 );
nand U10924 ( n1247, g6837, n1215 );
nand U10925 ( new_g30296_, n1224, n1225 );
nand U10926 ( n1224, g2264, n7113 );
nand U10927 ( n1225, g7084, n1215 );
nand U10928 ( new_g30304_, n1198, n1199 );
nand U10929 ( n1198, g2285, n7436 );
nand U10930 ( n1199, n7390, n1200 );
nand U10931 ( new_g30302_, n1203, n1204 );
nand U10932 ( n1203, g1591, n7448 );
nand U10933 ( n1204, n7400, n1205 );
nand U10934 ( new_g30301_, n1206, n1207 );
nand U10935 ( n1206, g2279, n7117 );
nand U10936 ( n1207, g6837, n1200 );
nand U10937 ( new_g30303_, n1201, n1202 );
nand U10938 ( n1201, g2282, n7113 );
nand U10939 ( n1202, g7084, n1200 );
nand U10940 ( new_g30295_, n1226, n1227 );
nand U10941 ( n1226, g1585, n7118 );
nand U10942 ( n1227, g6573, n1205 );
nand U10943 ( new_g30299_, n1216, n1217 );
nand U10944 ( n1216, g1588, n7114 );
nand U10945 ( n1217, g6782, n1205 );
nand U10946 ( new_g30245_, n1543, n1544 );
nand U10947 ( n1543, g213, n7120 );
nand U10948 ( n1544, g6231, n1501 );
nand U10949 ( new_g30246_, n1541, n1542 );
nand U10950 ( n1541, g216, n7116 );
nand U10951 ( n1542, g6313, n1501 );
nand U10952 ( n1266, n1334, n1335 );
nand U10953 ( n1334, n852, n1336 );
nand U10954 ( n1335, n1048, g785 );
xor U10955 ( n1336, n1337, n1022 );
nand U10956 ( n1306, n1370, n1371 );
nand U10957 ( n1370, n890, n1372 );
nand U10958 ( n1371, n1073, g97 );
xor U10959 ( n1372, n1373, n1059 );
nor U10960 ( n3716, g851, n7119 );
nor U10961 ( n3814, g163, n7120 );
nand U10962 ( n4238, n4239, n4240 );
or U10963 ( n4240, n7436, g2238 );
nor U10964 ( n4239, n4241, n4242 );
nor U10965 ( n4241, g2240, n7113 );
nand U10966 ( n3607, n3608, n3609 );
or U10967 ( n3609, n7448, g1544 );
nor U10968 ( n3608, n3610, n3612 );
nor U10969 ( n3610, g1546, n7114 );
nand U10970 ( n3712, n3713, n3714 );
or U10971 ( n3714, n7460, g850 );
nor U10972 ( n3713, n3715, n3716 );
nor U10973 ( n3715, g852, n7115 );
nand U10974 ( n3810, n3811, n3812 );
or U10975 ( n3812, n7472, g162 );
nor U10976 ( n3811, n3813, n3814 );
nor U10977 ( n3813, g164, n7116 );
nand U10978 ( new_g30300_, n1213, n1214 );
nand U10979 ( n1213, g2267, n7436 );
nand U10980 ( n1214, n7391, n1215 );
nand U10981 ( new_g30279_, n1286, n1287 );
nand U10982 ( n1286, g1567, n7118 );
nand U10983 ( n1287, g6573, n1235 );
nand U10984 ( new_g30287_, n1255, n1256 );
nand U10985 ( n1255, g1570, n7114 );
nand U10986 ( n1256, g6782, n1235 );
nand U10987 ( new_g30294_, n1233, n1234 );
nand U10988 ( n1233, g1573, n7448 );
nand U10989 ( n1234, n7401, n1235 );
nand U10990 ( new_g30277_, n1295, n1296 );
nand U10991 ( n1295, g876, n7115 );
nand U10992 ( n1296, g6518, n1266 );
nand U10993 ( new_g30267_, n1341, n1342 );
nand U10994 ( n1341, g189, n7116 );
nand U10995 ( n1342, g6313, n1306 );
nand U10996 ( new_g30298_, n1218, n1219 );
nand U10997 ( n1218, g897, n7460 );
nand U10998 ( n1219, n7410, n1220 );
nand U10999 ( new_g30285_, n1264, n1265 );
nand U11000 ( n1264, g879, n7460 );
nand U11001 ( n1265, n7411, n1266 );
nand U11002 ( new_g30292_, n1238, n1239 );
nand U11003 ( n1238, g210, n7472 );
nand U11004 ( n1239, n7420, n1240 );
nand U11005 ( new_g30275_, n1304, n1305 );
nand U11006 ( n1304, g192, n7472 );
nand U11007 ( n1305, n7421, n1306 );
nand U11008 ( new_g30286_, n1257, n1258 );
nand U11009 ( n1257, g891, n7119 );
nand U11010 ( n1258, g6368, n1220 );
nand U11011 ( new_g30293_, n1236, n1237 );
nand U11012 ( n1236, g894, n7115 );
nand U11013 ( n1237, g6518, n1220 );
nand U11014 ( new_g30269_, n1332, n1333 );
nand U11015 ( n1332, g873, n7119 );
nand U11016 ( n1333, g6368, n1266 );
nand U11017 ( new_g30276_, n1297, n1298 );
nand U11018 ( n1297, g204, n7120 );
nand U11019 ( n1298, g6231, n1240 );
nand U11020 ( new_g30284_, n1267, n1268 );
nand U11021 ( n1267, g207, n7116 );
nand U11022 ( n1268, g6313, n1240 );
nand U11023 ( new_g30261_, n1368, n1369 );
nand U11024 ( n1368, g186, n7120 );
nand U11025 ( n1369, g6231, n1306 );
nor U11026 ( n4247, g2245, n7117 );
nor U11027 ( n3617, g1551, n7118 );
nor U11028 ( n3721, g857, n7119 );
nor U11029 ( n3819, g169, n7120 );
and U11030 ( n1178, g2257, n2116 );
and U11031 ( n1196, g1563, n2157 );
and U11032 ( n1138, g869, n2196 );
and U11033 ( n1158, g181, n2230 );
nand U11034 ( n2116, n4244, n4245 );
or U11035 ( n4245, n7436, g2244 );
nor U11036 ( n4244, n4246, n4247 );
nor U11037 ( n4246, g2246, n7113 );
nand U11038 ( n2157, n3614, n3615 );
or U11039 ( n3615, n7448, g1550 );
nor U11040 ( n3614, n3616, n3617 );
nor U11041 ( n3616, g1552, n7114 );
nand U11042 ( n2196, n3718, n3719 );
or U11043 ( n3719, n7460, g856 );
nor U11044 ( n3718, n3720, n3721 );
nor U11045 ( n3720, g858, n7115 );
nand U11046 ( n2230, n3816, n3817 );
or U11047 ( n3817, n7472, g168 );
nor U11048 ( n3816, n3818, n3819 );
nor U11049 ( n3818, g170, n7116 );
or U11050 ( n4195, n7347, n7348 );
nor U11051 ( n7347, n7117, g2230 );
nor U11052 ( n7348, n7113, g2231 );
or U11053 ( n3561, n7349, n7350 );
nor U11054 ( n7349, n7118, g1536 );
nor U11055 ( n7350, n7114, g1537 );
or U11056 ( n3662, n7351, n7352 );
nor U11057 ( n7351, n7119, g842 );
nor U11058 ( n7352, n7115, g843 );
or U11059 ( n3761, n7353, n7354 );
nor U11060 ( n7353, n7120, g154 );
nor U11061 ( n7354, n7116, g155 );
xor U11062 ( n4211, g2185, n4212 );
nor U11063 ( n4212, n4213, n4214 );
nor U11064 ( n4213, g2223, n7435 );
nand U11065 ( n4214, n4215, n4216 );
xor U11066 ( n3577, g1491, n3578 );
nor U11067 ( n3578, n3579, n3580 );
nor U11068 ( n3579, g1529, n7447 );
nand U11069 ( n3580, n3581, n3582 );
or U11070 ( n4216, n7113, g2225 );
or U11071 ( n3582, n7114, g1531 );
xor U11072 ( n3680, g801, n3681 );
nor U11073 ( n3681, n3682, n3684 );
nor U11074 ( n3682, g835, n7459 );
nand U11075 ( n3684, n3685, n3686 );
xor U11076 ( n3779, g113, n3780 );
nor U11077 ( n3780, n3781, n3783 );
nor U11078 ( n3781, g147, n7471 );
nand U11079 ( n3783, n3784, n3785 );
or U11080 ( n3686, n7115, g837 );
or U11081 ( n3785, n7116, g149 );
or U11082 ( n4215, n7117, g2224 );
or U11083 ( n3581, n7118, g1530 );
or U11084 ( n3685, n7119, g836 );
or U11085 ( n3784, n7120, g148 );
nand U11086 ( n4346, g3233, n638 );
not U11087 ( n638, g3230 );
nor U11088 ( n4279, n4291, n4292 );
nand U11089 ( n4291, n4294, n4295 );
nand U11090 ( n4292, n637, n4293 );
nand U11091 ( n4294, g3113, n4297 );
nand U11092 ( n6175, n6176, n6177 );
nor U11093 ( n6177, n6178, n6179 );
nor U11094 ( n6176, n6180, n4346 );
and U11095 ( n6179, g3114, n4297 );
nand U11096 ( n4340, n4341, n4342 );
nor U11097 ( n4342, n4343, n4344 );
nor U11098 ( n4341, n4345, n4346 );
and U11099 ( n4344, g3120, n4297 );
nor U11100 ( n1173, n1174, n1175 );
nand U11101 ( n1175, g2384, n532 );
nor U11102 ( n1191, n1192, n1193 );
nand U11103 ( n1193, g1690, n421 );
nor U11104 ( n1133, n1134, n1135 );
nand U11105 ( n1135, g996, n312 );
nor U11106 ( n1153, n1154, n1155 );
nand U11107 ( n1155, g309, n191 );
nand U11108 ( new_g30341_, n1162, n1163 );
nand U11109 ( n1162, g2394, n7430 );
nand U11110 ( n1163, n1108, g7264 );
nand U11111 ( new_g30503_, n1109, n1110 );
nand U11112 ( n1109, g1700, n7442 );
nand U11113 ( n1110, n1111, g7014 );
nand U11114 ( new_g30485_, n1117, n1118 );
nand U11115 ( n1117, g1006, n7454 );
nand U11116 ( n1118, n1114, g6712 );
nand U11117 ( new_g30505_, n1106, n1107 );
nand U11118 ( n1106, g2393, n7433 );
nand U11119 ( n1107, n1108, g5555 );
nand U11120 ( new_g30487_, n1115, n1116 );
nand U11121 ( n1115, g1699, n7445 );
nand U11122 ( n1116, n1111, g5511 );
nand U11123 ( new_g30470_, n1122, n1123 );
nand U11124 ( n1122, g1005, n7457 );
nand U11125 ( n1123, n1114, g5472 );
nand U11126 ( new_g30455_, n1142, n1143 );
nand U11127 ( n1142, g318, n7469 );
nand U11128 ( n1143, n1121, g5437 );
nand U11129 ( new_g30468_, n1140, n1141 );
nand U11130 ( n1140, g319, n7466 );
nand U11131 ( n1141, n1121, g6447 );
nand U11132 ( new_g30356_, n1160, n1161 );
nand U11133 ( n1160, g2395, n7425 );
nand U11134 ( n1161, n1108, g2476 );
nand U11135 ( new_g30338_, n1180, n1181 );
nand U11136 ( n1180, g1701, n7437 );
nand U11137 ( n1181, n1111, g1782 );
nand U11138 ( new_g30500_, n1112, n1113 );
nand U11139 ( n1112, g1007, n7449 );
nand U11140 ( n1113, n1114, g1088 );
nand U11141 ( new_g30482_, n1119, n1120 );
nand U11142 ( n1119, g320, n7461 );
nand U11143 ( n1120, n1121, g401 );
nor U11144 ( new_g27315_, n2945, n2946 );
nor U11145 ( n2945, g1269, n342 );
nor U11146 ( n2946, n2904, n2901 );
nor U11147 ( new_g27332_, n2890, n2891 );
nor U11148 ( n2890, g1963, n451 );
nor U11149 ( n2891, n2866, n2863 );
nor U11150 ( new_g27321_, n2926, n2927 );
nor U11151 ( n2926, g1962, n449 );
nor U11152 ( n2927, n2866, n2889 );
nor U11153 ( new_g27338_, n2871, n2872 );
nor U11154 ( n2871, g2656, n564 );
nor U11155 ( n2872, n2844, n2851 );
nor U11156 ( new_g27281_, n3101, n3102 );
nor U11157 ( n3101, g582, n219 );
nor U11158 ( n3102, n2959, n3031 );
nor U11159 ( new_g27295_, n3032, n3033 );
nor U11160 ( n3032, g583, n221 );
nor U11161 ( n3033, n2959, n2956 );
nor U11162 ( new_g27311_, n2957, n2958 );
nor U11163 ( n2957, g581, n220 );
nor U11164 ( n2958, n2959, n2907 );
nor U11165 ( new_g27301_, n3013, n3014 );
nor U11166 ( n3013, g1268, n340 );
nor U11167 ( n3014, n2904, n2944 );
nor U11168 ( new_g27328_, n2902, n2903 );
nor U11169 ( n2902, g1267, n341 );
nor U11170 ( n2903, n2904, n2869 );
nor U11171 ( new_g27340_, n2864, n2865 );
nor U11172 ( n2864, g1961, n450 );
nor U11173 ( n2865, n2866, n2847 );
nor U11174 ( new_g27344_, n2852, n2853 );
nor U11175 ( n2852, g2657, n566 );
nor U11176 ( n2853, n2844, n2841 );
nor U11177 ( new_g27347_, n2842, n2843 );
nor U11178 ( n2842, g2655, n565 );
nor U11179 ( n2843, n2844, n2837 );
nor U11180 ( n7043, n6193, n4346 );
nor U11181 ( n6193, g3123, n4709 );
nor U11182 ( new_g27327_, n2905, n2906 );
nor U11183 ( n2905, g584, n220 );
nor U11184 ( n2906, n2907, n2908 );
nor U11185 ( new_g27339_, n2867, n2868 );
nor U11186 ( n2867, g1270, n341 );
nor U11187 ( n2868, n2869, n2870 );
nor U11188 ( new_g27346_, n2845, n2846 );
nor U11189 ( n2845, g1964, n450 );
nor U11190 ( n2846, n2847, n2848 );
nor U11191 ( new_g27354_, n2835, n2836 );
nor U11192 ( n2835, g2658, n565 );
nor U11193 ( n2836, n2837, n2838 );
nor U11194 ( new_g27329_, n2899, n2900 );
nor U11195 ( n2899, g1272, n342 );
nor U11196 ( n2900, n2870, n2901 );
nor U11197 ( new_g27341_, n2861, n2862 );
nor U11198 ( n2861, g1966, n451 );
nor U11199 ( n2862, n2848, n2863 );
nor U11200 ( new_g27333_, n2887, n2888 );
nor U11201 ( n2887, g1965, n449 );
nor U11202 ( n2888, n2848, n2889 );
nor U11203 ( new_g27345_, n2849, n2850 );
nor U11204 ( n2849, g2659, n564 );
nor U11205 ( n2850, n2838, n2851 );
nor U11206 ( new_g27296_, n3029, n3030 );
nor U11207 ( n3029, g585, n219 );
nor U11208 ( n3030, n2908, n3031 );
nor U11209 ( new_g27312_, n2954, n2955 );
nor U11210 ( n2954, g586, n221 );
nor U11211 ( n2955, n2908, n2956 );
nor U11212 ( new_g27316_, n2942, n2943 );
nor U11213 ( n2942, g1271, n340 );
nor U11214 ( n2943, n2870, n2944 );
nor U11215 ( new_g27348_, n2839, n2840 );
nor U11216 ( n2839, g2660, n566 );
nor U11217 ( n2840, n2838, n2841 );
nor U11218 ( new_g27269_, n3187, n3188 );
nor U11219 ( n3187, g579, n219 );
nor U11220 ( n3188, n3036, n3031 );
nor U11221 ( new_g27280_, n3106, n3107 );
nor U11222 ( n3106, g580, n221 );
nor U11223 ( n3107, n3036, n2956 );
nor U11224 ( new_g27300_, n3018, n3019 );
nor U11225 ( n3018, g1266, n342 );
nor U11226 ( n3019, n2949, n2901 );
nor U11227 ( new_g27320_, n2931, n2932 );
nor U11228 ( n2931, g1960, n451 );
nor U11229 ( n2932, n2894, n2863 );
nor U11230 ( new_g27306_, n2996, n2997 );
nor U11231 ( n2996, g1959, n449 );
nor U11232 ( n2997, n2894, n2889 );
nor U11233 ( new_g27326_, n2909, n2910 );
nor U11234 ( n2909, g2653, n564 );
nor U11235 ( n2910, n2856, n2851 );
nor U11236 ( new_g27294_, n3034, n3035 );
nor U11237 ( n3034, g578, n220 );
nor U11238 ( n3035, n3036, n2907 );
nor U11239 ( new_g27286_, n3084, n3085 );
nor U11240 ( n3084, g1265, n340 );
nor U11241 ( n3085, n2949, n2944 );
nor U11242 ( new_g27314_, n2947, n2948 );
nor U11243 ( n2947, g1264, n341 );
nor U11244 ( n2948, n2949, n2869 );
nor U11245 ( new_g27331_, n2892, n2893 );
nor U11246 ( n2892, g1958, n450 );
nor U11247 ( n2893, n2894, n2847 );
nor U11248 ( new_g27337_, n2876, n2877 );
nor U11249 ( n2876, g2654, n566 );
nor U11250 ( n2877, n2856, n2841 );
nor U11251 ( new_g27343_, n2854, n2855 );
nor U11252 ( n2854, g2652, n565 );
nor U11253 ( n2855, n2856, n2837 );
nand U11254 ( g25435, n6194, n637 );
nor U11255 ( n6194, n6195, n6196 );
and U11256 ( n6195, g3110, n4297 );
nor U11257 ( n6196, g3125, n4709 );
nor U11258 ( new_g27285_, n3088, n3089 );
nor U11259 ( n3088, g1263, n342 );
nor U11260 ( n3089, n3022, n2901 );
nor U11261 ( new_g27305_, n3000, n3001 );
nor U11262 ( n3000, g1957, n451 );
nor U11263 ( n3001, n2935, n2863 );
nor U11264 ( new_g27290_, n3048, n3049 );
nor U11265 ( n3048, g1956, n449 );
nor U11266 ( n3049, n2935, n2889 );
nor U11267 ( new_g27310_, n2960, n2961 );
nor U11268 ( n2960, g2650, n564 );
nor U11269 ( n2961, n2880, n2851 );
nor U11270 ( new_g27307_, n2992, n2993 );
nor U11271 ( n2992, g2421, n42 );
nor U11272 ( n2993, n2994, n2859 );
nor U11273 ( new_g27287_, n3080, n3081 );
nor U11274 ( n3080, g1727, n39 );
nor U11275 ( n3081, n3082, n2897 );
nor U11276 ( new_g27270_, n3181, n3183 );
nor U11277 ( n3181, g1033, n36 );
nor U11278 ( n3183, n3184, n2952 );
nor U11279 ( new_g27258_, n3270, n3271 );
nor U11280 ( n3270, g346, n33 );
nor U11281 ( n3271, n3272, n3039 );
nor U11282 ( new_g27268_, n3191, n3192 );
nor U11283 ( n3191, g577, n221 );
nor U11284 ( n3192, n3110, n2956 );
nor U11285 ( new_g27279_, n3108, n3109 );
nor U11286 ( n3108, g575, n220 );
nor U11287 ( n3109, n3110, n2907 );
nor U11288 ( new_g27261_, n3238, n3239 );
nor U11289 ( n3238, g576, n219 );
nor U11290 ( n3239, n3110, n3031 );
nor U11291 ( new_g27299_, n3020, n3021 );
nor U11292 ( n3020, g1261, n341 );
nor U11293 ( n3021, n3022, n2869 );
nor U11294 ( new_g27273_, n3149, n3150 );
nor U11295 ( n3149, g1262, n340 );
nor U11296 ( n3150, n3022, n2944 );
nor U11297 ( new_g27319_, n2933, n2934 );
nor U11298 ( n2933, g1955, n450 );
nor U11299 ( n2934, n2935, n2847 );
nor U11300 ( new_g27325_, n2913, n2914 );
nor U11301 ( n2913, g2651, n566 );
nor U11302 ( n2914, n2880, n2841 );
nor U11303 ( new_g27336_, n2878, n2879 );
nor U11304 ( n2878, g2649, n565 );
nor U11305 ( n2879, n2880, n2837 );
nor U11306 ( new_g27291_, n3046, n3047 );
nor U11307 ( n3046, g2418, n41 );
nor U11308 ( n3047, n2994, n2883 );
nor U11309 ( new_g27276_, n3117, n3118 );
nor U11310 ( n3117, g2429, n40 );
nor U11311 ( n3118, n2994, n2917 );
nor U11312 ( new_g27274_, n3147, n3148 );
nor U11313 ( n3147, g1724, n38 );
nor U11314 ( n3148, n3082, n2938 );
nor U11315 ( new_g27264_, n3206, n3207 );
nor U11316 ( n3206, g1735, n37 );
nor U11317 ( n3207, n3082, n3004 );
nor U11318 ( new_g27262_, n3236, n3237 );
nor U11319 ( n3236, g1030, n35 );
nor U11320 ( n3237, n3184, n3025 );
nor U11321 ( new_g27257_, n3274, n3275 );
nor U11322 ( n3274, g1041, n34 );
nor U11323 ( n3275, n3184, n3092 );
nor U11324 ( new_g27255_, n3304, n3305 );
nor U11325 ( n3304, g343, n32 );
nor U11326 ( n3305, n3272, n3113 );
nor U11327 ( new_g27253_, n3306, n3307 );
nor U11328 ( n3306, g354, n31 );
nor U11329 ( n3307, n3272, n3196 );
or U11330 ( g25420, n4346, n4706 );
nand U11331 ( n4706, n4707, n4708 );
nand U11332 ( n4708, g3112, n4297 );
nand U11333 ( n4707, g3126, n151 );
or U11334 ( g25442, n4346, n4703 );
nand U11335 ( n4703, n4704, n4705 );
nand U11336 ( n4705, g3111, n4297 );
nand U11337 ( n4704, g3124, n151 );
nor U11338 ( n6801, n6806, n6807 );
nand U11339 ( n6807, n6808, n6809 );
nand U11340 ( n6809, n6810, n6811 );
nand U11341 ( n6810, g2615, n7501 );
nor U11342 ( n6415, n6420, n6421 );
nand U11343 ( n6421, n6422, n6423 );
nand U11344 ( n6423, n6424, n6425 );
nand U11345 ( n6424, g1227, n7501 );
nand U11346 ( n6811, g2612, g3229 );
nand U11347 ( n6425, g1224, g3229 );
nand U11348 ( n7075, n6784, n6785 );
nand U11349 ( n6785, g2584, n6786 );
nor U11350 ( n6784, n6801, n6802 );
xor U11351 ( n6786, n6787, n6788 );
nand U11352 ( n7055, n6398, n6399 );
nand U11353 ( n6399, g1196, n6400 );
nor U11354 ( n6398, n6415, n6416 );
xor U11355 ( n6400, n6401, n6402 );
nor U11356 ( n6610, n6615, n6616 );
nand U11357 ( n6616, n6617, n6618 );
nand U11358 ( n6618, n6619, n6620 );
nand U11359 ( n6619, g1921, n7501 );
nand U11360 ( n6620, g1918, g3229 );
nand U11361 ( n7065, n6591, n6592 );
nand U11362 ( n6592, g1890, n6593 );
nor U11363 ( n6591, n6610, n6611 );
xor U11364 ( n6593, n6594, n6595 );
nor U11365 ( n6222, n6227, n6228 );
nand U11366 ( n6228, n6229, n6230 );
nand U11367 ( n6230, n6231, n6232 );
nand U11368 ( n6232, g541, n7501 );
nand U11369 ( n6231, g538, g3229 );
nand U11370 ( n7045, n6205, n6206 );
nand U11371 ( n6206, g510, n6207 );
nor U11372 ( n6205, n6222, n6223 );
xor U11373 ( n6207, n6208, n6209 );
nand U11374 ( new_g29182_, n1763, n1765 );
nand U11375 ( n1763, g2397, n1813 );
nand U11376 ( n1765, n121, n1751 );
not U11377 ( n121, n1813 );
nand U11378 ( new_g29181_, n1824, n1825 );
nand U11379 ( n1824, g1704, n1826 );
nand U11380 ( n1825, n56, n1760 );
not U11381 ( n56, n1826 );
nand U11382 ( new_g29178_, n1832, n1833 );
nand U11383 ( n1832, g1703, n1876 );
nand U11384 ( n1833, n55, n1760 );
not U11385 ( n55, n1876 );
nand U11386 ( new_g29185_, n1754, n1756 );
nand U11387 ( n1754, g2398, n1757 );
nand U11388 ( n1756, n122, n1751 );
not U11389 ( n122, n1757 );
nand U11390 ( new_g29173_, n1888, n1889 );
nand U11391 ( n1888, g1010, n1890 );
nand U11392 ( n1889, n78, n1829 );
not U11393 ( n78, n1890 );
nand U11394 ( new_g29170_, n1897, n1898 );
nand U11395 ( n1897, g1009, n1947 );
nand U11396 ( n1898, n77, n1829 );
not U11397 ( n77, n1947 );
nand U11398 ( new_g29169_, n1959, n1960 );
nand U11399 ( n1959, g323, n1961 );
nand U11400 ( n1960, n100, n1894 );
not U11401 ( n100, n1961 );
nand U11402 ( new_g29167_, n1962, n1963 );
nand U11403 ( n1962, g322, n2013 );
nand U11404 ( n1963, n99, n1894 );
not U11405 ( n99, n2013 );
nand U11406 ( new_g29187_, n1749, n1750 );
nand U11407 ( n1749, g2396, n1752 );
nand U11408 ( n1750, n1751, n123 );
not U11409 ( n123, n1752 );
nand U11410 ( new_g29184_, n1758, n1759 );
nand U11411 ( n1758, g1702, n1761 );
nand U11412 ( n1759, n1760, n57 );
not U11413 ( n57, n1761 );
nand U11414 ( new_g29179_, n1827, n1828 );
nand U11415 ( n1827, g1008, n1830 );
nand U11416 ( n1828, n1829, n79 );
not U11417 ( n79, n1830 );
nand U11418 ( new_g29172_, n1891, n1893 );
nand U11419 ( n1891, g321, n1895 );
nand U11420 ( n1893, n1894, n101 );
not U11421 ( n101, n1895 );
or U11422 ( n1093, n2116, n7355 );
or U11423 ( n681, n2157, n7356 );
or U11424 ( n718, n2196, n7357 );
or U11425 ( n752, n2230, n7358 );
nand U11426 ( n1251, n3906, n3907 );
nand U11427 ( n3907, g2267, n7389 );
nor U11428 ( n3906, n3908, n3909 );
and U11429 ( n3908, n7474, g2264 );
nand U11430 ( n1291, n3979, n3980 );
nand U11431 ( n3980, g1573, n7399 );
nor U11432 ( n3979, n3981, n3982 );
and U11433 ( n3981, n7480, g1570 );
nand U11434 ( n1337, n4049, n4050 );
nand U11435 ( n4050, g879, n7409 );
nor U11436 ( n4049, n4051, n4052 );
and U11437 ( n4051, n7486, g876 );
nand U11438 ( n1373, n4120, n4121 );
nand U11439 ( n4121, g192, n7419 );
nor U11440 ( n4120, n4122, n4123 );
and U11441 ( n4122, n7492, g189 );
and U11442 ( n3909, n7477, g2261 );
and U11443 ( n3982, n7483, g1567 );
and U11444 ( n4052, n7489, g873 );
and U11445 ( n4123, n7495, g186 );
nand U11446 ( n801, n3910, n3911 );
nand U11447 ( n3911, g2348, n7388 );
nor U11448 ( n3910, n3912, n3913 );
and U11449 ( n3912, n7474, g2345 );
nand U11450 ( n837, n3983, n3984 );
nand U11451 ( n3984, g1654, n7398 );
nor U11452 ( n3983, n3985, n3986 );
and U11453 ( n3985, n7480, g1651 );
nand U11454 ( n875, n4053, n4054 );
nand U11455 ( n4054, g960, n7408 );
nor U11456 ( n4053, n4055, n4056 );
and U11457 ( n4055, n7486, g957 );
nand U11458 ( n921, n4124, n4125 );
nand U11459 ( n4125, g273, n7418 );
nor U11460 ( n4124, n4126, n4127 );
and U11461 ( n4126, n7492, g270 );
and U11462 ( n3913, n7477, g2342 );
and U11463 ( n3986, n7483, g1648 );
and U11464 ( n4056, n7489, g954 );
and U11465 ( n4127, n7495, g267 );
nand U11466 ( n934, n3928, n3929 );
nand U11467 ( n3929, g2312, n7393 );
nor U11468 ( n3928, n3930, n3931 );
nand U11469 ( n978, n3999, n4000 );
nand U11470 ( n4000, g1618, n7403 );
nor U11471 ( n3999, n4001, n4002 );
nand U11472 ( n1019, n4069, n4070 );
nand U11473 ( n4070, g924, n7413 );
nor U11474 ( n4069, n4071, n4072 );
nand U11475 ( n1055, n4140, n4141 );
nand U11476 ( n4141, g237, n7423 );
nor U11477 ( n4140, n4142, n4143 );
and U11478 ( n3931, n7477, g2306 );
and U11479 ( n4002, n7483, g1612 );
and U11480 ( n4072, n7489, g918 );
and U11481 ( n4143, n7495, g231 );
nand U11482 ( n1083, n4937, n4938 );
or U11483 ( n4938, n7426, g2395 );
nor U11484 ( n4937, n4939, n4940 );
nor U11485 ( n4939, g2394, n7429 );
nand U11486 ( n671, n4954, n4955 );
or U11487 ( n4955, n7438, g1701 );
nor U11488 ( n4954, n4956, n4957 );
nor U11489 ( n4956, g1700, n7441 );
nand U11490 ( n707, n4971, n4972 );
or U11491 ( n4972, n7450, g1007 );
nor U11492 ( n4971, n4973, n4974 );
nor U11493 ( n4973, g1006, n7453 );
nand U11494 ( n742, n4986, n4987 );
or U11495 ( n4987, n7462, g320 );
nor U11496 ( n4986, n4988, n4989 );
nor U11497 ( n4988, g319, n7466 );
nor U11498 ( n4940, g2393, n7432 );
nor U11499 ( n4957, g1699, n7444 );
nor U11500 ( n4974, g1005, n7456 );
nor U11501 ( n4989, g318, n7468 );
and U11502 ( n3930, n7474, g2309 );
and U11503 ( n4001, n7480, g1615 );
and U11504 ( n4071, n7486, g921 );
and U11505 ( n4142, n7492, g234 );
buf U11506 ( n7431, n542 );
not U11507 ( n542, g5555 );
buf U11508 ( n7443, n430 );
not U11509 ( n430, g5511 );
buf U11510 ( n7455, n321 );
not U11511 ( n321, g5472 );
buf U11512 ( n7467, n200 );
not U11513 ( n200, g5437 );
buf U11514 ( n7452, n324 );
not U11515 ( n324, g6712 );
buf U11516 ( n7428, n546 );
not U11517 ( n546, g7264 );
nand U11518 ( n805, n3949, n3950 );
nand U11519 ( n3950, g2303, n7391 );
nor U11520 ( n3949, n3951, n3952 );
and U11521 ( n3951, g7084, g2300 );
nand U11522 ( n841, n4019, n4020 );
nand U11523 ( n4020, g1609, n7401 );
nor U11524 ( n4019, n4021, n4022 );
and U11525 ( n4021, g6782, g1606 );
nand U11526 ( n879, n4089, n4090 );
nand U11527 ( n4090, g915, n7411 );
nor U11528 ( n4089, n4091, n4092 );
and U11529 ( n4091, g6518, g912 );
nand U11530 ( n925, n4160, n4161 );
nand U11531 ( n4161, g228, n7421 );
nor U11532 ( n4160, n4162, n4163 );
and U11533 ( n4162, g6313, g225 );
and U11534 ( n3952, g6837, g2297 );
and U11535 ( n4022, g6573, g1603 );
and U11536 ( n4092, g6368, g909 );
and U11537 ( n4163, g6231, g222 );
buf U11538 ( n7464, n204 );
not U11539 ( n204, g6447 );
nor U11540 ( new_g28774_, n2077, n2078 );
nor U11541 ( n2078, n7432, n2064 );
nor U11542 ( n2077, g2502, n2080 );
nor U11543 ( n2080, n118, n7432 );
nor U11544 ( new_g28783_, n2066, n2067 );
nor U11545 ( n2067, n7429, n2064 );
nor U11546 ( n2066, g2503, n2068 );
nor U11547 ( n2068, n118, n7429 );
nor U11548 ( new_g28761_, n2122, n2123 );
nor U11549 ( n2123, n7444, n2075 );
nor U11550 ( n2122, g1808, n2125 );
nor U11551 ( n2125, n52, n7444 );
nor U11552 ( new_g28772_, n2086, n2087 );
nor U11553 ( n2087, n7441, n2075 );
nor U11554 ( n2086, g1809, n2088 );
nor U11555 ( n2088, n52, n7441 );
nor U11556 ( new_g28747_, n2163, n2164 );
nor U11557 ( n2164, n7456, n2095 );
nor U11558 ( n2163, g1114, n2166 );
nor U11559 ( n2166, n74, n7456 );
nor U11560 ( new_g28759_, n2130, n2131 );
nor U11561 ( n2131, n7453, n2095 );
nor U11562 ( n2130, g1115, n2132 );
nor U11563 ( n2132, n74, n7453 );
nor U11564 ( new_g28736_, n2203, n2204 );
nor U11565 ( n2204, n7468, n2138 );
nor U11566 ( n2203, g427, n2206 );
nor U11567 ( n2206, n96, n7468 );
nor U11568 ( new_g28745_, n2171, n2172 );
nor U11569 ( n2172, n7465, n2138 );
nor U11570 ( n2171, g428, n2173 );
nor U11571 ( n2173, n96, n7465 );
nor U11572 ( new_g28788_, n2061, n2062 );
nor U11573 ( n2062, n7425, n2064 );
nor U11574 ( n2061, g2501, n2065 );
nor U11575 ( n2065, n118, n7425 );
nor U11576 ( new_g28778_, n2073, n2074 );
nor U11577 ( n2074, n7437, n2075 );
nor U11578 ( n2073, g1807, n2076 );
nor U11579 ( n2076, n52, n7437 );
nor U11580 ( new_g28767_, n2093, n2094 );
nor U11581 ( n2094, n7449, n2095 );
nor U11582 ( n2093, g1113, n2096 );
nor U11583 ( n2096, n74, n7449 );
nor U11584 ( new_g28754_, n2136, n2137 );
nor U11585 ( n2137, n7461, n2138 );
nor U11586 ( n2136, g426, n2139 );
nor U11587 ( n2139, n96, n7461 );
buf U11588 ( n7440, n433 );
not U11589 ( n433, g7014 );
nand U11590 ( n1211, n3923, n3925 );
nand U11591 ( n3925, g2285, n7394 );
nor U11592 ( n3923, n3926, n3927 );
nand U11593 ( n1231, n3995, n3996 );
nand U11594 ( n3996, g1591, n7404 );
nor U11595 ( n3995, n3997, n3998 );
nand U11596 ( n1262, n4065, n4066 );
nand U11597 ( n4066, g897, n7414 );
nor U11598 ( n4065, n4067, n4068 );
nand U11599 ( n1302, n4136, n4137 );
nand U11600 ( n4137, g210, n7424 );
nor U11601 ( n4136, n4138, n4139 );
and U11602 ( n3927, n7477, g2279 );
and U11603 ( n3998, n7483, g1585 );
and U11604 ( n4068, n7489, g891 );
and U11605 ( n4139, n7495, g204 );
and U11606 ( n3926, n7474, g2282 );
and U11607 ( n3997, n7480, g1588 );
and U11608 ( n4067, n7486, g894 );
and U11609 ( n4138, n7492, g207 );
nand U11610 ( n900, n3932, n3933 );
nand U11611 ( n3933, g2321, n7393 );
nor U11612 ( n3932, n3934, n3935 );
and U11613 ( n3934, n7474, g2318 );
nand U11614 ( n947, n4003, n4004 );
nand U11615 ( n4004, g1627, n7403 );
nor U11616 ( n4003, n4005, n4006 );
and U11617 ( n4005, n7480, g1624 );
nand U11618 ( n991, n4073, n4074 );
nand U11619 ( n4074, g933, n7413 );
nor U11620 ( n4073, n4075, n4076 );
and U11621 ( n4075, n7486, g930 );
nand U11622 ( n1032, n4144, n4145 );
nand U11623 ( n4145, g246, n7423 );
nor U11624 ( n4144, n4146, n4147 );
and U11625 ( n4146, n7492, g243 );
and U11626 ( n3935, n7477, g2315 );
and U11627 ( n4006, n7483, g1621 );
and U11628 ( n4076, n7489, g927 );
and U11629 ( n4147, n7495, g240 );
nand U11630 ( n784, n3914, n3916 );
nand U11631 ( n3916, g2276, n7389 );
nor U11632 ( n3914, n3917, n3918 );
and U11633 ( n3917, n7474, g2273 );
nand U11634 ( n817, n3987, n3988 );
nand U11635 ( n3988, g1582, n7399 );
nor U11636 ( n3987, n3989, n3990 );
and U11637 ( n3989, n7480, g1579 );
nand U11638 ( n853, n4057, n4058 );
nand U11639 ( n4058, g888, n7409 );
nor U11640 ( n4057, n4059, n4060 );
and U11641 ( n4059, n7486, g885 );
nand U11642 ( n891, n4128, n4129 );
nand U11643 ( n4129, g201, n7419 );
nor U11644 ( n4128, n4130, n4131 );
and U11645 ( n4130, n7492, g198 );
and U11646 ( n3918, n7477, g2270 );
and U11647 ( n3990, n7483, g1576 );
and U11648 ( n4060, n7489, g882 );
and U11649 ( n4131, n7495, g195 );
nor U11650 ( n4931, g2388, n7430 );
nor U11651 ( n4948, g1694, n7442 );
nor U11652 ( n4965, g1000, n7454 );
nand U11653 ( n1277, n3957, n3958 );
nand U11654 ( n3958, g2294, n7389 );
nor U11655 ( n3957, n3959, n3960 );
and U11656 ( n3959, g7084, g2291 );
nand U11657 ( n1323, n4027, n4028 );
nand U11658 ( n4028, g1600, n7399 );
nor U11659 ( n4027, n4029, n4030 );
and U11660 ( n4029, g6782, g1597 );
nand U11661 ( n1359, n4097, n4098 );
nand U11662 ( n4098, g906, n7409 );
nor U11663 ( n4097, n4099, n4100 );
and U11664 ( n4099, g6518, g903 );
nand U11665 ( n1393, n4168, n4169 );
nand U11666 ( n4169, g219, n7419 );
nor U11667 ( n4168, n4170, n4171 );
and U11668 ( n4170, g6313, g216 );
nand U11669 ( n1082, n4929, n4930 );
or U11670 ( n4930, n7425, g2389 );
nor U11671 ( n4929, n4931, n4932 );
nor U11672 ( n4932, g2387, n7433 );
nand U11673 ( n670, n4946, n4947 );
or U11674 ( n4947, n7437, g1695 );
nor U11675 ( n4946, n4948, n4949 );
nor U11676 ( n4949, g1693, n7445 );
nand U11677 ( n706, n4963, n4964 );
or U11678 ( n4964, n7449, g1001 );
nor U11679 ( n4963, n4965, n4966 );
nor U11680 ( n4966, g999, n7457 );
nand U11681 ( n741, n4978, n4979 );
or U11682 ( n4979, n7461, g314 );
nor U11683 ( n4978, n4980, n4981 );
nor U11684 ( n4980, g313, n7465 );
and U11685 ( n3960, g6837, g2288 );
and U11686 ( n4030, g6573, g1594 );
and U11687 ( n4100, g6368, g900 );
and U11688 ( n4171, g6231, g213 );
nor U11689 ( n4981, g312, n7469 );
nand U11690 ( n1312, n3953, n3954 );
nand U11691 ( n3954, g2330, n7390 );
nor U11692 ( n3953, n3955, n3956 );
and U11693 ( n3955, g7084, g2327 );
nand U11694 ( n1348, n4023, n4024 );
nand U11695 ( n4024, g1636, n7400 );
nor U11696 ( n4023, n4025, n4026 );
and U11697 ( n4025, g6782, g1633 );
nand U11698 ( n1382, n4093, n4094 );
nand U11699 ( n4094, g942, n7410 );
nor U11700 ( n4093, n4095, n4096 );
and U11701 ( n4095, g6518, g939 );
nand U11702 ( n1407, n4164, n4165 );
nand U11703 ( n4165, g255, n7420 );
nor U11704 ( n4164, n4166, n4167 );
and U11705 ( n4166, g6313, g252 );
and U11706 ( n3956, g6837, g2324 );
and U11707 ( n4026, g6573, g1630 );
and U11708 ( n4096, g6368, g936 );
and U11709 ( n4167, g6231, g249 );
nand U11710 ( n1274, n3941, n3942 );
nand U11711 ( n3942, g2339, n7392 );
nor U11712 ( n3941, n3943, n3944 );
and U11713 ( n3943, g7084, g2336 );
nand U11714 ( n1320, n4011, n4012 );
nand U11715 ( n4012, g1645, n7402 );
nor U11716 ( n4011, n4013, n4014 );
and U11717 ( n4013, g6782, g1642 );
nand U11718 ( n1356, n4081, n4082 );
nand U11719 ( n4082, g951, n7412 );
nor U11720 ( n4081, n4083, n4084 );
and U11721 ( n4083, g6518, g948 );
nand U11722 ( n1390, n4152, n4153 );
nand U11723 ( n4153, g264, n7422 );
nor U11724 ( n4152, n4154, n4155 );
and U11725 ( n4154, g6313, g261 );
and U11726 ( n3944, g6837, g2333 );
and U11727 ( n4014, g6573, g1639 );
and U11728 ( n4084, g6368, g945 );
and U11729 ( n4155, g6231, g258 );
nand U11730 ( new_g29621_, n1602, n1603 );
nand U11731 ( n1602, g2388, n7430 );
nand U11732 ( n1603, n1601, g7264 );
nand U11733 ( new_g29612_, n1624, n1625 );
nand U11734 ( n1624, g1000, n7454 );
nand U11735 ( n1625, n1617, g6712 );
nand U11736 ( new_g29618_, n1607, n1608 );
nand U11737 ( n1607, g2387, n7433 );
nand U11738 ( n1608, n1601, g5555 );
nand U11739 ( new_g29613_, n1618, n1619 );
nand U11740 ( n1618, g1693, n7445 );
nand U11741 ( n1619, n1606, g5511 );
nand U11742 ( new_g29617_, n1613, n1614 );
nand U11743 ( n1613, g1694, n7442 );
nand U11744 ( n1614, n1606, g7014 );
nand U11745 ( new_g29609_, n1629, n1630 );
nand U11746 ( n1629, g999, n7457 );
nand U11747 ( n1630, n1617, g5472 );
nand U11748 ( new_g29606_, n1637, n1638 );
nand U11749 ( n1637, g312, n7469 );
nand U11750 ( n1638, n1628, g5437 );
nand U11751 ( new_g29608_, n1635, n1636 );
nand U11752 ( n1635, g313, n7466 );
nand U11753 ( n1636, n1628, g6447 );
nand U11754 ( new_g29623_, n1599, n1600 );
nand U11755 ( n1599, g2389, n7425 );
nand U11756 ( n1600, n1601, g2476 );
nand U11757 ( new_g29620_, n1604, n1605 );
nand U11758 ( n1604, g1695, n7437 );
nand U11759 ( n1605, n1606, g1782 );
nand U11760 ( new_g29616_, n1615, n1616 );
nand U11761 ( n1615, g1001, n7449 );
nand U11762 ( n1616, n1617, g1088 );
nand U11763 ( new_g29611_, n1626, n1627 );
nand U11764 ( n1626, g314, n7461 );
nand U11765 ( n1627, n1628, g401 );
nand U11766 ( new_g28773_, n2084, n2085 );
nand U11767 ( n2084, g2486, n7430 );
nand U11768 ( n2085, g7264, n2071 );
nand U11769 ( new_g28746_, n2169, n2170 );
nand U11770 ( n2169, g1098, n7454 );
nand U11771 ( n2170, g6712, n2135 );
nand U11772 ( new_g28763_, n2097, n2098 );
nand U11773 ( n2097, g2483, n7433 );
nand U11774 ( n2098, g5555, n2071 );
nand U11775 ( new_g28749_, n2140, n2141 );
nand U11776 ( n2140, g1789, n7445 );
nand U11777 ( n2141, g5511, n2092 );
nand U11778 ( new_g28760_, n2128, n2129 );
nand U11779 ( n2128, g1792, n7442 );
nand U11780 ( n2129, g7014, n2092 );
nand U11781 ( new_g28738_, n2177, n2178 );
nand U11782 ( n2177, g1095, n7457 );
nand U11783 ( n2178, g5472, n2135 );
nand U11784 ( new_g28732_, n2211, n2212 );
nand U11785 ( n2211, g408, n7469 );
nand U11786 ( n2212, g5437, n2176 );
nand U11787 ( new_g28735_, n2209, n2210 );
nand U11788 ( n2209, g411, n7466 );
nand U11789 ( n2210, g6447, n2176 );
nand U11790 ( new_g28782_, n2069, n2070 );
nand U11791 ( n2069, g2489, n7425 );
nand U11792 ( n2070, g2476, n2071 );
nand U11793 ( new_g28771_, n2089, n2091 );
nand U11794 ( n2089, g1795, n7437 );
nand U11795 ( n2091, g1782, n2092 );
nand U11796 ( new_g28758_, n2133, n2134 );
nand U11797 ( n2133, g1101, n7449 );
nand U11798 ( n2134, g1088, n2135 );
nand U11799 ( new_g28744_, n2174, n2175 );
nand U11800 ( n2174, g414, n7461 );
nand U11801 ( n2175, g401, n2176 );
nand U11802 ( n1084, n4933, n4934 );
or U11803 ( n4934, n7425, g2392 );
nor U11804 ( n4933, n4935, n4936 );
nor U11805 ( n4936, g2390, n7433 );
nor U11806 ( n4935, g2391, n7430 );
nor U11807 ( n4969, g1003, n7454 );
nand U11808 ( n708, n4967, n4968 );
or U11809 ( n4968, n7449, g1004 );
nor U11810 ( n4967, n4969, n4970 );
nor U11811 ( n4970, g1002, n7457 );
nand U11812 ( n672, n4950, n4951 );
or U11813 ( n4951, n7437, g1698 );
nor U11814 ( n4950, n4952, n4953 );
nor U11815 ( n4953, g1696, n7445 );
nor U11816 ( n4952, g1697, n7442 );
nand U11817 ( n743, n4982, n4983 );
or U11818 ( n4983, n7461, g317 );
nor U11819 ( n4982, n4984, n4985 );
nor U11820 ( n4985, g315, n7469 );
nor U11821 ( n4984, g316, n7466 );
nand U11822 ( new_g29221_, n1662, n1663 );
nand U11823 ( n1662, g2495, n7430 );
nand U11824 ( n1663, g7264, n1661 );
nand U11825 ( new_g29204_, n1706, n1707 );
nand U11826 ( n1706, g1107, n7454 );
nand U11827 ( n1707, g6712, n1688 );
nand U11828 ( new_g29213_, n1667, n1668 );
nand U11829 ( n1667, g2492, n7433 );
nand U11830 ( n1668, g5555, n1661 );
nand U11831 ( new_g29205_, n1689, n1690 );
nand U11832 ( n1689, g1798, n7445 );
nand U11833 ( n1690, g5511, n1666 );
nand U11834 ( new_g29212_, n1684, n1685 );
nand U11835 ( n1684, g1801, n7442 );
nand U11836 ( n1685, g7014, n1666 );
nand U11837 ( new_g29198_, n1711, n1712 );
nand U11838 ( n1711, g1104, n7457 );
nand U11839 ( n1712, g5472, n1688 );
nand U11840 ( new_g29194_, n1730, n1731 );
nand U11841 ( n1730, g417, n7469 );
nand U11842 ( n1731, g5437, n1710 );
nand U11843 ( new_g29197_, n1728, n1729 );
nand U11844 ( n1728, g420, n7466 );
nand U11845 ( n1729, g6447, n1710 );
nand U11846 ( new_g29226_, n1659, n1660 );
nand U11847 ( n1659, g2498, n7425 );
nand U11848 ( n1660, g2476, n1661 );
nand U11849 ( new_g29218_, n1664, n1665 );
nand U11850 ( n1664, g1804, n7437 );
nand U11851 ( n1665, g1782, n1666 );
nand U11852 ( new_g29209_, n1686, n1687 );
nand U11853 ( n1686, g1110, n7449 );
nand U11854 ( n1687, g1088, n1688 );
nand U11855 ( new_g29201_, n1708, n1709 );
nand U11856 ( n1708, g423, n7461 );
nand U11857 ( n1709, g401, n1710 );
buf U11858 ( n7427, n547 );
not U11859 ( n547, g2476 );
buf U11860 ( n7439, n434 );
not U11861 ( n434, g1782 );
buf U11862 ( n7451, n325 );
not U11863 ( n325, g1088 );
buf U11864 ( n7463, n205 );
not U11865 ( n205, g401 );
buf U11866 ( n7434, n519 );
not U11867 ( n519, g2241 );
buf U11868 ( n7446, n409 );
not U11869 ( n409, g1547 );
buf U11870 ( n7458, n300 );
not U11871 ( n300, g853 );
buf U11872 ( n7470, n179 );
not U11873 ( n179, g165 );
nand U11874 ( new_g24059_, n4920, n4921 );
nand U11875 ( n4920, g305, n7501 );
nand U11876 ( n4921, g3229, n7288 );
nand U11877 ( new_g24083_, n4916, n4917 );
nand U11878 ( n4916, g1686, n7501 );
nand U11879 ( n4917, g3229, n7289 );
nand U11880 ( new_g24092_, n4914, n4915 );
nand U11881 ( n4914, g2380, n7501 );
nand U11882 ( n4915, g3229, n7291 );
nand U11883 ( new_g24072_, n4918, n4919 );
nand U11884 ( n4919, g992, n7501 );
nand U11885 ( n4918, g3229, n7292 );
nand U11886 ( n1752, n1753, g2476 );
nand U11887 ( n1761, n1762, g1782 );
nand U11888 ( n1830, n1831, g1088 );
nand U11889 ( n1895, n1896, g401 );
nor U11890 ( new_g26672_, n3532, n3533 );
nor U11891 ( n3532, g2478, n3534 );
nor U11892 ( n3533, n7432, n3526 );
nor U11893 ( n3534, n7432, n7215 );
nor U11894 ( new_g26676_, n3524, n3525 );
nor U11895 ( n3524, g2479, n3527 );
nor U11896 ( n3525, n7429, n3526 );
nor U11897 ( n3527, n7429, n7215 );
nor U11898 ( new_g26667_, n3546, n3547 );
nor U11899 ( n3546, g1784, n3632 );
nor U11900 ( n3547, n7444, n3530 );
nor U11901 ( n3632, n7444, n7216 );
nor U11902 ( new_g26670_, n3539, n3540 );
nor U11903 ( n3539, g1785, n3541 );
nor U11904 ( n3540, n7441, n3530 );
nor U11905 ( n3541, n7441, n7216 );
nor U11906 ( new_g26661_, n3645, n3646 );
nor U11907 ( n3645, g1090, n3735 );
nor U11908 ( n3646, n7456, n3544 );
nor U11909 ( n3735, n7456, n7214 );
nor U11910 ( new_g26665_, n3637, n3639 );
nor U11911 ( n3637, g1091, n3640 );
nor U11912 ( n3639, n7453, n3544 );
nor U11913 ( n3640, n7453, n7214 );
nor U11914 ( new_g26655_, n3744, n3745 );
nor U11915 ( n3744, g403, n3832 );
nor U11916 ( n3745, n7468, n3643 );
nor U11917 ( n3832, n7468, n7217 );
nor U11918 ( new_g26659_, n3741, n3742 );
nor U11919 ( n3741, g404, n3743 );
nor U11920 ( n3742, n7465, n3643 );
nor U11921 ( n3743, n7465, n7217 );
nor U11922 ( new_g26025_, n4179, n4180 );
nor U11923 ( n4179, g2477, n4260 );
nor U11924 ( n4180, n7425, n3526 );
nor U11925 ( n4260, n7425, n7215 );
nor U11926 ( new_g26675_, n3528, n3529 );
nor U11927 ( n3528, g1783, n3531 );
nor U11928 ( n3529, n7437, n3530 );
nor U11929 ( n3531, n7437, n7216 );
nor U11930 ( new_g26669_, n3542, n3543 );
nor U11931 ( n3542, g1089, n3545 );
nor U11932 ( n3543, n7449, n3544 );
nor U11933 ( n3545, n7449, n7214 );
nor U11934 ( new_g26664_, n3641, n3642 );
nor U11935 ( n3641, g402, n3644 );
nor U11936 ( n3642, n7461, n3643 );
nor U11937 ( n3644, n7461, n7217 );
nand U11938 ( n1890, n1831, g6712 );
nand U11939 ( n1757, n1753, g7264 );
nand U11940 ( n1813, n1753, g5555 );
nand U11941 ( n1826, n1762, g7014 );
nand U11942 ( n1876, n1762, g5511 );
nand U11943 ( n1947, n1831, g5472 );
nand U11944 ( n1961, n1896, g6447 );
nand U11945 ( n2013, n1896, g5437 );
nor U11946 ( n4225, g2205, n7435 );
nor U11947 ( n3592, g1511, n7447 );
nor U11948 ( n3697, g817, n7459 );
nor U11949 ( n3795, g129, n7471 );
nor U11950 ( n4194, g2229, n7435 );
nor U11951 ( n3560, g1535, n7447 );
nor U11952 ( n3661, g841, n7459 );
nor U11953 ( n3760, g153, n7471 );
nand U11954 ( n2750, n120, n3390 );
nand U11955 ( n3390, n3391, n3392 );
or U11956 ( n3392, n7117, g2254 );
nor U11957 ( n3391, n3393, n3394 );
nand U11958 ( n2773, n54, n3427 );
nand U11959 ( n3427, n3428, n3429 );
or U11960 ( n3429, n7118, g1560 );
nor U11961 ( n3428, n3430, n3431 );
nand U11962 ( n2794, n76, n3464 );
nand U11963 ( n3464, n3466, n3467 );
or U11964 ( n3467, n7119, g866 );
nor U11965 ( n3466, n3468, n3469 );
nand U11966 ( n2810, n98, n3497 );
nand U11967 ( n3497, n3498, n3499 );
or U11968 ( n3499, n7120, g178 );
nor U11969 ( n3498, n3500, n3502 );
nor U11970 ( n3393, g2255, n7113 );
nor U11971 ( n3430, g1561, n7114 );
nor U11972 ( n3468, g867, n7115 );
nor U11973 ( n3500, g179, n7116 );
nand U11974 ( new_g26826_, n3355, n3356 );
nand U11975 ( n3355, g2516, n7430 );
nand U11976 ( n3356, n3354, g7264 );
nand U11977 ( new_g26814_, n3415, n3416 );
nand U11978 ( n3415, g1128, n7454 );
nand U11979 ( n3416, n3385, g6712 );
nand U11980 ( new_g26823_, n3363, n3364 );
nand U11981 ( n3363, g2513, n7433 );
nand U11982 ( n3364, n3354, g5555 );
nand U11983 ( new_g26816_, n3400, n3401 );
nand U11984 ( n3400, g1819, n7445 );
nand U11985 ( n3401, n3362, g5511 );
nand U11986 ( new_g26821_, n3378, n3379 );
nand U11987 ( n3378, g1822, n7442 );
nand U11988 ( n3379, n3362, g7014 );
nand U11989 ( new_g26810_, n3437, n3439 );
nand U11990 ( n3437, g1125, n7457 );
nand U11991 ( n3439, n3385, g5472 );
nand U11992 ( new_g26805_, n3476, n3477 );
nand U11993 ( n3476, g438, n7469 );
nand U11994 ( n3477, n3422, g5437 );
nand U11995 ( new_g26808_, n3454, n3455 );
nand U11996 ( n3454, g441, n7466 );
nand U11997 ( n3455, n3422, g6447 );
nand U11998 ( new_g26827_, n3352, n3353 );
nand U11999 ( n3352, g2519, n7425 );
nand U12000 ( n3353, n3354, g2476 );
nand U12001 ( new_g26824_, n3360, n3361 );
nand U12002 ( n3360, g1825, n7437 );
nand U12003 ( n3361, n3362, g1782 );
nand U12004 ( new_g26818_, n3383, n3384 );
nand U12005 ( n3383, g1131, n7449 );
nand U12006 ( n3384, n3385, g1088 );
nand U12007 ( new_g26812_, n3420, n3421 );
nand U12008 ( n3420, g444, n7461 );
nand U12009 ( n3421, n3422, g401 );
or U12010 ( n2729, n7359, n2743 );
nand U12011 ( n7359, n2744, g2384 );
or U12012 ( n2737, n7360, n2766 );
nand U12013 ( n7360, n2767, g1690 );
or U12014 ( n2758, n7361, n2787 );
nand U12015 ( n7361, n2788, g996 );
or U12016 ( n2781, n7362, n2803 );
nand U12017 ( n7362, n2804, g309 );
nor U12018 ( new_g27767_, n2740, n2741 );
nor U12019 ( n2740, g2523, n2745 );
nor U12020 ( n2741, n7432, n2729 );
nor U12021 ( n2745, n7432, n2731 );
nor U12022 ( new_g27769_, n2732, n2733 );
nor U12023 ( n2732, g2524, n2734 );
nor U12024 ( n2733, n7429, n2729 );
nor U12025 ( n2734, n7429, n2731 );
nor U12026 ( new_g27764_, n2762, n2764 );
nor U12027 ( n2762, g1829, n2768 );
nor U12028 ( n2764, n7444, n2737 );
nor U12029 ( n2768, n7444, n2739 );
nor U12030 ( new_g27766_, n2753, n2754 );
nor U12031 ( n2753, g1830, n2755 );
nor U12032 ( n2754, n7441, n2737 );
nor U12033 ( n2755, n7441, n2739 );
nor U12034 ( new_g27761_, n2784, n2785 );
nor U12035 ( n2784, g1135, n2789 );
nor U12036 ( n2785, n7456, n2758 );
nor U12037 ( n2789, n7456, n2761 );
nor U12038 ( new_g27763_, n2776, n2777 );
nor U12039 ( n2776, g1136, n2778 );
nor U12040 ( n2777, n7453, n2758 );
nor U12041 ( n2778, n7453, n2761 );
nor U12042 ( new_g27759_, n2800, n2801 );
nor U12043 ( n2800, g448, n2805 );
nor U12044 ( n2801, n7468, n2781 );
nor U12045 ( n2805, n7468, n2783 );
nor U12046 ( new_g27760_, n2797, n2798 );
nor U12047 ( n2797, g449, n2799 );
nor U12048 ( n2798, n7465, n2781 );
nor U12049 ( n2799, n7465, n2783 );
nor U12050 ( new_g27771_, n2727, n2728 );
nor U12051 ( n2727, g2522, n2730 );
nor U12052 ( n2728, n7425, n2729 );
nor U12053 ( n2730, n7425, n2731 );
nor U12054 ( new_g27768_, n2735, n2736 );
nor U12055 ( n2735, g1828, n2738 );
nor U12056 ( n2736, n7437, n2737 );
nor U12057 ( n2738, n7437, n2739 );
nor U12058 ( new_g27765_, n2756, n2757 );
nor U12059 ( n2756, g1134, n2760 );
nor U12060 ( n2757, n7449, n2758 );
nor U12061 ( n2760, n7449, n2761 );
nor U12062 ( new_g27762_, n2779, n2780 );
nor U12063 ( n2779, g447, n2782 );
nor U12064 ( n2780, n7461, n2781 );
nor U12065 ( n2782, n7461, n2783 );
nand U12066 ( n2731, g2384, n2746 );
nand U12067 ( n2746, n2747, n2748 );
nand U12068 ( n2747, n2752, n2750 );
nand U12069 ( n2748, n2749, n543 );
nand U12070 ( n2739, g1690, n2769 );
nand U12071 ( n2769, n2770, n2771 );
nand U12072 ( n2770, n2775, n2773 );
nand U12073 ( n2771, n2772, n431 );
nand U12074 ( n2761, g996, n2790 );
nand U12075 ( n2790, n2791, n2792 );
nand U12076 ( n2791, n2796, n2794 );
nand U12077 ( n2792, n2793, n322 );
nand U12078 ( n2783, g309, n2806 );
nand U12079 ( n2806, n2807, n2808 );
nand U12080 ( n2807, n2812, n2810 );
nand U12081 ( n2808, n2809, n201 );
or U12082 ( n4235, n7436, g2235 );
or U12083 ( n3604, n7448, g1541 );
or U12084 ( n3708, n7460, g847 );
or U12085 ( n3807, n7472, g159 );
nor U12086 ( new_g27334_, n2884, n2885 );
nor U12087 ( n2884, g2451, n42 );
nor U12088 ( n2885, n2886, n2859 );
nor U12089 ( new_g27317_, n2939, n2940 );
nor U12090 ( n2939, g1757, n39 );
nor U12091 ( n2940, n2941, n2897 );
nor U12092 ( new_g27297_, n3026, n3027 );
nor U12093 ( n3026, g1063, n36 );
nor U12094 ( n3027, n3028, n2952 );
nor U12095 ( new_g27277_, n3114, n3115 );
nor U12096 ( n3114, g376, n33 );
nor U12097 ( n3115, n3116, n3039 );
nor U12098 ( new_g27309_, n2983, n2984 );
nor U12099 ( n2983, g2459, n40 );
nor U12100 ( n2984, n2886, n2917 );
nor U12101 ( new_g27323_, n2921, n2922 );
nor U12102 ( n2921, g2448, n41 );
nor U12103 ( n2922, n2886, n2883 );
nor U12104 ( new_g27289_, n3071, n3072 );
nor U12105 ( n3071, g1765, n37 );
nor U12106 ( n3072, n2941, n3004 );
nor U12107 ( new_g27303_, n3008, n3009 );
nor U12108 ( n3008, g1754, n38 );
nor U12109 ( n3009, n2941, n2938 );
nor U12110 ( new_g27272_, n3172, n3173 );
nor U12111 ( n3172, g1071, n34 );
nor U12112 ( n3173, n3028, n3092 );
nor U12113 ( new_g27283_, n3096, n3097 );
nor U12114 ( n3096, g1060, n35 );
nor U12115 ( n3097, n3028, n3025 );
nor U12116 ( new_g27260_, n3261, n3262 );
nor U12117 ( n3261, g384, n31 );
nor U12118 ( n3262, n3116, n3196 );
nor U12119 ( new_g27266_, n3201, n3202 );
nor U12120 ( n3201, g373, n32 );
nor U12121 ( n3202, n3116, n3113 );
nand U12122 ( n6125, n6191, n6192 );
nor U12123 ( n6192, g3198, g3194 );
nor U12124 ( n6191, g3191, n7108 );
nor U12125 ( n6173, n6125, g3204 );
nand U12126 ( n4321, n4329, n4330 );
nor U12127 ( n4330, n4331, n4332 );
nor U12128 ( n4329, n4336, n4337 );
and U12129 ( n4331, n4308, g3136 );
and U12130 ( n4336, n146, g3210 );
nand U12131 ( n4339, n4347, n4348 );
nor U12132 ( n4347, n4353, n4354 );
nor U12133 ( n4348, n4349, n4350 );
and U12134 ( n4354, n4286, g3086 );
nand U12135 ( n4350, n4351, n4352 );
nand U12136 ( n4351, g3096, n4289 );
nand U12137 ( n4352, g3094, n4314 );
and U12138 ( n6154, n6173, g3201 );
nand U12139 ( n6174, n6181, n6182 );
nor U12140 ( n6181, n6187, n6188 );
nor U12141 ( n6182, n6183, n6184 );
and U12142 ( n6188, g3101, n4286 );
nand U12143 ( n6184, n6185, n6186 );
nand U12144 ( n6185, n4289, g3108 );
nand U12145 ( n6186, n4314, g3106 );
nor U12146 ( new_g27342_, n2857, n2858 );
nor U12147 ( n2857, g2466, n42 );
nor U12148 ( n2858, n2859, n2860 );
nor U12149 ( new_g27330_, n2895, n2896 );
nor U12150 ( n2895, g1772, n39 );
nor U12151 ( n2896, n2897, n2898 );
nor U12152 ( new_g27313_, n2950, n2951 );
nor U12153 ( n2950, g1078, n36 );
nor U12154 ( n2951, n2952, n2953 );
nor U12155 ( new_g27293_, n3037, n3038 );
nor U12156 ( n3037, g391, n33 );
nor U12157 ( n3038, n3039, n3040 );
nand U12158 ( n6144, n6145, n6146 );
nor U12159 ( n6145, n6151, n6152 );
nor U12160 ( n6146, n6147, n6148 );
and U12161 ( n6152, g3104, n4313 );
and U12162 ( n6148, g3100, n4317 );
nor U12163 ( new_g27324_, n2915, n2916 );
nor U12164 ( n2915, g2473, n40 );
nor U12165 ( n2916, n2860, n2917 );
nor U12166 ( new_g27304_, n3002, n3003 );
nor U12167 ( n3002, g1779, n37 );
nor U12168 ( n3003, n2898, n3004 );
nor U12169 ( new_g27318_, n2936, n2937 );
nor U12170 ( n2936, g1769, n38 );
nor U12171 ( n2937, n2898, n2938 );
nor U12172 ( new_g27284_, n3090, n3091 );
nor U12173 ( n3090, g1085, n34 );
nor U12174 ( n3091, n2953, n3092 );
nor U12175 ( new_g27267_, n3193, n3194 );
nor U12176 ( n3193, g398, n31 );
nor U12177 ( n3194, n3040, n3196 );
nor U12178 ( new_g27278_, n3111, n3112 );
nor U12179 ( n3111, g388, n32 );
nor U12180 ( n3112, n3040, n3113 );
nor U12181 ( new_g27335_, n2881, n2882 );
nor U12182 ( n2881, g2463, n41 );
nor U12183 ( n2882, n2860, n2883 );
nor U12184 ( new_g27298_, n3023, n3024 );
nor U12185 ( n3023, g1075, n35 );
nor U12186 ( n3024, n2953, n3025 );
and U12187 ( n4324, n7363, n7364 );
nand U12188 ( n7363, n4305, g3211 );
nand U12189 ( n7364, n4317, g3085 );
and U12190 ( n6147, n4305, g3098 );
nor U12191 ( n6156, n6170, n6171 );
nor U12192 ( n6170, n4338, n7091 );
and U12193 ( n6171, n4304, g3099 );
nor U12194 ( n4299, n4300, n4301 );
nand U12195 ( n4301, n4302, n4303 );
nand U12196 ( n4300, n4306, n4307 );
nand U12197 ( n4302, g3158, n4305 );
nand U12198 ( n4306, g3155, n146 );
and U12199 ( n6151, g3105, n4318 );
and U12200 ( n4337, n4304, g3084 );
and U12201 ( n4323, n7365, n7366 );
nand U12202 ( n7365, n4318, g3093 );
nand U12203 ( n7366, n4313, g3092 );
nand U12204 ( n4709, n6197, n6167 );
nor U12205 ( n6197, g3204, n6168 );
nor U12206 ( n6172, n7109, g3188 );
and U12207 ( n6167, n6172, g3201 );
and U12208 ( n4345, g3132, n151 );
nand U12209 ( n6168, n6199, n6200 );
nor U12210 ( n6199, g3194, g3191 );
nor U12211 ( n6200, g3198, g3197 );
nor U12212 ( new_g27322_, n2923, n2924 );
nor U12213 ( n2923, g2436, n42 );
nor U12214 ( n2924, n2925, n2859 );
nor U12215 ( new_g27302_, n3010, n3011 );
nor U12216 ( n3010, g1742, n39 );
nor U12217 ( n3011, n3012, n2897 );
nor U12218 ( new_g27282_, n3098, n3099 );
nor U12219 ( n3098, g1048, n36 );
nor U12220 ( n3099, n3100, n2952 );
nor U12221 ( new_g27265_, n3203, n3204 );
nor U12222 ( n3203, g361, n33 );
nor U12223 ( n3204, n3205, n3039 );
nand U12224 ( n6129, n6163, n6164 );
nor U12225 ( n6164, g3204, g3201 );
and U12226 ( n6163, n6155, n149 );
nor U12227 ( n6157, n6158, n6159 );
and U12228 ( n6158, g3134, n4308 );
nand U12229 ( n6159, n6160, n6162 );
nand U12230 ( n6160, g3147, n4335 );
nor U12231 ( new_g27292_, n3041, n3042 );
nor U12232 ( n3041, g2444, n40 );
nor U12233 ( n3042, n2925, n2917 );
nor U12234 ( new_g27308_, n2990, n2991 );
nor U12235 ( n2990, g2433, n41 );
nor U12236 ( n2991, n2925, n2883 );
nor U12237 ( new_g27275_, n3142, n3143 );
nor U12238 ( n3142, g1750, n37 );
nor U12239 ( n3143, n3012, n3004 );
nor U12240 ( new_g27288_, n3078, n3079 );
nor U12241 ( n3078, g1739, n38 );
nor U12242 ( n3079, n3012, n2938 );
nor U12243 ( new_g27263_, n3231, n3232 );
nor U12244 ( n3231, g1056, n34 );
nor U12245 ( n3232, n3100, n3092 );
nor U12246 ( new_g27271_, n3179, n3180 );
nor U12247 ( n3179, g1045, n35 );
nor U12248 ( n3180, n3100, n3025 );
nor U12249 ( new_g27256_, n3299, n3300 );
nor U12250 ( n3299, g369, n31 );
nor U12251 ( n3300, n3205, n3196 );
nor U12252 ( new_g27259_, n3268, n3269 );
nor U12253 ( n3268, g358, n32 );
nor U12254 ( n3269, n3205, n3113 );
nand U12255 ( n4332, n4333, n4334 );
nand U12256 ( n4333, g3142, n4335 );
nand U12257 ( n4334, n148, n49 );
nand U12258 ( n4303, g3161, n4304 );
nand U12259 ( n4309, n4315, n4316 );
nand U12260 ( n4315, g3179, n4318 );
nand U12261 ( n4316, g3164, n4317 );
nor U12262 ( n4280, n4281, n4282 );
nand U12263 ( n4282, n4283, n4284 );
nand U12264 ( n4281, n4287, n4288 );
nand U12265 ( n4284, g3170, n4285 );
nand U12266 ( n4293, g3127, n151 );
nand U12267 ( n4288, g3088, n4289 );
nand U12268 ( n4310, n4311, n4312 );
nand U12269 ( n4312, g3176, n4313 );
nand U12270 ( n4311, g3182, n4314 );
and U12271 ( n6153, n6190, n145 );
nor U12272 ( n6190, g3201, n7112 );
and U12273 ( n6178, g3103, n4296 );
nand U12274 ( n6132, g3204, n6155 );
nor U12275 ( n6155, g3207, g3188 );
and U12276 ( n4308, n6169, g3201 );
nor U12277 ( n6169, n6168, n6132 );
and U12278 ( n6187, g3102, n4285 );
and U12279 ( n4343, n4296, g3091 );
and U12280 ( n4353, n4285, g3087 );
nor U12281 ( n6180, g3128, n4709 );
nand U12282 ( n6901, n6981, n1582 );
nor U12283 ( n6981, g2637, g2633 );
nand U12284 ( n6703, n6781, n2024 );
nor U12285 ( n6781, g1943, g1939 );
nand U12286 ( n6508, n6587, n3869 );
nor U12287 ( n6587, g1249, g1245 );
and U12288 ( n4286, n6189, n145 );
nor U12289 ( n6189, g3201, n6132 );
nand U12290 ( n6315, n6393, n6394 );
nor U12291 ( n6393, new_g21851_, n6395 );
nor U12292 ( n6394, g563, g559 );
nor U12293 ( n6395, g499, n7162 );
nor U12294 ( n1442, g2397, n7432 );
nor U12295 ( n1488, g1703, n7444 );
nor U12296 ( n1534, g1009, n7456 );
nor U12297 ( n1575, g322, n7468 );
nand U12298 ( n1434, n1439, n1440 );
or U12299 ( n1440, n7425, g2396 );
nor U12300 ( n1439, n1441, n1442 );
nor U12301 ( n1441, g2398, n7429 );
nand U12302 ( n1478, n1484, n1486 );
or U12303 ( n1486, n7437, g1702 );
nor U12304 ( n1484, n1487, n1488 );
nor U12305 ( n1487, g1704, n7441 );
nand U12306 ( n1526, n1531, n1532 );
or U12307 ( n1532, n7449, g1008 );
nor U12308 ( n1531, n1533, n1534 );
nor U12309 ( n1533, g1010, n7453 );
nand U12310 ( n1567, n1572, n1573 );
or U12311 ( n1573, n7461, g321 );
nor U12312 ( n1572, n1574, n1575 );
nor U12313 ( n1574, g323, n7465 );
nand U12314 ( n4283, g3167, n4286 );
and U12315 ( n6183, g3107, n4290 );
nand U12316 ( n4295, g3173, n4296 );
nand U12317 ( n4307, g3135, n4308 );
and U12318 ( n4349, n4290, g3095 );
nand U12319 ( new_g21851_, n6999, n7000 );
nand U12320 ( n6999, g544, g499 );
nand U12321 ( n7000, n7001, g548 );
nor U12322 ( n7001, g6485, g499 );
nand U12323 ( n3869, n6993, n6994 );
or U12324 ( n6993, g1230, n7156 );
nand U12325 ( n6994, n6996, n6997 );
nand U12326 ( n6997, g1234, n7122 );
nand U12327 ( n2024, n6988, n6989 );
or U12328 ( n6988, g1924, n7182 );
nand U12329 ( n6989, n6990, n6991 );
nand U12330 ( n6991, g1928, n7155 );
nor U12331 ( n6990, g1880, n6992 );
nor U12332 ( n6992, n3869, n7155 );
nor U12333 ( n6984, g2574, n6987 );
nor U12334 ( n6987, n2024, n7160 );
nor U12335 ( n6996, g1186, n6998 );
and U12336 ( n6998, new_g21851_, g6750 );
nand U12337 ( n1582, n6982, n6983 );
or U12338 ( n6982, g2618, n7183 );
nand U12339 ( n6983, n6984, n6985 );
nand U12340 ( n6985, g2622, n7160 );
nand U12341 ( n4287, g3185, n4290 );
nand U12342 ( n6138, n7367, n7368 );
nand U12343 ( n7367, n4308, g3139 );
or U12344 ( n7368, g3133, n4709 );
nand U12345 ( n6126, g3188, n7109 );
and U12346 ( n3419, n3462, n3463 );
nand U12347 ( n3462, n306, n7214 );
nand U12348 ( n3463, g996, n2794 );
and U12349 ( n3359, n3388, n3389 );
nand U12350 ( n3388, n525, n7215 );
nand U12351 ( n3389, g2384, n2750 );
and U12352 ( n3382, n3425, n3426 );
nand U12353 ( n3425, n415, n7216 );
nand U12354 ( n3426, g1690, n2773 );
and U12355 ( n3459, n3495, n3496 );
nand U12356 ( n3495, n185, n7217 );
nand U12357 ( n3496, g309, n2810 );
nand U12358 ( new_g26822_, n3376, n3377 );
nand U12359 ( n3376, g2507, n7430 );
nand U12360 ( n3377, n3359, g7264 );
nand U12361 ( new_g26809_, n3452, n3453 );
nand U12362 ( n3452, g1119, n7454 );
nand U12363 ( n3453, n3419, g6712 );
nand U12364 ( new_g26817_, n3386, n3387 );
nand U12365 ( n3386, g2504, n7433 );
nand U12366 ( n3387, n3359, g5555 );
nand U12367 ( new_g26811_, n3423, n3424 );
nand U12368 ( n3423, g1810, n7445 );
nand U12369 ( n3424, n3382, g5511 );
nand U12370 ( new_g26815_, n3413, n3414 );
nand U12371 ( n3413, g1813, n7442 );
nand U12372 ( n3414, n3382, g7014 );
nand U12373 ( new_g26806_, n3460, n3461 );
nand U12374 ( n3460, g1116, n7457 );
nand U12375 ( n3461, n3419, g5472 );
nand U12376 ( new_g26803_, n3493, n3494 );
nand U12377 ( n3493, g429, n7469 );
nand U12378 ( n3494, n3459, g5437 );
nand U12379 ( new_g26804_, n3490, n3491 );
nand U12380 ( n3490, g432, n7466 );
nand U12381 ( n3491, n3459, g6447 );
nand U12382 ( new_g26825_, n3357, n3358 );
nand U12383 ( n3357, g2510, n7425 );
nand U12384 ( n3358, n3359, g2476 );
nand U12385 ( new_g26820_, n3380, n3381 );
nand U12386 ( n3380, g1816, n7437 );
nand U12387 ( n3381, n3382, g1782 );
nand U12388 ( new_g26813_, n3417, n3418 );
nand U12389 ( n3417, g1122, n7449 );
nand U12390 ( n3418, n3419, g1088 );
nand U12391 ( new_g26807_, n3457, n3458 );
nand U12392 ( n3457, g435, n7461 );
nand U12393 ( n3458, n3459, g401 );
nand U12394 ( n6117, n6118, n6119 );
nand U12395 ( n6118, g3151, n4335 );
nand U12396 ( n6119, g3201, n6120 );
nand U12397 ( n6120, n6121, n6122 );
nand U12398 ( n6122, n6123, n6124 );
nor U12399 ( n6124, g185, n7112 );
nor U12400 ( n6123, n6125, n6126 );
nor U12401 ( n3651, g1091, n7454 );
and U12402 ( n1632, n3649, n3650 );
or U12403 ( n3650, n7449, g1089 );
nor U12404 ( n3649, n3651, n3652 );
nor U12405 ( n3652, g1090, n7457 );
nor U12406 ( n4185, g2479, n7429 );
and U12407 ( n1610, n4183, n4184 );
or U12408 ( n4184, n7425, g2477 );
nor U12409 ( n4183, n4185, n4186 );
nor U12410 ( n4186, g2478, n7432 );
nor U12411 ( new_g22173_, n5147, n5149 );
nor U12412 ( n5147, g2239, n515 );
nor U12413 ( n5149, n511, n5133 );
nor U12414 ( new_g22185_, n5127, n5128 );
nor U12415 ( n5127, g2240, n518 );
nor U12416 ( n5128, n511, n5121 );
nor U12417 ( new_g22152_, n5194, n5195 );
nor U12418 ( n5194, g1545, n406 );
nor U12419 ( n5195, n402, n5168 );
nor U12420 ( new_g22169_, n5161, n5162 );
nor U12421 ( n5161, g1546, n408 );
nor U12422 ( n5162, n402, n5141 );
nor U12423 ( new_g22129_, n5240, n5241 );
nor U12424 ( n5240, g851, n297 );
nor U12425 ( n5241, n293, n5214 );
nor U12426 ( new_g22148_, n5207, n5208 );
nor U12427 ( n5207, g852, n299 );
nor U12428 ( n5208, n293, n5176 );
nor U12429 ( new_g22103_, n5283, n5284 );
nor U12430 ( n5283, g163, n176 );
nor U12431 ( n5284, n172, n5258 );
nor U12432 ( new_g22125_, n5252, n5253 );
nor U12433 ( n5252, g164, n178 );
nor U12434 ( n5253, n172, n5221 );
nor U12435 ( new_g22194_, n5117, n5118 );
nor U12436 ( n5117, g2238, n520 );
nor U12437 ( n5118, n511, n5116 );
nor U12438 ( new_g22180_, n5136, n5137 );
nor U12439 ( n5136, g1544, n410 );
nor U12440 ( n5137, n402, n5126 );
nor U12441 ( new_g22164_, n5171, n5172 );
nor U12442 ( n5171, g850, n301 );
nor U12443 ( n5172, n293, n5146 );
nor U12444 ( new_g22143_, n5217, n5218 );
nor U12445 ( n5217, g162, n180 );
nor U12446 ( n5218, n172, n5181 );
nor U12447 ( n3552, g1784, n7445 );
nor U12448 ( n3751, g403, n7469 );
and U12449 ( n1621, n3549, n3550 );
or U12450 ( n3550, n7437, g1783 );
nor U12451 ( n3549, n3551, n3552 );
nor U12452 ( n3551, g1785, n7441 );
and U12453 ( n1640, n3748, n3749 );
or U12454 ( n3749, n7461, g402 );
nor U12455 ( n3748, n3750, n3751 );
nor U12456 ( n3750, g404, n7466 );
nor U12457 ( new_g22155_, n5182, n5183 );
nor U12458 ( n5182, g2236, n515 );
nor U12459 ( n5183, n510, n5133 );
nor U12460 ( new_g22172_, n5154, n5155 );
nor U12461 ( n5154, g2237, n518 );
nor U12462 ( n5155, n510, n5121 );
nor U12463 ( new_g22132_, n5230, n5231 );
nor U12464 ( n5230, g1542, n406 );
nor U12465 ( n5231, n401, n5168 );
nor U12466 ( new_g22151_, n5200, n5201 );
nor U12467 ( n5200, g1543, n408 );
nor U12468 ( n5201, n401, n5141 );
nor U12469 ( new_g22106_, n5273, n5274 );
nor U12470 ( n5273, g848, n297 );
nor U12471 ( n5274, n292, n5214 );
nor U12472 ( new_g22128_, n5246, n5247 );
nor U12473 ( n5246, g849, n299 );
nor U12474 ( n5247, n292, n5176 );
nor U12475 ( new_g22081_, n5317, n5318 );
nor U12476 ( n5317, g160, n176 );
nor U12477 ( n5318, n171, n5258 );
nor U12478 ( new_g22102_, n5290, n5291 );
nor U12479 ( n5290, g161, n178 );
nor U12480 ( n5291, n171, n5221 );
nor U12481 ( new_g22184_, n5129, n5130 );
nor U12482 ( n5129, g2235, n520 );
nor U12483 ( n5130, n510, n5116 );
nor U12484 ( new_g22168_, n5163, n5164 );
nor U12485 ( n5163, g1541, n410 );
nor U12486 ( n5164, n401, n5126 );
nor U12487 ( new_g22147_, n5209, n5210 );
nor U12488 ( n5209, g847, n301 );
nor U12489 ( n5210, n292, n5146 );
nor U12490 ( new_g22124_, n5254, n5255 );
nor U12491 ( n5254, g159, n180 );
nor U12492 ( n5255, n171, n5181 );
nand U12493 ( n6121, n6127, n149 );
nor U12494 ( n6127, g3207, g3204 );
nand U12495 ( n2883, n2995, g7264 );
nand U12496 ( n3025, n3185, g6712 );
nand U12497 ( n2917, n2995, g5555 );
nand U12498 ( n2938, n3083, g7014 );
nand U12499 ( n3004, n3083, g5511 );
nand U12500 ( n3092, n3185, g5472 );
nand U12501 ( n3113, n3273, g6447 );
nand U12502 ( n3196, n3273, g5437 );
nand U12503 ( n2859, n2995, g2476 );
nand U12504 ( n2897, n3083, g1782 );
nand U12505 ( n2952, n3185, g1088 );
nand U12506 ( n3039, n3273, g401 );
and U12507 ( n6149, g3207, g3188 );
nand U12508 ( n7052, n6250, n6296 );
nand U12509 ( n6296, n6297, n247 );
nor U12510 ( n6297, n6298, n6299 );
nor U12511 ( n6298, g533, n226 );
nand U12512 ( n7053, n6269, n6304 );
nand U12513 ( n6304, n6305, n247 );
nor U12514 ( n6305, n6306, n6307 );
nor U12515 ( n6306, g531, n226 );
nand U12516 ( n7050, n6269, n6270 );
nand U12517 ( n6270, n6271, n247 );
nor U12518 ( n6271, n6272, n6273 );
nor U12519 ( n6272, g530, n226 );
nand U12520 ( n7054, n6260, n6316 );
nand U12521 ( n6316, n6317, n247 );
nor U12522 ( n6317, n6318, n6319 );
nor U12523 ( n6318, g529, n226 );
nand U12524 ( n7047, n6250, n6251 );
nand U12525 ( n6251, n6252, n247 );
nor U12526 ( n6252, n6253, n6254 );
nor U12527 ( n6253, g534, n226 );
nand U12528 ( n7048, n6260, n6261 );
nand U12529 ( n6261, n6262, n247 );
nor U12530 ( n6262, n6263, n6264 );
nor U12531 ( n6263, g532, n226 );
nor U12532 ( n6284, g536, n226 );
nor U12533 ( n6236, g537, n226 );
nand U12534 ( n7077, n6812, n6813 );
nand U12535 ( n6813, n6814, n581 );
nor U12536 ( n6814, n6815, n6816 );
nor U12537 ( n6815, g2607, n233 );
nand U12538 ( n7066, n6621, n6622 );
nand U12539 ( n6622, n6623, n464 );
nor U12540 ( n6623, n6624, n6625 );
nor U12541 ( n6624, g1913, n236 );
nand U12542 ( n7056, n6426, n6427 );
nand U12543 ( n6427, n6428, n355 );
nor U12544 ( n6428, n6429, n6430 );
nor U12545 ( n6429, g1219, n239 );
nand U12546 ( n7061, n6471, n6472 );
nand U12547 ( n6472, n6473, n355 );
nor U12548 ( n6473, n6474, n6475 );
nor U12549 ( n6474, g1217, n239 );
nand U12550 ( n7082, n6812, n6874 );
nand U12551 ( n6874, n6875, n581 );
nor U12552 ( n6875, n6877, n6878 );
nor U12553 ( n6877, g2608, n233 );
nand U12554 ( n7083, n6860, n6886 );
nand U12555 ( n6886, n6887, n581 );
nor U12556 ( n6887, n6888, n6889 );
nor U12557 ( n6888, g2604, n233 );
nand U12558 ( n7081, n6860, n6861 );
nand U12559 ( n6861, n6862, n581 );
nor U12560 ( n6862, n6863, n6864 );
nor U12561 ( n6863, g2605, n233 );
nand U12562 ( n7072, n6621, n6679 );
nand U12563 ( n6679, n6680, n464 );
nor U12564 ( n6680, n6681, n6682 );
nor U12565 ( n6681, g1914, n236 );
nand U12566 ( n7073, n6666, n6689 );
nand U12567 ( n6689, n6690, n464 );
nor U12568 ( n6690, n6691, n6692 );
nor U12569 ( n6691, g1910, n236 );
nand U12570 ( n7071, n6666, n6667 );
nand U12571 ( n6667, n6668, n464 );
nor U12572 ( n6668, n6669, n6670 );
nor U12573 ( n6669, g1911, n236 );
nand U12574 ( n7070, n6633, n6657 );
nand U12575 ( n6657, n6658, n464 );
nor U12576 ( n6658, n6659, n6660 );
nor U12577 ( n6659, g1909, n236 );
nand U12578 ( n7068, n6633, n6634 );
nand U12579 ( n6634, n6635, n464 );
nor U12580 ( n6635, n6636, n6637 );
nor U12581 ( n6636, g1912, n236 );
nand U12582 ( n7060, n6438, n6462 );
nand U12583 ( n6462, n6463, n355 );
nor U12584 ( n6463, n6464, n6465 );
nor U12585 ( n6464, g1215, n239 );
nand U12586 ( n7057, n6438, n6439 );
nand U12587 ( n6439, n6440, n355 );
nor U12588 ( n6440, n6441, n6442 );
nor U12589 ( n6441, g1218, n239 );
nand U12590 ( n7080, n6824, n6850 );
nand U12591 ( n6850, n6851, n581 );
nor U12592 ( n6851, n6852, n6853 );
nor U12593 ( n6852, g2603, n233 );
nand U12594 ( n7078, n6824, n6825 );
nand U12595 ( n6825, n6826, n581 );
nor U12596 ( n6826, n6827, n6828 );
nor U12597 ( n6827, g2606, n233 );
nand U12598 ( n7062, n6426, n6484 );
nand U12599 ( n6484, n6485, n355 );
nor U12600 ( n6485, n6486, n6487 );
nor U12601 ( n6486, g1220, n239 );
nand U12602 ( n7063, n6471, n6494 );
nand U12603 ( n6494, n6495, n355 );
nor U12604 ( n6495, n6496, n6497 );
nor U12605 ( n6496, g1216, n239 );
nor U12606 ( n6906, g2611, n233 );
nor U12607 ( n6836, g2610, n233 );
nor U12608 ( n6707, g1917, n236 );
nor U12609 ( n6645, g1916, n236 );
nor U12610 ( n6512, g1223, n239 );
nor U12611 ( n6450, g1222, n239 );
nor U12612 ( n6136, g2984, g2985 );
nand U12613 ( n6135, g3120, n49 );
nand U12614 ( new_g28349_, n2503, n2504 );
nand U12615 ( n2503, g617, n7171 );
nand U12616 ( n2504, g6642, n2395 );
nor U12617 ( n3256, g582, n7162 );
nand U12618 ( n2639, n3253, n3254 );
or U12619 ( n3254, n7169, g581 );
nor U12620 ( n3253, n3255, n3256 );
nor U12621 ( n3255, g583, n7171 );
nand U12622 ( new_g28345_, n2597, n2598 );
nand U12623 ( n2597, g614, n7162 );
nand U12624 ( n2598, g6485, n2395 );
nand U12625 ( new_g28353_, n2393, n2394 );
nand U12626 ( n2393, g620, n7169 );
nand U12627 ( n2394, g550, n2395 );
nand U12628 ( new_g28342_, n2612, n2613 );
nand U12629 ( n2612, g605, n7162 );
nand U12630 ( n2613, n2507, g6485 );
nand U12631 ( new_g28344_, n2610, n2611 );
nand U12632 ( n2610, g608, n7171 );
nand U12633 ( n2611, n2507, g6642 );
nand U12634 ( new_g28348_, n2505, n2506 );
nand U12635 ( n2505, g611, n7169 );
nand U12636 ( n2506, n2507, g550 );
nand U12637 ( n2535, n3164, n3165 );
or U12638 ( n3165, n7167, g1267 );
nor U12639 ( n3164, n3166, n3167 );
nor U12640 ( n3166, g1269, n7159 );
nand U12641 ( n2424, n3063, n3064 );
or U12642 ( n3064, n7168, g1961 );
nor U12643 ( n3063, n3065, n3066 );
nor U12644 ( n3065, g1963, n7158 );
nor U12645 ( n3066, g1962, n7155 );
nor U12646 ( n3167, g1268, n7122 );
nand U12647 ( new_g28357_, n2373, n2374 );
nand U12648 ( n2373, g1994, n7155 );
nand U12649 ( n2374, g7052, n2259 );
nand U12650 ( new_g28360_, n2281, n2282 );
nand U12651 ( n2281, g1306, n7167 );
nand U12652 ( n2282, g1236, n2283 );
nand U12653 ( new_g28366_, n2257, n2258 );
nand U12654 ( n2257, g2000, n7168 );
nand U12655 ( n2258, g1930, n2259 );
nand U12656 ( new_g28351_, n2488, n2489 );
nand U12657 ( n2488, g1300, n7122 );
nand U12658 ( n2489, g6750, n2283 );
nand U12659 ( new_g28355_, n2388, n2389 );
nand U12660 ( n2388, g1303, n7159 );
nand U12661 ( n2389, g6944, n2283 );
nand U12662 ( new_g28362_, n2276, n2277 );
nand U12663 ( n2276, g1997, n7158 );
nand U12664 ( n2277, g7194, n2259 );
nand U12665 ( n6137, n7369, n7370 );
nand U12666 ( n6134, g3114, n6137 );
nand U12667 ( n2311, n2975, n2976 );
or U12668 ( n2976, n7179, g2655 );
nor U12669 ( n2975, n2977, n2978 );
nor U12670 ( n2977, g2657, n7161 );
nor U12671 ( n2978, g2656, n7160 );
nand U12672 ( new_g28371_, n2249, n2250 );
nand U12673 ( n2249, g2694, n7179 );
nand U12674 ( n2250, g2624, n2251 );
nand U12675 ( new_g28368_, n2252, n2253 );
nand U12676 ( n2252, g2691, n7161 );
nand U12677 ( n2253, g7390, n2251 );
nand U12678 ( new_g28364_, n2260, n2261 );
nand U12679 ( n2260, g2688, n7160 );
nand U12680 ( n2261, g7302, n2251 );
nand U12681 ( new_g28350_, n2501, n2502 );
nand U12682 ( n2501, g1294, n7159 );
nand U12683 ( n2502, n2392, g6944 );
nand U12684 ( new_g28354_, n2390, n2391 );
nand U12685 ( n2390, g1297, n7167 );
nand U12686 ( n2391, n2392, g1236 );
nand U12687 ( new_g28361_, n2278, n2279 );
nand U12688 ( n2278, g1991, n7168 );
nand U12689 ( n2279, n2280, g1930 );
nand U12690 ( new_g28346_, n2508, n2509 );
nand U12691 ( n2508, g1291, n7122 );
nand U12692 ( n2509, n2392, g6750 );
nand U12693 ( new_g28356_, n2386, n2387 );
nand U12694 ( n2386, g1988, n7158 );
nand U12695 ( n2387, n2280, g7194 );
nand U12696 ( new_g28352_, n2396, n2397 );
nand U12697 ( n2396, g1985, n7155 );
nand U12698 ( n2397, n2280, g7052 );
nand U12699 ( new_g28367_, n2254, n2255 );
nand U12700 ( n2254, g2685, n7179 );
nand U12701 ( n2255, n2256, g2624 );
nand U12702 ( new_g28363_, n2274, n2275 );
nand U12703 ( n2274, g2682, n7161 );
nand U12704 ( n2275, n2256, g7390 );
nand U12705 ( new_g28358_, n2284, n2285 );
nand U12706 ( n2284, g2679, n7160 );
nand U12707 ( n2285, n2256, g7302 );
nand U12708 ( n2632, n3249, n3250 );
or U12709 ( n3250, n7169, g578 );
nor U12710 ( n3249, n3251, n3252 );
nor U12711 ( n3251, g580, n7171 );
nor U12712 ( n3252, g579, n7162 );
nor U12713 ( n3260, g585, n7162 );
nand U12714 ( n2651, n3257, n3258 );
or U12715 ( n3258, n7169, g584 );
nor U12716 ( n3257, n3259, n3260 );
nor U12717 ( n3259, g586, n7171 );
nand U12718 ( n2029, g2138, n2713 );
nand U12719 ( n2714, g2147, n3338 );
nand U12720 ( n2035, g1444, n2717 );
nand U12721 ( n2718, g1453, n3342 );
nand U12722 ( n2041, g758, n2721 );
nand U12723 ( n2722, g767, n3346 );
nand U12724 ( n2047, g70, n2725 );
nand U12725 ( n2726, g79, n3350 );
nand U12726 ( n3339, g2156, n4263 );
nand U12727 ( n3343, g1462, n4267 );
nand U12728 ( n3347, g776, n4271 );
nand U12729 ( n3351, g88, n4275 );
nand U12730 ( n1645, g2129, n2028 );
nand U12731 ( n1648, g1435, n2034 );
nand U12732 ( n1651, g749, n2040 );
nand U12733 ( n1654, g61, n2046 );
nor U12734 ( new_g29582_, n29, n1643 );
xor U12735 ( n1643, n1644, g2120 );
nand U12736 ( n1644, g2124, n30 );
not U12737 ( n30, n1645 );
nor U12738 ( new_g29581_, n27, n1646 );
xor U12739 ( n1646, n1647, g1426 );
nand U12740 ( n1647, g1430, n28 );
not U12741 ( n28, n1648 );
nor U12742 ( new_g29580_, n25, n1649 );
xor U12743 ( n1649, n1650, g740 );
nand U12744 ( n1650, g744, n26 );
not U12745 ( n26, n1651 );
nor U12746 ( new_g29579_, n23, n1652 );
xor U12747 ( n1652, n1653, g52 );
nand U12748 ( n1653, g56, n24 );
not U12749 ( n24, n1654 );
and U12750 ( n4263, g2160, n4264 );
and U12751 ( n4267, g1466, n4268 );
and U12752 ( n4271, g780, n4272 );
and U12753 ( n4275, g92, n4276 );
nand U12754 ( n2528, n3160, n3161 );
or U12755 ( n3161, n7167, g1264 );
nor U12756 ( n3160, n3162, n3163 );
nor U12757 ( n3162, g1266, n7159 );
nand U12758 ( n2416, n3059, n3060 );
or U12759 ( n3060, n7168, g1958 );
nor U12760 ( n3059, n3061, n3062 );
nor U12761 ( n3061, g1960, n7158 );
nor U12762 ( n3062, g1959, n7155 );
nor U12763 ( n3163, g1265, n7122 );
nand U12764 ( n2547, n3168, n3169 );
or U12765 ( n3169, n7167, g1270 );
nor U12766 ( n3168, n3170, n3171 );
nor U12767 ( n3170, g1272, n7159 );
nand U12768 ( n2436, n3067, n3068 );
or U12769 ( n3068, n7168, g1964 );
nor U12770 ( n3067, n3069, n3070 );
nor U12771 ( n3069, g1966, n7158 );
nor U12772 ( n3070, g1965, n7155 );
nor U12773 ( n3171, g1271, n7122 );
nand U12774 ( n2304, n2971, n2972 );
or U12775 ( n2972, n7179, g2652 );
nor U12776 ( n2971, n2973, n2974 );
nor U12777 ( n2973, g2654, n7161 );
nor U12778 ( n2974, g2653, n7160 );
nand U12779 ( n2323, n2979, n2980 );
or U12780 ( n2980, n7179, g2658 );
nor U12781 ( n2979, n2981, n2982 );
nor U12782 ( n2981, g2660, n7161 );
nor U12783 ( n2982, g2659, n7160 );
nand U12784 ( n4830, n621, n5427 );
nand U12785 ( n5427, n5428, n640 );
nand U12786 ( n5428, n5429, n5430 );
and U12787 ( n5429, g3018, g3032 );
nor U12788 ( n4461, n5426, g3234 );
nor U12789 ( new_g23359_, n619, n4990 );
xor U12790 ( n4990, n4832, g3028 );
nor U12791 ( new_g25202_, n619, n4683 );
xor U12792 ( n4683, n4684, g3032 );
nand U12793 ( n2060, n3880, n3881 );
nand U12794 ( n3880, g985, n7228 );
nand U12795 ( n3881, n3882, g986 );
nand U12796 ( n1590, n1591, n1592 );
nand U12797 ( n1591, g2380, n7430 );
nand U12798 ( n1592, new_g28903_, g7264 );
nor U12799 ( n2057, n2058, n2059 );
and U12800 ( n2059, n7442, g1686 );
nor U12801 ( n2058, n7441, n2060 );
and U12802 ( n3882, n7371, n7372 );
nand U12803 ( n7371, new_g21346_, g6712 );
nand U12804 ( n7372, n7454, g992 );
nand U12805 ( new_g21346_, n5494, n5495 );
or U12806 ( n5494, g299, g298 );
nand U12807 ( n5495, n5496, g305 );
and U12808 ( n5496, n7466, g299 );
and U12809 ( new_g28903_, n2055, n2056 );
nand U12810 ( n2055, g1679, n7247 );
nand U12811 ( n2056, n2057, g1680 );
nand U12812 ( n7036, n7039, n7041 );
nand U12813 ( n7041, n6137, n7121 );
nor U12814 ( n7039, g3147, n7042 );
nor U12815 ( n7042, g3142, n6136 );
nor U12816 ( new_g30055_, n1588, n1589 );
and U12817 ( n1589, g2373, n7287 );
nor U12818 ( n1588, n7287, n1590 );
nand U12819 ( g25489, n7032, n7033 );
nand U12820 ( n7033, n7034, n7035 );
nand U12821 ( n7032, n7036, n7035 );
nor U12822 ( n7034, g3151, g3142 );
nor U12823 ( n2110, g2503, n7429 );
nor U12824 ( n2189, g1115, n7453 );
nand U12825 ( n1680, n2108, n2109 );
or U12826 ( n2109, n7426, g2501 );
nor U12827 ( n2108, n2110, n2111 );
nor U12828 ( n2111, g2502, n7432 );
nand U12829 ( n1724, n2186, n2188 );
or U12830 ( n2188, n7450, g1113 );
nor U12831 ( n2186, n2189, n2190 );
nor U12832 ( n2190, g1114, n7456 );
nand U12833 ( n2624, n3245, n3246 );
or U12834 ( n3246, n7169, g575 );
nor U12835 ( n3245, n3247, n3248 );
nor U12836 ( n3247, g577, n7171 );
nor U12837 ( n3248, g576, n7162 );
nor U12838 ( new_g24446_, n4828, n4829 );
nor U12839 ( n4828, g3036, n4831 );
nand U12840 ( n4829, n4684, n4830 );
nand U12841 ( n1702, n2149, n2150 );
or U12842 ( n2150, n7438, g1807 );
nor U12843 ( n2149, n2151, n2152 );
nor U12844 ( n2151, g1809, n7441 );
nand U12845 ( n1744, n2221, n2222 );
or U12846 ( n2222, n7462, g426 );
nor U12847 ( n2221, n2224, n2225 );
nor U12848 ( n2224, g428, n7465 );
nor U12849 ( n2152, g1808, n7444 );
nor U12850 ( n2225, g427, n7468 );
nor U12851 ( new_g29355_, n27, n1656 );
xor U12852 ( n1656, g1430, n1648 );
nor U12853 ( new_g29354_, n25, n1657 );
xor U12854 ( n1657, g744, n1651 );
nor U12855 ( new_g29353_, n23, n1658 );
xor U12856 ( n1658, g56, n1654 );
nor U12857 ( new_g29357_, n29, n1655 );
xor U12858 ( n1655, g2124, n1645 );
nand U12859 ( n7035, g3147, n7037 );
nand U12860 ( n7037, n7038, g3142 );
nor U12861 ( n7038, n7121, n7091 );
nand U12862 ( n2520, n3156, n3157 );
or U12863 ( n3157, n7167, g1261 );
nor U12864 ( n3156, n3158, n3159 );
nor U12865 ( n3158, g1263, n7159 );
nand U12866 ( n2408, n3055, n3056 );
or U12867 ( n3056, n7168, g1955 );
nor U12868 ( n3055, n3057, n3058 );
nor U12869 ( n3057, g1957, n7158 );
nor U12870 ( n3058, g1956, n7155 );
nor U12871 ( n3159, g1262, n7122 );
nand U12872 ( n2296, n2967, n2968 );
or U12873 ( n2968, n7179, g2649 );
nor U12874 ( n2967, n2969, n2970 );
nor U12875 ( n2969, g2651, n7161 );
nor U12876 ( n2970, g2650, n7160 );
nor U12877 ( new_g26048_, n620, n4172 );
nor U12878 ( n4172, n621, n4173 );
not U12879 ( n620, n4175 );
xor U12880 ( n4173, g2998, n4174 );
nor U12881 ( n6934, g2782, n7163 );
nor U12882 ( n6734, g2088, n7164 );
nor U12883 ( n6539, g1394, n7165 );
and U12884 ( n4398, n6931, n6932 );
or U12885 ( n6932, n7178, g2781 );
nor U12886 ( n6931, n6933, n6934 );
nor U12887 ( n6933, g2783, n7172 );
and U12888 ( n4441, n6731, n6732 );
or U12889 ( n6732, n7177, g2087 );
nor U12890 ( n6731, n6733, n6734 );
nor U12891 ( n6733, g2089, n7173 );
and U12892 ( n4490, n6536, n6537 );
or U12893 ( n6537, n7176, g1393 );
nor U12894 ( n6536, n6538, n6539 );
nor U12895 ( n6538, g1395, n7174 );
nor U12896 ( n6938, g2776, n7163 );
nor U12897 ( n6947, g2800, n7163 );
nor U12898 ( n6738, g2082, n7164 );
nor U12899 ( n6747, g2106, n7164 );
nor U12900 ( n6543, g1388, n7165 );
nor U12901 ( n6552, g1412, n7165 );
and U12902 ( n4404, n6935, n6936 );
or U12903 ( n6936, n7178, g2775 );
nor U12904 ( n6935, n6937, n6938 );
nor U12905 ( n6937, g2777, n7172 );
and U12906 ( n4447, n6735, n6736 );
or U12907 ( n6736, n7177, g2081 );
nor U12908 ( n6735, n6737, n6738 );
nor U12909 ( n6737, g2083, n7173 );
and U12910 ( n4496, n6540, n6541 );
or U12911 ( n6541, n7176, g1387 );
nor U12912 ( n6540, n6542, n6543 );
nor U12913 ( n6542, g1389, n7174 );
and U12914 ( n4387, n6944, n6945 );
or U12915 ( n6945, n7178, g2799 );
nor U12916 ( n6944, n6946, n6947 );
nor U12917 ( n6946, g2801, n7172 );
and U12918 ( n4430, n6744, n6745 );
or U12919 ( n6745, n7177, g2105 );
nor U12920 ( n6744, n6746, n6747 );
nor U12921 ( n6746, g2107, n7173 );
and U12922 ( n4479, n6549, n6550 );
or U12923 ( n6550, n7176, g1411 );
nor U12924 ( n6549, n6551, n6552 );
nor U12925 ( n6551, g1413, n7174 );
nor U12926 ( n6951, g2797, n7163 );
nor U12927 ( n6751, g2103, n7164 );
nor U12928 ( n6556, g1409, n7165 );
and U12929 ( n4386, n6948, n6949 );
or U12930 ( n6949, n7178, g2796 );
nor U12931 ( n6948, n6950, n6951 );
nor U12932 ( n6950, g2798, n7172 );
and U12933 ( n4429, n6748, n6749 );
or U12934 ( n6749, n7177, g2102 );
nor U12935 ( n6748, n6750, n6751 );
nor U12936 ( n6750, g2104, n7173 );
and U12937 ( n4478, n6553, n6554 );
or U12938 ( n6554, n7176, g1408 );
nor U12939 ( n6553, n6555, n6556 );
nor U12940 ( n6555, g1410, n7174 );
nor U12941 ( n6344, g708, n7170 );
and U12942 ( n4529, n6341, n6342 );
or U12943 ( n6342, n7181, g707 );
nor U12944 ( n6341, n6343, n6344 );
nor U12945 ( n6343, g709, n7180 );
nor U12946 ( n6348, g702, n7170 );
nor U12947 ( n6357, g726, n7170 );
and U12948 ( n4535, n6345, n6346 );
or U12949 ( n6346, n7181, g701 );
nor U12950 ( n6345, n6347, n6348 );
nor U12951 ( n6347, g703, n7180 );
and U12952 ( n4518, n6354, n6355 );
or U12953 ( n6355, n7181, g725 );
nor U12954 ( n6354, n6356, n6357 );
nor U12955 ( n6356, g727, n7180 );
nor U12956 ( n6361, g723, n7170 );
and U12957 ( n4517, n6358, n6359 );
or U12958 ( n6359, n7181, g722 );
nor U12959 ( n6358, n6360, n6361 );
nor U12960 ( n6360, g724, n7180 );
nand U12961 ( n4393, n6973, n6974 );
or U12962 ( n6974, n7178, g2790 );
nor U12963 ( n6973, n6975, n6976 );
nor U12964 ( n6975, g2792, n7172 );
nand U12965 ( n4436, n6773, n6774 );
or U12966 ( n6774, n7177, g2096 );
nor U12967 ( n6773, n6775, n6776 );
nor U12968 ( n6775, g2098, n7173 );
nand U12969 ( n4485, n6578, n6579 );
or U12970 ( n6579, n7176, g1402 );
nor U12971 ( n6578, n6580, n6581 );
nor U12972 ( n6580, g1404, n7174 );
nor U12973 ( n6976, g2791, n7163 );
nor U12974 ( n6776, g2097, n7164 );
nor U12975 ( n6581, g1403, n7165 );
nor U12976 ( n6269, n227, n6312 );
and U12977 ( n6312, n6313, n6243 );
not U12978 ( n227, n6250 );
and U12979 ( n6313, n6314, g499 );
nand U12980 ( n6952, n6967, n596 );
nor U12981 ( n6967, n6972, n4393 );
nor U12982 ( n6972, n6977, n6978 );
nor U12983 ( n6977, g2812, n7163 );
nand U12984 ( n6752, n6767, n478 );
nor U12985 ( n6767, n6772, n4436 );
nor U12986 ( n6772, n6777, n6778 );
nor U12987 ( n6777, g2118, n7164 );
nand U12988 ( n6557, n6572, n370 );
nor U12989 ( n6572, n6577, n4485 );
nor U12990 ( n6577, n6582, n6583 );
nor U12991 ( n6582, g1424, n7165 );
nor U12992 ( n6860, n234, n6893 );
and U12993 ( n6893, n6895, n6843 );
not U12994 ( n234, n6812 );
and U12995 ( n6895, n6859, g2574 );
nor U12996 ( n6666, n237, n6696 );
and U12997 ( n6696, n6697, n6651 );
not U12998 ( n237, n6621 );
and U12999 ( n6697, n6665, g1880 );
nor U13000 ( n6471, n240, n6501 );
and U13001 ( n6501, n6502, n6456 );
not U13002 ( n240, n6426 );
and U13003 ( n6502, n6470, g1186 );
nand U13004 ( n4524, n6383, n6384 );
or U13005 ( n6384, n7181, g716 );
nor U13006 ( n6383, n6385, n6386 );
nor U13007 ( n6385, g718, n7180 );
nor U13008 ( n6386, g717, n7170 );
nand U13009 ( n6362, n6377, n261 );
nor U13010 ( n6377, n6382, n4524 );
nor U13011 ( n6382, n6387, n6388 );
nor U13012 ( n6387, g738, n7170 );
nor U13013 ( n6962, g2773, n7163 );
nor U13014 ( n6762, g2079, n7164 );
nor U13015 ( n6567, g1385, n7165 );
nand U13016 ( n6911, n6959, n6960 );
or U13017 ( n6960, n7178, g2772 );
nor U13018 ( n6959, n6961, n6962 );
nor U13019 ( n6961, g2774, n7172 );
nand U13020 ( n6712, n6759, n6760 );
or U13021 ( n6760, n7177, g2078 );
nor U13022 ( n6759, n6761, n6762 );
nor U13023 ( n6761, g2080, n7173 );
nand U13024 ( n6517, n6564, n6565 );
or U13025 ( n6565, n7176, g1384 );
nor U13026 ( n6564, n6566, n6567 );
nor U13027 ( n6566, g1386, n7174 );
nand U13028 ( n6869, n6963, n6964 );
or U13029 ( n6964, n7178, g2787 );
nor U13030 ( n6963, n6965, n6966 );
nor U13031 ( n6965, g2789, n7172 );
nand U13032 ( n6674, n6763, n6764 );
or U13033 ( n6764, n7177, g2093 );
nor U13034 ( n6763, n6765, n6766 );
nor U13035 ( n6765, g2095, n7173 );
nand U13036 ( n6479, n6568, n6569 );
or U13037 ( n6569, n7176, g1399 );
nor U13038 ( n6568, n6570, n6571 );
nor U13039 ( n6570, g1401, n7174 );
nor U13040 ( n6966, g2788, n7163 );
nor U13041 ( n6766, g2094, n7164 );
nor U13042 ( n6571, g1400, n7165 );
nand U13043 ( n6242, n6369, n6370 );
or U13044 ( n6370, n7181, g698 );
nor U13045 ( n6369, n6371, n6372 );
nor U13046 ( n6371, g700, n7180 );
nor U13047 ( n6372, g699, n7170 );
nand U13048 ( n3077, n3217, n3218 );
or U13049 ( n3218, n7438, g1742 );
nor U13050 ( n3217, n3219, n3220 );
nor U13051 ( n3220, g1750, n7444 );
nor U13052 ( n3130, g2433, n7429 );
nor U13053 ( n3219, g1739, n7442 );
nor U13054 ( n3287, g1045, n7453 );
nand U13055 ( n2989, n3128, n3129 );
or U13056 ( n3129, n7426, g2436 );
nor U13057 ( n3128, n3130, n3131 );
nor U13058 ( n3131, g2444, n7432 );
nand U13059 ( n3178, n3285, n3286 );
or U13060 ( n3286, n7450, g1048 );
nor U13061 ( n3285, n3287, n3288 );
nor U13062 ( n3288, g1056, n7456 );
nand U13063 ( n6311, n6373, n6374 );
or U13064 ( n6374, n7181, g713 );
nor U13065 ( n6373, n6375, n6376 );
nor U13066 ( n6375, g715, n7180 );
nor U13067 ( n6376, g714, n7170 );
nor U13068 ( n3320, g369, n7468 );
nand U13069 ( n3267, n3317, n3318 );
or U13070 ( n3318, n7462, g361 );
nor U13071 ( n3317, n3319, n3320 );
nor U13072 ( n3319, g358, n7465 );
nor U13073 ( new_g29111_, n2030, n2031 );
nor U13074 ( n2030, g1435, n2034 );
nand U13075 ( n2031, n1648, n2033 );
nor U13076 ( new_g29110_, n2037, n2038 );
nor U13077 ( n2037, g749, n2040 );
nand U13078 ( n2038, n1651, n2039 );
nor U13079 ( new_g29109_, n2042, n2043 );
nor U13080 ( n2042, g61, n2046 );
nand U13081 ( n2043, n1654, n2044 );
nor U13082 ( new_g29112_, n2025, n2026 );
nor U13083 ( n2025, g2129, n2028 );
nand U13084 ( n2026, n1645, n2027 );
nand U13085 ( n4392, n6968, n6969 );
or U13086 ( n6969, n7178, g2793 );
nor U13087 ( n6968, n6970, n6971 );
nor U13088 ( n6970, g2795, n7172 );
nand U13089 ( n4435, n6768, n6769 );
or U13090 ( n6769, n7177, g2099 );
nor U13091 ( n6768, n6770, n6771 );
nor U13092 ( n6770, g2101, n7173 );
nand U13093 ( n4484, n6573, n6574 );
or U13094 ( n6574, n7176, g1405 );
nor U13095 ( n6573, n6575, n6576 );
nor U13096 ( n6575, g1407, n7174 );
nor U13097 ( n6971, g2794, n7163 );
nor U13098 ( n6771, g2100, n7164 );
nor U13099 ( n6576, g1406, n7165 );
nor U13100 ( n6958, g2785, n7163 );
nor U13101 ( n6758, g2091, n7164 );
nor U13102 ( n6563, g1397, n7165 );
nand U13103 ( n6832, n6955, n6956 );
or U13104 ( n6956, n7178, g2784 );
nor U13105 ( n6955, n6957, n6958 );
nor U13106 ( n6957, g2786, n7172 );
nand U13107 ( n6641, n6755, n6756 );
or U13108 ( n6756, n7177, g2090 );
nor U13109 ( n6755, n6757, n6758 );
nor U13110 ( n6757, g2092, n7173 );
nand U13111 ( n6446, n6560, n6561 );
or U13112 ( n6561, n7176, g1396 );
nor U13113 ( n6560, n6562, n6563 );
nor U13114 ( n6562, g1398, n7174 );
nand U13115 ( new_g22002_, n4830, n5424 );
nand U13116 ( n5424, n5425, n4832 );
or U13117 ( n5425, g3018, n5426 );
nand U13118 ( n4523, n6378, n6379 );
or U13119 ( n6379, n7181, g719 );
nor U13120 ( n6378, n6380, n6381 );
nor U13121 ( n6380, g721, n7180 );
nor U13122 ( n6381, g720, n7170 );
nor U13123 ( n6368, g711, n7170 );
nand U13124 ( n6268, n6365, n6366 );
or U13125 ( n6366, n7181, g710 );
nor U13126 ( n6365, n6367, n6368 );
nor U13127 ( n6367, g712, n7180 );
nand U13128 ( new_g25265_, n4175, n4458 );
nand U13129 ( n4458, n4459, n4461 );
nor U13130 ( n4459, n4174, n4462 );
nor U13131 ( n4462, g3080, g2993 );
nor U13132 ( n3126, g2418, n7429 );
nor U13133 ( n3283, g1030, n7453 );
nand U13134 ( n3045, n3124, n3125 );
or U13135 ( n3125, n7426, g2421 );
nor U13136 ( n3124, n3126, n3127 );
nor U13137 ( n3127, g2429, n7432 );
nand U13138 ( n3235, n3281, n3282 );
or U13139 ( n3282, n7450, g1033 );
nor U13140 ( n3281, n3283, n3284 );
nor U13141 ( n3284, g1041, n7456 );
or U13142 ( n6978, n7373, n7374 );
nor U13143 ( n7373, n7178, g2811 );
nor U13144 ( n7374, n7172, g2813 );
or U13145 ( n6778, n7375, n7376 );
nor U13146 ( n7375, n7177, g2117 );
nor U13147 ( n7376, n7173, g2119 );
or U13148 ( n6583, n7377, n7378 );
nor U13149 ( n7377, n7176, g1423 );
nor U13150 ( n7378, n7174, g1425 );
nand U13151 ( n5470, g3139, n639 );
not U13152 ( n639, g3231 );
nand U13153 ( new_g21882_, n5461, n5462 );
nand U13154 ( n5461, g2878, n7244 );
nand U13155 ( n5462, n7384, n5463 );
nand U13156 ( n3940, n6077, n6078 );
nor U13157 ( n6077, g2896, g2892 );
nor U13158 ( n6078, g2900, n6079 );
or U13159 ( n6079, g2903, g2908 );
not U13160 ( n640, g3234 );
nand U13161 ( new_g21878_, n5468, n5469 );
nand U13162 ( n5468, g7519, n7382 );
nand U13163 ( n5469, n5463, n7244 );
nand U13164 ( new_g21880_, n5464, n5466 );
nand U13165 ( n5464, g2877, n7244 );
nand U13166 ( n5466, n5467, n7382 );
nand U13167 ( new_g20874_, n5808, n5809 );
nand U13168 ( n5808, g8096, n7382 );
nand U13169 ( n5809, n5467, n7244 );
nor U13170 ( n3216, g1735, n7444 );
nor U13171 ( n3316, g354, n7468 );
nand U13172 ( n3146, n3213, n3214 );
or U13173 ( n3214, n7438, g1727 );
nor U13174 ( n3213, n3215, n3216 );
nor U13175 ( n3215, g1724, n7441 );
nand U13176 ( n3303, n3313, n3314 );
or U13177 ( n3314, n7462, g346 );
nor U13178 ( n3313, n3315, n3316 );
nor U13179 ( n3315, g343, n7465 );
nor U13180 ( n3394, g2253, n7435 );
nor U13181 ( n3469, g865, n7459 );
nor U13182 ( new_g26031_, n4178, n621 );
xor U13183 ( n4178, n3517, g3010 );
nor U13184 ( new_g24445_, n4833, n621 );
xor U13185 ( n4833, n622, g3002 );
nor U13186 ( n3431, g1559, n7447 );
nor U13187 ( n3502, g177, n7471 );
or U13188 ( n6388, n7379, n7380 );
nor U13189 ( n7379, n7181, g737 );
nor U13190 ( n7380, n7180, g739 );
nand U13191 ( n2638, n2692, n2693 );
nand U13192 ( n2693, g368, g337 );
and U13193 ( n2692, n2694, n2695 );
nand U13194 ( n2694, g5629, g364 );
nand U13195 ( n2534, n2588, n2589 );
nand U13196 ( n2589, g1055, g1024 );
and U13197 ( n2588, n2590, n2591 );
nand U13198 ( n2590, g5657, g1051 );
nand U13199 ( n2423, n2478, n2479 );
nand U13200 ( n2479, g1749, g1718 );
and U13201 ( n2478, n2481, n2482 );
nand U13202 ( n2481, g5695, g1745 );
nand U13203 ( n2695, g5648, g366 );
nand U13204 ( n2591, g5686, g1053 );
nand U13205 ( n2482, g5738, g1747 );
nand U13206 ( n4403, n6940, n6941 );
or U13207 ( n6941, n7178, g2778 );
nor U13208 ( n6940, n6942, n6943 );
nor U13209 ( n6942, g2780, n7172 );
nand U13210 ( n4446, n6740, n6741 );
or U13211 ( n6741, n7177, g2084 );
nor U13212 ( n6740, n6742, n6743 );
nor U13213 ( n6742, g2086, n7173 );
nand U13214 ( n4495, n6545, n6546 );
or U13215 ( n6546, n7176, g1390 );
nor U13216 ( n6545, n6547, n6548 );
nor U13217 ( n6547, g1392, n7174 );
nor U13218 ( n6943, g2779, n7163 );
nor U13219 ( n6743, g2085, n7164 );
nor U13220 ( n6548, g1391, n7165 );
nand U13221 ( n4406, n6927, n6928 );
or U13222 ( n6928, n7178, g2805 );
nor U13223 ( n6927, n6929, n6930 );
nor U13224 ( n6929, g2807, n7172 );
nand U13225 ( n4449, n6727, n6728 );
or U13226 ( n6728, n7177, g2111 );
nor U13227 ( n6727, n6729, n6730 );
nor U13228 ( n6729, g2113, n7173 );
nand U13229 ( n4498, n6532, n6533 );
or U13230 ( n6533, n7176, g1417 );
nor U13231 ( n6532, n6534, n6535 );
nor U13232 ( n6534, g1419, n7174 );
nor U13233 ( n6930, g2806, n7163 );
nor U13234 ( n6730, g2112, n7164 );
nor U13235 ( n6535, g1418, n7165 );
nand U13236 ( n4534, n6350, n6351 );
or U13237 ( n6351, n7181, g704 );
nor U13238 ( n6350, n6352, n6353 );
nor U13239 ( n6352, g706, n7180 );
nor U13240 ( n6353, g705, n7170 );
nor U13241 ( n3134, g2448, n7430 );
nand U13242 ( n2919, n3132, n3133 );
or U13243 ( n3133, n7426, g2451 );
nor U13244 ( n3132, n3134, n3135 );
nor U13245 ( n3135, g2459, n7433 );
nand U13246 ( n4537, n6337, n6338 );
or U13247 ( n6338, n7181, g731 );
nor U13248 ( n6337, n6339, n6340 );
nor U13249 ( n6339, g733, n7180 );
nor U13250 ( n6340, g732, n7170 );
nand U13251 ( n3006, n3221, n3222 );
or U13252 ( n3222, n7438, g1757 );
nor U13253 ( n3221, n3223, n3224 );
nor U13254 ( n3224, g1765, n7444 );
nor U13255 ( n3223, g1754, n7442 );
nor U13256 ( n3291, g1060, n7453 );
nand U13257 ( n3094, n3289, n3290 );
or U13258 ( n3290, n7450, g1063 );
nor U13259 ( n3289, n3291, n3292 );
nor U13260 ( n3292, g1071, n7456 );
nand U13261 ( n3198, n3321, n3322 );
or U13262 ( n3322, n7462, g376 );
nor U13263 ( n3321, n3323, n3324 );
nor U13264 ( n3323, g373, n7465 );
nor U13265 ( n3324, g384, n7468 );
nand U13266 ( g16496, g2987, n6113 );
nand U13267 ( n6113, g5388, n7123 );
nand U13268 ( n2686, g396, g5648 );
nand U13269 ( n2582, g1083, g5686 );
nand U13270 ( n2471, g1777, g5738 );
nand U13271 ( n2668, n2683, n2684 );
nand U13272 ( n2684, g324, g337 );
and U13273 ( n2683, n2685, n2686 );
nand U13274 ( n2685, g394, g5629 );
nand U13275 ( n2564, n2579, n2580 );
nand U13276 ( n2580, g1011, g1024 );
and U13277 ( n2579, n2581, n2582 );
nand U13278 ( n2581, g1081, g5657 );
nand U13279 ( n2453, n2468, n2469 );
nand U13280 ( n2469, g1705, g1718 );
and U13281 ( n2468, n2470, n2471 );
nand U13282 ( n2470, g1775, g5695 );
nand U13283 ( n2310, n2364, n2365 );
nand U13284 ( n2365, g2443, g2412 );
and U13285 ( n2364, n2366, n2367 );
nand U13286 ( n2366, g5747, g2439 );
nand U13287 ( n2367, g5796, g2441 );
nand U13288 ( new_g24226_, n4866, n4867 );
nand U13289 ( n4866, g2553, n7262 );
nand U13290 ( n4867, g8167, n528 );
nand U13291 ( new_g24214_, n4882, n4884 );
nand U13292 ( n4882, g2552, n7263 );
nand U13293 ( n4884, g8087, n528 );
nand U13294 ( new_g24213_, n4886, n4888 );
nand U13295 ( n4886, g1165, n7264 );
nand U13296 ( n4888, g8007, n308 );
nand U13297 ( new_g24181_, n4904, n4905 );
nand U13298 ( n4904, g1164, n7265 );
nand U13299 ( n4905, g7961, n308 );
nand U13300 ( new_g24238_, n4854, n4855 );
nand U13301 ( n4854, g2554, n7271 );
nand U13302 ( n4855, g2560, n528 );
nand U13303 ( new_g24223_, n4870, n4871 );
nand U13304 ( n4870, g1166, n7270 );
nand U13305 ( n4871, g1172, n308 );
nand U13306 ( new_g24207_, n4897, n4898 );
nand U13307 ( n4897, g478, n7268 );
nand U13308 ( n4898, g7956, n187 );
nand U13309 ( new_g24178_, n4909, n4910 );
nand U13310 ( n4909, g477, n7269 );
nand U13311 ( n4910, g7909, n187 );
nand U13312 ( new_g24216_, n4878, n4879 );
nand U13313 ( n4878, g479, n7273 );
nand U13314 ( n4879, g485, n187 );
nand U13315 ( new_g24219_, n4874, n4875 );
nand U13316 ( n4874, g1859, n7266 );
nand U13317 ( n4875, g8082, n417 );
nand U13318 ( new_g24208_, n4893, n4894 );
nand U13319 ( n4893, g1858, n7267 );
nand U13320 ( n4894, g8012, n417 );
nand U13321 ( new_g24231_, n4860, n4861 );
nand U13322 ( n4860, g1860, n7272 );
nand U13323 ( n4861, g1866, n417 );
nand U13324 ( n2358, g2471, g5796 );
nand U13325 ( n2340, n2355, n2356 );
nand U13326 ( n2356, g2399, g2412 );
and U13327 ( n2355, n2357, n2358 );
nand U13328 ( n2357, g2469, g5747 );
nor U13329 ( new_g28637_, n29, n2239 );
xor U13330 ( n2239, g2133, n2029 );
nor U13331 ( new_g28636_, n27, n2240 );
xor U13332 ( n2240, g1439, n2035 );
nor U13333 ( new_g28635_, n25, n2241 );
xor U13334 ( n2241, g753, n2041 );
nor U13335 ( new_g28634_, n23, n2242 );
xor U13336 ( n2242, g65, n2047 );
nand U13337 ( new_g23418_, n4922, n4923 );
nand U13338 ( n4922, g2533, n7262 );
nand U13339 ( n4923, n527, g8167 );
nand U13340 ( new_g23407_, n4926, n4927 );
nand U13341 ( n4926, g2530, n7263 );
nand U13342 ( n4927, n527, g8087 );
nand U13343 ( new_g23406_, n4941, n4942 );
nand U13344 ( n4941, g1145, n7264 );
nand U13345 ( n4942, n307, g8007 );
nand U13346 ( new_g23392_, n4960, n4961 );
nand U13347 ( n4960, g1142, n7265 );
nand U13348 ( n4961, n307, g7961 );
nand U13349 ( new_g24209_, n4891, n4892 );
nand U13350 ( n4891, g2536, n7271 );
nand U13351 ( n4892, n527, g2560 );
nand U13352 ( new_g24179_, n4907, n4908 );
nand U13353 ( n4907, g1148, n7270 );
nand U13354 ( n4908, n307, g1172 );
nand U13355 ( new_g23413_, n4924, n4925 );
nand U13356 ( n4924, g1839, n7266 );
nand U13357 ( n4925, n416, g8082 );
nand U13358 ( new_g23400_, n4943, n4944 );
nand U13359 ( n4943, g1836, n7267 );
nand U13360 ( n4944, n416, g8012 );
nand U13361 ( new_g24182_, n4902, n4903 );
nand U13362 ( n4902, g1842, n7272 );
nand U13363 ( n4903, n416, g1866 );
nand U13364 ( new_g23399_, n4958, n4959 );
nand U13365 ( n4958, g458, n7268 );
nand U13366 ( n4959, n186, g7956 );
nand U13367 ( new_g23385_, n4975, n4976 );
nand U13368 ( n4975, g455, n7269 );
nand U13369 ( n4976, n186, g7909 );
nand U13370 ( new_g24174_, n4912, n4913 );
nand U13371 ( n4912, g461, n7273 );
nand U13372 ( n4913, n186, g485 );
and U13373 ( n5933, g3136, n639 );
nand U13374 ( new_g24237_, n4856, n4857 );
nand U13375 ( n4856, g2543, n7262 );
nand U13376 ( n4857, g8167, n3887 );
nand U13377 ( new_g24225_, n4868, n4869 );
nand U13378 ( n4868, g2540, n7263 );
nand U13379 ( n4869, g8087, n3887 );
nand U13380 ( new_g24230_, n4862, n4863 );
nand U13381 ( n4862, g1849, n7266 );
nand U13382 ( n4863, g8082, n3963 );
nand U13383 ( new_g24218_, n4876, n4877 );
nand U13384 ( n4876, g1846, n7267 );
nand U13385 ( n4877, g8012, n3963 );
nand U13386 ( new_g24222_, n4872, n4873 );
nand U13387 ( n4872, g1155, n7264 );
nand U13388 ( n4873, g8007, n4033 );
nand U13389 ( new_g24212_, n4889, n4890 );
nand U13390 ( n4889, g1152, n7265 );
nand U13391 ( n4890, g7961, n4033 );
nand U13392 ( new_g24215_, n4880, n4881 );
nand U13393 ( n4880, g468, n7268 );
nand U13394 ( n4881, g7956, n4103 );
nand U13395 ( new_g24206_, n4899, n4901 );
nand U13396 ( n4899, g465, n7269 );
nand U13397 ( n4901, g7909, n4103 );
nand U13398 ( new_g24250_, n4850, n4851 );
nand U13399 ( n4850, g2546, n7271 );
nand U13400 ( n4851, g2560, n3887 );
nand U13401 ( new_g24243_, n4852, n4853 );
nand U13402 ( n4852, g1852, n7272 );
nand U13403 ( n4853, g1866, n3963 );
nand U13404 ( new_g24235_, n4858, n4859 );
nand U13405 ( n4858, g1158, n7270 );
nand U13406 ( n4859, g1172, n4033 );
nand U13407 ( new_g24228_, n4864, n4865 );
nand U13408 ( n4864, g471, n7273 );
nand U13409 ( n4865, g485, n4103 );
nand U13410 ( n2363, g2456, g5796 );
nand U13411 ( n2328, n2360, n2361 );
nand U13412 ( n2361, g2458, g2412 );
and U13413 ( n2360, n2362, n2363 );
nand U13414 ( n2362, g2454, g5747 );
nand U13415 ( n2691, g381, g5648 );
nand U13416 ( n2587, g1068, g5686 );
nand U13417 ( n2477, g1762, g5738 );
nand U13418 ( n2656, n2688, n2689 );
nand U13419 ( n2689, g383, g337 );
and U13420 ( n2688, n2690, n2691 );
nand U13421 ( n2690, g379, g5629 );
nand U13422 ( n2552, n2584, n2585 );
nand U13423 ( n2585, g1070, g1024 );
and U13424 ( n2584, n2586, n2587 );
nand U13425 ( n2586, g1066, g5657 );
nand U13426 ( n2441, n2473, n2474 );
nand U13427 ( n2474, g1764, g1718 );
and U13428 ( n2473, n2475, n2477 );
nand U13429 ( n2475, g1760, g5695 );
nand U13430 ( new_g30801_, n641, n642 );
nand U13431 ( n641, g3108, n7245 );
nand U13432 ( n642, g3109, n235 );
nand U13433 ( new_g30796_, n646, n647 );
nand U13434 ( n646, g3106, n7242 );
nand U13435 ( n647, g8106, n235 );
nand U13436 ( new_g30798_, n644, n645 );
nand U13437 ( n644, g3107, n7243 );
nand U13438 ( n645, g8030, n235 );
nand U13439 ( n3177, n3293, n3294 );
or U13440 ( n3294, n7450, g1078 );
nor U13441 ( n3293, n3295, n3296 );
nor U13442 ( n3296, g1085, n7457 );
nor U13443 ( n3138, g2463, n7430 );
nor U13444 ( n3295, g1075, n7454 );
nand U13445 ( n2988, n3136, n3137 );
or U13446 ( n3137, n7426, g2466 );
nor U13447 ( n3136, n3138, n3139 );
nor U13448 ( n3139, g2473, n7433 );
nor U13449 ( new_g28147_, n2715, n2716 );
nor U13450 ( n2715, g1444, n2717 );
nand U13451 ( n2716, n2035, n2033 );
nor U13452 ( new_g28146_, n2719, n2720 );
nor U13453 ( n2719, g758, n2721 );
nand U13454 ( n2720, n2041, n2039 );
nor U13455 ( new_g28145_, n2723, n2724 );
nor U13456 ( n2723, g70, n2725 );
nand U13457 ( n2724, n2047, n2044 );
nand U13458 ( n3076, n3225, n3226 );
or U13459 ( n3226, n7438, g1772 );
nor U13460 ( n3225, n3227, n3228 );
nor U13461 ( n3228, g1779, n7445 );
nor U13462 ( new_g28148_, n2711, n2712 );
nor U13463 ( n2711, g2138, n2713 );
nand U13464 ( n2712, n2029, n2027 );
nor U13465 ( n3227, g1769, n7442 );
xor U13466 ( n3905, g2160, n498 );
xor U13467 ( n3978, g1466, n390 );
xor U13468 ( n4048, g780, n281 );
xor U13469 ( n4119, g92, n160 );
nand U13470 ( n3266, n3325, n3326 );
or U13471 ( n3326, n7462, g391 );
nor U13472 ( n3325, n3327, n3328 );
nor U13473 ( n3328, g398, n7469 );
xor U13474 ( n3921, g2156, n502 );
xor U13475 ( n3993, g1462, n394 );
xor U13476 ( n4063, g776, n285 );
xor U13477 ( n4134, g88, n164 );
nor U13478 ( n3327, g388, n7466 );
nor U13479 ( n3900, n3902, n3903 );
xor U13480 ( n3902, n7189, n501 );
nand U13481 ( n3903, n3904, n3905 );
xor U13482 ( n3904, g2120, n500 );
nor U13483 ( n3974, n3975, n3976 );
xor U13484 ( n3975, n7190, n393 );
nand U13485 ( n3976, n3977, n3978 );
xor U13486 ( n3977, g1426, n392 );
nor U13487 ( n4044, n4045, n4046 );
xor U13488 ( n4045, n7191, n284 );
nand U13489 ( n4046, n4047, n4048 );
xor U13490 ( n4047, g740, n283 );
nor U13491 ( n4114, n4115, n4116 );
xor U13492 ( n4115, n7192, n163 );
nand U13493 ( n4116, n4117, n4119 );
xor U13494 ( n4117, g52, n162 );
nor U13495 ( n3899, n3919, n3920 );
xor U13496 ( n3919, g2147, n900 );
nand U13497 ( n3920, n3921, n3922 );
xor U13498 ( n3922, n7210, n1211 );
nor U13499 ( n3973, n3991, n3992 );
xor U13500 ( n3991, g1453, n947 );
nand U13501 ( n3992, n3993, n3994 );
xor U13502 ( n3994, n7211, n1231 );
nor U13503 ( n4043, n4061, n4062 );
xor U13504 ( n4061, g767, n991 );
nand U13505 ( n4062, n4063, n4064 );
xor U13506 ( n4064, n7212, n1262 );
nor U13507 ( n4113, n4132, n4133 );
xor U13508 ( n4132, g79, n1032 );
nand U13509 ( n4133, n4134, n4135 );
xor U13510 ( n4135, n7213, n1302 );
nor U13511 ( n3370, g2524, n7430 );
nor U13512 ( n3445, g1136, n7454 );
nand U13513 ( n2743, n3368, n3369 );
or U13514 ( n3369, n7426, g2522 );
nor U13515 ( n3368, n3370, n3371 );
nor U13516 ( n3371, g2523, n7433 );
nand U13517 ( n2787, n3443, n3444 );
or U13518 ( n3444, n7450, g1134 );
nor U13519 ( n3443, n3445, n3446 );
nor U13520 ( n3446, g1135, n7457 );
nor U13521 ( n3407, g1830, n7442 );
nand U13522 ( n2766, n3405, n3406 );
or U13523 ( n3406, n7438, g1828 );
nor U13524 ( n3405, n3407, n3408 );
nor U13525 ( n3408, g1829, n7445 );
nor U13526 ( n3484, g449, n7466 );
nand U13527 ( n2803, n3481, n3482 );
or U13528 ( n3482, n7462, g447 );
nor U13529 ( n3481, n3484, n3485 );
nor U13530 ( n3485, g448, n7469 );
and U13531 ( new_g20884_, g3054, n640 );
nand U13532 ( n2830, g672, n3739 );
nand U13533 ( n3740, g646, n4848 );
nand U13534 ( n2825, g1358, n3635 );
nand U13535 ( n3636, g1332, n4844 );
nand U13536 ( n2820, g2052, n3537 );
nand U13537 ( n3538, g2026, n4840 );
nand U13538 ( n3335, g2746, n3522 );
nand U13539 ( n3523, g2720, n4836 );
nand U13540 ( n2238, g679, n2829 );
nand U13541 ( n2709, g1365, n2824 );
nand U13542 ( n2706, g2059, n2819 );
nand U13543 ( n2703, g2753, n3334 );
nand U13544 ( n4849, g633, n5007 );
nand U13545 ( n4845, g1319, n5459 );
nand U13546 ( n4841, g2013, n5448 );
nand U13547 ( n4837, g2707, n5443 );
nor U13548 ( n5008, n7181, g659 );
nor U13549 ( n5460, n7176, g1345 );
nor U13550 ( n5449, n7177, g2039 );
nor U13551 ( n5444, n7178, g2733 );
and U13552 ( n5007, g640, n5008 );
and U13553 ( n5459, g1326, n5460 );
and U13554 ( n5448, g2020, n5449 );
and U13555 ( n5443, g2714, n5444 );
nand U13556 ( n3946, n3947, n3948 );
xor U13557 ( n3947, g2138, n507 );
xor U13558 ( n3948, g2124, n506 );
nand U13559 ( n4016, n4017, n4018 );
xor U13560 ( n4017, g1444, n399 );
xor U13561 ( n4018, g1430, n398 );
nand U13562 ( n4086, n4087, n4088 );
xor U13563 ( n4087, g758, n290 );
xor U13564 ( n4088, g744, n289 );
nand U13565 ( n4157, n4158, n4159 );
xor U13566 ( n4158, g70, n169 );
xor U13567 ( n4159, g56, n168 );
or U13568 ( new_g20497_, g3079, g3234 );
or U13569 ( new_g19152_, g2933, g51 );
nor U13570 ( new_g16823_, n7295, g51 );
nor U13571 ( new_g20877_, g3234, n7187 );
nor U13572 ( new_g16802_, g51, n7253 );
nor U13573 ( new_g27621_, n29, n2831 );
xor U13574 ( n2831, g2142, n2714 );
nor U13575 ( new_g27612_, n27, n2832 );
xor U13576 ( n2832, g1448, n2718 );
nor U13577 ( new_g27603_, n25, n2833 );
xor U13578 ( n2833, g762, n2722 );
nor U13579 ( new_g27594_, n23, n2834 );
xor U13580 ( n2834, g74, n2726 );
nand U13581 ( new_g18975_, n5867, n5868 );
nand U13582 ( n5867, n7384, g2981 );
nand U13583 ( n5868, g2195, n7244 );
nand U13584 ( new_g18781_, n5911, n5912 );
nand U13585 ( n5911, g2956, n7384 );
nand U13586 ( n5912, g1501, n7498 );
nand U13587 ( new_g18968_, n5869, n5870 );
nand U13588 ( n5869, n7384, g2978 );
nand U13589 ( n5870, g2190, n7244 );
nand U13590 ( new_g18803_, n5905, n5906 );
nand U13591 ( n5905, g2953, n7383 );
nand U13592 ( n5906, g1496, n7498 );
buf U13593 ( n7497, g2879 );
nand U13594 ( new_g18942_, n5873, n5874 );
nand U13595 ( n5873, n7384, g2975 );
nand U13596 ( n5874, g2185, n7244 );
nand U13597 ( new_g20417_, n5824, n5825 );
nand U13598 ( n5824, g7334, n7382 );
nand U13599 ( n5825, g2963, n7244 );
nand U13600 ( new_g20343_, n5832, n5833 );
nand U13601 ( n5832, g6442, n7382 );
nand U13602 ( n5833, g2969, n7244 );
nand U13603 ( new_g19184_, n5843, n5844 );
nand U13604 ( n5843, g4590, n7382 );
nand U13605 ( n5844, g2975, n7244 );
nand U13606 ( new_g19163_, n5853, n5854 );
nand U13607 ( n5853, g4090, n7382 );
nand U13608 ( n5854, g2981, n7244 );
nand U13609 ( new_g19154_, n5859, n5860 );
nand U13610 ( n5859, g8251, n7383 );
nand U13611 ( n5860, g2874, n7244 );
nand U13612 ( new_g18867_, n5887, n5888 );
nand U13613 ( n5887, n7384, g2969 );
nand U13614 ( n5888, g2175, n7498 );
nand U13615 ( new_g18852_, n5891, n5892 );
nand U13616 ( n5891, g2941, n7383 );
nand U13617 ( n5892, g1481, n7498 );
nand U13618 ( new_g18821_, n5899, n5900 );
nand U13619 ( n5899, g2947, n7384 );
nand U13620 ( n5900, g1491, n7498 );
nand U13621 ( new_g18836_, n5895, n5896 );
nand U13622 ( n5895, n7384, g2966 );
nand U13623 ( n5896, g2170, n7498 );
nand U13624 ( new_g18906_, n5877, n5879 );
nand U13625 ( n5877, n7384, g2972 );
nand U13626 ( n5879, g2180, n7498 );
nand U13627 ( new_g18885_, n5880, n5881 );
nand U13628 ( n5880, n7384, g2874 );
nand U13629 ( n5881, g2200, n7498 );
nand U13630 ( new_g18866_, n5889, n5890 );
nand U13631 ( n5889, g2938, n7383 );
nand U13632 ( n5890, g1476, n7498 );
nand U13633 ( new_g18835_, n5897, n5898 );
nand U13634 ( n5897, g2944, n7383 );
nand U13635 ( n5898, g1486, n7498 );
nand U13636 ( new_g18754_, n5919, n5920 );
nand U13637 ( n5919, g2959, n7384 );
nand U13638 ( n5920, g1506, n7498 );
nand U13639 ( new_g18957_, n5871, n5872 );
nand U13640 ( n5871, n7384, g2963 );
nand U13641 ( n5872, g2165, n7244 );
nand U13642 ( new_g18883_, n5883, n5884 );
nand U13643 ( n5883, g2935, n7383 );
nand U13644 ( n5884, g1471, n7498 );
nand U13645 ( new_g19167_, n5851, n5852 );
nand U13646 ( n5851, g4200, n7382 );
nand U13647 ( n5852, g2938, n7244 );
nand U13648 ( new_g20376_, n5826, n5827 );
nand U13649 ( n5826, g6895, n7382 );
nand U13650 ( n5827, g2966, n7244 );
nand U13651 ( new_g20310_, n5841, n5842 );
nand U13652 ( n5841, g6225, n7382 );
nand U13653 ( n5842, g2972, n7244 );
nand U13654 ( new_g19173_, n5847, n5848 );
nand U13655 ( n5847, g4323, n7383 );
nand U13656 ( n5848, g2978, n7244 );
nand U13657 ( new_g19157_, n5857, n5858 );
nand U13658 ( n5857, g3993, n7383 );
nand U13659 ( n5858, g2941, n7244 );
nand U13660 ( new_g19149_, n5863, n5864 );
nand U13661 ( n5863, g8175, n7383 );
nand U13662 ( n5864, g2944, n7244 );
nand U13663 ( new_g19144_, n5865, n5866 );
nand U13664 ( n5865, g8023, n7383 );
nand U13665 ( n5866, g2947, n7244 );
nand U13666 ( new_g19172_, n5849, n5850 );
nand U13667 ( n5849, g4321, n7382 );
nand U13668 ( n5850, g2953, n7244 );
nand U13669 ( new_g19162_, n5855, n5856 );
nand U13670 ( n5855, g4088, n7383 );
nand U13671 ( n5856, g2956, n7244 );
nand U13672 ( new_g19153_, n5861, n5862 );
nand U13673 ( n5861, g8249, n7383 );
nand U13674 ( n5862, g2959, n7244 );
nand U13675 ( new_g19178_, n5845, n5846 );
nand U13676 ( n5845, g4450, n7382 );
nand U13677 ( n5846, g2935, n7244 );
nor U13678 ( new_g28199_, n267, n2710 );
xor U13679 ( n2710, n2238, g686 );
nor U13680 ( new_g27718_, n376, n2815 );
xor U13681 ( n2815, n2709, g1372 );
nor U13682 ( new_g27722_, n484, n2814 );
xor U13683 ( n2814, n2706, g2066 );
nor U13684 ( new_g27724_, n603, n2813 );
xor U13685 ( n2813, n2703, g2760 );
nor U13686 ( new_g25260_, n4503, n4504 );
nor U13687 ( n4503, g735, n4538 );
nor U13688 ( n4504, n4456, n255 );
nor U13689 ( new_g25262_, n4500, n4501 );
nor U13690 ( n4500, g736, n4502 );
nor U13691 ( n4501, n4456, n256 );
nor U13692 ( new_g25266_, n4454, n4455 );
nor U13693 ( n4454, g734, n4457 );
nor U13694 ( n4455, n4456, n257 );
nor U13695 ( new_g25272_, n4372, n4373 );
nor U13696 ( n4372, g2809, n4407 );
nor U13697 ( n4373, n4363, n590 );
nor U13698 ( new_g25280_, n4365, n4366 );
nor U13699 ( n4365, g2810, n4367 );
nor U13700 ( n4366, n4363, n591 );
nor U13701 ( new_g25288_, n4361, n4362 );
nor U13702 ( n4361, g2808, n4364 );
nor U13703 ( n4362, n4363, n592 );
nor U13704 ( new_g25268_, n4415, n4416 );
nor U13705 ( n4415, g2115, n4450 );
nor U13706 ( n4416, n4370, n472 );
nor U13707 ( new_g25271_, n4408, n4409 );
nor U13708 ( n4408, g2116, n4410 );
nor U13709 ( n4409, n4370, n473 );
nor U13710 ( new_g25279_, n4368, n4369 );
nor U13711 ( n4368, g2114, n4371 );
nor U13712 ( n4369, n4370, n474 );
nor U13713 ( new_g25263_, n4463, n4465 );
nor U13714 ( n4463, g1421, n4499 );
nor U13715 ( n4465, n4413, n364 );
nor U13716 ( new_g25267_, n4451, n4452 );
nor U13717 ( n4451, g1422, n4453 );
nor U13718 ( n4452, n4413, n365 );
nor U13719 ( new_g25270_, n4411, n4412 );
nor U13720 ( n4411, g1420, n4414 );
nor U13721 ( n4412, n4413, n366 );
and U13722 ( n4456, n4505, n4506 );
nor U13723 ( n4505, n4536, n4537 );
nor U13724 ( n4506, n4507, n4508 );
nor U13725 ( n4536, g728, n7181 );
and U13726 ( n4363, n4374, n4375 );
nor U13727 ( n4374, n4405, n4406 );
nor U13728 ( n4375, n4376, n4377 );
nor U13729 ( n4405, g2802, n7178 );
and U13730 ( n4370, n4417, n4418 );
nor U13731 ( n4417, n4448, n4449 );
nor U13732 ( n4418, n4419, n4420 );
nor U13733 ( n4448, g2108, n7177 );
and U13734 ( n4413, n4466, n4467 );
nor U13735 ( n4466, n4497, n4498 );
nor U13736 ( n4467, n4468, n4469 );
nor U13737 ( n4497, g1414, n7176 );
nor U13738 ( n4511, n4525, n4526 );
nand U13739 ( n4526, n4527, n4528 );
nand U13740 ( n4525, n4530, n4531 );
xor U13741 ( n4528, g646, n4529 );
nor U13742 ( n4380, n4394, n4395 );
nand U13743 ( n4395, n4396, n4397 );
nand U13744 ( n4394, n4399, n4400 );
xor U13745 ( n4397, g2720, n4398 );
nor U13746 ( n4423, n4437, n4438 );
nand U13747 ( n4438, n4439, n4440 );
nand U13748 ( n4437, n4442, n4443 );
xor U13749 ( n4440, g2026, n4441 );
nor U13750 ( n4472, n4486, n4487 );
nand U13751 ( n4487, n4488, n4489 );
nand U13752 ( n4486, n4491, n4492 );
xor U13753 ( n4489, g1332, n4490 );
nand U13754 ( n4508, n4509, n4510 );
or U13755 ( n4509, n7180, g730 );
nand U13756 ( n4510, n4511, n4512 );
nor U13757 ( n4512, n4513, n4514 );
nand U13758 ( n4377, n4378, n4379 );
or U13759 ( n4378, n7172, g2804 );
nand U13760 ( n4379, n4380, n4381 );
nor U13761 ( n4381, n4382, n4383 );
nand U13762 ( n4420, n4421, n4422 );
or U13763 ( n4421, n7173, g2110 );
nand U13764 ( n4422, n4423, n4424 );
nor U13765 ( n4424, n4425, n4426 );
nand U13766 ( n4469, n4470, n4471 );
or U13767 ( n4470, n7174, g1416 );
nand U13768 ( n4471, n4472, n4473 );
nor U13769 ( n4473, n4474, n4475 );
nor U13770 ( n4530, n4532, n4533 );
xor U13771 ( n4533, n4534, g653 );
xor U13772 ( n4532, n4535, n7203 );
nor U13773 ( n4399, n4401, n4402 );
xor U13774 ( n4402, n4403, g2727 );
xor U13775 ( n4401, n4404, n7199 );
nor U13776 ( n4442, n4444, n4445 );
xor U13777 ( n4445, n4446, g2033 );
xor U13778 ( n4444, n4447, n7200 );
nor U13779 ( n4491, n4493, n4494 );
xor U13780 ( n4494, n4495, g1339 );
xor U13781 ( n4493, n4496, n7201 );
nand U13782 ( n5088, n6480, n6481 );
nand U13783 ( n6481, g1297, g1236 );
nor U13784 ( n6480, n6482, n6483 );
and U13785 ( n6482, g6944, g1294 );
and U13786 ( n6483, g6750, g1291 );
nand U13787 ( n5070, n6870, n6871 );
nand U13788 ( n6871, g2685, g2624 );
nor U13789 ( n6870, n6872, n6873 );
and U13790 ( n6873, g7302, g2679 );
and U13791 ( n6872, g7390, g2682 );
nand U13792 ( n6314, n6329, n6330 );
nor U13793 ( n6329, n6391, n6392 );
nor U13794 ( n6330, n260, n6331 );
nor U13795 ( n6391, g735, n7170 );
nand U13796 ( n6859, n6896, n6897 );
nor U13797 ( n6896, n6899, n6900 );
nor U13798 ( n6897, n595, n6898 );
nor U13799 ( n6899, g2809, n7163 );
nand U13800 ( n6665, n6698, n6699 );
nor U13801 ( n6698, n6701, n6702 );
nor U13802 ( n6699, n477, n6700 );
nor U13803 ( n6701, g2115, n7164 );
nand U13804 ( n6470, n6503, n6504 );
nor U13805 ( n6503, n6506, n6507 );
nor U13806 ( n6504, n369, n6505 );
nor U13807 ( n6506, g1421, n7165 );
nand U13808 ( n5097, n6323, n6324 );
nand U13809 ( n6324, g611, g550 );
nor U13810 ( n6323, n6325, n6326 );
and U13811 ( n6325, g6642, g608 );
and U13812 ( n6326, g6485, g605 );
xor U13813 ( n4521, n4524, g666 );
xor U13814 ( n4390, n4393, g2740 );
xor U13815 ( n4433, n4436, g2046 );
xor U13816 ( n4482, n4485, g1352 );
nand U13817 ( n4513, n4519, n4520 );
xor U13818 ( n4520, g672, n262 );
nor U13819 ( n4519, n4521, n4522 );
xor U13820 ( n4522, n4523, g679 );
nand U13821 ( n4382, n4388, n4389 );
xor U13822 ( n4389, g2746, n597 );
nor U13823 ( n4388, n4390, n4391 );
xor U13824 ( n4391, n4392, g2753 );
nand U13825 ( n4425, n4431, n4432 );
xor U13826 ( n4432, g2052, n479 );
nor U13827 ( n4431, n4433, n4434 );
xor U13828 ( n4434, n4435, g2059 );
nand U13829 ( n4474, n4480, n4481 );
xor U13830 ( n4481, g1358, n371 );
nor U13831 ( n4480, n4482, n4483 );
xor U13832 ( n4483, n4484, g1365 );
nand U13833 ( n5079, n6675, n6676 );
nand U13834 ( n6676, g1991, g1930 );
nor U13835 ( n6675, n6677, n6678 );
and U13836 ( n6678, g7052, g1985 );
and U13837 ( n6677, g7194, g1988 );
nor U13838 ( new_g27131_, n3336, n3337 );
nor U13839 ( n3336, g2147, n3338 );
nand U13840 ( n3337, n2714, n2027 );
nor U13841 ( new_g27129_, n3340, n3341 );
nor U13842 ( n3340, g1453, n3342 );
nand U13843 ( n3341, n2718, n2033 );
nor U13844 ( new_g27123_, n3344, n3345 );
nor U13845 ( n3344, g767, n3346 );
nand U13846 ( n3345, n2722, n2039 );
nor U13847 ( new_g27120_, n3348, n3349 );
nor U13848 ( n3348, g79, n3350 );
nand U13849 ( n3349, n2726, n2044 );
xor U13850 ( n3938, g2129, n1274 );
xor U13851 ( n4009, g1435, n1320 );
xor U13852 ( n4079, g749, n1356 );
xor U13853 ( n4150, g61, n1390 );
nand U13854 ( n2273, n6918, n6919 );
nand U13855 ( n6919, g2694, g2624 );
nor U13856 ( n6918, n6920, n6921 );
and U13857 ( n6921, g7302, g2688 );
and U13858 ( n6920, g7390, g2691 );
nand U13859 ( n2609, n6277, n6278 );
nand U13860 ( n6278, g620, g550 );
nor U13861 ( n6277, n6279, n6280 );
and U13862 ( n6279, g6642, g617 );
and U13863 ( n6280, g6485, g614 );
nand U13864 ( n2385, n6718, n6719 );
nand U13865 ( n6719, g2000, g1930 );
nor U13866 ( n6718, n6720, n6721 );
and U13867 ( n6721, g7052, g1994 );
and U13868 ( n6720, g7194, g1997 );
nor U13869 ( new_g27672_, n2826, n2827 );
nor U13870 ( n2826, g679, n2829 );
nand U13871 ( n2827, n2238, n2828 );
nor U13872 ( new_g27678_, n2821, n2822 );
nor U13873 ( n2821, g1365, n2824 );
nand U13874 ( n2822, n2709, n2823 );
nor U13875 ( new_g27682_, n2816, n2817 );
nor U13876 ( n2816, g2059, n2819 );
nand U13877 ( n2817, n2706, n2818 );
nor U13878 ( new_g27243_, n3331, n3332 );
nor U13879 ( n3331, g2753, n3334 );
nand U13880 ( n3332, n2703, n3333 );
xor U13881 ( n4531, g640, n263 );
xor U13882 ( n4400, g2714, n599 );
xor U13883 ( n4443, g2020, n480 );
xor U13884 ( n4492, g1326, n372 );
nand U13885 ( n5133, g2257, n7477 );
nand U13886 ( n5121, g2257, n7474 );
nand U13887 ( n5168, g1563, n7483 );
nand U13888 ( n5141, g1563, n7480 );
nand U13889 ( n5214, g869, n7489 );
nand U13890 ( n5176, g869, n7486 );
nand U13891 ( n5258, g181, n7495 );
nand U13892 ( n5221, g181, n7492 );
nor U13893 ( new_g22045_, n5380, n5381 );
nor U13894 ( n5381, n7128, n5133 );
nor U13895 ( n5380, g2218, n515 );
nor U13896 ( new_g22061_, n5355, n5356 );
nor U13897 ( n5356, n7132, n5133 );
nor U13898 ( n5355, g2221, n515 );
nor U13899 ( new_g22078_, n5328, n5329 );
nor U13900 ( n5329, n7092, n5133 );
nor U13901 ( n5328, g2224, n515 );
nor U13902 ( new_g22099_, n5297, n5298 );
nor U13903 ( n5298, n7149, n5133 );
nor U13904 ( n5297, g2227, n515 );
nor U13905 ( new_g22117_, n5261, n5262 );
nor U13906 ( n5262, n7144, n5133 );
nor U13907 ( n5261, g2230, n515 );
nor U13908 ( new_g22140_, n5224, n5225 );
nor U13909 ( n5225, n7142, n5133 );
nor U13910 ( n5224, g2233, n515 );
nor U13911 ( new_g22170_, n5159, n5160 );
nor U13912 ( n5160, n7130, n5133 );
nor U13913 ( n5159, g2206, n515 );
nor U13914 ( new_g22183_, n5131, n5132 );
nor U13915 ( n5132, n7124, n5133 );
nor U13916 ( n5131, g2209, n515 );
nor U13917 ( new_g22060_, n5358, n5359 );
nor U13918 ( n5359, n7128, n5121 );
nor U13919 ( n5358, g2219, n518 );
nor U13920 ( new_g22077_, n5331, n5332 );
nor U13921 ( n5332, n7132, n5121 );
nor U13922 ( n5331, g2222, n518 );
nor U13923 ( new_g22098_, n5299, n5300 );
nor U13924 ( n5300, n7092, n5121 );
nor U13925 ( n5299, g2225, n518 );
nor U13926 ( new_g22116_, n5263, n5264 );
nor U13927 ( n5264, n7149, n5121 );
nor U13928 ( n5263, g2228, n518 );
nor U13929 ( new_g22139_, n5226, n5227 );
nor U13930 ( n5227, n7144, n5121 );
nor U13931 ( n5226, g2231, n518 );
nor U13932 ( new_g22154_, n5189, n5190 );
nor U13933 ( n5190, n7142, n5121 );
nor U13934 ( n5189, g2234, n518 );
nor U13935 ( new_g22182_, n5134, n5135 );
nor U13936 ( n5135, n7130, n5121 );
nor U13937 ( n5134, g2207, n518 );
nor U13938 ( new_g22193_, n5119, n5120 );
nor U13939 ( n5120, n7124, n5121 );
nor U13940 ( n5119, g2210, n518 );
nor U13941 ( new_g22035_, n5401, n5402 );
nor U13942 ( n5402, n7129, n5168 );
nor U13943 ( n5401, g1524, n406 );
nor U13944 ( new_g22044_, n5382, n5383 );
nor U13945 ( n5383, n7133, n5168 );
nor U13946 ( n5382, g1527, n406 );
nor U13947 ( new_g22059_, n5360, n5361 );
nor U13948 ( n5361, n7093, n5168 );
nor U13949 ( n5360, g1530, n406 );
nor U13950 ( new_g22075_, n5335, n5336 );
nor U13951 ( n5336, n7150, n5168 );
nor U13952 ( n5335, g1533, n406 );
nor U13953 ( new_g22092_, n5304, n5305 );
nor U13954 ( n5305, n7145, n5168 );
nor U13955 ( n5304, g1536, n406 );
nor U13956 ( new_g22114_, n5267, n5268 );
nor U13957 ( n5268, n7143, n5168 );
nor U13958 ( n5267, g1539, n406 );
nor U13959 ( new_g22149_, n5205, n5206 );
nor U13960 ( n5206, n7131, n5168 );
nor U13961 ( n5205, g1512, n406 );
nor U13962 ( new_g22167_, n5165, n5167 );
nor U13963 ( n5167, n7125, n5168 );
nor U13964 ( n5165, g1515, n406 );
nor U13965 ( new_g22043_, n5385, n5386 );
nor U13966 ( n5386, n7129, n5141 );
nor U13967 ( n5385, g1525, n408 );
nor U13968 ( new_g22058_, n5362, n5363 );
nor U13969 ( n5363, n7133, n5141 );
nor U13970 ( n5362, g1528, n408 );
nor U13971 ( new_g22074_, n5337, n5338 );
nor U13972 ( n5338, n7093, n5141 );
nor U13973 ( n5337, g1531, n408 );
nor U13974 ( new_g22091_, n5306, n5307 );
nor U13975 ( n5307, n7150, n5141 );
nor U13976 ( n5306, g1534, n408 );
nor U13977 ( new_g22113_, n5269, n5270 );
nor U13978 ( n5270, n7145, n5141 );
nor U13979 ( n5269, g1537, n408 );
nor U13980 ( new_g22131_, n5236, n5237 );
nor U13981 ( n5237, n7143, n5141 );
nor U13982 ( n5236, g1540, n408 );
nor U13983 ( new_g22166_, n5169, n5170 );
nor U13984 ( n5170, n7131, n5141 );
nor U13985 ( n5169, g1513, n408 );
nor U13986 ( new_g22179_, n5138, n5140 );
nor U13987 ( n5140, n7125, n5141 );
nor U13988 ( n5138, g1516, n408 );
nor U13989 ( new_g22029_, n5415, n5416 );
nor U13990 ( n5416, n7134, n5214 );
nor U13991 ( n5415, g830, n297 );
nor U13992 ( new_g22034_, n5403, n5404 );
nor U13993 ( n5404, n7140, n5214 );
nor U13994 ( n5403, g833, n297 );
nor U13995 ( new_g22042_, n5387, n5388 );
nor U13996 ( n5388, n7095, n5214 );
nor U13997 ( n5387, g836, n297 );
nor U13998 ( new_g22056_, n5367, n5368 );
nor U13999 ( n5368, n7153, n5214 );
nor U14000 ( n5367, g839, n297 );
nor U14001 ( new_g22068_, n5342, n5343 );
nor U14002 ( n5343, n7151, n5214 );
nor U14003 ( n5342, g842, n297 );
nor U14004 ( new_g22089_, n5310, n5311 );
nor U14005 ( n5311, n7146, n5214 );
nor U14006 ( n5310, g845, n297 );
nor U14007 ( new_g22126_, n5250, n5251 );
nor U14008 ( n5251, n7137, n5214 );
nor U14009 ( n5250, g818, n297 );
nor U14010 ( new_g22146_, n5212, n5213 );
nor U14011 ( n5213, n7126, n5214 );
nor U14012 ( n5212, g821, n297 );
nor U14013 ( new_g22033_, n5405, n5407 );
nor U14014 ( n5407, n7134, n5176 );
nor U14015 ( n5405, g831, n299 );
nor U14016 ( new_g22041_, n5389, n5390 );
nor U14017 ( n5390, n7140, n5176 );
nor U14018 ( n5389, g834, n299 );
nor U14019 ( new_g22055_, n5369, n5370 );
nor U14020 ( n5370, n7095, n5176 );
nor U14021 ( n5369, g837, n299 );
nor U14022 ( new_g22067_, n5344, n5345 );
nor U14023 ( n5345, n7153, n5176 );
nor U14024 ( n5344, g840, n299 );
nor U14025 ( new_g22088_, n5313, n5314 );
nor U14026 ( n5314, n7151, n5176 );
nor U14027 ( n5313, g843, n299 );
nor U14028 ( new_g22105_, n5279, n5280 );
nor U14029 ( n5280, n7146, n5176 );
nor U14030 ( n5279, g846, n299 );
nor U14031 ( new_g22145_, n5215, n5216 );
nor U14032 ( n5216, n7137, n5176 );
nor U14033 ( n5215, g819, n299 );
nor U14034 ( new_g22163_, n5173, n5174 );
nor U14035 ( n5174, n7126, n5176 );
nor U14036 ( n5173, g822, n299 );
nor U14037 ( new_g22025_, n5422, n5423 );
nor U14038 ( n5423, n7136, n5258 );
nor U14039 ( n5422, g142, n176 );
nor U14040 ( new_g22028_, n5417, n5418 );
nor U14041 ( n5418, n7141, n5258 );
nor U14042 ( n5417, g145, n176 );
nor U14043 ( new_g22032_, n5408, n5409 );
nor U14044 ( n5409, n7096, n5258 );
nor U14045 ( n5408, g148, n176 );
nor U14046 ( new_g22039_, n5394, n5395 );
nor U14047 ( n5395, n7154, n5258 );
nor U14048 ( n5394, g151, n176 );
nor U14049 ( new_g22049_, n5373, n5374 );
nor U14050 ( n5374, n7152, n5258 );
nor U14051 ( n5373, g154, n176 );
nor U14052 ( new_g22065_, n5349, n5350 );
nor U14053 ( n5350, n7147, n5258 );
nor U14054 ( n5349, g157, n176 );
nor U14055 ( new_g22100_, n5295, n5296 );
nor U14056 ( n5296, n7138, n5258 );
nor U14057 ( n5295, g130, n176 );
nor U14058 ( new_g22123_, n5256, n5257 );
nor U14059 ( n5257, n7127, n5258 );
nor U14060 ( n5256, g133, n176 );
nor U14061 ( new_g22027_, n5419, n5420 );
nor U14062 ( n5420, n7136, n5221 );
nor U14063 ( n5419, g143, n178 );
nor U14064 ( new_g22031_, n5411, n5412 );
nor U14065 ( n5412, n7141, n5221 );
nor U14066 ( n5411, g146, n178 );
nor U14067 ( new_g22038_, n5396, n5398 );
nor U14068 ( n5398, n7096, n5221 );
nor U14069 ( n5396, g149, n178 );
nor U14070 ( new_g22048_, n5376, n5377 );
nor U14071 ( n5377, n7154, n5221 );
nor U14072 ( n5376, g152, n178 );
nor U14073 ( new_g22064_, n5351, n5352 );
nor U14074 ( n5352, n7152, n5221 );
nor U14075 ( n5351, g155, n178 );
nor U14076 ( new_g22080_, n5324, n5325 );
nor U14077 ( n5325, n7147, n5221 );
nor U14078 ( n5324, g158, n178 );
nor U14079 ( new_g22122_, n5259, n5260 );
nor U14080 ( n5260, n7138, n5221 );
nor U14081 ( n5259, g131, n178 );
nor U14082 ( new_g22142_, n5219, n5220 );
nor U14083 ( n5220, n7127, n5221 );
nor U14084 ( n5219, g134, n178 );
nand U14085 ( n2500, n6523, n6524 );
nand U14086 ( n6524, g1306, g1236 );
nor U14087 ( n6523, n6525, n6526 );
and U14088 ( n6525, g6944, g1303 );
and U14089 ( n6526, g6750, g1300 );
xor U14090 ( n4527, g660, n264 );
xor U14091 ( n4396, g2734, n600 );
xor U14092 ( n4439, g2040, n481 );
xor U14093 ( n4488, g1346, n373 );
nand U14094 ( n4514, n4515, n4516 );
xor U14095 ( n4515, g692, n4518 );
xor U14096 ( n4516, g686, n4517 );
nand U14097 ( n4383, n4384, n4385 );
xor U14098 ( n4384, g2766, n4387 );
xor U14099 ( n4385, g2760, n4386 );
nand U14100 ( n4426, n4427, n4428 );
xor U14101 ( n4427, g2072, n4430 );
xor U14102 ( n4428, g2066, n4429 );
nand U14103 ( n4475, n4476, n4477 );
xor U14104 ( n4476, g1378, n4479 );
xor U14105 ( n4477, g1372, n4478 );
nor U14106 ( n3876, g1192, n3878 );
nor U14107 ( n3878, n3879, n7159 );
nor U14108 ( n2050, g1886, n2052 );
nor U14109 ( n2052, n2053, n7158 );
nand U14110 ( n1586, n1587, n7274 );
nand U14111 ( n1587, g7390, new_g28990_ );
nand U14112 ( n3879, n5490, n5491 );
or U14113 ( n5490, g507, n7188 );
nand U14114 ( n5491, n5493, n7188 );
nand U14115 ( n2053, n3874, n3875 );
nand U14116 ( n3874, n7229, g1192 );
nand U14117 ( n3875, n3876, n3877 );
nor U14118 ( n5493, g16297, g6642 );
and U14119 ( new_g28990_, n2048, n2049 );
nand U14120 ( n2048, n7248, g1886 );
nand U14121 ( n2049, n2050, n2051 );
nor U14122 ( new_g30061_, n1583, n1584 );
nor U14123 ( n1584, g2581, n7274 );
nor U14124 ( n1583, n1585, n1586 );
and U14125 ( n1585, g16437, n7161 );
nand U14126 ( new_g29936_, n1597, n1598 );
nand U14127 ( n1597, g3103, n7242 );
nand U14128 ( n1598, g8106, n238 );
nand U14129 ( new_g29939_, n1595, n1596 );
nand U14130 ( n1595, g3104, n7243 );
nand U14131 ( n1596, g8030, n238 );
nand U14132 ( new_g29941_, n1593, n1594 );
nand U14133 ( n1593, g3105, n7245 );
nand U14134 ( n1594, g3109, n238 );
nand U14135 ( n3395, n4553, n4554 );
nor U14136 ( n4553, n4557, n4558 );
nor U14137 ( n4554, n4555, n4556 );
nand U14138 ( n4557, g2175, g2180 );
nand U14139 ( n3432, n4581, n4582 );
nor U14140 ( n4581, n4585, n4586 );
nor U14141 ( n4582, n4583, n4584 );
nand U14142 ( n4585, g1481, g1486 );
nand U14143 ( n4556, g2185, g2190 );
nand U14144 ( n4584, g1491, g1496 );
nand U14145 ( n4555, g2195, g2200 );
nand U14146 ( n4583, g1501, g1506 );
nor U14147 ( new_g26532_, n29, n3870 );
xor U14148 ( n3870, n3339, g2151 );
nor U14149 ( new_g26531_, n27, n3871 );
xor U14150 ( n3871, n3343, g1457 );
nor U14151 ( new_g26530_, n25, n3872 );
xor U14152 ( n3872, n3347, g771 );
nor U14153 ( new_g26529_, n23, n3873 );
xor U14154 ( n3873, n3351, g83 );
and U14155 ( n2628, n2697, n2698 );
nand U14156 ( n2698, g353, g337 );
and U14157 ( n2697, n2699, n2700 );
nand U14158 ( n2699, g349, g5629 );
and U14159 ( n2524, n2593, n2594 );
nand U14160 ( n2594, g1040, g1024 );
and U14161 ( n2593, n2595, n2596 );
nand U14162 ( n2595, g1036, g5657 );
and U14163 ( n2412, n2484, n2485 );
nand U14164 ( n2485, g1734, g1718 );
and U14165 ( n2484, n2486, n2487 );
nand U14166 ( n2486, g1730, g5695 );
nand U14167 ( n2700, g351, g5648 );
nand U14168 ( n2596, g1038, g5686 );
nand U14169 ( n2487, g1732, g5738 );
nand U14170 ( n3470, n4613, n4614 );
nor U14171 ( n4613, n4617, n4618 );
nor U14172 ( n4614, n4615, n4616 );
nand U14173 ( n4617, g793, g797 );
nand U14174 ( n3503, n4646, n4647 );
nor U14175 ( n4646, n4650, n4651 );
nor U14176 ( n4647, n4648, n4649 );
nand U14177 ( n4650, g105, g109 );
nand U14178 ( n4616, g801, g805 );
nand U14179 ( n4649, g113, g117 );
nand U14180 ( n4615, g809, g813 );
nand U14181 ( n4648, g121, g125 );
nand U14182 ( n2956, g6642, new_g22578_ );
nand U14183 ( n3031, g6485, new_g22578_ );
nand U14184 ( new_g22578_, n5093, n5094 );
nand U14185 ( n5093, n5096, n5069 );
nand U14186 ( n5094, n5095, g510 );
nand U14187 ( n5096, n5097, n3868 );
nand U14188 ( n2907, g550, new_g22578_ );
and U14189 ( n2300, n2369, n2370 );
nand U14190 ( n2370, g2428, g2412 );
and U14191 ( n2369, n2371, n2372 );
nand U14192 ( n2371, g2424, g5747 );
nand U14193 ( n2372, g2426, g5796 );
nand U14194 ( n4558, g2165, g2170 );
nand U14195 ( n4586, g1471, g1476 );
nand U14196 ( n2944, g6750, new_g22615_ );
nand U14197 ( new_g22615_, n5084, n5085 );
nand U14198 ( n5084, n5087, n5069 );
nand U14199 ( n5085, n5086, g1196 );
nand U14200 ( n5087, n5088, n3862 );
nand U14201 ( n2869, g1236, new_g22615_ );
nand U14202 ( n2901, g6944, new_g22615_ );
nand U14203 ( n2841, g7390, new_g22687_ );
nand U14204 ( new_g22687_, n5065, n5066 );
nand U14205 ( n5065, n5068, n5069 );
nand U14206 ( n5066, n5067, g2584 );
nand U14207 ( n5068, n5070, n3844 );
nand U14208 ( n2837, g2624, new_g22687_ );
nand U14209 ( n2851, g7302, new_g22687_ );
and U14210 ( new_g13110_, n6072, n6073 );
nor U14211 ( n6073, n6074, n6075 );
nor U14212 ( n6072, n7218, n6076 );
or U14213 ( n6074, g2917, g2920 );
nand U14214 ( n6076, g2883, n43 );
nor U14215 ( new_g25259_, n4539, n4540 );
nor U14216 ( n4540, n3395, n4541 );
nor U14217 ( n4539, g2253, n10 );
nor U14218 ( new_g25257_, n4542, n4543 );
nor U14219 ( n4543, n3395, n4544 );
nor U14220 ( n4542, g2255, n11 );
nor U14221 ( new_g25253_, n4550, n4551 );
nor U14222 ( n4551, n3395, n4552 );
nor U14223 ( n4550, g2254, n13 );
nor U14224 ( new_g25256_, n4545, n4546 );
nor U14225 ( n4546, n7130, n4541 );
nor U14226 ( n4545, g2250, n10 );
nor U14227 ( new_g25252_, n4559, n4560 );
nor U14228 ( n4560, n7130, n4544 );
nor U14229 ( n4559, g2252, n11 );
nor U14230 ( new_g25247_, n4571, n4572 );
nor U14231 ( n4572, n7130, n4552 );
nor U14232 ( n4571, g2251, n13 );
nor U14233 ( new_g25251_, n4561, n4562 );
nor U14234 ( n4562, n7124, n4541 );
nor U14235 ( n4561, g2247, n10 );
nor U14236 ( new_g25246_, n4573, n4574 );
nor U14237 ( n4574, n7124, n4544 );
nor U14238 ( n4573, g2249, n11 );
nor U14239 ( new_g25237_, n4599, n4600 );
nor U14240 ( n4600, n7124, n4552 );
nor U14241 ( n4599, g2248, n13 );
nor U14242 ( new_g25245_, n4575, n4576 );
nor U14243 ( n4576, n4577, n4541 );
nor U14244 ( n4575, g2244, n10 );
nor U14245 ( new_g25236_, n4601, n4602 );
nor U14246 ( n4602, n4577, n4544 );
nor U14247 ( n4601, g2246, n11 );
nor U14248 ( new_g25227_, n4628, n4629 );
nor U14249 ( n4629, n4577, n4552 );
nor U14250 ( n4628, g2245, n13 );
nor U14251 ( new_g25255_, n4547, n4548 );
nor U14252 ( n4548, n3432, n4549 );
nor U14253 ( n4547, g1559, n12 );
nor U14254 ( new_g25250_, n4563, n4564 );
nor U14255 ( n4564, n3432, n4565 );
nor U14256 ( n4563, g1561, n14 );
nor U14257 ( new_g25244_, n4578, n4579 );
nor U14258 ( n4579, n3432, n4580 );
nor U14259 ( n4578, g1560, n16 );
nor U14260 ( new_g25249_, n4566, n4567 );
nor U14261 ( n4567, n7131, n4549 );
nor U14262 ( n4566, g1556, n12 );
nor U14263 ( new_g25243_, n4587, n4588 );
nor U14264 ( n4588, n7131, n4565 );
nor U14265 ( n4587, g1558, n14 );
nor U14266 ( new_g25235_, n4603, n4604 );
nor U14267 ( n4604, n7131, n4580 );
nor U14268 ( n4603, g1557, n16 );
nor U14269 ( new_g25242_, n4589, n4590 );
nor U14270 ( n4590, n7125, n4549 );
nor U14271 ( n4589, g1553, n12 );
nor U14272 ( new_g25234_, n4605, n4606 );
nor U14273 ( n4606, n7125, n4565 );
nor U14274 ( n4605, g1555, n14 );
nor U14275 ( new_g25225_, n4632, n4633 );
nor U14276 ( n4633, n7125, n4580 );
nor U14277 ( n4632, g1554, n16 );
nor U14278 ( new_g25233_, n4607, n4608 );
nor U14279 ( n4608, n4609, n4549 );
nor U14280 ( n4607, g1550, n12 );
nor U14281 ( new_g25224_, n4634, n4635 );
nor U14282 ( n4635, n4609, n4565 );
nor U14283 ( n4634, g1552, n14 );
nor U14284 ( new_g25217_, n4656, n4657 );
nor U14285 ( n4657, n4609, n4580 );
nor U14286 ( n4656, g1551, n16 );
nor U14287 ( new_g25248_, n4568, n4569 );
nor U14288 ( n4569, n3470, n4570 );
nor U14289 ( n4568, g865, n15 );
nor U14290 ( new_g25241_, n4591, n4592 );
nor U14291 ( n4592, n3470, n4593 );
nor U14292 ( n4591, g867, n17 );
nor U14293 ( new_g25232_, n4610, n4611 );
nor U14294 ( n4611, n3470, n4612 );
nor U14295 ( n4610, g866, n19 );
nor U14296 ( new_g25240_, n4594, n4595 );
nor U14297 ( n4595, n7137, n4570 );
nor U14298 ( n4594, g862, n15 );
nor U14299 ( new_g25231_, n4619, n4620 );
nor U14300 ( n4620, n7137, n4593 );
nor U14301 ( n4619, g864, n17 );
nor U14302 ( new_g25223_, n4636, n4637 );
nor U14303 ( n4637, n7137, n4612 );
nor U14304 ( n4636, g863, n19 );
nor U14305 ( new_g25230_, n4621, n4622 );
nor U14306 ( n4622, n7126, n4570 );
nor U14307 ( n4621, g859, n15 );
nor U14308 ( new_g25222_, n4638, n4639 );
nor U14309 ( n4639, n7126, n4593 );
nor U14310 ( n4638, g861, n17 );
nor U14311 ( new_g25215_, n4660, n4661 );
nor U14312 ( n4661, n7126, n4612 );
nor U14313 ( n4660, g860, n19 );
nor U14314 ( new_g25221_, n4640, n4641 );
nor U14315 ( n4641, n4642, n4570 );
nor U14316 ( n4640, g856, n15 );
nor U14317 ( new_g25214_, n4662, n4663 );
nor U14318 ( n4663, n4642, n4593 );
nor U14319 ( n4662, g858, n17 );
nor U14320 ( new_g25209_, n4671, n4672 );
nor U14321 ( n4672, n4642, n4612 );
nor U14322 ( n4671, g857, n19 );
nor U14323 ( new_g25239_, n4596, n4597 );
nor U14324 ( n4597, n3503, n4598 );
nor U14325 ( n4596, g177, n18 );
nor U14326 ( new_g25229_, n4623, n4624 );
nor U14327 ( n4624, n3503, n4625 );
nor U14328 ( n4623, g179, n20 );
nor U14329 ( new_g25220_, n4643, n4644 );
nor U14330 ( n4644, n3503, n4645 );
nor U14331 ( n4643, g178, n21 );
nor U14332 ( new_g25228_, n4626, n4627 );
nor U14333 ( n4627, n7138, n4598 );
nor U14334 ( n4626, g174, n18 );
nor U14335 ( new_g25219_, n4652, n4653 );
nor U14336 ( n4653, n7138, n4625 );
nor U14337 ( n4652, g176, n20 );
nor U14338 ( new_g25213_, n4664, n4665 );
nor U14339 ( n4665, n7138, n4645 );
nor U14340 ( n4664, g175, n21 );
nor U14341 ( new_g25218_, n4654, n4655 );
nor U14342 ( n4655, n7127, n4598 );
nor U14343 ( n4654, g171, n18 );
nor U14344 ( new_g25212_, n4666, n4667 );
nor U14345 ( n4667, n7127, n4625 );
nor U14346 ( n4666, g173, n20 );
nor U14347 ( new_g25207_, n4675, n4676 );
nor U14348 ( n4676, n7127, n4645 );
nor U14349 ( n4675, g172, n21 );
nor U14350 ( new_g25211_, n4668, n4669 );
nor U14351 ( n4669, n4670, n4598 );
nor U14352 ( n4668, g168, n18 );
nor U14353 ( new_g25206_, n4677, n4678 );
nor U14354 ( n4678, n4670, n4625 );
nor U14355 ( n4677, g170, n20 );
nor U14356 ( new_g25204_, n4679, n4680 );
nor U14357 ( n4680, n4670, n4645 );
nor U14358 ( n4679, g169, n21 );
nand U14359 ( n2271, n4742, n4743 );
nor U14360 ( n4742, n4747, n4748 );
and U14361 ( n4743, n4744, n4745 );
and U14362 ( n4747, g7302, g2661 );
nand U14363 ( n6083, g2645, g7390 );
nand U14364 ( n4745, n4746, g2598 );
nor U14365 ( n4746, new_g12539_, n7198 );
and U14366 ( new_g12539_, n6080, n6081 );
nand U14367 ( n6081, g2647, g2624 );
and U14368 ( n6080, n6082, n6083 );
nand U14369 ( n6082, g2643, g7302 );
nand U14370 ( n2847, g1930, new_g22651_ );
nand U14371 ( n2863, g7194, new_g22651_ );
nand U14372 ( n2889, g7052, new_g22651_ );
nand U14373 ( new_g22651_, n5075, n5076 );
nand U14374 ( n5075, n5078, n5069 );
nand U14375 ( n5076, n5077, g1890 );
nand U14376 ( n5078, n5079, n3853 );
nand U14377 ( n2608, n4815, n4816 );
nor U14378 ( n4815, n4820, n4821 );
and U14379 ( n4816, n4817, n4818 );
and U14380 ( n4821, g550, g593 );
nand U14381 ( n6099, g571, g6642 );
nand U14382 ( n4618, g785, g789 );
nand U14383 ( n4651, g97, g101 );
nand U14384 ( n4818, n4819, g524 );
nor U14385 ( n4819, new_g12487_, n7198 );
and U14386 ( new_g12487_, n6096, n6097 );
nand U14387 ( n6097, g573, g550 );
and U14388 ( n6096, n6098, n6099 );
nand U14389 ( n6098, g569, g6485 );
and U14390 ( n2607, n4804, n4805 );
nor U14391 ( n4804, n4809, n4810 );
and U14392 ( n4805, n4806, n4807 );
and U14393 ( n4809, g6485, g596 );
nand U14394 ( n6111, g567, g6642 );
nand U14395 ( n4807, n4808, g542 );
nor U14396 ( n4808, new_g12457_, n7198 );
and U14397 ( new_g12457_, n6108, n6109 );
nand U14398 ( n6109, g489, g550 );
and U14399 ( n6108, n6110, n6111 );
nand U14400 ( n6110, g565, g6485 );
nor U14401 ( new_g26776_, n267, n3519 );
xor U14402 ( n3519, n2830, g666 );
nor U14403 ( new_g26781_, n376, n3518 );
xor U14404 ( n3518, n2825, g1352 );
nor U14405 ( new_g26789_, n484, n3514 );
xor U14406 ( n3514, n2820, g2046 );
nor U14407 ( new_g26795_, n603, n3513 );
xor U14408 ( n3513, n3335, g2740 );
and U14409 ( n2270, n4723, n4724 );
nor U14410 ( n4723, n4728, n4729 );
and U14411 ( n4724, n4725, n4726 );
and U14412 ( n4728, g7302, g2670 );
nand U14413 ( n6095, g2641, g7390 );
nand U14414 ( n4726, n4727, g2616 );
nor U14415 ( n4727, new_g12499_, n7198 );
and U14416 ( new_g12499_, n6092, n6093 );
nand U14417 ( n6093, g2564, g2624 );
and U14418 ( n6092, n6094, n6095 );
nand U14419 ( n6094, g2639, g7302 );
nand U14420 ( n2499, n4795, n4796 );
nor U14421 ( n4795, n4800, n4801 );
and U14422 ( n4796, n4797, n4798 );
and U14423 ( n4800, g6750, g1273 );
nand U14424 ( n6090, g1255, g6750 );
nand U14425 ( n4798, n4799, g1210 );
nor U14426 ( n4799, new_g12507_, n7198 );
and U14427 ( new_g12507_, n6088, n6089 );
nand U14428 ( n6089, g1259, g1236 );
and U14429 ( n6088, n6090, n6091 );
nand U14430 ( n6091, g1257, g6944 );
nand U14431 ( n2384, n4770, n4771 );
nor U14432 ( n4770, n4775, n4776 );
and U14433 ( n4771, n4772, n4773 );
and U14434 ( n4775, g7052, g1967 );
and U14435 ( n2498, n4779, n4780 );
nor U14436 ( n4779, n4784, n4785 );
and U14437 ( n4780, n4781, n4782 );
and U14438 ( n4785, g6944, g1285 );
nand U14439 ( n6106, g1251, g6750 );
nand U14440 ( n6087, g1951, g7194 );
nand U14441 ( n4782, n4783, g1228 );
nor U14442 ( n4783, new_g12467_, n7198 );
nand U14443 ( n4773, n4774, g1904 );
nor U14444 ( n4774, new_g12524_, n7198 );
and U14445 ( new_g12524_, n6084, n6085 );
nand U14446 ( n6085, g1953, g1930 );
and U14447 ( n6084, n6086, n6087 );
nand U14448 ( n6086, g1949, g7052 );
and U14449 ( new_g12467_, n6104, n6105 );
nand U14450 ( n6105, g1176, g1236 );
and U14451 ( n6104, n6106, n6107 );
nand U14452 ( n6107, g1253, g6944 );
and U14453 ( n2383, n4751, n4752 );
nor U14454 ( n4751, n4756, n4757 );
and U14455 ( n4752, n4753, n4754 );
and U14456 ( n4756, g7052, g1976 );
nand U14457 ( n6103, g1947, g7194 );
nand U14458 ( n4754, n4755, g1922 );
nor U14459 ( n4755, new_g12482_, n7198 );
and U14460 ( new_g12482_, n6100, n6101 );
nand U14461 ( n6101, g1870, g1930 );
and U14462 ( n6100, n6102, n6103 );
nand U14463 ( n6102, g1945, g7052 );
nor U14464 ( new_g25940_, n4261, n4262 );
nor U14465 ( n4261, g2156, n4263 );
nand U14466 ( n4262, n3339, n2027 );
nor U14467 ( new_g25938_, n4265, n4266 );
nor U14468 ( n4265, g1462, n4267 );
nand U14469 ( n4266, n3343, n2033 );
nor U14470 ( new_g25935_, n4269, n4270 );
nor U14471 ( n4269, g776, n4271 );
nand U14472 ( n4270, n3347, n2039 );
nor U14473 ( new_g25932_, n4273, n4274 );
nor U14474 ( n4273, g88, n4275 );
nand U14475 ( n4274, n3351, n2044 );
nand U14476 ( n7088, n7014, n7015 );
nand U14477 ( n7015, g2498, g2476 );
nor U14478 ( n7014, n7016, n7017 );
and U14479 ( n7017, g5555, g2492 );
nand U14480 ( n7086, n7005, n7006 );
nand U14481 ( n7006, g1110, g1088 );
nor U14482 ( n7005, n7007, n7008 );
and U14483 ( n7008, g5472, g1104 );
and U14484 ( n7007, g6712, g1107 );
and U14485 ( n7016, g7264, g2495 );
nand U14486 ( n7087, n7009, n7010 );
nand U14487 ( n7010, g1804, g1782 );
nor U14488 ( n7009, n7011, n7012 );
and U14489 ( n7011, g7014, g1801 );
nand U14490 ( n7044, n6201, n6202 );
nand U14491 ( n6202, g423, g401 );
nor U14492 ( n6201, n6203, n6204 );
and U14493 ( n6203, g6447, g420 );
and U14494 ( n7012, g5511, g1798 );
and U14495 ( n6204, g5437, g417 );
nand U14496 ( n3877, g16355, n7159 );
nor U14497 ( new_g26660_, n3736, n3738 );
nor U14498 ( n3736, g672, n3739 );
nand U14499 ( n3738, n2830, n2828 );
nor U14500 ( new_g26666_, n3633, n3634 );
nor U14501 ( n3633, g1358, n3635 );
nand U14502 ( n3634, n2825, n2823 );
nor U14503 ( new_g26671_, n3535, n3536 );
nor U14504 ( n3535, g2052, n3537 );
nand U14505 ( n3536, n2820, n2818 );
nor U14506 ( new_g26677_, n3520, n3521 );
nor U14507 ( n3520, g2746, n3522 );
nand U14508 ( n3521, n3335, n3333 );
nand U14509 ( n2751, n3396, n3397 );
nand U14510 ( n3397, g2510, g2476 );
nor U14511 ( n3396, n3398, n3399 );
and U14512 ( n3399, g5555, g2504 );
nand U14513 ( n2795, n3471, n3472 );
nand U14514 ( n3472, g1122, g1088 );
nor U14515 ( n3471, n3473, n3475 );
and U14516 ( n3475, g5472, g1116 );
and U14517 ( n3473, g6712, g1119 );
and U14518 ( n3398, g7264, g2507 );
nand U14519 ( new_g12433_, n7384, n6112 );
nand U14520 ( n6112, g8021, n7293 );
nand U14521 ( n2774, n3433, n3434 );
nand U14522 ( n3434, g1816, g1782 );
nor U14523 ( n3433, n3435, n3436 );
and U14524 ( n3435, g7014, g1813 );
nand U14525 ( n2811, n3504, n3505 );
nand U14526 ( n3505, g435, g401 );
nor U14527 ( n3504, n3506, n3507 );
and U14528 ( n3506, g6447, g432 );
and U14529 ( n3436, g5511, g1810 );
and U14530 ( n3507, g5437, g429 );
nand U14531 ( n3868, n5098, n5099 );
nand U14532 ( n5099, g496, g550 );
nor U14533 ( n5098, n5100, n5101 );
and U14534 ( n5100, g6642, g493 );
and U14535 ( n5101, g6485, g490 );
nand U14536 ( n3365, n5452, n5453 );
nand U14537 ( n5453, g2519, g2476 );
nor U14538 ( n5452, n5454, n5455 );
and U14539 ( n5455, g5555, g2513 );
nand U14540 ( n3440, n5039, n5040 );
nand U14541 ( n5040, g1131, g1088 );
nor U14542 ( n5039, n5041, n5042 );
and U14543 ( n5042, g5472, g1125 );
and U14544 ( n5041, g6712, g1128 );
and U14545 ( n5454, g7264, g2516 );
nand U14546 ( n3862, n5089, n5090 );
nand U14547 ( n5090, g1183, g1236 );
nor U14548 ( n5089, n5091, n5092 );
and U14549 ( n5091, g6944, g1180 );
and U14550 ( n5092, g6750, g1177 );
nand U14551 ( n3844, n5071, n5072 );
nand U14552 ( n5072, g2571, g2624 );
nor U14553 ( n5071, n5073, n5074 );
and U14554 ( n5074, g7302, g2565 );
and U14555 ( n5073, g7390, g2568 );
nand U14556 ( n3402, n5029, n5030 );
nand U14557 ( n5030, g1825, g1782 );
nor U14558 ( n5029, n5031, n5032 );
and U14559 ( n5031, g7014, g1822 );
nand U14560 ( n3478, n5047, n5048 );
nand U14561 ( n5048, g444, g401 );
nor U14562 ( n5047, n5049, n5050 );
and U14563 ( n5049, g6447, g441 );
and U14564 ( n5032, g5511, g1819 );
and U14565 ( n5050, g5437, g438 );
nand U14566 ( n3853, n5080, n5081 );
nand U14567 ( n5081, g1877, g1930 );
nor U14568 ( n5080, n5082, n5083 );
and U14569 ( n5083, g7052, g1871 );
and U14570 ( n5082, g7194, g1874 );
nor U14571 ( new_g25067_, n29, n4699 );
xnor U14572 ( n4699, n4264, g2160 );
nor U14573 ( new_g25056_, n27, n4700 );
xnor U14574 ( n4700, n4268, g1466 );
nor U14575 ( new_g25042_, n25, n4701 );
xnor U14576 ( n4701, n4272, g780 );
nor U14577 ( new_g25027_, n23, n4702 );
xnor U14578 ( n4702, n4276, g92 );
and U14579 ( n5481, g3018, g3028 );
nor U14580 ( n5482, n5431, n5484 );
or U14581 ( n5484, g3032, g3036 );
nand U14582 ( n5431, n5485, n5486 );
nor U14583 ( n5485, n7100, n5489 );
nor U14584 ( n5486, n5487, n5488 );
nand U14585 ( n5489, g3013, g3002 );
nand U14586 ( n5488, g2998, n7099 );
nand U14587 ( n2101, n2118, n2119 );
nand U14588 ( n2119, g2489, g2476 );
nor U14589 ( n2118, n2120, n2121 );
and U14590 ( n2121, g5555, g2483 );
nand U14591 ( n2180, n2198, n2199 );
nand U14592 ( n2199, g1101, g1088 );
nor U14593 ( n2198, n2201, n2202 );
and U14594 ( n2202, g5472, g1095 );
and U14595 ( n2201, g6712, g1098 );
and U14596 ( n2120, g7264, g2486 );
nand U14597 ( new_g24499_, n4802, n4803 );
nand U14598 ( n4802, g596, n7162 );
nand U14599 ( n4803, n4767, g6485 );
nand U14600 ( new_g24508_, n4788, n4789 );
nand U14601 ( n4788, g599, n7171 );
nand U14602 ( n4789, n4767, g6642 );
nand U14603 ( new_g24519_, n4765, n4766 );
nand U14604 ( n4765, g602, n7169 );
nand U14605 ( n4766, n4767, g550 );
nand U14606 ( new_g24532_, n4737, n4738 );
nand U14607 ( n4737, g1288, n7167 );
nand U14608 ( n4738, n4739, g1236 );
nand U14609 ( new_g24545_, n4718, n4719 );
nand U14610 ( n4718, g1982, n7168 );
nand U14611 ( n4719, n4720, g1930 );
nand U14612 ( new_g24547_, n4715, n4716 );
nand U14613 ( n4715, g2667, n7179 );
nand U14614 ( n4716, n4717, g2624 );
nand U14615 ( new_g24557_, n4710, n4711 );
nand U14616 ( n4710, g2676, n7179 );
nand U14617 ( n4711, n4712, g2624 );
nand U14618 ( new_g24511_, n4777, n4778 );
nand U14619 ( n4777, g1282, n7122 );
nand U14620 ( n4778, n4739, g6750 );
nand U14621 ( new_g24537_, n4730, n4731 );
nand U14622 ( n4730, g2664, n7161 );
nand U14623 ( n4731, n4717, g7390 );
nand U14624 ( new_g24548_, n4713, n4714 );
nand U14625 ( n4713, g2673, n7161 );
nand U14626 ( n4714, n4712, g7390 );
nand U14627 ( new_g24522_, n4760, n4761 );
nand U14628 ( n4760, g1285, n7159 );
nand U14629 ( n4761, n4739, g6944 );
nand U14630 ( new_g24535_, n4732, n4733 );
nand U14631 ( n4732, g1979, n7158 );
nand U14632 ( n4733, n4720, g7194 );
nand U14633 ( new_g24525_, n4749, n4750 );
nand U14634 ( n4749, g1976, n7155 );
nand U14635 ( n4750, n4720, g7052 );
nand U14636 ( new_g24527_, n4740, n4741 );
nand U14637 ( n4740, g2661, n7160 );
nand U14638 ( n4741, n4717, g7302 );
nand U14639 ( new_g24538_, n4721, n4722 );
nand U14640 ( n4721, g2670, n7160 );
nand U14641 ( n4722, n4712, g7302 );
nand U14642 ( n2143, n2159, n2160 );
nand U14643 ( n2160, g1795, g1782 );
nor U14644 ( n2159, n2161, n2162 );
and U14645 ( n2161, g7014, g1792 );
nand U14646 ( n2215, n2232, n2233 );
nand U14647 ( n2233, g414, g401 );
nor U14648 ( n2232, n2234, n2235 );
and U14649 ( n2234, g6447, g411 );
and U14650 ( n2162, g5511, g1789 );
and U14651 ( n2235, g5437, g408 );
nand U14652 ( n5000, n4174, g2998 );
nand U14653 ( n4695, n4696, g3002 );
nor U14654 ( new_g25185_, n267, n4698 );
xor U14655 ( n4698, n3740, g660 );
nor U14656 ( new_g25189_, n376, n4697 );
xor U14657 ( n4697, n3636, g1346 );
nor U14658 ( new_g25194_, n484, n4692 );
xor U14659 ( n4692, n3538, g2040 );
nor U14660 ( new_g25197_, n603, n4691 );
xor U14661 ( n4691, n3523, g2734 );
nand U14662 ( n5691, n5750, g2612 );
nor U14663 ( n5750, g2733, n7101 );
nand U14664 ( n5731, n5776, g1918 );
nor U14665 ( n5776, g2039, n7102 );
nand U14666 ( n5765, n5796, g1224 );
nor U14667 ( n5796, g1345, n7103 );
nand U14668 ( n5791, n5807, g538 );
nor U14669 ( n5807, g659, n7104 );
nor U14670 ( new_g20939_, n5721, n5722 );
nor U14671 ( n5721, g2774, n4367 );
nor U14672 ( n5722, n7254, n591 );
nor U14673 ( new_g20941_, n5717, n5718 );
nor U14674 ( n5717, g2801, n4367 );
nor U14675 ( n5718, n7258, n591 );
nor U14676 ( new_g20963_, n5687, n5688 );
nor U14677 ( n5687, g2777, n4367 );
nor U14678 ( n5688, n7199, n591 );
nor U14679 ( new_g20982_, n5650, n5651 );
nor U14680 ( n5650, g2780, n4367 );
nor U14681 ( n5651, n7194, n591 );
nor U14682 ( new_g21005_, n5612, n5613 );
nor U14683 ( n5612, g2783, n4367 );
nor U14684 ( n5613, n7279, n591 );
nor U14685 ( new_g21026_, n5576, n5577 );
nor U14686 ( n5576, g2786, n4367 );
nor U14687 ( n5577, n7219, n591 );
nor U14688 ( new_g21044_, n5546, n5547 );
nor U14689 ( n5546, g2789, n4367 );
nor U14690 ( n5547, n7280, n591 );
nor U14691 ( new_g21061_, n5524, n5525 );
nor U14692 ( n5524, g2792, n4367 );
nor U14693 ( n5525, n7234, n591 );
nor U14694 ( new_g21074_, n5509, n5510 );
nor U14695 ( n5509, g2795, n4367 );
nor U14696 ( n5510, n7275, n591 );
nor U14697 ( new_g21082_, n5499, n5500 );
nor U14698 ( n5499, g2798, n4367 );
nor U14699 ( n5500, n7249, n591 );
nor U14700 ( new_g20962_, n5689, n5690 );
nor U14701 ( n5689, g2772, n4364 );
nor U14702 ( n5690, n7254, n592 );
nor U14703 ( new_g20965_, n5683, n5684 );
nor U14704 ( n5683, g2799, n4364 );
nor U14705 ( n5684, n7258, n592 );
nor U14706 ( new_g20981_, n5652, n5653 );
nor U14707 ( n5652, g2775, n4364 );
nor U14708 ( n5653, n7199, n592 );
nor U14709 ( new_g21004_, n5614, n5615 );
nor U14710 ( n5614, g2778, n4364 );
nor U14711 ( n5615, n7194, n592 );
nor U14712 ( new_g21025_, n5578, n5579 );
nor U14713 ( n5578, g2781, n4364 );
nor U14714 ( n5579, n7279, n592 );
nor U14715 ( new_g21043_, n5548, n5549 );
nor U14716 ( n5548, g2784, n4364 );
nor U14717 ( n5549, n7219, n592 );
nor U14718 ( new_g21060_, n5526, n5527 );
nor U14719 ( n5526, g2787, n4364 );
nor U14720 ( n5527, n7280, n592 );
nor U14721 ( new_g21073_, n5511, n5512 );
nor U14722 ( n5511, g2790, n4364 );
nor U14723 ( n5512, n7234, n592 );
nor U14724 ( new_g21081_, n5502, n5503 );
nor U14725 ( n5502, g2793, n4364 );
nor U14726 ( n5503, n7275, n592 );
nor U14727 ( new_g21094_, n5497, n5498 );
nor U14728 ( n5497, g2796, n4364 );
nor U14729 ( n5498, n7249, n592 );
nor U14730 ( new_g20915_, n5755, n5756 );
nor U14731 ( n5755, g2080, n4410 );
nor U14732 ( n5756, n7255, n473 );
nor U14733 ( new_g20917_, n5751, n5752 );
nor U14734 ( n5751, g2107, n4410 );
nor U14735 ( n5752, n7259, n473 );
nor U14736 ( new_g20935_, n5727, n5728 );
nor U14737 ( n5727, g2083, n4410 );
nor U14738 ( n5728, n7200, n473 );
nor U14739 ( new_g20954_, n5694, n5695 );
nor U14740 ( n5694, g2086, n4410 );
nor U14741 ( n5695, n7195, n473 );
nor U14742 ( new_g20978_, n5658, n5659 );
nor U14743 ( n5658, g2089, n4410 );
nor U14744 ( n5659, n7281, n473 );
nor U14745 ( new_g21000_, n5624, n5626 );
nor U14746 ( n5624, g2092, n4410 );
nor U14747 ( n5626, n7220, n473 );
nor U14748 ( new_g21020_, n5586, n5587 );
nor U14749 ( n5586, g2095, n4410 );
nor U14750 ( n5587, n7282, n473 );
nor U14751 ( new_g21040_, n5555, n5556 );
nor U14752 ( n5555, g2098, n4410 );
nor U14753 ( n5556, n7235, n473 );
nor U14754 ( new_g21055_, n5530, n5531 );
nor U14755 ( n5530, g2101, n4410 );
nor U14756 ( n5531, n7276, n473 );
nor U14757 ( new_g21072_, n5513, n5514 );
nor U14758 ( n5513, g2104, n4410 );
nor U14759 ( n5514, n7250, n473 );
nor U14760 ( new_g20934_, n5729, n5730 );
nor U14761 ( n5729, g2078, n4371 );
nor U14762 ( n5730, n7255, n474 );
nor U14763 ( new_g20937_, n5723, n5724 );
nor U14764 ( n5723, g2105, n4371 );
nor U14765 ( n5724, n7259, n474 );
nor U14766 ( new_g20953_, n5696, n5697 );
nor U14767 ( n5696, g2081, n4371 );
nor U14768 ( n5697, n7200, n474 );
nor U14769 ( new_g20977_, n5660, n5661 );
nor U14770 ( n5660, g2084, n4371 );
nor U14771 ( n5661, n7195, n474 );
nor U14772 ( new_g20999_, n5627, n5628 );
nor U14773 ( n5627, g2087, n4371 );
nor U14774 ( n5628, n7281, n474 );
nor U14775 ( new_g21019_, n5588, n5590 );
nor U14776 ( n5588, g2090, n4371 );
nor U14777 ( n5590, n7220, n474 );
nor U14778 ( new_g21039_, n5557, n5558 );
nor U14779 ( n5557, g2093, n4371 );
nor U14780 ( n5558, n7282, n474 );
nor U14781 ( new_g21054_, n5532, n5533 );
nor U14782 ( n5532, g2096, n4371 );
nor U14783 ( n5533, n7235, n474 );
nor U14784 ( new_g21071_, n5515, n5516 );
nor U14785 ( n5515, g2099, n4371 );
nor U14786 ( n5516, n7276, n474 );
nor U14787 ( new_g21080_, n5504, n5506 );
nor U14788 ( n5504, g2102, n4371 );
nor U14789 ( n5506, n7250, n474 );
nor U14790 ( new_g20896_, n5781, n5782 );
nor U14791 ( n5781, g1386, n4453 );
nor U14792 ( n5782, n7256, n365 );
nor U14793 ( new_g20898_, n5777, n5778 );
nor U14794 ( n5777, g1413, n4453 );
nor U14795 ( n5778, n7260, n365 );
nor U14796 ( new_g20911_, n5761, n5762 );
nor U14797 ( n5761, g1389, n4453 );
nor U14798 ( n5762, n7201, n365 );
nor U14799 ( new_g20926_, n5734, n5735 );
nor U14800 ( n5734, g1392, n4453 );
nor U14801 ( n5735, n7196, n365 );
nor U14802 ( new_g20950_, n5702, n5703 );
nor U14803 ( n5702, g1395, n4453 );
nor U14804 ( n5703, n7283, n365 );
nor U14805 ( new_g20973_, n5669, n5670 );
nor U14806 ( n5669, g1398, n4453 );
nor U14807 ( n5670, n7221, n365 );
nor U14808 ( new_g20994_, n5635, n5636 );
nor U14809 ( n5635, g1401, n4453 );
nor U14810 ( n5636, n7284, n365 );
nor U14811 ( new_g21016_, n5597, n5598 );
nor U14812 ( n5597, g1404, n4453 );
nor U14813 ( n5598, n7236, n365 );
nor U14814 ( new_g21034_, n5561, n5562 );
nor U14815 ( n5561, g1407, n4453 );
nor U14816 ( n5562, n7277, n365 );
nor U14817 ( new_g21053_, n5534, n5535 );
nor U14818 ( n5534, g1410, n4453 );
nor U14819 ( n5535, n7251, n365 );
nor U14820 ( new_g20910_, n5763, n5764 );
nor U14821 ( n5763, g1384, n4414 );
nor U14822 ( n5764, n7256, n366 );
nor U14823 ( new_g20913_, n5757, n5758 );
nor U14824 ( n5757, g1411, n4414 );
nor U14825 ( n5758, n7260, n366 );
nor U14826 ( new_g20925_, n5736, n5737 );
nor U14827 ( n5736, g1387, n4414 );
nor U14828 ( n5737, n7201, n366 );
nor U14829 ( new_g20949_, n5704, n5705 );
nor U14830 ( n5704, g1390, n4414 );
nor U14831 ( n5705, n7196, n366 );
nor U14832 ( new_g20972_, n5671, n5672 );
nor U14833 ( n5671, g1393, n4414 );
nor U14834 ( n5672, n7283, n366 );
nor U14835 ( new_g20993_, n5637, n5638 );
nor U14836 ( n5637, g1396, n4414 );
nor U14837 ( n5638, n7221, n366 );
nor U14838 ( new_g21015_, n5599, n5600 );
nor U14839 ( n5599, g1399, n4414 );
nor U14840 ( n5600, n7284, n366 );
nor U14841 ( new_g21033_, n5563, n5564 );
nor U14842 ( n5563, g1402, n4414 );
nor U14843 ( n5564, n7236, n366 );
nor U14844 ( new_g21052_, n5536, n5537 );
nor U14845 ( n5536, g1405, n4414 );
nor U14846 ( n5537, n7277, n366 );
nor U14847 ( new_g21070_, n5517, n5518 );
nor U14848 ( n5517, g1408, n4414 );
nor U14849 ( n5518, n7251, n366 );
nor U14850 ( new_g20879_, n5801, n5802 );
nor U14851 ( n5801, g700, n4502 );
nor U14852 ( n5802, n7257, n256 );
nor U14853 ( new_g20881_, n5797, n5798 );
nor U14854 ( n5797, g727, n4502 );
nor U14855 ( n5798, n7261, n256 );
nor U14856 ( new_g20892_, n5787, n5788 );
nor U14857 ( n5787, g703, n4502 );
nor U14858 ( n5788, n7203, n256 );
nor U14859 ( new_g20902_, n5768, n5769 );
nor U14860 ( n5768, g706, n4502 );
nor U14861 ( n5769, n7197, n256 );
nor U14862 ( new_g20922_, n5742, n5743 );
nor U14863 ( n5742, g709, n4502 );
nor U14864 ( n5743, n7285, n256 );
nor U14865 ( new_g20945_, n5713, n5714 );
nor U14866 ( n5713, g712, n4502 );
nor U14867 ( n5714, n7222, n256 );
nor U14868 ( new_g20967_, n5679, n5680 );
nor U14869 ( n5679, g715, n4502 );
nor U14870 ( n5680, n7286, n256 );
nor U14871 ( new_g20990_, n5644, n5645 );
nor U14872 ( n5644, g718, n4502 );
nor U14873 ( n5645, n7237, n256 );
nor U14874 ( new_g21010_, n5604, n5605 );
nor U14875 ( n5604, g721, n4502 );
nor U14876 ( n5605, n7278, n256 );
nor U14877 ( new_g21032_, n5565, n5566 );
nor U14878 ( n5565, g724, n4502 );
nor U14879 ( n5566, n7252, n256 );
nor U14880 ( new_g20891_, n5789, n5790 );
nor U14881 ( n5789, g698, n4457 );
nor U14882 ( n5790, n7257, n257 );
nor U14883 ( new_g20894_, n5783, n5784 );
nor U14884 ( n5783, g725, n4457 );
nor U14885 ( n5784, n7261, n257 );
nor U14886 ( new_g20901_, n5770, n5771 );
nor U14887 ( n5770, g701, n4457 );
nor U14888 ( n5771, n7203, n257 );
nor U14889 ( new_g20921_, n5744, n5745 );
nor U14890 ( n5744, g704, n4457 );
nor U14891 ( n5745, n7197, n257 );
nor U14892 ( new_g20944_, n5715, n5716 );
nor U14893 ( n5715, g707, n4457 );
nor U14894 ( n5716, n7285, n257 );
nor U14895 ( new_g20966_, n5681, n5682 );
nor U14896 ( n5681, g710, n4457 );
nor U14897 ( n5682, n7222, n257 );
nor U14898 ( new_g20989_, n5646, n5647 );
nor U14899 ( n5646, g713, n4457 );
nor U14900 ( n5647, n7286, n257 );
nor U14901 ( new_g21009_, n5606, n5607 );
nor U14902 ( n5606, g716, n4457 );
nor U14903 ( n5607, n7237, n257 );
nor U14904 ( new_g21031_, n5567, n5568 );
nor U14905 ( n5567, g719, n4457 );
nor U14906 ( n5568, n7278, n257 );
nor U14907 ( new_g21051_, n5538, n5539 );
nor U14908 ( n5538, g722, n4457 );
nor U14909 ( n5539, n7252, n257 );
and U14910 ( n4748, g2624, g2667 );
nand U14911 ( n1672, g2384, n2101 );
nand U14912 ( n1716, g996, n2180 );
and U14913 ( n4820, g6485, g587 );
nor U14914 ( new_g20918_, n5748, n5749 );
nor U14915 ( n5748, g2773, n4407 );
nor U14916 ( n5749, n7254, n590 );
nor U14917 ( new_g20919_, n5746, n5747 );
nor U14918 ( n5746, g2800, n4407 );
nor U14919 ( n5747, n7258, n590 );
nor U14920 ( new_g20940_, n5719, n5720 );
nor U14921 ( n5719, g2776, n4407 );
nor U14922 ( n5720, n7199, n590 );
nor U14923 ( new_g20964_, n5685, n5686 );
nor U14924 ( n5685, g2779, n4407 );
nor U14925 ( n5686, n7194, n590 );
nor U14926 ( new_g20983_, n5648, n5649 );
nor U14927 ( n5648, g2782, n4407 );
nor U14928 ( n5649, n7279, n590 );
nor U14929 ( new_g21006_, n5610, n5611 );
nor U14930 ( n5610, g2785, n4407 );
nor U14931 ( n5611, n7219, n590 );
nor U14932 ( new_g21027_, n5574, n5575 );
nor U14933 ( n5574, g2788, n4407 );
nor U14934 ( n5575, n7280, n590 );
nor U14935 ( new_g21045_, n5544, n5545 );
nor U14936 ( n5544, g2791, n4407 );
nor U14937 ( n5545, n7234, n590 );
nor U14938 ( new_g21062_, n5522, n5523 );
nor U14939 ( n5522, g2794, n4407 );
nor U14940 ( n5523, n7275, n590 );
nor U14941 ( new_g21075_, n5507, n5508 );
nor U14942 ( n5507, g2797, n4407 );
nor U14943 ( n5508, n7249, n590 );
nor U14944 ( new_g20899_, n5774, n5775 );
nor U14945 ( n5774, g2079, n4450 );
nor U14946 ( n5775, n7255, n472 );
nor U14947 ( new_g20900_, n5772, n5773 );
nor U14948 ( n5772, g2106, n4450 );
nor U14949 ( n5773, n7259, n472 );
nor U14950 ( new_g20916_, n5753, n5754 );
nor U14951 ( n5753, g2082, n4450 );
nor U14952 ( n5754, n7200, n472 );
nor U14953 ( new_g20936_, n5725, n5726 );
nor U14954 ( n5725, g2085, n4450 );
nor U14955 ( n5726, n7195, n472 );
nor U14956 ( new_g20955_, n5692, n5693 );
nor U14957 ( n5692, g2088, n4450 );
nor U14958 ( n5693, n7281, n472 );
nor U14959 ( new_g20979_, n5656, n5657 );
nor U14960 ( n5656, g2091, n4450 );
nor U14961 ( n5657, n7220, n472 );
nor U14962 ( new_g21001_, n5622, n5623 );
nor U14963 ( n5622, g2094, n4450 );
nor U14964 ( n5623, n7282, n472 );
nor U14965 ( new_g21021_, n5584, n5585 );
nor U14966 ( n5584, g2097, n4450 );
nor U14967 ( n5585, n7235, n472 );
nor U14968 ( new_g21041_, n5553, n5554 );
nor U14969 ( n5553, g2100, n4450 );
nor U14970 ( n5554, n7276, n472 );
nor U14971 ( new_g21056_, n5528, n5529 );
nor U14972 ( n5528, g2103, n4450 );
nor U14973 ( n5529, n7250, n472 );
nor U14974 ( new_g20882_, n5794, n5795 );
nor U14975 ( n5794, g1385, n4499 );
nor U14976 ( n5795, n7256, n364 );
nor U14977 ( new_g20883_, n5792, n5793 );
nor U14978 ( n5792, g1412, n4499 );
nor U14979 ( n5793, n7260, n364 );
nor U14980 ( new_g20897_, n5779, n5780 );
nor U14981 ( n5779, g1388, n4499 );
nor U14982 ( n5780, n7201, n364 );
nor U14983 ( new_g20912_, n5759, n5760 );
nor U14984 ( n5759, g1391, n4499 );
nor U14985 ( n5760, n7196, n364 );
nor U14986 ( new_g20927_, n5732, n5733 );
nor U14987 ( n5732, g1394, n4499 );
nor U14988 ( n5733, n7283, n364 );
nor U14989 ( new_g20951_, n5700, n5701 );
nor U14990 ( n5700, g1397, n4499 );
nor U14991 ( n5701, n7221, n364 );
nor U14992 ( new_g20974_, n5667, n5668 );
nor U14993 ( n5667, g1400, n4499 );
nor U14994 ( n5668, n7284, n364 );
nor U14995 ( new_g20995_, n5633, n5634 );
nor U14996 ( n5633, g1403, n4499 );
nor U14997 ( n5634, n7236, n364 );
nor U14998 ( new_g21017_, n5595, n5596 );
nor U14999 ( n5595, g1406, n4499 );
nor U15000 ( n5596, n7277, n364 );
nor U15001 ( new_g21035_, n5559, n5560 );
nor U15002 ( n5559, g1409, n4499 );
nor U15003 ( n5560, n7251, n364 );
nor U15004 ( new_g20875_, n5805, n5806 );
nor U15005 ( n5805, g699, n4538 );
nor U15006 ( n5806, n7257, n255 );
nor U15007 ( new_g20876_, n5803, n5804 );
nor U15008 ( n5803, g726, n4538 );
nor U15009 ( n5804, n7261, n255 );
nor U15010 ( new_g20880_, n5799, n5800 );
nor U15011 ( n5799, g702, n4538 );
nor U15012 ( n5800, n7203, n255 );
nor U15013 ( new_g20893_, n5785, n5786 );
nor U15014 ( n5785, g705, n4538 );
nor U15015 ( n5786, n7197, n255 );
nor U15016 ( new_g20903_, n5766, n5767 );
nor U15017 ( n5766, g708, n4538 );
nor U15018 ( n5767, n7285, n255 );
nor U15019 ( new_g20923_, n5740, n5741 );
nor U15020 ( n5740, g711, n4538 );
nor U15021 ( n5741, n7222, n255 );
nor U15022 ( new_g20946_, n5711, n5712 );
nor U15023 ( n5711, g714, n4538 );
nor U15024 ( n5712, n7286, n255 );
nor U15025 ( new_g20968_, n5677, n5678 );
nor U15026 ( n5677, g717, n4538 );
nor U15027 ( n5678, n7237, n255 );
nor U15028 ( new_g20991_, n5642, n5643 );
nor U15029 ( n5642, g720, n4538 );
nor U15030 ( n5643, n7278, n255 );
nor U15031 ( new_g21011_, n5601, n5603 );
nor U15032 ( n5601, g723, n4538 );
nor U15033 ( n5603, n7252, n255 );
nand U15034 ( n4832, n5426, g3018 );
nor U15035 ( n4831, n4832, n7240 );
nand U15036 ( n4684, g3036, n4831 );
and U15037 ( n4810, g6642, g599 );
and U15038 ( n4801, g1236, g1279 );
and U15039 ( n4776, g1930, g1973 );
nand U15040 ( n1694, g1690, n2143 );
nand U15041 ( n1735, g309, n2215 );
nand U15042 ( new_g28420_, n2247, n2248 );
nand U15043 ( n2247, g3100, n7242 );
nand U15044 ( n2248, g8106, n241 );
nand U15045 ( new_g28421_, n2245, n2246 );
nand U15046 ( n2245, g3101, n7243 );
nand U15047 ( n2246, g8030, n241 );
and U15048 ( n4729, g7390, g2673 );
nand U15049 ( new_g28425_, n2243, n2244 );
nand U15050 ( n2243, g3102, n7245 );
nand U15051 ( n2244, g3109, n241 );
and U15052 ( n4784, g6750, g1282 );
and U15053 ( n4757, g7194, g1979 );
nand U15054 ( n4744, g2664, g7390 );
nand U15055 ( n4817, g590, g6642 );
nand U15056 ( n4806, g602, g550 );
nand U15057 ( n4781, g1288, g1236 );
nand U15058 ( n4753, g1982, g1930 );
nand U15059 ( n4725, g2676, g2624 );
nor U15060 ( new_g24426_, n4846, n4847 );
nor U15061 ( n4846, g646, n4848 );
nand U15062 ( n4847, n3740, n2828 );
nor U15063 ( new_g24430_, n4842, n4843 );
nor U15064 ( n4842, g1332, n4844 );
nand U15065 ( n4843, n3636, n2823 );
nor U15066 ( new_g24434_, n4838, n4839 );
nor U15067 ( n4838, g2026, n4840 );
nand U15068 ( n4839, n3538, n2818 );
nor U15069 ( new_g24438_, n4834, n4835 );
nor U15070 ( n4834, g2720, n4836 );
nand U15071 ( n4835, n3523, n3333 );
nand U15072 ( n5126, g1563, n7400 );
nand U15073 ( n5146, g869, n7410 );
nand U15074 ( n5181, g181, n7420 );
nand U15075 ( n4797, g1276, g6944 );
nand U15076 ( n4772, g1970, g7194 );
nand U15077 ( n5116, g2257, n7390 );
nand U15078 ( n4994, g2883, g2950 );
or U15079 ( n4993, n4994, n7381 );
nand U15080 ( n4687, n4688, g2892 );
nor U15081 ( new_g26798_, n3508, n3509 );
xnor U15082 ( n3508, g2908, n3511 );
nor U15083 ( n3511, n3512, n7223 );
nand U15084 ( n5069, n5838, n5839 );
nor U15085 ( n5838, g3006, g3002 );
nor U15086 ( n5839, g3010, n5840 );
nand U15087 ( n5840, n7204, n7100 );
nand U15088 ( new_g24491_, n4813, n4814 );
nand U15089 ( n4813, g587, n7162 );
nand U15090 ( n4814, n4792, g6485 );
nand U15091 ( new_g24498_, n4811, n4812 );
nand U15092 ( n4811, g590, n7171 );
nand U15093 ( n4812, n4792, g6642 );
nand U15094 ( new_g24507_, n4790, n4791 );
nand U15095 ( n4790, g593, n7169 );
nand U15096 ( n4791, n4792, g550 );
nand U15097 ( new_g24521_, n4762, n4763 );
nand U15098 ( n4762, g1279, n7167 );
nand U15099 ( n4763, n4764, g1236 );
nand U15100 ( new_g24501_, n4793, n4794 );
nand U15101 ( n4793, g1273, n7122 );
nand U15102 ( n4794, n4764, g6750 );
nand U15103 ( new_g24510_, n4786, n4787 );
nand U15104 ( n4786, g1276, n7159 );
nand U15105 ( n4787, n4764, g6944 );
nand U15106 ( new_g24534_, n4734, n4735 );
nand U15107 ( n4734, g1973, n7168 );
nand U15108 ( n4735, n4736, g1930 );
nand U15109 ( new_g24524_, n4758, n4759 );
nand U15110 ( n4758, g1970, n7158 );
nand U15111 ( n4759, n4736, g7194 );
nand U15112 ( new_g24513_, n4768, n4769 );
nand U15113 ( n4768, g1967, n7155 );
nand U15114 ( n4769, n4736, g7052 );
nand U15115 ( n2051, g16399, n7158 );
nand U15116 ( n4690, n4825, g2924 );
nand U15117 ( n5818, g2950, g2908 );
and U15118 ( n4825, g2917, n4826 );
nor U15119 ( new_g25199_, n2, n4689 );
xor U15120 ( n4689, n4690, g2920 );
nor U15121 ( n6331, g734, n7181 );
nor U15122 ( n6898, g2808, n7178 );
nor U15123 ( n6700, g2114, n7177 );
nor U15124 ( n6505, g1420, n7176 );
nor U15125 ( new_g26037_, n4176, n3509 );
xor U15126 ( n4176, n3512, g2900 );
nand U15127 ( n5816, g2888, n7105 );
nor U15128 ( n6392, g736, n7180 );
nor U15129 ( n6900, g2810, n7172 );
nor U15130 ( n6702, g2116, n7173 );
nor U15131 ( n6507, g1422, n7174 );
or U15132 ( n6075, g2888, g2912 );
nand U15133 ( n5817, g2903, g2892 );
nand U15134 ( n4824, n3509, n5436 );
nand U15135 ( n5436, n5437, n7246 );
nand U15136 ( n5437, n5439, n5440 );
and U15137 ( n5439, g2912, g2920 );
nor U15138 ( new_g23357_, n2, n4995 );
xor U15139 ( n4995, n7, g2917 );
nand U15140 ( new_g26541_, n3865, n3866 );
nand U15141 ( n3865, g490, n7162 );
nand U15142 ( n3866, n3858, g6485 );
nand U15143 ( new_g26545_, n3863, n3864 );
nand U15144 ( n3863, g493, n7171 );
nand U15145 ( n3864, n3858, g6642 );
nand U15146 ( new_g26553_, n3856, n3857 );
nand U15147 ( n3856, g496, n7169 );
nand U15148 ( n3857, n3858, g550 );
nand U15149 ( new_g26569_, n3847, n3848 );
nand U15150 ( n3847, g1183, n7167 );
nand U15151 ( n3848, n3849, g1236 );
nand U15152 ( new_g26547_, n3859, n3860 );
nand U15153 ( n3859, g1177, n7122 );
nand U15154 ( n3860, n3849, g6750 );
nand U15155 ( new_g26557_, n3854, n3855 );
nand U15156 ( n3854, g1180, n7159 );
nand U15157 ( n3855, n3849, g6944 );
nor U15158 ( new_g23324_, n267, n5002 );
xor U15159 ( n5002, n4849, g653 );
nor U15160 ( new_g23329_, n376, n5001 );
xor U15161 ( n5001, n4845, g1339 );
nor U15162 ( new_g23339_, n484, n4997 );
xor U15163 ( n4997, n4841, g2033 );
nor U15164 ( new_g23348_, n603, n4996 );
xor U15165 ( n4996, n4837, g2727 );
nand U15166 ( new_g26616_, n3833, n3834 );
nand U15167 ( n3833, g2571, n7179 );
nand U15168 ( n3834, n3835, g2624 );
nand U15169 ( new_g26596_, n3836, n3837 );
nand U15170 ( n3836, g2568, n7161 );
nand U15171 ( n3837, n3835, g7390 );
nand U15172 ( new_g26575_, n3841, n3842 );
nand U15173 ( n3841, g2565, n7160 );
nand U15174 ( n3842, n3835, g7302 );
nor U15175 ( new_g20924_, n5738, n5739 );
nor U15176 ( n5738, g729, n259 );
nor U15177 ( n5739, n223, n5708 );
nor U15178 ( new_g20969_, n5675, n5676 );
nor U15179 ( n5675, g728, n269 );
nor U15180 ( n5676, n223, n5641 );
nor U15181 ( new_g20947_, n5709, n5710 );
nor U15182 ( n5709, g730, n267 );
nor U15183 ( n5710, n223, n2828 );
nor U15184 ( new_g24476_, n4822, n4823 );
nor U15185 ( n4822, g2924, n4825 );
nand U15186 ( n4823, n4690, n4824 );
nor U15187 ( new_g20952_, n5698, n5699 );
nor U15188 ( n5698, g1415, n368 );
nor U15189 ( n5699, n346, n5664 );
nor U15190 ( new_g20996_, n5631, n5632 );
nor U15191 ( n5631, g1414, n378 );
nor U15192 ( n5632, n346, n5594 );
nor U15193 ( new_g20975_, n5665, n5666 );
nor U15194 ( n5665, g1416, n376 );
nor U15195 ( n5666, n346, n2823 );
nand U15196 ( new_g26592_, n3838, n3839 );
nand U15197 ( n3838, g1877, n7168 );
nand U15198 ( n3839, n3840, g1930 );
nand U15199 ( new_g26573_, n3845, n3846 );
nand U15200 ( n3845, g1874, n7158 );
nand U15201 ( n3846, n3840, g7194 );
nand U15202 ( new_g26559_, n3850, n3851 );
nand U15203 ( n3850, g1871, n7155 );
nand U15204 ( n3851, n3840, g7052 );
nor U15205 ( new_g21007_, n5608, n5609 );
nor U15206 ( n5608, g2803, n594 );
nor U15207 ( n5609, n570, n5571 );
nor U15208 ( new_g21046_, n5542, n5543 );
nor U15209 ( n5542, g2802, n605 );
nor U15210 ( n5543, n570, n5521 );
nor U15211 ( new_g21028_, n5572, n5573 );
nor U15212 ( n5572, g2804, n603 );
nor U15213 ( n5573, n570, n3333 );
nor U15214 ( new_g22284_, n603, n5103 );
nor U15215 ( n5103, n4367, g2813 );
nor U15216 ( new_g22267_, n484, n5106 );
nor U15217 ( n5106, n4410, g2119 );
nor U15218 ( new_g22247_, n376, n5109 );
nor U15219 ( n5109, n4453, g1425 );
nor U15220 ( new_g22231_, n267, n5112 );
nor U15221 ( n5112, n4502, g739 );
nor U15222 ( new_g22299_, n605, n5102 );
nor U15223 ( n5102, n4364, g2811 );
nor U15224 ( new_g22280_, n486, n5104 );
nor U15225 ( n5104, n4371, g2117 );
nor U15226 ( new_g22263_, n378, n5107 );
nor U15227 ( n5107, n4414, g1423 );
nor U15228 ( new_g22242_, n269, n5110 );
nor U15229 ( n5110, n4457, g737 );
nor U15230 ( new_g20948_, n5706, n5707 );
nor U15231 ( n5706, g732, n259 );
nor U15232 ( n5707, n224, n5708 );
nor U15233 ( new_g20992_, n5639, n5640 );
nor U15234 ( n5639, g731, n269 );
nor U15235 ( n5640, n224, n5641 );
nor U15236 ( new_g20970_, n5673, n5674 );
nor U15237 ( n5673, g733, n267 );
nor U15238 ( n5674, n224, n2828 );
nor U15239 ( new_g20980_, n5654, n5655 );
nor U15240 ( n5654, g2109, n476 );
nor U15241 ( n5655, n455, n5619 );
nor U15242 ( new_g21022_, n5582, n5583 );
nor U15243 ( n5582, g2108, n486 );
nor U15244 ( n5583, n455, n5552 );
nor U15245 ( new_g21002_, n5620, n5621 );
nor U15246 ( n5620, g2110, n484 );
nor U15247 ( n5621, n455, n2818 );
nor U15248 ( new_g20976_, n5662, n5663 );
nor U15249 ( n5662, g1418, n368 );
nor U15250 ( n5663, n343, n5664 );
nor U15251 ( new_g21018_, n5591, n5592 );
nor U15252 ( n5591, g1417, n378 );
nor U15253 ( n5592, n343, n5594 );
nor U15254 ( new_g20997_, n5629, n5630 );
nor U15255 ( n5629, g1419, n376 );
nor U15256 ( n5630, n343, n2823 );
nor U15257 ( new_g21029_, n5569, n5570 );
nor U15258 ( n5569, g2806, n594 );
nor U15259 ( n5570, n567, n5571 );
nor U15260 ( new_g21063_, n5519, n5520 );
nor U15261 ( n5519, g2805, n605 );
nor U15262 ( n5520, n567, n5521 );
nor U15263 ( new_g21047_, n5540, n5541 );
nor U15264 ( n5540, g2807, n603 );
nor U15265 ( n5541, n567, n3333 );
nand U15266 ( new_g21842_, n5479, n5480 );
nand U15267 ( n5479, g554, n7169 );
nand U15268 ( n5480, g550, n2272 );
nand U15269 ( new_g21843_, n5477, n5478 );
nand U15270 ( n5477, g1240, n7167 );
nand U15271 ( n5478, g1236, n2272 );
nand U15272 ( new_g21845_, n5475, n5476 );
nand U15273 ( n5475, g1934, n7168 );
nand U15274 ( n5476, g1930, n2272 );
nand U15275 ( new_g21847_, n5472, n5473 );
nand U15276 ( n5472, g2628, n7179 );
nand U15277 ( n5473, g2624, n2272 );
nor U15278 ( new_g22269_, n594, n5105 );
nor U15279 ( n5105, n4407, g2812 );
nor U15280 ( new_g22249_, n476, n5108 );
nor U15281 ( n5108, n4450, g2118 );
nor U15282 ( new_g22234_, n368, n5111 );
nor U15283 ( n5111, n4499, g1424 );
nor U15284 ( new_g22218_, n259, n5113 );
nor U15285 ( n5113, n4538, g738 );
nor U15286 ( new_g21003_, n5617, n5618 );
nor U15287 ( n5617, g2112, n476 );
nor U15288 ( n5618, n452, n5619 );
nor U15289 ( new_g21042_, n5550, n5551 );
nor U15290 ( n5550, g2111, n486 );
nor U15291 ( n5551, n452, n5552 );
nor U15292 ( new_g21023_, n5580, n5581 );
nor U15293 ( n5580, g2113, n484 );
nor U15294 ( n5581, n452, n2818 );
nor U15295 ( n4507, g729, n7170 );
nor U15296 ( n4376, g2803, n7163 );
nor U15297 ( n4419, g2109, n7164 );
nor U15298 ( n4468, g1415, n7165 );
nor U15299 ( new_g22076_, n5333, n5334 );
nor U15300 ( n5334, n7128, n5116 );
nor U15301 ( n5333, g2217, n520 );
nor U15302 ( new_g22097_, n5301, n5302 );
nor U15303 ( n5302, n7132, n5116 );
nor U15304 ( n5301, g2220, n520 );
nor U15305 ( new_g22115_, n5265, n5266 );
nor U15306 ( n5266, n7092, n5116 );
nor U15307 ( n5265, g2223, n520 );
nor U15308 ( new_g22138_, n5228, n5229 );
nor U15309 ( n5229, n7149, n5116 );
nor U15310 ( n5228, g2226, n520 );
nor U15311 ( new_g22153_, n5191, n5192 );
nor U15312 ( n5192, n7144, n5116 );
nor U15313 ( n5191, g2229, n520 );
nor U15314 ( new_g22171_, n5156, n5158 );
nor U15315 ( n5158, n7142, n5116 );
nor U15316 ( n5156, g2232, n520 );
nor U15317 ( new_g22192_, n5122, n5123 );
nor U15318 ( n5123, n7130, n5116 );
nor U15319 ( n5122, g2205, n520 );
nor U15320 ( new_g22200_, n5114, n5115 );
nor U15321 ( n5115, n7124, n5116 );
nor U15322 ( n5114, g2208, n520 );
nor U15323 ( new_g22057_, n5364, n5365 );
nor U15324 ( n5365, n7129, n5126 );
nor U15325 ( n5364, g1523, n410 );
nor U15326 ( new_g22073_, n5340, n5341 );
nor U15327 ( n5341, n7133, n5126 );
nor U15328 ( n5340, g1526, n410 );
nor U15329 ( new_g22090_, n5308, n5309 );
nor U15330 ( n5309, n7093, n5126 );
nor U15331 ( n5308, g1529, n410 );
nor U15332 ( new_g22112_, n5271, n5272 );
nor U15333 ( n5272, n7150, n5126 );
nor U15334 ( n5271, g1532, n410 );
nor U15335 ( new_g22130_, n5238, n5239 );
nor U15336 ( n5239, n7145, n5126 );
nor U15337 ( n5238, g1535, n410 );
nor U15338 ( new_g22150_, n5203, n5204 );
nor U15339 ( n5204, n7143, n5126 );
nor U15340 ( n5203, g1538, n410 );
nor U15341 ( new_g22178_, n5142, n5143 );
nor U15342 ( n5143, n7131, n5126 );
nor U15343 ( n5142, g1511, n410 );
nor U15344 ( new_g22191_, n5124, n5125 );
nor U15345 ( n5125, n7125, n5126 );
nor U15346 ( n5124, g1514, n410 );
nor U15347 ( new_g22040_, n5391, n5392 );
nor U15348 ( n5392, n7134, n5146 );
nor U15349 ( n5391, g829, n301 );
nor U15350 ( new_g22054_, n5371, n5372 );
nor U15351 ( n5372, n7140, n5146 );
nor U15352 ( n5371, g832, n301 );
nor U15353 ( new_g22066_, n5346, n5347 );
nor U15354 ( n5347, n7095, n5146 );
nor U15355 ( n5346, g835, n301 );
nor U15356 ( new_g22087_, n5315, n5316 );
nor U15357 ( n5316, n7153, n5146 );
nor U15358 ( n5315, g838, n301 );
nor U15359 ( new_g22104_, n5281, n5282 );
nor U15360 ( n5282, n7151, n5146 );
nor U15361 ( n5281, g841, n301 );
nor U15362 ( new_g22127_, n5248, n5249 );
nor U15363 ( n5249, n7146, n5146 );
nor U15364 ( n5248, g844, n301 );
nor U15365 ( new_g22162_, n5177, n5178 );
nor U15366 ( n5178, n7137, n5146 );
nor U15367 ( n5177, g817, n301 );
nor U15368 ( new_g22177_, n5144, n5145 );
nor U15369 ( n5145, n7126, n5146 );
nor U15370 ( n5144, g820, n301 );
nor U15371 ( new_g22030_, n5413, n5414 );
nor U15372 ( n5414, n7136, n5181 );
nor U15373 ( n5413, g141, n180 );
nor U15374 ( new_g22037_, n5399, n5400 );
nor U15375 ( n5400, n7141, n5181 );
nor U15376 ( n5399, g144, n180 );
nor U15377 ( new_g22047_, n5378, n5379 );
nor U15378 ( n5379, n7096, n5181 );
nor U15379 ( n5378, g147, n180 );
nor U15380 ( new_g22063_, n5353, n5354 );
nor U15381 ( n5354, n7154, n5181 );
nor U15382 ( n5353, g150, n180 );
nor U15383 ( new_g22079_, n5326, n5327 );
nor U15384 ( n5327, n7152, n5181 );
nor U15385 ( n5326, g153, n180 );
nor U15386 ( new_g22101_, n5292, n5293 );
nor U15387 ( n5293, n7147, n5181 );
nor U15388 ( n5292, g156, n180 );
nor U15389 ( new_g22141_, n5222, n5223 );
nor U15390 ( n5223, n7138, n5181 );
nor U15391 ( n5222, g129, n180 );
nor U15392 ( new_g22161_, n5179, n5180 );
nor U15393 ( n5180, n7127, n5181 );
nor U15394 ( n5179, g132, n180 );
nor U15395 ( new_g24473_, n4827, n3509 );
xor U15396 ( n4827, n5, g2892 );
nor U15397 ( new_g23136_, n5005, n5006 );
nor U15398 ( n5005, g633, n5007 );
nand U15399 ( n5006, n4849, n2828 );
nor U15400 ( new_g21969_, n5457, n5458 );
nor U15401 ( n5457, g1319, n5459 );
nand U15402 ( n5458, n4845, n2823 );
nor U15403 ( new_g21972_, n5445, n5446 );
nor U15404 ( n5445, g2013, n5448 );
nand U15405 ( n5446, n4841, n2818 );
nor U15406 ( new_g21974_, n5441, n5442 );
nor U15407 ( n5441, g2707, n5443 );
nand U15408 ( n5442, n4837, n3333 );
nand U15409 ( new_g23047_, n5053, n5054 );
nand U15410 ( n5053, g2559, n7262 );
nand U15411 ( n5054, g8167, n545 );
nand U15412 ( new_g23132_, n5011, n5012 );
nand U15413 ( n5011, g2555, n7263 );
nand U15414 ( n5012, g8087, n545 );
nand U15415 ( new_g23014_, n5061, n5062 );
nand U15416 ( n5061, g1171, n7264 );
nand U15417 ( n5062, g8007, n323 );
nand U15418 ( new_g23110_, n5025, n5026 );
nand U15419 ( n5025, g1167, n7265 );
nand U15420 ( n5026, g7961, n323 );
nand U15421 ( new_g23076_, n5043, n5044 );
nand U15422 ( n5043, g2539, n7271 );
nand U15423 ( n5044, g2560, n545 );
nand U15424 ( new_g23039_, n5055, n5056 );
nand U15425 ( n5055, g1151, n7270 );
nand U15426 ( n5056, g1172, n323 );
xnor U15427 ( n5471, n6018, n6019 );
xor U15428 ( n6018, n6022, n6023 );
xor U15429 ( n6019, n6020, n6021 );
xnor U15430 ( n6022, g2874, g2963 );
xor U15431 ( n6020, g2981, g2978 );
xor U15432 ( n6021, g2975, g2972 );
nand U15433 ( new_g23030_, n5057, n5058 );
nand U15434 ( n5057, g1865, n7266 );
nand U15435 ( n5058, g8082, n432 );
nand U15436 ( new_g23123_, n5017, n5018 );
nand U15437 ( n5017, g1861, n7267 );
nand U15438 ( n5018, g8012, n432 );
nand U15439 ( new_g23000_, n5063, n5064 );
nand U15440 ( n5063, g484, n7268 );
nand U15441 ( n5064, g7956, n202 );
nand U15442 ( new_g23092_, n5035, n5036 );
nand U15443 ( n5035, g480, n7269 );
nand U15444 ( n5036, g7909, n202 );
nand U15445 ( new_g23058_, n5051, n5052 );
nand U15446 ( n5051, g1845, n7272 );
nand U15447 ( n5052, g1866, n432 );
nand U15448 ( new_g23022_, n5059, n5060 );
nand U15449 ( n5059, g464, n7273 );
nand U15450 ( n5060, g485, n202 );
xnor U15451 ( n5810, n6012, n6013 );
xor U15452 ( n6012, n6016, n6017 );
xor U15453 ( n6013, n6014, n6015 );
xnor U15454 ( n6016, g2935, g2938 );
xor U15455 ( n6014, g2959, g2956 );
xor U15456 ( n6015, g2953, g2947 );
xor U15457 ( n6023, g2969, g2966 );
xor U15458 ( n6017, g2944, g2941 );
nor U15459 ( new_g22026_, n5421, n3509 );
xor U15460 ( n5421, n4994, g2888 );
nor U15461 ( new_g13143_, n6056, n6057 );
nor U15462 ( n6056, g2539, n7160 );
nand U15463 ( n6057, n6058, n6059 );
or U15464 ( n6058, n7161, g2555 );
nor U15465 ( new_g13175_, n6032, n6033 );
nor U15466 ( n6032, g2554, n7160 );
nand U15467 ( n6033, n6034, n6035 );
or U15468 ( n6034, n7161, g2552 );
nor U15469 ( new_g13194_, n6024, n6025 );
nor U15470 ( n6024, g2563, n7160 );
nand U15471 ( n6025, n6026, n6027 );
or U15472 ( n6026, n7161, g2561 );
nor U15473 ( new_g13135_, n6060, n6061 );
nor U15474 ( n6060, g1845, n7155 );
nand U15475 ( n6061, n6062, n6063 );
or U15476 ( n6062, n7158, g1861 );
nor U15477 ( new_g13164_, n6040, n6041 );
nor U15478 ( n6040, g1860, n7155 );
nand U15479 ( n6041, n6042, n6043 );
or U15480 ( n6042, n7158, g1858 );
nor U15481 ( new_g13182_, n6028, n6029 );
nor U15482 ( n6028, g1869, n7155 );
nand U15483 ( n6029, n6030, n6031 );
or U15484 ( n6030, n7158, g1867 );
nor U15485 ( new_g13124_, n6064, n6065 );
nor U15486 ( n6064, g1151, n7122 );
nand U15487 ( n6065, n6066, n6067 );
or U15488 ( n6066, n7159, g1167 );
nor U15489 ( new_g13155_, n6048, n6049 );
nor U15490 ( n6048, g1166, n7122 );
nand U15491 ( n6049, n6050, n6051 );
or U15492 ( n6050, n7159, g1164 );
nor U15493 ( new_g13171_, n6036, n6037 );
nor U15494 ( n6036, g1175, n7122 );
nand U15495 ( n6037, n6038, n6039 );
or U15496 ( n6038, n7159, g1173 );
nor U15497 ( new_g13111_, n6068, n6069 );
nor U15498 ( n6068, g464, n7162 );
nand U15499 ( n6069, n6070, n6071 );
or U15500 ( n6070, n7171, g480 );
nor U15501 ( new_g13149_, n6052, n6053 );
nor U15502 ( n6052, g479, n7162 );
nand U15503 ( n6053, n6054, n6055 );
or U15504 ( n6054, n7171, g477 );
nor U15505 ( new_g13160_, n6044, n6045 );
nor U15506 ( n6044, g488, n7162 );
nand U15507 ( n6045, n6046, n6047 );
or U15508 ( n6046, n7171, g486 );
or U15509 ( n6059, n7179, g2559 );
or U15510 ( n6035, n7179, g2553 );
or U15511 ( n6027, n7179, g2562 );
or U15512 ( n6063, n7168, g1865 );
or U15513 ( n6043, n7168, g1859 );
or U15514 ( n6031, n7168, g1868 );
or U15515 ( n6067, n7167, g1171 );
or U15516 ( n6051, n7167, g1165 );
or U15517 ( n6039, n7167, g1174 );
or U15518 ( n6071, n7169, g484 );
or U15519 ( n6055, n7169, g478 );
or U15520 ( n6047, n7169, g487 );
and U15521 ( n4577, n4630, n4631 );
nor U15522 ( n4631, g2195, g2190 );
nor U15523 ( n4630, n7142, n7092 );
and U15524 ( n4609, n4658, n4659 );
nor U15525 ( n4659, g1501, g1496 );
nor U15526 ( n4658, n7143, n7093 );
nand U15527 ( n2828, g6911, g630 );
nand U15528 ( n2823, g7161, g1316 );
nand U15529 ( n2818, g7357, g2010 );
nand U15530 ( n3333, g7487, g2704 );
nand U15531 ( new_g25452_, n4355, n4356 );
nand U15532 ( n4355, g3099, n7245 );
nand U15533 ( n4356, g3109, new_g21851_ );
nand U15534 ( new_g25450_, n4359, n4360 );
nand U15535 ( n4359, g3097, n7242 );
nand U15536 ( n4360, g8106, new_g21851_ );
nand U15537 ( new_g25451_, n4357, n4358 );
nand U15538 ( n4357, g3098, n7243 );
nand U15539 ( n4358, g8030, new_g21851_ );
nand U15540 ( new_g23133_, n5009, n5010 );
nand U15541 ( n5009, g2562, n7262 );
nand U15542 ( n5010, g8167, n3365 );
nand U15543 ( new_g23114_, n5021, n5022 );
nand U15544 ( n5021, g2561, n7263 );
nand U15545 ( n5022, g8087, n3365 );
nand U15546 ( new_g23111_, n5023, n5024 );
nand U15547 ( n5023, g1174, n7264 );
nand U15548 ( n5024, g8007, n3440 );
nand U15549 ( new_g23081_, n5037, n5038 );
nand U15550 ( n5037, g1173, n7265 );
nand U15551 ( n5038, g7961, n3440 );
nand U15552 ( new_g23126_, n5013, n5014 );
nand U15553 ( n5013, g1175, n7270 );
nand U15554 ( n5014, g1172, n3440 );
nand U15555 ( new_g21970_, n5450, n5451 );
nand U15556 ( n5450, g2563, n7271 );
nand U15557 ( n5451, g2560, n3365 );
and U15558 ( n4642, n4673, n4674 );
nor U15559 ( n4674, g809, g805 );
nor U15560 ( n4673, n7146, n7095 );
and U15561 ( n4670, n4681, n4682 );
nor U15562 ( n4682, g121, g117 );
nor U15563 ( n4681, n7147, n7096 );
nand U15564 ( new_g23124_, n5015, n5016 );
nand U15565 ( n5015, g1868, n7266 );
nand U15566 ( n5016, g8082, n3402 );
nand U15567 ( new_g23097_, n5027, n5028 );
nand U15568 ( n5027, g1867, n7267 );
nand U15569 ( n5028, g8012, n3402 );
nand U15570 ( new_g23093_, n5033, n5034 );
nand U15571 ( n5033, g487, n7268 );
nand U15572 ( n5034, g7956, n3478 );
nand U15573 ( new_g23067_, n5045, n5046 );
nand U15574 ( n5045, g486, n7269 );
nand U15575 ( n5046, g7909, n3478 );
nand U15576 ( new_g23137_, n5003, n5004 );
nand U15577 ( n5003, g1869, n7272 );
nand U15578 ( n5004, g1866, n3402 );
nand U15579 ( new_g23117_, n5019, n5020 );
nand U15580 ( n5019, g488, n7273 );
nand U15581 ( n5020, g485, n3478 );
xor U15582 ( new_g16132_, g2962, n5471 );
xor U15583 ( new_g16181_, g2934, n5810 );
nand U15584 ( new_g16803_, n6001, n6002 );
nand U15585 ( n6001, g3066, g2987 );
nand U15586 ( n6002, g3047, n7239 );
nand U15587 ( new_g16866_, n5979, n5980 );
nand U15588 ( n5979, g3070, g2987 );
nand U15589 ( n5980, g3051, n7239 );
nand U15590 ( new_g16851_, n5991, n5992 );
nand U15591 ( n5991, g3068, g2987 );
nand U15592 ( n5992, g3049, n7239 );
nand U15593 ( new_g16824_, n5999, n6000 );
nand U15594 ( n5999, g3062, g2987 );
nand U15595 ( n6000, g3043, n7239 );
nand U15596 ( new_g16853_, n5989, n5990 );
nand U15597 ( n5989, g3064, g2987 );
nand U15598 ( n5990, g3045, n7239 );
nand U15599 ( new_g16844_, n5995, n5996 );
nand U15600 ( n5995, g3063, g2987 );
nand U15601 ( n5996, g3044, n7239 );
nand U15602 ( new_g16835_, n5997, n5998 );
nand U15603 ( n5997, g3067, g2987 );
nand U15604 ( n5998, g3048, n7239 );
nand U15605 ( new_g16857_, n5985, n5986 );
nand U15606 ( n5985, g3069, g2987 );
nand U15607 ( n5986, g3050, n7239 );
nand U15608 ( new_g16860_, n5983, n5984 );
nand U15609 ( n5983, g3065, g2987 );
nand U15610 ( n5984, g3046, n7239 );
nand U15611 ( new_g18868_, n5885, n5886 );
nand U15612 ( n5885, g3078, g2987 );
nand U15613 ( n5886, g3060, n7239 );
nand U15614 ( new_g18804_, n5903, n5904 );
nand U15615 ( n5903, g3076, g2987 );
nand U15616 ( n5904, g3058, n7239 );
nand U15617 ( new_g18755_, n5917, n5918 );
nand U15618 ( n5917, g3075, g2987 );
nand U15619 ( n5918, g3057, n7239 );
nand U15620 ( new_g16854_, n5987, n5988 );
nand U15621 ( n5987, g3072, g2987 );
nand U15622 ( n5988, g3053, n7239 );
nand U15623 ( new_g16861_, n5981, n5982 );
nand U15624 ( n5981, g3073, g2987 );
nand U15625 ( n5982, g3055, n7239 );
nand U15626 ( new_g16845_, n5993, n5994 );
nand U15627 ( n5993, g3071, g2987 );
nand U15628 ( n5994, g3052, n7239 );
nand U15629 ( new_g16880_, n5977, n5978 );
nand U15630 ( n5977, g3074, g2987 );
nand U15631 ( n5978, g3056, n7239 );
nand U15632 ( new_g18837_, n5893, n5894 );
nand U15633 ( n5893, g3077, g2987 );
nand U15634 ( n5894, g3059, n7239 );
nand U15635 ( new_g18907_, n5875, n5876 );
nand U15636 ( n5875, g2997, g2987 );
nand U15637 ( n5876, g3061, n7239 );
nand U15638 ( new_g20314_, n5836, n5837 );
nand U15639 ( n5836, g659, n7181 );
nand U15640 ( n5837, n628, g629 );
nand U15641 ( new_g20333_, n5834, n5835 );
nand U15642 ( n5834, g1345, n7176 );
nand U15643 ( n5835, n628, g1315 );
nand U15644 ( new_g20353_, n5830, n5831 );
nand U15645 ( n5830, g2039, n7177 );
nand U15646 ( n5831, n628, g2009 );
nand U15647 ( new_g20375_, n5828, n5829 );
nand U15648 ( n5828, g2733, n7178 );
nand U15649 ( n5829, n628, g2703 );
xnor U15650 ( n6011, n7018, n7019 );
xor U15651 ( n7019, n7020, n7021 );
xor U15652 ( n7018, n7023, n7024 );
xnor U15653 ( n7020, g8275, g8274 );
xnor U15654 ( n5934, n7025, n7026 );
xor U15655 ( n7026, n7027, n7028 );
xor U15656 ( n7025, n7029, n7030 );
xnor U15657 ( n7027, g8261, g8260 );
xor U15658 ( n7024, g8271, g8270 );
xor U15659 ( n7030, g8259, g8264 );
xor U15660 ( n7089, g3083, n6011 );
xor U15661 ( n7090, g2990, n5934 );
nor U15662 ( n5440, g2924, g2917 );
nor U15663 ( n5430, g3036, g3028 );
xnor U15664 ( n7021, g8273, g8272 );
xnor U15665 ( n7028, g8266, g8265 );
nand U15666 ( new_g18678_, n5929, n5930 );
nand U15667 ( n5930, g557, n7169 );
or U15668 ( n5929, n7169, g554 );
nand U15669 ( new_g18707_, n5927, n5928 );
nand U15670 ( n5928, g1243, n7167 );
or U15671 ( n5927, n7167, g1240 );
nand U15672 ( new_g18743_, n5921, n5922 );
nand U15673 ( n5922, g1937, n7168 );
or U15674 ( n5921, n7168, g1934 );
nand U15675 ( new_g18780_, n5913, n5914 );
nand U15676 ( n5914, g2631, n7179 );
or U15677 ( n5913, n7179, g2628 );
xnor U15678 ( n7023, g8269, g8268 );
xnor U15679 ( n7029, g8263, g8262 );
nand U15680 ( new_g18726_, n5923, n5924 );
nand U15681 ( n5923, g557, g550 );
nand U15682 ( n5924, g510, n7169 );
nand U15683 ( new_g18763_, n5915, n5916 );
nand U15684 ( n5915, g1243, g1236 );
nand U15685 ( n5916, g1196, n7167 );
nand U15686 ( new_g18794_, n5907, n5908 );
nand U15687 ( n5907, g1937, g1930 );
nand U15688 ( n5908, g1890, n7168 );
nand U15689 ( new_g18820_, n5901, n5902 );
nand U15690 ( n5901, g2631, g2624 );
nand U15691 ( n5902, g2584, n7179 );
nand U15692 ( n5641, g629, g630 );
nand U15693 ( n5594, g1315, g1316 );
nand U15694 ( n5552, g2009, g2010 );
nand U15695 ( n5521, g2703, g2704 );
nand U15696 ( n5708, g6677, g630 );
nand U15697 ( n5664, g6979, g1316 );
nand U15698 ( n5619, g7229, g2010 );
nand U15699 ( n5571, g7425, g2704 );
nand U15700 ( new_g17229_, n5965, n5966 );
nand U15701 ( n5965, g8106, g499 );
nand U15702 ( n5966, g3155, n7242 );
nand U15703 ( new_g17247_, n5955, n5956 );
nand U15704 ( n5955, g8030, g499 );
nand U15705 ( n5956, g3158, n7243 );
nand U15706 ( new_g18669_, n5931, n5932 );
nand U15707 ( n5931, g559, g8106 );
nand U15708 ( n5932, g3210, n7242 );
nand U15709 ( new_g18719_, n5925, n5926 );
nand U15710 ( n5925, g559, g8030 );
nand U15711 ( n5926, g3211, n7243 );
nand U15712 ( new_g17236_, n5959, n5960 );
nand U15713 ( n5960, g8106, g1186 );
nand U15714 ( n5959, g3164, n7242 );
nand U15715 ( new_g17248_, n5953, n5954 );
nand U15716 ( n5954, g8106, g1880 );
nand U15717 ( n5953, g3173, n7242 );
nand U15718 ( new_g17271_, n5947, n5948 );
nand U15719 ( n5948, g8106, g2574 );
nand U15720 ( n5947, g3182, n7242 );
nand U15721 ( new_g17270_, n5949, n5950 );
nand U15722 ( n5950, g8030, g1186 );
nand U15723 ( n5949, g3167, n7243 );
nand U15724 ( new_g17303_, n5943, n5944 );
nand U15725 ( n5944, g8030, g1880 );
nand U15726 ( n5943, g3176, n7243 );
nand U15727 ( new_g17341_, n5939, n5940 );
nand U15728 ( n5940, g8030, g2574 );
nand U15729 ( n5939, g3185, n7243 );
nand U15730 ( new_g17222_, n5975, n5976 );
nand U15731 ( n5976, g1245, g8106 );
nand U15732 ( n5975, g3085, n7242 );
nand U15733 ( new_g17224_, n5973, n5974 );
nand U15734 ( n5974, g1939, g8106 );
nand U15735 ( n5973, g3091, n7242 );
nand U15736 ( new_g17226_, n5969, n5970 );
nand U15737 ( n5970, g2633, g8106 );
nand U15738 ( n5969, g3094, n7242 );
nand U15739 ( new_g17225_, n5971, n5972 );
nand U15740 ( n5972, g1245, g8030 );
nand U15741 ( n5971, g3086, n7243 );
nand U15742 ( new_g17228_, n5967, n5968 );
nand U15743 ( n5968, g1939, g8030 );
nand U15744 ( n5967, g3092, n7243 );
nand U15745 ( new_g17235_, n5961, n5962 );
nand U15746 ( n5962, g2633, g8030 );
nand U15747 ( n5961, g3095, n7243 );
nand U15748 ( new_g17302_, n5945, n5946 );
nand U15749 ( n5945, g3109, g499 );
nand U15750 ( n5946, g3161, n7245 );
nand U15751 ( new_g18782_, n5909, n5910 );
nand U15752 ( n5909, g559, g3109 );
nand U15753 ( n5910, g3084, n7245 );
nand U15754 ( new_g17340_, n5941, n5942 );
nand U15755 ( n5942, g3109, g1186 );
nand U15756 ( n5941, g3170, n7245 );
nand U15757 ( new_g17383_, n5937, n5938 );
nand U15758 ( n5938, g3109, g1880 );
nand U15759 ( n5937, g3179, n7245 );
nand U15760 ( new_g17429_, n5935, n5936 );
nand U15761 ( n5936, g3109, g2574 );
nand U15762 ( n5935, g3088, n7245 );
nand U15763 ( new_g17234_, n5963, n5964 );
nand U15764 ( n5964, g1245, g3109 );
nand U15765 ( n5963, g3087, n7245 );
nand U15766 ( new_g17246_, n5957, n5958 );
nand U15767 ( n5958, g1939, g3109 );
nand U15768 ( n5957, g3093, n7245 );
nand U15769 ( new_g17269_, n5951, n5952 );
nand U15770 ( n5952, g2633, g3109 );
nand U15771 ( n5951, g3096, n7245 );
nand U15772 ( new_g16654_, n6009, n6010 );
nand U15773 ( n6010, g510, g629 );
nand U15774 ( n6009, g630, n7181 );
nand U15775 ( new_g16671_, n6007, n6008 );
nand U15776 ( n6008, g1196, g1315 );
nand U15777 ( n6007, g1316, n7176 );
nand U15778 ( new_g16692_, n6005, n6006 );
nand U15779 ( n6006, g1890, g2009 );
nand U15780 ( n6005, g2010, n7177 );
nand U15781 ( new_g16718_, n6003, n6004 );
nand U15782 ( n6004, g2584, g2703 );
nand U15783 ( n6003, g2704, n7178 );
not U15784 ( n7385, g2241 );
not U15785 ( n7386, g2241 );
not U15786 ( n7387, g2241 );
not U15787 ( n7388, n7385 );
not U15788 ( n7389, n7385 );
not U15789 ( n7390, n7385 );
not U15790 ( n7391, n7386 );
not U15791 ( n7392, n7387 );
not U15792 ( n7393, n7387 );
not U15793 ( n7394, n7387 );
not U15794 ( n7395, g1547 );
not U15795 ( n7396, g1547 );
not U15796 ( n7397, g1547 );
not U15797 ( n7398, n7395 );
not U15798 ( n7399, n7395 );
not U15799 ( n7400, n7395 );
not U15800 ( n7401, n7396 );
not U15801 ( n7402, n7397 );
not U15802 ( n7403, n7397 );
not U15803 ( n7404, n7397 );
not U15804 ( n7405, g853 );
not U15805 ( n7406, g853 );
not U15806 ( n7407, g853 );
not U15807 ( n7408, n7405 );
not U15808 ( n7409, n7405 );
not U15809 ( n7410, n7405 );
not U15810 ( n7411, n7406 );
not U15811 ( n7412, n7407 );
not U15812 ( n7413, n7407 );
not U15813 ( n7414, n7407 );
not U15814 ( n7415, g165 );
not U15815 ( n7416, g165 );
not U15816 ( n7417, g165 );
not U15817 ( n7418, n7415 );
not U15818 ( n7419, n7415 );
not U15819 ( n7420, n7415 );
not U15820 ( n7421, n7416 );
not U15821 ( n7422, n7417 );
not U15822 ( n7423, n7417 );
not U15823 ( n7424, n7417 );
endmodule

