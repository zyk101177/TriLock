module dff (clk, reset, Q, D);
input wire clk, reset, D;
output reg Q;

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      Q <= 1'b0;
    end
    else begin
      Q <= D;
    end
  end

endmodule


module s13207_ori ( clk, reset, g43, g49, g633, g634, g635, g645, g647, g648, g690,
g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757,
g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554,
g786, g1206, g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196,
g29, g22, g28, g10, g23, g37, g26, g1, g27, g42, g11, g32, g41, g31,
g45, g9, g44, g21, g30, g25, g206, g291, g372, g453, g534, g594, g785,
g1006, g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817,
g1824, g1829, g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888,
g3077, g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316,
g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663, g4664,
g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687, g5729, g6207,
g6212, g6223, g6236, g6269, g6425, g6648, g6653, g6675, g6849, g6850,
g6895, g6909, g7048, g7063, g7103, g7283, g7284, g7285, g7286, g7287,
g7288, g7289, g7290, g7291, g7292, g7293, g7294, g7295, g7298, g7423,
g7424, g7425, g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729,
g7730, g7731, g7732, g8216, g8217, g8218, g8219, g8234, g8661, g8663,
g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308,
g9310, g9312, g9314, g9378, g7763, g1205, g3856, g3857, g3854, g1193,
g1197, g1201, g6294, g6376, g1195, g6300, g6292, g6298, g6291, g6293,
g6304, g6296, g6289, g6297, g6306, g6290, g6303, g6305, g6302, g6308,
g6288, g6307, g6299, g6301, g6295 );
input clk, reset, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698,
g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781,
g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786,
g1206, g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29,
g22, g28, g10, g23, g37, g26, g1, g27, g42, g11, g32, g41, g31, g45,
g9, g44, g21, g30, g25;
output g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246,
g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871,
g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159,
g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373,
g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669,
g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269,
g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063,
g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291,
g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504,
g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216,
g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132,
g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378,
g7763, g1205, g3856, g3857, g3854, g1193, g1197, g1201, g6294, g6376,
g1195, g6300, g6292, g6298, g6291, g6293, g6304, g6296, g6289, g6297,
g6306, g6290, g6303, g6305, g6302, g6308, g6288, g6307, g6299, g6301,
g6295;
wire g49, g1000, g1008, g1554, g24, g29, g22, g28, g10, g23, g37, g26, ex_wire0, ex_wire1, ex_wire2, ex_wire3, ex_wire4, ex_wire5, ex_wire6, ex_wire7, ex_wire8, ex_wire9, ex_wire10, ex_wire11, ex_wire12, ex_wire13, ex_wire14, ex_wire15, ex_wire16, ex_wire17, ex_wire18, ex_wire19, ex_wire20, ex_wire21, ex_wire22, ex_wire23, ex_wire24, g1,
g27, g42, g11, g32, g41, g31, g9, g44, g21, g30, g25, g1313, g611, g4,
g100, new_g9354_, new_g5242_, g1158, new_g8895_, g1514, new_g6169_,
new_g9007_, g1327, g600, g628, new_g5214_, new_g6091_, new_g4264_,
new_g9000_, new_g7238_, g459, g976, g681, g162, g114, g483, g706,
new_g8897_, g1018, new_g6164_, g138, new_g4812_, g995, g1450, g597,
g759, g1499, new_g7788_, g940, new_g6577_, g83, g1211, new_g8155_,
g985, new_g6123_, g1486, new_g5201_, new_g7677_, g874, g809,
new_g5255_, g228, new_g4354_, g673, new_g6181_, g330, g1345,
new_g7825_, g297, g134, g489, new_g9387_, new_g6579_, new_g6275_,
new_g3237_, new_g9008_, new_g4878_, g775, g371, new_g7007_, g62, g560,
new_g5489_, g74, new_g5203_, g603, new_g6284_, new_g6718_, new_g8998_,
new_g9010_, new_g5234_, g390, g480, new_g6170_, g623, new_g6282_, g5,
new_g4256_, new_g7027_, g1354, g606, new_g4232_, new_g8992_,
new_g5440_, new_g6912_, g1339, new_g5220_, g1322, new_g6740_, g243,
g625, g518, new_g7029_, g1519, new_g5208_, g999, new_g8985_, g746,
g1207, new_g5256_, g321, g1325, g629, new_g5254_, new_g5563_,
new_g7086_, g1416, g685, g1013, new_g8893_, g770, g225, g86,
new_g8894_, g1351, new_g5236_, new_g4825_, new_g9006_, new_g6287_,
g110, new_g4868_, g5669, new_g8981_, new_g5657_, new_g5231_, g1226,
new_g7235_, g942, new_g5441_, new_g8978_, g8, new_g6590_, new_g5559_,
new_g8607_, g618, new_g8987_, new_g8068_, new_g7406_, g601, g945,
g6207, new_g6277_, new_g7605_, g168, g1424, g714, g1342, g626,
new_g6460_, g1462, g12, new_g8901_, new_g4263_, g45, new_g6966_,
new_g5216_, new_g5223_, g219, g48, g855, new_g5576_, new_g4284_,
g1217, new_g4349_, g1494, new_g6611_, g632, new_g8641_, new_g6273_,
new_g6445_, g1092, new_g6280_, g669, new_g8994_, g1229, g762,
new_g8980_, new_g5188_, new_g5572_, new_g4819_, g758, g324, g7505,
g614, g80, new_g8896_, new_g8976_, g1412, new_g6180_, new_g5210_,
new_g5715_, g926, new_g4364_, g767, new_g5202_, new_g7679_, g1330,
g765, new_g7242_, g1176, g1296, g1397, g452, g1360, g1504, new_g9009_,
g1300, new_g5233_, new_g9004_, g607, new_g7328_, g598, g1284, g774,
g677, g68, new_g7021_, g661, g544, g866, new_g5235_, new_g8983_,
g1304, g889, g1269, new_g6188_, new_g8989_, g584, new_g4705_,
new_g3515_, new_g5193_, g174, g612, new_g7480_, g1357, g741,
new_g7220_, new_g8902_, g1467, new_g5218_, new_g8986_, g1323,
new_g7041_, new_g5748_, g1439, g130, g1220, g859, new_g7025_, g621,
g990, new_g5624_, g1319, g8216, new_g4272_, new_g7080_, new_g5708_,
g710, new_g6585_, g237, g1097, g973, g1318, g465, new_g7033_, g222,
new_g7312_, g384, g249, g1227, new_g5222_, g828, g7507, new_g8911_,
new_g7449_, g9128, new_g7791_, new_g5560_, g1214, g1336, g1260,
new_g7697_, new_g5227_, g1224, g300, g7731, new_g7228_, new_g7031_,
g89, new_g9355_, g1392, g1400, g613, g1317, new_g5722_, new_g8899_,
g1405, g1292, g1321, g718, new_g7240_, g1333, new_g4681_, g306,
new_g9002_, new_g7177_, g318, g1435, new_g6571_, g883, g408, g825,
new_g7227_, g309, new_g7002_, g6425, g979, new_g9356_, new_g5215_,
g609, g437, new_g5211_, new_g7324_, g871, new_g9080_, g1328, g77,
new_g6735_, g1225, g333, g1148, new_g5706_, g3829, g595, g9132, g105,
g65, new_g5753_, g387, new_g5241_, g615, new_g6285_, g1329,
new_g6664_, new_g8584_, new_g8991_, g462, new_g5213_, new_g7832_,
g468, g6653, g630, g495, g610, new_g5204_, new_g9003_, g1348, g822,
g1432, g278, g1017, new_g7020_, g378, new_g8982_, g761, new_g3339_,
g1007, new_g7596_, new_g4374_, g7506, g984, new_g5195_, g764,
new_g5243_, g773, new_g4297_, new_g4317_, new_g6685_, new_g8995_,
new_g5513_, new_g8629_, new_g7128_, new_g6457_, new_g5200_,
new_g5237_, g803, new_g8801_, g202, g1443, g617, new_g7314_, g1230,
g1243, g6, g126, g944, new_g8990_, g216, g440, g471, g627, new_g5707_,
new_g8988_, new_g7030_, g887, new_g4327_, new_g8997_, new_g4840_,
new_g7271_, new_g5052_, g605, g252, g1025, new_g6739_, g959, g154,
new_g6120_, new_g3259_, new_g7783_, new_g6159_, new_g4720_, g580,
new_g5228_, g933, g356, g619, g1444, new_g5452_, new_g5711_, g7063,
g1320, new_g5672_, g760, g158, g819, g1268, new_g9358_, g1223,
new_g7197_, g402, new_g8984_, g246, g769, new_g8999_, g596,
new_g5212_, new_g5194_, g187, g290, new_g5704_, new_g7209_,
new_g5716_, new_g4879_, new_g5205_, new_g7321_, g71, new_g5475_, g772,
new_g5537_, g599, g2, new_g4837_, new_g7089_, new_g7017_, g240, g207,
new_g7087_, new_g7827_, new_g5686_, new_g6459_, new_g9338_, g1253,
new_g5538_, g1033, new_g5260_, g631, new_g8793_, new_g9005_,
new_g4688_, new_g4747_, g1324, new_g6115_, g533, g381, new_g6274_,
new_g9337_, g1272, g1021, new_g5747_, g1394, g47, new_g8900_, g540,
g275, new_g5238_, g778, g1087, new_g9357_, g95, new_g6954_, g604,
new_g8076_, g7, new_g5245_, new_g5196_, g1280, new_g7318_, new_g6165_,
new_g5545_, g1477, new_g6686_, new_g8996_, new_g4711_, g414,
new_g7782_, g768, new_g6458_, new_g5479_, g536, new_g5259_, g359,
g557, new_g4676_, g1454, g771, new_g5253_, g6212, new_g5265_, g486,
new_g5710_, new_g4299_, new_g7254_, new_g7810_, g1489, g1288, g620,
g998, g534, new_g6283_, g730, new_g8993_, g665, g327, new_g7826_,
new_g7837_, new_g7787_, new_g6949_, new_g7232_, new_g7036_, g734,
new_g5244_, new_g5230_, new_g5209_, g5687, new_g5264_, new_g3429_,
new_g4280_, g1307, new_g5751_, new_g8779_, g492, new_g5752_, g763,
new_g7217_, g766, g1267, new_g5566_, g399, new_g6286_, new_g5219_,
new_g4728_, new_g7426_, new_g6276_, new_g7415_, g1276, g602,
new_g4236_, g142, new_g9001_, new_g7008_, new_g6643_, new_g5232_,
g567, new_g7833_, g1231, new_g5698_, g303, new_g6602_, g1481, g652,
new_g7443_, g616, g1228, new_g7537_, g3, new_g5221_, new_g8979_, g521,
g405, new_g9339_, g608, new_g6262_, g411, new_g4249_, new_g5229_,
g1247, g118, new_g5217_, new_g8059_, g122, new_g6281_, g196,
new_g6951_, g1057, g591, g1126, g1114, g1149, g423, g952, g573, g264,
g579, g840, g951, g516, g846, g348, g417, g426, g1110, g429, g553,
g535, g443, g1142, g587, g117, g267, g180, g1179, g507, g377, g513,
g456, g837, g362, g342, g420, g236, g432, g498, g274, g953, g295,
g234, g834, g258, g949, g365, g141, g527, g345, g1509, g103, g281,
g1130, g1061, g255, g129, g184, g339, g212, g1106, g351, g474, g524,
g312, g1077, g570, g261, g354, g133, g843, g293, g397, g284, g108,
g183, g563, g815, g446, g233, g55, g1102, g137, g539, g395, g501,
g550, g394, g799, g1138, g232, g454, g477, g1045, g1053, g849, g588,
g214, g179, g396, g1098, g1122, g556, g270, g213, g355, g583, g852,
g1041, g435, g375, g504, g547, g313, g1134, g185, g1049, g376, g1118,
g1069, g1037, g215, g150, g316, g476, g315, g296, g950, g273, g93,
g235, g292, g510, g566, g948, g336, g121, g146, g182, g1065, g231,
g374, g436, g393, g125, g455, g458, g475, g98, g543, g517, g398, g831,
g314, g145, g478, g373, g211, g457, g181, g317, g954, g294, g113,
g479, g1379, g1378, g1376, g1377, g1374, g1373, g1371, g1372, g1030,
g1366, g1365, g1363, g1364, g1383, g1382, g1380, g1381, g1166, g1370,
g1369, g1367, g1368, g943, g1387, g1386, g1384, g1385, g972, g971,
g1263, g1257, g1415, g186, g205, g210, g195, g1513, g1266, g1408,
g1388, g1459, g1375, g875, n610, n629, n709, n794, n983, n1023, n1042,
n1092, n1122, n1300, n1374, n1566, n1585, n1669, n1768, n1822, n1860,
n2014, n2107, n2252, n2403, n2423, n2467, n2478, n2566, n2638, n2722,
n2775, n2784, n2824, n2837, n2896, n2991, n3035, n3043, n3055, n3069,
n3202, n3211, n3282, n3329, n3338, n3482, n1, n3, n4, n5, n6, n7, n8,
n12, n15, n16, n17, n18, n23, n24, n26, n27, n28, n29, n30, n31, n32,
n34, n36, n38, n39, n40, n41, n44, n45, n47, n48, n56, n58, n59, n60,
n66, n68, n69, n79, n80, n81, n82, n84, n87, n89, n95, n96, n101,
n106, n107, n108, n116, n117, n119, n121, n127, n128, n140, n141,
n156, n167, n184, n188, n189, n190, n191, n192, n193, n196, n197,
n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
n220, n221, n222, n225, n226, n227, n228, n229, n230, n231, n232,
n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
n266, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
n301, n302, n303, n306, n307, n308, n309, n310, n311, n312, n313,
n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
n336, n337, n338, n339, n340, n341, n342, n343, n346, n347, n348,
n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
n382, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n407,
n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
n443, n444, n445, n446, n447, n448, n449, n451, n452, n453, n454,
n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
n556, n557, n558, n559, n560, n561, n564, n565, n566, n567, n568,
n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
n580, n581, n582, n583, n584, n586, n587, n588, n589, n590, n591,
n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
n603, n604, n605, n606, n607, n608, n609, n611, n612, n613, n614,
n615, n616, n617, n618, n619, n620, n621, n622, n623, n625, n626,
n627, n628, n630, n631, n632, n633, n634, n635, n636, n637, n638,
n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
n672, n673, n676, n677, n678, n679, n682, n683, n684, n685, n686,
n687, n688, n689, n690, n691, n692, n693, n695, n696, n697, n698,
n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n710,
n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
n733, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
n756, n757, n758, n760, n761, n762, n763, n764, n765, n766, n767,
n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
n790, n791, n792, n793, n795, n796, n797, n798, n799, n800, n801,
n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
n879, n880, n881, n882, n883, n884, n885, n886, n889, n890, n891,
n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
n982, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1045,
n1046, n1050, n1051, n1052, n1053, n1054, n1055, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1177, n1180, n1183, n1184, n1185, n1186, n1187, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442, n1444, n1445, n1446, n1447,
n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
n1468, n1469, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
n1510, n1511, n1512, n1513, n1514, n1515, n1517, n1518, n1519, n1520,
n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
n1561, n1562, n1563, n1564, n1565, n1567, n1568, n1569, n1570, n1571,
n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
n1582, n1583, n1584, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1612, n1613,
n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1623, n1624,
n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
n1666, n1667, n1668, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
n1687, n1688, n1689, n1690, n1692, n1693, n1694, n1695, n1696, n1697,
n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, g6675, g6223,
n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1769,
n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
n1820, n1821, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
n1851, n1852;
assign g5729 = g49;
assign g6269 = g1000;
assign g6909 = g1008;
assign g5143 = g1554;
assign g6294 = g24;
assign g6300 = g29;
assign g6292 = g22;
assign g6298 = g28;
assign g6291 = g10;
assign g6293 = g23;
assign g6304 = g37;
assign g6296 = g26;
assign g6289 = g1;
assign g6297 = g27;
assign g6306 = g42;
assign g6290 = g11;
assign g6303 = g32;
assign g6305 = g41;
assign g6302 = g31;
assign g6288 = g9;
assign g6307 = g44;
assign g6299 = g21;
assign g6301 = g30;
assign g6376 = g25;
assign g6295 = g25;
assign g7291 = 1'b1;
assign g7290 = 1'b1;
assign g7504 = g5669;
assign g7295 = 1'b1;
assign g7294 = 1'b1;
assign g7284 = 1'b1;
assign g7729 = g6207;
assign g6308 = g45;
assign g7287 = 1'b1;
assign g7289 = 1'b1;
assign g5678 = g7505;
assign g7286 = 1'b1;
assign g7293 = 1'b1;
assign g6648 = g8216;
assign g5684 = g7507;
assign g9204 = g9128;
assign g7292 = 1'b1;
assign g6236 = g7731;
assign g8218 = g6425;
assign g3859 = g3829;
assign g3860 = g3829;
assign g8234 = g9132;
assign g8217 = g6653;
assign g3077 = g1017;
assign g5682 = g7506;
assign g8663 = g7063;
assign g7288 = 1'b1;
assign g7730 = g6212;
assign g372 = g534;
assign g291 = g534;
assign g594 = g534;
assign g206 = g534;
assign g453 = g534;
assign g7285 = 1'b1;
assign g7508 = g5687;
assign g7283 = 1'b1;
assign g8661 = 1'b0;
assign g8219 = g6675;
assign g7732 = g6223;

dff g183_reg ( clk, reset, g183, g10 );
dff g1012_reg ( clk, reset, n709, g43 );
dff g1014_reg ( clk, reset, n1860, n709 );
dff g186_reg ( clk, reset, g186, g1198 );
dff g959_reg ( clk, reset, g959, n1688 );
not U_inv0 ( n1781, g959 );
dff g449_reg ( clk, reset, g3159, g1206 );
not U_inv1 ( n1839, g3159 );
dff g452_reg ( clk, reset, g452, g3159 );
dff g1197_reg ( clk, reset, g1197, g1196 );
dff g1397_reg ( clk, reset, g1397, g28 );
dff g1400_reg ( clk, reset, g1400, g29 );
dff g1240_reg ( clk, reset, g1894, g1234 );
dff g530_reg ( clk, reset, g3191, g1202 );
not U_inv2 ( n1838, g3191 );
dff g533_reg ( clk, reset, g533, g3191 );
dff g1013_reg ( clk, reset, g1013, n1860 );
dff g815_reg ( clk, reset, g815, n1785 );
not U_inv3 ( n1785, g815 );
dff g819_reg ( clk, reset, g819, new_g7328_ );
dff g287_reg ( clk, reset, g3096, g1194 );
not U_inv4 ( n1840, g3096 );
dff g290_reg ( clk, reset, g290, g3096 );
dff g933_reg ( clk, reset, g933, n1690 );
dff g368_reg ( clk, reset, g3130, g1198 );
not U_inv5 ( n1841, g3130 );
dff g371_reg ( clk, reset, g371, g3130 );
dff g1236_reg ( clk, reset, g5571, g1894 );
dff g1231_reg ( clk, reset, g1231, g5571 );
not U_inv6 ( n1766, g1231 );
dff g1244_reg ( clk, reset, n2566, g1231 );
dff g1429_reg ( clk, reset, ex_wire0, g5571 );
not U_inv7 ( n1845, ex_wire0 );
dff g1394_reg ( clk, reset, g1394, g27 );
dff g942_reg ( clk, reset, g942, g941 );
dff g828_reg ( clk, reset, g828, new_g7318_ );
not U_inv8 ( n1723, g828 );
dff g822_reg ( clk, reset, g822, n1686 );
dff g825_reg ( clk, reset, g825, n1685 );
not U_inv9 ( n1698, g825 );
dff g1392_reg ( clk, reset, g1392, g26 );
dff g195_reg ( clk, reset, g195, g1194 );
dff g1199_reg ( clk, reset, n3035, g24 );
dff g1245_reg ( clk, reset, g1246, n2566 );
dff g1207_reg ( clk, reset, g1207, new_g4249_ );
not U_inv10 ( n1704, g1207 );
dff g517_reg ( clk, reset, g517, g1207 );
dff g355_reg ( clk, reset, g355, g1207 );
dff g359_reg ( clk, reset, g359, new_g5253_ );
dff g436_reg ( clk, reset, g436, g1207 );
dff g65_reg ( clk, reset, g65, g65 );
not U_inv11 ( n1699, g65 );
dff g945_reg ( clk, reset, g945, n1687 );
dff g940_reg ( clk, reset, g940, new_g4676_ );
dff g936_reg ( clk, reset, ex_wire1, new_g4349_ );
not U_inv12 ( n1722, ex_wire1 );
dff g809_reg ( clk, reset, g809, n1684 );
dff g778_reg ( clk, reset, g778, new_g7029_ );
dff g799_reg ( clk, reset, g799, new_g7321_ );
dff g803_reg ( clk, reset, g803, new_g7324_ );
dff g806_reg ( clk, reset, ex_wire2, n1683 );
not U_inv13 ( n1742, ex_wire2 );
dff g775_reg ( clk, reset, g775, new_g7314_ );
dff g812_reg ( clk, reset, ex_wire3, new_g7312_ );
not U_inv14 ( n1756, ex_wire3 );
dff g1195_reg ( clk, reset, g1195, g23 );
dff g274_reg ( clk, reset, g274, g1207 );
dff g278_reg ( clk, reset, g278, new_g5241_ );
dff g871_reg ( clk, reset, g871, n1689 );
dff g874_reg ( clk, reset, g874, n127 );
dff g440_reg ( clk, reset, g440, new_g5259_ );
dff g184_reg ( clk, reset, g184, g1 );
dff g210_reg ( clk, reset, g210, g1206 );
dff g1524_reg ( clk, reset, g1911, g37 );
dff g1513_reg ( clk, reset, g1513, g1911 );
dff g1211_reg ( clk, reset, g1211, new_g4297_ );
not U_inv15 ( n1734, g1211 );
dff g273_reg ( clk, reset, g273, g1211 );
dff g275_reg ( clk, reset, g275, new_g5233_ );
dff g354_reg ( clk, reset, g354, g1211 );
dff g356_reg ( clk, reset, g356, new_g5242_ );
dff g516_reg ( clk, reset, g516, g1211 );
dff g518_reg ( clk, reset, g518, new_g5260_ );
dff g1200_reg ( clk, reset, n1023, n3035 );
dff g1201_reg ( clk, reset, g1201, n1023 );
dff g1191_reg ( clk, reset, n2403, g22 );
dff g1192_reg ( clk, reset, n3282, n2403 );
dff g1223_reg ( clk, reset, g1223, new_g5545_ );
not U_inv16 ( n1733, g1223 );
dff g314_reg ( clk, reset, g314, g1223 );
dff g476_reg ( clk, reset, g476, g1223 );
dff g486_reg ( clk, reset, g486, new_g5232_ );
dff g233_reg ( clk, reset, g233, g1223 );
dff g243_reg ( clk, reset, g243, new_g5201_ );
dff g1254_reg ( clk, reset, g2662, new_g5559_ );
dff g1214_reg ( clk, reset, g1214, new_g4868_ );
not U_inv17 ( n1702, g1214 );
dff g398_reg ( clk, reset, g398, g1214 );
dff g317_reg ( clk, reset, g317, g1214 );
dff g333_reg ( clk, reset, g333, new_g5234_ );
dff g479_reg ( clk, reset, g479, g1214 );
dff g495_reg ( clk, reset, g495, new_g5255_ );
dff g1217_reg ( clk, reset, g1217, new_g5566_ );
not U_inv18 ( n1732, g1217 );
dff g478_reg ( clk, reset, g478, g1217 );
dff g492_reg ( clk, reset, g492, new_g5244_ );
dff g316_reg ( clk, reset, g316, g1217 );
dff g330_reg ( clk, reset, g330, new_g5228_ );
dff g235_reg ( clk, reset, g235, g1217 );
dff g249_reg ( clk, reset, g249, new_g5216_ );
dff g397_reg ( clk, reset, g397, g1217 );
dff g1220_reg ( clk, reset, g1220, new_g5537_ );
not U_inv19 ( n1744, g1220 );
dff g315_reg ( clk, reset, g315, g1220 );
dff g327_reg ( clk, reset, g327, new_g5218_ );
dff g477_reg ( clk, reset, g477, g1220 );
dff g489_reg ( clk, reset, g489, new_g5237_ );
dff g234_reg ( clk, reset, g234, g1220 );
dff g246_reg ( clk, reset, g246, new_g5209_ );
dff g396_reg ( clk, reset, g396, g1220 );
dff g408_reg ( clk, reset, g408, new_g5230_ );
dff g312_reg ( clk, reset, g312, g1225 );
dff g318_reg ( clk, reset, g318, new_g5195_ );
dff g393_reg ( clk, reset, g393, g1225 );
dff g399_reg ( clk, reset, g399, new_g5204_ );
dff g231_reg ( clk, reset, g231, g1225 );
dff g237_reg ( clk, reset, g237, new_g5188_ );
dff g474_reg ( clk, reset, g474, g1225 );
dff g480_reg ( clk, reset, g480, new_g5214_ );
dff g1224_reg ( clk, reset, g1224, new_g6115_ );
not U_inv20 ( n1703, g1224 );
dff g313_reg ( clk, reset, g313, g1224 );
dff g394_reg ( clk, reset, g394, g1224 );
dff g402_reg ( clk, reset, g402, new_g5213_ );
dff g232_reg ( clk, reset, g232, g1224 );
dff g240_reg ( clk, reset, g240, new_g5194_ );
dff g475_reg ( clk, reset, g475, g1224 );
dff g483_reg ( clk, reset, g483, new_g5222_ );
dff g1257_reg ( clk, reset, g1257, new_g4837_ );
dff g1263_reg ( clk, reset, g1263, new_g4819_ );
dff g1247_reg ( clk, reset, g1247, new_g5686_ );
not U_inv21 ( n1759, g1247 );
dff g1226_reg ( clk, reset, g1226, new_g6123_ );
not U_inv22 ( n1737, g1226 );
dff g458_reg ( clk, reset, g458, g1226 );
dff g471_reg ( clk, reset, g471, new_g5722_ );
dff g377_reg ( clk, reset, g377, g1226 );
dff g390_reg ( clk, reset, g390, new_g5715_ );
dff g296_reg ( clk, reset, g296, g1226 );
dff g309_reg ( clk, reset, g309, new_g5710_ );
dff g215_reg ( clk, reset, g215, g1226 );
dff g228_reg ( clk, reset, g228, new_g5706_ );
dff g1227_reg ( clk, reset, g1227, new_g6585_ );
not U_inv23 ( n1765, g1227 );
dff g457_reg ( clk, reset, g457, g1227 );
dff g468_reg ( clk, reset, g468, new_g5716_ );
dff g295_reg ( clk, reset, g295, g1227 );
dff g214_reg ( clk, reset, g214, g1227 );
dff g225_reg ( clk, reset, g225, new_g5704_ );
dff g1228_reg ( clk, reset, g1228, new_g6590_ );
not U_inv24 ( n1707, g1228 );
dff g294_reg ( clk, reset, g294, g1228 );
dff g303_reg ( clk, reset, g303, new_g5217_ );
dff g375_reg ( clk, reset, g375, g1228 );
dff g456_reg ( clk, reset, g456, g1228 );
dff g465_reg ( clk, reset, g465, new_g5236_ );
dff g213_reg ( clk, reset, g213, g1228 );
dff g222_reg ( clk, reset, g222, new_g5208_ );
dff g1229_reg ( clk, reset, g1229, new_g6577_ );
not U_inv25 ( n1755, g1229 );
dff g212_reg ( clk, reset, g212, g1229 );
dff g219_reg ( clk, reset, g219, new_g5200_ );
dff g374_reg ( clk, reset, g374, g1229 );
dff g455_reg ( clk, reset, g455, g1229 );
dff g293_reg ( clk, reset, g293, g1229 );
dff g1230_reg ( clk, reset, g1230, new_g7020_ );
not U_inv26 ( n1708, g1230 );
dff g454_reg ( clk, reset, g454, g1230 );
dff g292_reg ( clk, reset, g292, g1230 );
dff g297_reg ( clk, reset, g297, new_g5202_ );
dff g211_reg ( clk, reset, g211, g1230 );
dff g373_reg ( clk, reset, g373, g1230 );
dff g378_reg ( clk, reset, g378, new_g5212_ );
dff g1266_reg ( clk, reset, g1266, new_g4878_ );
dff g1269_reg ( clk, reset, g1269, new_g4879_ );
dff g1268_reg ( clk, reset, g1268, new_g4280_ );
dff g1267_reg ( clk, reset, g1267, new_g3259_ );
dff g1329_reg ( clk, reset, g1329, g1267 );
not U_inv27 ( n1770, g1329 );
dff g395_reg ( clk, reset, g395, g1223 );
dff g405_reg ( clk, reset, g405, new_g5220_ );
dff g1251_reg ( clk, reset, g8216, n68 );
not U_inv28 ( n1749, g8216 );
dff g1390_reg ( clk, reset, n3055, g8216 );
dff g1391_reg ( clk, reset, ex_wire4, n3055 );
not U_inv29 ( n1827, ex_wire4 );
dff g216_reg ( clk, reset, g216, new_g5193_ );
dff g236_reg ( clk, reset, g236, g1214 );
dff g252_reg ( clk, reset, g252, new_g5227_ );
dff g205_reg ( clk, reset, g205, g1202 );
dff g576_reg ( clk, reset, g2844, g1206 );
not U_inv30 ( n1844, g2844 );
dff g595_reg ( clk, reset, g595, g2844 );
dff g1243_reg ( clk, reset, g1243, g1894 );
dff g1431_reg ( clk, reset, ex_wire5, g1243 );
not U_inv31 ( n1847, ex_wire5 );
dff g1330_reg ( clk, reset, g1330, new_g5475_ );
not U_inv32 ( n1731, g1330 );
dff g1333_reg ( clk, reset, g1333, new_g5479_ );
not U_inv33 ( n1701, g1333 );
dff g1336_reg ( clk, reset, g1336, new_g5489_ );
dff g1339_reg ( clk, reset, g1339, new_g5513_ );
not U_inv34 ( n1735, g1339 );
dff g1342_reg ( clk, reset, g1342, new_g6091_ );
dff g1345_reg ( clk, reset, g1345, new_g7002_ );
not U_inv35 ( n1738, g1345 );
dff g1348_reg ( clk, reset, g1348, new_g7007_ );
not U_inv36 ( n1772, g1348 );
dff g1260_reg ( clk, reset, g1260, new_g5538_ );
not U_inv37 ( n1789, g1260 );
dff g1252_reg ( clk, reset, ex_wire6, g1260 );
not U_inv38 ( n1791, ex_wire6 );
dff g1430_reg ( clk, reset, ex_wire7, n1791 );
not U_inv39 ( n1848, ex_wire7 );
dff g1415_reg ( clk, reset, g1415, n56 );
dff g1412_reg ( clk, reset, g1412, new_g4840_ );
dff g1443_reg ( clk, reset, g1443, n1791 );
not U_inv40 ( n1711, g1443 );
dff g1432_reg ( clk, reset, g1432, new_g4236_ );
not U_inv41 ( g6675, g1432 );
dff g1435_reg ( clk, reset, g1435, new_g4263_ );
dff g1439_reg ( clk, reset, g1439, new_g4284_ );
dff g33_reg ( clk, reset, g7507, new_g4264_ );
dff g38_reg ( clk, reset, g5687, new_g4812_ );
not U_inv42 ( n1773, g5687 );
dff g1459_reg ( clk, reset, g1459, n1789 );
dff g1424_reg ( clk, reset, g1424, n1789 );
not U_inv43 ( n1713, g1424 );
dff g1428_reg ( clk, reset, ex_wire8, g1424 );
not U_inv44 ( n1846, ex_wire8 );
dff g1408_reg ( clk, reset, g1408, n59 );
dff g1405_reg ( clk, reset, g1405, new_g4825_ );
dff g1416_reg ( clk, reset, g1416, new_g3339_ );
not U_inv45 ( n1712, g1416 );
dff g1421_reg ( clk, reset, ex_wire9, new_g4354_ );
not U_inv46 ( n1786, ex_wire9 );
dff g1409_reg ( clk, reset, g1724, new_g4364_ );
dff g1307_reg ( clk, reset, g1307, n1789 );
not U_inv47 ( n1710, g1307 );
dff g521_reg ( clk, reset, g521, new_g5264_ );
dff g300_reg ( clk, reset, g300, new_g5210_ );
dff g376_reg ( clk, reset, g376, g1227 );
dff g387_reg ( clk, reset, g387, new_g5711_ );
dff g1193_reg ( clk, reset, g1193, n3282 );
dff g324_reg ( clk, reset, g324, new_g5211_ );
dff g321_reg ( clk, reset, g321, new_g5203_ );
dff g414_reg ( clk, reset, g414, new_g5243_ );
dff g306_reg ( clk, reset, g306, new_g5707_ );
dff g411_reg ( clk, reset, g411, new_g5235_ );
dff g1204_reg ( clk, reset, n610, g1203 );
dff g1205_reg ( clk, reset, g1205, n610 );
dff g384_reg ( clk, reset, g384, new_g5229_ );
dff g459_reg ( clk, reset, g459, new_g5221_ );
dff g381_reg ( clk, reset, g381, new_g5219_ );
dff g1351_reg ( clk, reset, g1351, new_g7008_ );
not U_inv48 ( n1748, g1351 );
dff g1354_reg ( clk, reset, g1354, new_g7197_ );
dff g1357_reg ( clk, reset, g1357, new_g7677_ );
not U_inv49 ( n1753, g1357 );
dff g435_reg ( clk, reset, g435, g1211 );
dff g437_reg ( clk, reset, g437, new_g5254_ );
dff g995_reg ( clk, reset, g995, new_g6954_ );
dff g985_reg ( clk, reset, g985, new_g6949_ );
dff g990_reg ( clk, reset, g990, new_g6951_ );
dff g462_reg ( clk, reset, g462, new_g5231_ );
dff g1360_reg ( clk, reset, g1360, new_g7679_ );
not U_inv50 ( n1771, g1360 );
dff g1450_reg ( clk, reset, g1450, new_g4272_ );
not U_inv51 ( n1754, g1450 );
dff g1444_reg ( clk, reset, g1444, new_g4256_ );
not U_inv52 ( n1779, g1444 );
dff g1454_reg ( clk, reset, g1454, new_g4299_ );
not U_inv53 ( n1709, g1454 );
dff g1461_reg ( clk, reset, g3829, new_g3429_ );
dff g1460_reg ( clk, reset, g534, new_g3237_ );
dff g1179_reg ( clk, reset, g1179, g4373 );
dff g1176_reg ( clk, reset, g1176, new_g4374_ );
dff g1081_reg ( clk, reset, g1944, new_g4747_ );
not U_inv54 ( n1776, g1944 );
dff g1156_reg ( clk, reset, n2014, g1944 );
dff g1157_reg ( clk, reset, n3069, n2014 );
dff g1159_reg ( clk, reset, n3329, n3069 );
dff g1158_reg ( clk, reset, g1158, n3329 );
not U_inv55 ( n1705, g1158 );
dff g646_reg ( clk, reset, n1669, n1705 );
dff g652_reg ( clk, reset, g652, n1669 );
not U_inv56 ( n1761, g652 );
dff g1153_reg ( clk, reset, n2784, new_g5708_ );
dff g1154_reg ( clk, reset, n3211, n2784 );
dff g1155_reg ( clk, reset, n1122, n3211 );
dff g1185_reg ( clk, reset, n2775, n1122 );
dff g1097_reg ( clk, reset, g1097, n2775 );
not U_inv57 ( n1778, g1097 );
dff g1098_reg ( clk, reset, g1098, new_g5441_ );
dff g1102_reg ( clk, reset, g1102, new_g5452_ );
dff g1106_reg ( clk, reset, g1106, new_g6602_ );
dff g1110_reg ( clk, reset, g1110, new_g7025_ );
not U_inv58 ( n1741, g1110 );
dff g1114_reg ( clk, reset, g1114, new_g7227_ );
dff g1118_reg ( clk, reset, g1118, new_g7443_ );
dff g1173_reg ( clk, reset, g7425, new_g7217_ );
dff g1170_reg ( clk, reset, g7424, g7425 );
dff g1167_reg ( clk, reset, g7423, g7424 );
dff g1166_reg ( clk, reset, g1166, g7423 );
dff g1077_reg ( clk, reset, g1077, new_g7426_ );
dff g1084_reg ( clk, reset, g2888, new_g6571_ );
not U_inv59 ( n1780, g2888 );
dff g1146_reg ( clk, reset, n1822, g2888 );
dff g1147_reg ( clk, reset, n3202, n1822 );
dff g1148_reg ( clk, reset, g1148, n3202 );
not U_inv60 ( n1750, g1148 );
dff g1122_reg ( clk, reset, g1122, new_g7697_ );
not U_inv61 ( n1769, g1122 );
dff g1126_reg ( clk, reset, g1126, new_g8155_ );
dff g1142_reg ( clk, reset, g1142, new_g8076_ );
dff g1087_reg ( clk, reset, g1087, new_g5624_ );
dff g1092_reg ( clk, reset, g1092, new_g7087_ );
not U_inv62 ( n1729, g1092 );
dff g1130_reg ( clk, reset, g1130, new_g7030_ );
not U_inv63 ( n1700, g1130 );
dff g1134_reg ( clk, reset, g1134, new_g7033_ );
dff g1138_reg ( clk, reset, g1138, new_g7036_ );
not U_inv64 ( n1820, g1138 );
dff g1149_reg ( clk, reset, g1149, new_g7041_ );
dff g1037_reg ( clk, reset, g1037, new_g6966_ );
not U_inv65 ( n1730, g1037 );
dff g1041_reg ( clk, reset, g1041, new_g7177_ );
not U_inv66 ( n1823, g1041 );
dff g1045_reg ( clk, reset, g1045, new_g7415_ );
not U_inv67 ( n1736, g1045 );
dff g1049_reg ( clk, reset, g1049, new_g7605_ );
dff g1053_reg ( clk, reset, g1053, new_g8068_ );
not U_inv68 ( n1821, g1053 );
dff g1057_reg ( clk, reset, g1057, new_g8607_ );
not U_inv69 ( n1743, g1057 );
dff g1061_reg ( clk, reset, g1061, new_g8793_ );
dff g1065_reg ( clk, reset, g1065, new_g8901_ );
not U_inv70 ( n1758, g1065 );
dff g1069_reg ( clk, reset, g1069, new_g8978_ );
dff g1073_reg ( clk, reset, g4267, new_g9080_ );
dff g1163_reg ( clk, reset, g4371, g4267 );
dff g1160_reg ( clk, reset, g4370, g4371 );
dff g1182_reg ( clk, reset, g4372, g4370 );
dff g1186_reg ( clk, reset, g4373, g4372 );
dff g71_reg ( clk, reset, g71, g3 );
not U_inv71 ( n1716, g71 );
dff g632_reg ( clk, reset, g632, g48 );
dff g766_reg ( clk, reset, g766, g48 );
dff g142_reg ( clk, reset, g142, g48 );
dff g145_reg ( clk, reset, g145, g142 );
dff g1313_reg ( clk, reset, g1313, new_g4688_ );
dff g624_reg ( clk, reset, ex_wire10, g48 );
not U_inv72 ( n1720, ex_wire10 );
dff g758_reg ( clk, reset, g758, g48 );
not U_inv73 ( n1718, g758 );
dff g774_reg ( clk, reset, g774, g48 );
dff g109_reg ( clk, reset, n1374, g48 );
dff g110_reg ( clk, reset, g110, n1374 );
dff g113_reg ( clk, reset, g113, g110 );
dff g68_reg ( clk, reset, g68, g48 );
not U_inv74 ( n1693, g68 );
dff g621_reg ( clk, reset, g621, g48 );
dff g1388_reg ( clk, reset, g1388, new_g6181_ );
dff g613_reg ( clk, reset, g613, g48 );
dff g1383_reg ( clk, reset, g1383, new_g6283_ );
dff g600_reg ( clk, reset, g600, g48 );
dff g1370_reg ( clk, reset, g1370, new_g6280_ );
dff g608_reg ( clk, reset, g608, g48 );
dff g1375_reg ( clk, reset, g1375, new_g6169_ );
dff g47_reg ( clk, reset, g47, new_g9387_ );
dff g741_reg ( clk, reset, g741, n196 );
not U_inv75 ( n1783, g741 );
dff g104_reg ( clk, reset, n1585, g3 );
dff g105_reg ( clk, reset, g105, n1585 );
dff g108_reg ( clk, reset, g108, g105 );
dff g599_reg ( clk, reset, g599, g3 );
dff g1363_reg ( clk, reset, g1363, new_g6276_ );
dff g765_reg ( clk, reset, g765, g3 );
dff g607_reg ( clk, reset, g607, g3 );
dff g1371_reg ( clk, reset, g1371, new_g6164_ );
dff g631_reg ( clk, reset, g631, g3 );
dff g620_reg ( clk, reset, g620, g3 );
dff g1384_reg ( clk, reset, g1384, new_g6170_ );
dff g773_reg ( clk, reset, g773, g3 );
dff g612_reg ( clk, reset, g612, g3 );
dff g1376_reg ( clk, reset, g1376, new_g6281_ );
dff g138_reg ( clk, reset, g138, g3 );
dff g141_reg ( clk, reset, g141, g138 );
dff g1317_reg ( clk, reset, g1317, new_g5052_ );
dff g623_reg ( clk, reset, g623, g3 );
not U_inv76 ( n1719, g623 );
dff g162_reg ( clk, reset, g162, g162 );
dff g1004_reg ( clk, reset, n2467, new_g6643_ );
dff g1005_reg ( clk, reset, n1566, n2467 );
dff g998_reg ( clk, reset, g998, n1566 );
dff g1007_reg ( clk, reset, g1007, new_g8641_ );
dff g1034_reg ( clk, reset, g6425, new_g8801_ );
not U_inv77 ( n1725, g6425 );
dff g185_reg ( clk, reset, g185, g6425 );
dff g971_reg ( clk, reset, g971, n1725 );
dff g976_reg ( clk, reset, g976, new_g7827_ );
dff g963_reg ( clk, reset, g1870, new_g7406_ );
dff g970_reg ( clk, reset, ex_wire11, g1870 );
not U_inv78 ( n1814, ex_wire11 );
dff g973_reg ( clk, reset, g973, new_g7537_ );
dff g966_reg ( clk, reset, g1871, n66 );
dff g969_reg ( clk, reset, ex_wire12, g1871 );
not U_inv79 ( n1815, ex_wire12 );
dff g984_reg ( clk, reset, g984, new_g8976_ );
dff g979_reg ( clk, reset, g979, new_g6664_ );
dff g972_reg ( clk, reset, g972, g979 );
dff g1271_reg ( clk, reset, n2478, new_g4232_ );
dff g1270_reg ( clk, reset, n1092, n2478 );
dff g172_reg ( clk, reset, ex_wire13, n1092 );
not U_inv80 ( n1849, ex_wire13 );
dff g1308_reg ( clk, reset, n983, new_g5572_ );
dff g1309_reg ( clk, reset, n2252, n983 );
dff g1310_reg ( clk, reset, n3338, n2252 );
dff g1311_reg ( clk, reset, n2824, n3338 );
dff g1312_reg ( clk, reset, n629, n2824 );
dff g1304_reg ( clk, reset, g1304, n629 );
dff g1272_reg ( clk, reset, g1272, new_g5560_ );
dff g543_reg ( clk, reset, g543, g1272 );
dff g544_reg ( clk, reset, g544, new_g5256_ );
dff g1276_reg ( clk, reset, g1276, new_g5563_ );
not U_inv81 ( n1764, g1276 );
dff g539_reg ( clk, reset, g539, g1276 );
dff g540_reg ( clk, reset, g540, new_g5245_ );
dff g1280_reg ( clk, reset, g1280, new_g6611_ );
not U_inv82 ( n1831, g1280 );
dff g535_reg ( clk, reset, g535, g1280 );
dff g536_reg ( clk, reset, g536, new_g5238_ );
dff g1284_reg ( clk, reset, g1284, new_g7017_ );
dff g587_reg ( clk, reset, g587, g1284 );
dff g560_reg ( clk, reset, g560, new_g5215_ );
dff g1292_reg ( clk, reset, g1292, new_g7021_ );
not U_inv83 ( n1746, g1292 );
dff g579_reg ( clk, reset, g579, g1292 );
dff g580_reg ( clk, reset, g580, new_g5196_ );
dff g1300_reg ( clk, reset, g1300, new_g7027_ );
dff g566_reg ( clk, reset, g566, g1300 );
dff g567_reg ( clk, reset, g567, new_g5223_ );
dff g1253_reg ( clk, reset, g1253, new_g4681_ );
dff g1250_reg ( clk, reset, g6653, new_g6579_ );
dff g1396_reg ( clk, reset, n2896, g6653 );
dff g1398_reg ( clk, reset, ex_wire14, n2896 );
not U_inv84 ( n1825, ex_wire14 );
dff g1288_reg ( clk, reset, g1288, new_g7220_ );
dff g583_reg ( clk, reset, g583, g1288 );
dff g584_reg ( clk, reset, g584, new_g5205_ );
dff g1296_reg ( clk, reset, g1296, new_g7031_ );
dff g556_reg ( clk, reset, g556, g1296 );
dff g557_reg ( clk, reset, g557, new_g5265_ );
dff g563_reg ( clk, reset, g563, new_g8899_ );
dff g625_reg ( clk, reset, g625, g8 );
dff g614_reg ( clk, reset, g614, g8 );
dff g1382_reg ( clk, reset, g1382, new_g6285_ );
dff g767_reg ( clk, reset, g767, g8 );
dff g601_reg ( clk, reset, g601, g8 );
dff g1369_reg ( clk, reset, g1369, new_g6282_ );
dff g114_reg ( clk, reset, g114, g8 );
dff g117_reg ( clk, reset, g117, g114 );
dff g759_reg ( clk, reset, g759, g8 );
dff g52_reg ( clk, reset, ex_wire15, g8 );
not U_inv85 ( n1692, ex_wire15 );
dff g948_reg ( clk, reset, g948, new_g7825_ );
dff g55_reg ( clk, reset, g55, new_g7480_ );
dff g62_reg ( clk, reset, g62, n106 );
not U_inv86 ( n1724, g62 );
dff g527_reg ( clk, reset, g527, new_g9010_ );
dff g524_reg ( clk, reset, g524, new_g9009_ );
dff g513_reg ( clk, reset, g513, new_g9003_ );
dff g510_reg ( clk, reset, g510, new_g9001_ );
dff g507_reg ( clk, reset, g507, new_g8999_ );
dff g504_reg ( clk, reset, g504, new_g8996_ );
dff g501_reg ( clk, reset, g501, new_g8992_ );
dff g118_reg ( clk, reset, g118, g7 );
dff g121_reg ( clk, reset, g121, g118 );
dff g760_reg ( clk, reset, g760, g7 );
dff g768_reg ( clk, reset, g768, g7 );
dff g86_reg ( clk, reset, g86, g7 );
dff g626_reg ( clk, reset, g626, g7 );
dff g602_reg ( clk, reset, g602, g7 );
dff g1368_reg ( clk, reset, g1368, new_g6284_ );
dff g615_reg ( clk, reset, g615, g7 );
dff g1381_reg ( clk, reset, g1381, new_g6287_ );
dff g949_reg ( clk, reset, g949, new_g7782_ );
dff g950_reg ( clk, reset, g950, new_g7787_ );
dff g951_reg ( clk, reset, g951, new_g7791_ );
dff g952_reg ( clk, reset, g952, new_g7810_ );
dff g953_reg ( clk, reset, g953, new_g7826_ );
dff g954_reg ( clk, reset, g954, new_g7783_ );
dff g943_reg ( clk, reset, g943, new_g7788_ );
dff g944_reg ( clk, reset, g944, new_g5657_ );
dff g12_reg ( clk, reset, g12, g7048 );
dff g890_reg ( clk, reset, n794, new_g6445_ );
dff g878_reg ( clk, reset, g4316, n794 );
not U_inv87 ( n1787, g4316 );
dff g926_reg ( clk, reset, g926, g4316 );
not U_inv88 ( n1763, g926 );
dff g891_reg ( clk, reset, g1783, g926 );
dff g896_reg ( clk, reset, g1829, g1783 );
dff g901_reg ( clk, reset, g1824, g1829 );
dff g906_reg ( clk, reset, g1817, g1824 );
dff g911_reg ( clk, reset, g1810, g1817 );
dff g916_reg ( clk, reset, g1804, g1810 );
dff g921_reg ( clk, reset, g1798, g1804 );
dff g883_reg ( clk, reset, g883, g1798 );
dff g852_reg ( clk, reset, g852, g883 );
dff g849_reg ( clk, reset, g849, g1798 );
dff g846_reg ( clk, reset, g846, g1804 );
dff g843_reg ( clk, reset, g843, g1810 );
dff g840_reg ( clk, reset, g840, g1817 );
dff g837_reg ( clk, reset, g837, g1824 );
dff g834_reg ( clk, reset, g834, g1829 );
dff g831_reg ( clk, reset, g831, g1783 );
dff g866_reg ( clk, reset, g866, new_g4327_ );
not U_inv89 ( n1752, g866 );
dff g863_reg ( clk, reset, ex_wire16, n1774 );
not U_inv90 ( n1696, ex_wire16 );
dff g598_reg ( clk, reset, g598, g2 );
dff g1364_reg ( clk, reset, g1364, new_g6274_ );
dff g619_reg ( clk, reset, g619, g2 );
dff g1385_reg ( clk, reset, g1385, new_g6165_ );
dff g134_reg ( clk, reset, g134, g2 );
dff g137_reg ( clk, reset, g137, g134 );
dff g1318_reg ( clk, reset, g1318, new_g6262_ );
dff g622_reg ( clk, reset, ex_wire17, g2 );
not U_inv91 ( n1721, ex_wire17 );
dff g606_reg ( clk, reset, g606, g2 );
dff g1372_reg ( clk, reset, g1372, new_g6159_ );
dff g630_reg ( clk, reset, g630, g2 );
dff g772_reg ( clk, reset, g772, g2 );
dff g74_reg ( clk, reset, g74, g2 );
not U_inv92 ( n1715, g74 );
dff g764_reg ( clk, reset, g764, g2 );
dff g99_reg ( clk, reset, n2638, g2 );
dff g100_reg ( clk, reset, g100, n2638 );
dff g103_reg ( clk, reset, g103, g100 );
dff g611_reg ( clk, reset, g611, g2 );
dff g1377_reg ( clk, reset, g1377, new_g6277_ );
dff g158_reg ( clk, reset, g158, g158 );
not U_inv93 ( n1790, g158 );
dff g199_reg ( clk, reset, n1042, n1790 );
dff g200_reg ( clk, reset, n2991, n1042 );
dff g201_reg ( clk, reset, n3482, n2991 );
dff g190_reg ( clk, reset, ex_wire18, n3482 );
not U_inv94 ( n1788, ex_wire18 );
dff g207_reg ( clk, reset, g207, new_g4728_ );
dff g182_reg ( clk, reset, g182, g207 );
dff g187_reg ( clk, reset, g187, new_g4720_ );
dff g180_reg ( clk, reset, g180, g187 );
dff g196_reg ( clk, reset, g196, new_g4711_ );
dff g179_reg ( clk, reset, g179, g196 );
dff g617_reg ( clk, reset, g617, g5 );
dff g1387_reg ( clk, reset, g1387, new_g5752_ );
dff g609_reg ( clk, reset, g609, g5 );
dff g1379_reg ( clk, reset, g1379, new_g6188_ );
dff g762_reg ( clk, reset, g762, g5 );
dff g770_reg ( clk, reset, g770, g5 );
dff g604_reg ( clk, reset, g604, g5 );
dff g1374_reg ( clk, reset, g1374, new_g5747_ );
dff g80_reg ( clk, reset, g80, g5 );
not U_inv95 ( n1714, g80 );
dff g365_reg ( clk, reset, g365, new_g9006_ );
dff g362_reg ( clk, reset, g362, new_g9005_ );
dff g351_reg ( clk, reset, g351, new_g8997_ );
dff g348_reg ( clk, reset, g348, new_g8994_ );
dff g345_reg ( clk, reset, g345, new_g8990_ );
dff g342_reg ( clk, reset, g342, new_g8986_ );
dff g339_reg ( clk, reset, g339, new_g8983_ );
dff g336_reg ( clk, reset, g336, new_g8981_ );
dff g284_reg ( clk, reset, g284, new_g9004_ );
dff g281_reg ( clk, reset, g281, new_g9002_ );
dff g270_reg ( clk, reset, g270, new_g8993_ );
dff g267_reg ( clk, reset, g267, new_g8989_ );
dff g264_reg ( clk, reset, g264, new_g8985_ );
dff g261_reg ( clk, reset, g261, new_g8982_ );
dff g258_reg ( clk, reset, g258, new_g8980_ );
dff g255_reg ( clk, reset, g255, new_g8979_ );
dff g168_reg ( clk, reset, g168, g168 );
dff g1029_reg ( clk, reset, g1017, g168 );
not U_inv96 ( n1782, g1017 );
dff g1018_reg ( clk, reset, g1018, new_g7832_ );
dff g1025_reg ( clk, reset, g1025, new_g7837_ );
dff g1021_reg ( clk, reset, g1021, new_g7833_ );
dff g1033_reg ( clk, reset, g1033, new_g8911_ );
dff g150_reg ( clk, reset, g150, g150 );
dff g603_reg ( clk, reset, g603, g6 );
dff g1367_reg ( clk, reset, g1367, new_g6286_ );
dff g83_reg ( clk, reset, g83, g6 );
dff g714_reg ( clk, reset, g714, g714 );
dff g718_reg ( clk, reset, g718, g718 );
dff g710_reg ( clk, reset, g710, g710 );
dff g685_reg ( clk, reset, g685, g685 );
dff g597_reg ( clk, reset, g597, g4 );
dff g1365_reg ( clk, reset, g1365, new_g6273_ );
dff g130_reg ( clk, reset, g130, g4 );
dff g133_reg ( clk, reset, g133, g130 );
dff g1319_reg ( clk, reset, g1319, new_g6685_ );
not U_inv97 ( n1775, g1319 );
dff g77_reg ( clk, reset, g77, g4 );
not U_inv98 ( n1717, g77 );
dff g746_reg ( clk, reset, g746, n889 );
not U_inv99 ( n1784, g746 );
dff g446_reg ( clk, reset, g446, new_g9008_ );
dff g443_reg ( clk, reset, g443, new_g9007_ );
dff g432_reg ( clk, reset, g432, new_g9000_ );
dff g429_reg ( clk, reset, g429, new_g8998_ );
dff g426_reg ( clk, reset, g426, new_g8995_ );
dff g423_reg ( clk, reset, g423, new_g8991_ );
dff g420_reg ( clk, reset, g420, new_g8987_ );
dff g417_reg ( clk, reset, g417, new_g8984_ );
dff g570_reg ( clk, reset, g570, new_g8902_ );
dff g573_reg ( clk, reset, g573, new_g8900_ );
dff g591_reg ( clk, reset, g591, new_g8897_ );
dff g588_reg ( clk, reset, g588, new_g8896_ );
dff g553_reg ( clk, reset, g553, new_g8895_ );
dff g550_reg ( clk, reset, g550, new_g8894_ );
dff g547_reg ( clk, reset, g547, new_g8893_ );
dff g859_reg ( clk, reset, g859, g859 );
not U_inv100 ( n1694, g859 );
dff g855_reg ( clk, reset, g855, g855 );
not U_inv101 ( n1695, g855 );
dff g605_reg ( clk, reset, g605, g4 );
dff g1373_reg ( clk, reset, g1373, new_g5751_ );
dff g94_reg ( clk, reset, n2423, g4 );
dff g95_reg ( clk, reset, g95, n2423 );
dff g98_reg ( clk, reset, g98, g95 );
dff g763_reg ( clk, reset, g763, g4 );
dff g610_reg ( clk, reset, g610, g4 );
dff g1378_reg ( clk, reset, g1378, new_g6275_ );
dff g771_reg ( clk, reset, g771, g4 );
dff g629_reg ( clk, reset, g629, g4 );
dff g618_reg ( clk, reset, g618, g4 );
dff g1386_reg ( clk, reset, g1386, new_g5753_ );
dff g154_reg ( clk, reset, g154, new_g7128_ );
dff g734_reg ( clk, reset, g734, g734 );
dff g673_reg ( clk, reset, g673, g673 );
dff g761_reg ( clk, reset, g761, g6 );
dff g1402_reg ( clk, reset, n3043, new_g5672_ );
dff g1403_reg ( clk, reset, n2107, n3043 );
dff g1404_reg ( clk, reset, n1300, n2107 );
dff g16_reg ( clk, reset, g7505, n1300 );
not U_inv102 ( n1829, g7505 );
dff g1393_reg ( clk, reset, n2722, g7505 );
dff g1395_reg ( clk, reset, ex_wire19, n2722 );
not U_inv103 ( n1826, ex_wire19 );
dff g769_reg ( clk, reset, g769, g6 );
dff g616_reg ( clk, reset, g616, g6 );
dff g1380_reg ( clk, reset, g1380, new_g5748_ );
dff g1389_reg ( clk, reset, g6212, new_g3515_ );
dff g627_reg ( clk, reset, g627, g6 );
dff g122_reg ( clk, reset, g122, g6 );
dff g125_reg ( clk, reset, g125, g122 );
dff g665_reg ( clk, reset, g665, g665 );
dff g628_reg ( clk, reset, g628, g5 );
dff g20_reg ( clk, reset, g7506, new_g5576_ );
dff g126_reg ( clk, reset, g126, g5 );
dff g129_reg ( clk, reset, g129, g126 );
dff g1320_reg ( clk, reset, g1320, new_g6735_ );
not U_inv104 ( n1745, g1320 );
dff g1321_reg ( clk, reset, g1321, new_g6718_ );
dff g1323_reg ( clk, reset, g1323, new_g6739_ );
dff g1322_reg ( clk, reset, g1322, new_g6686_ );
not U_inv105 ( n1762, g1322 );
dff g1324_reg ( clk, reset, g1324, new_g6740_ );
not U_inv106 ( n1740, g1324 );
dff g1325_reg ( clk, reset, g1325, new_g7086_ );
not U_inv107 ( n1777, g1325 );
dff g1326_reg ( clk, reset, ex_wire20, new_g7080_ );
not U_inv108 ( n1751, ex_wire20 );
dff g1327_reg ( clk, reset, g1327, new_g7089_ );
dff g92_reg ( clk, reset, n1768, g5 );
dff g89_reg ( clk, reset, g89, n1768 );
dff g93_reg ( clk, reset, g93, g89 );
dff g1328_reg ( clk, reset, g1328, new_g6912_ );
dff g13_reg ( clk, reset, g5669, new_g6460_ );
dff g596_reg ( clk, reset, g596, g5 );
dff g1366_reg ( clk, reset, g1366, new_g6180_ );
dff g174_reg ( clk, reset, g174, g174 );
not U_inv109 ( n1706, g174 );
dff g1486_reg ( clk, reset, g1486, new_g7254_ );
not U_inv110 ( g6223, g1486 );
dff g1481_reg ( clk, reset, g1481, new_g7271_ );
dff g1489_reg ( clk, reset, g1489, new_g7228_ );
dff g1494_reg ( clk, reset, g1494, new_g7232_ );
not U_inv111 ( n1767, g1494 );
dff g1499_reg ( clk, reset, g1499, new_g7235_ );
dff g1504_reg ( clk, reset, g1504, new_g7238_ );
not U_inv112 ( n1739, g1504 );
dff g1509_reg ( clk, reset, g1509, new_g7240_ );
dff g1514_reg ( clk, reset, g1514, new_g7242_ );
dff g1519_reg ( clk, reset, g1519, new_g7449_ );
not U_inv113 ( n1760, g1519 );
dff g1462_reg ( clk, reset, g1462, new_g7596_ );
dff g1467_reg ( clk, reset, g1467, new_g8059_ );
dff g1472_reg ( clk, reset, ex_wire21, new_g8584_ );
not U_inv114 ( n1757, ex_wire21 );
dff g1477_reg ( clk, reset, g1477, new_g8779_ );
dff g669_reg ( clk, reset, g669, g669 );
dff g730_reg ( clk, reset, g730, g730 );
dff g202_reg ( clk, reset, g202, new_g4705_ );
dff g181_reg ( clk, reset, g181, g202 );
dff g677_reg ( clk, reset, g677, g677 );
dff g888_reg ( clk, reset, g785, new_g6458_ );
not U_inv115 ( n1817, g785 );
dff g889_reg ( clk, reset, g889, new_g6459_ );
dff g887_reg ( clk, reset, g887, new_g6457_ );
not U_inv116 ( n1747, g887 );
dff g875_reg ( clk, reset, g875, new_g4317_ );
dff g661_reg ( clk, reset, g661, g661 );
dff g173_reg ( clk, reset, g6207, g6207 );
dff g498_reg ( clk, reset, g498, new_g8988_ );
dff g706_reg ( clk, reset, g706, g706 );
dff g146_reg ( clk, reset, g146, g146 );
not U_inv117 ( n1697, g146 );
dff g1030_reg ( clk, reset, g1030, new_g7209_ );
dff g1189_reg ( clk, reset, ex_wire22, new_g5698_ );
not U_inv118 ( n1828, ex_wire22 );
dff g1399_reg ( clk, reset, n2837, g7731 );
dff g1401_reg ( clk, reset, ex_wire23, n2837 );
not U_inv119 ( n1824, ex_wire23 );
dff g999_reg ( clk, reset, g999, new_g8629_ );
dff g681_reg ( clk, reset, g681, g681 );
dff g689_reg ( clk, reset, ex_wire24, new_g5440_ );
not U_inv120 ( g6895, ex_wire24 );
dff g1225_reg ( clk, reset, g1225, new_g6120_ );
dff g8_reg ( clk, reset, g8, new_g9358_ );
dff g6_reg ( clk, reset, g6, new_g9356_ );
dff g5_reg ( clk, reset, g5, new_g9355_ );
dff g7_reg ( clk, reset, g7, new_g9357_ );
dff g2_reg ( clk, reset, g2, new_g9339_ );
dff g4_reg ( clk, reset, g4, new_g9354_ );
dff g3_reg ( clk, reset, g3, new_g9338_ );
dff g48_reg ( clk, reset, g48, new_g9337_ );
nand U2043 ( n1774, n1752, n1696 );
nor U2044 ( n631, g68, g71 );
nor U2045 ( n616, n1693, g71 );
not U2046 ( n31, n373 );
not U2047 ( n29, n710 );
not U2048 ( n27, n720 );
not U2049 ( n28, n715 );
not U2050 ( n34, n644 );
not U2051 ( n23, n328 );
not U2052 ( n24, n676 );
not U2053 ( n140, n797 );
xor U2054 ( n206, new_g9337_, new_g9338_ );
xor U2055 ( n202, n203, n204 );
xor U2056 ( n203, n207, n208 );
xor U2057 ( n204, n205, n206 );
xnor U2058 ( n207, new_g9355_, new_g9356_ );
nand U2059 ( n656, n663, n664 );
nand U2060 ( n373, n651, n652 );
nor U2061 ( n652, n653, n654 );
nor U2062 ( n651, n656, n657 );
nand U2063 ( n654, n655, n645 );
xor U2064 ( n205, new_g9339_, new_g9354_ );
xor U2065 ( n208, new_g9357_, new_g9358_ );
and U2066 ( n239, n31, n321 );
not U2067 ( n39, n663 );
not U2068 ( n40, n664 );
not U2069 ( n41, n650 );
nand U2070 ( n710, n817, n106 );
nor U2071 ( n817, n119, n587 );
nand U2072 ( n720, n620, n106 );
nand U2073 ( n715, n106, n621 );
nand U2074 ( n653, n644, n648 );
nand U2075 ( n644, n1180, n590 );
not U2076 ( n47, n849 );
not U2077 ( n32, n648 );
not U2078 ( n36, n645 );
nand U2079 ( n328, n607, n608 );
nor U2080 ( n607, n622, n623 );
nor U2081 ( n608, n609, n611 );
nand U2082 ( n623, n625, n587 );
not U2083 ( n26, n219 );
nand U2084 ( n609, n618, n619 );
nor U2085 ( n618, n621, n222 );
nor U2086 ( n619, n26, n620 );
nand U2087 ( n676, n590, n632 );
nand U2088 ( n611, n612, n613 );
nor U2089 ( n612, n264, n252 );
nor U2090 ( n613, n226, n341 );
nand U2091 ( n622, n627, n628 );
and U2092 ( n627, n472, n630 );
nor U2093 ( n628, n225, n392 );
and U2094 ( n222, n615, n590 );
nor U2095 ( n625, n255, n391 );
not U2096 ( n38, n655 );
not U2097 ( n30, n630 );
not U2098 ( g7103, n936 );
nor U2099 ( n218, n587, n116 );
nor U2100 ( n215, n587, n117 );
not U2101 ( n117, n590 );
nor U2102 ( n797, n167, n141 );
nand U2103 ( n1419, n1433, n1310 );
not U2104 ( n81, n1245 );
not U2105 ( n82, n1318 );
not U2106 ( n4, g4655 );
nor U2107 ( n661, n359, n1715 );
nor U2108 ( n540, n541, n328 );
nor U2109 ( n541, n542, n543 );
nand U2110 ( n542, n564, n565 );
nand U2111 ( n543, n544, n545 );
not U2112 ( n3, new_g9387_ );
nand U2113 ( n663, n669, n670 );
and U2114 ( n670, n1717, n614 );
nor U2115 ( n669, n671, n107 );
not U2116 ( n107, n661 );
nand U2117 ( new_g9338_, n514, n515 );
nor U2118 ( n515, n516, n517 );
nor U2119 ( n514, n534, n535 );
or U2120 ( n516, n526, n527 );
nand U2121 ( n545, n321, n546 );
nand U2122 ( n546, n547, n548 );
nor U2123 ( n547, n556, n557 );
nor U2124 ( n548, n549, n550 );
nor U2125 ( n605, n606, n328 );
nor U2126 ( n606, n633, n634 );
nand U2127 ( n633, n682, n683 );
nand U2128 ( n634, n635, n636 );
nand U2129 ( new_g9337_, n576, n577 );
nor U2130 ( n577, n578, n579 );
nor U2131 ( n576, n599, n600 );
or U2132 ( n578, n591, n592 );
nand U2133 ( n636, n321, n637 );
nand U2134 ( n637, n638, n639 );
nor U2135 ( n638, n665, n666 );
nor U2136 ( n639, n640, n641 );
nand U2137 ( n664, n754, n661 );
nor U2138 ( n754, n119, n662 );
nand U2139 ( n650, n660, n661 );
nor U2140 ( n660, n116, n662 );
nand U2141 ( n657, n650, n658 );
nand U2142 ( n658, n659, n631 );
nor U2143 ( n419, n420, n328 );
nor U2144 ( n420, n421, n422 );
nand U2145 ( n421, n439, n440 );
nand U2146 ( n422, n423, n424 );
nand U2147 ( new_g9354_, n395, n396 );
and U2148 ( n396, n397, n398 );
nor U2149 ( n395, n413, n414 );
nor U2150 ( n397, n407, n408 );
nand U2151 ( n423, n321, n425 );
nand U2152 ( n425, n426, n427 );
nor U2153 ( n426, n433, n434 );
nor U2154 ( n427, n428, n429 );
nor U2155 ( n479, n480, n328 );
nor U2156 ( n480, n481, n482 );
nand U2157 ( n481, n501, n502 );
nand U2158 ( n482, n483, n484 );
nand U2159 ( new_g9339_, n452, n453 );
nor U2160 ( n453, n454, n455 );
nor U2161 ( n452, n473, n474 );
or U2162 ( n454, n464, n465 );
nand U2163 ( n484, n321, n485 );
nand U2164 ( n485, n486, n487 );
nor U2165 ( n486, n493, n494 );
nor U2166 ( n487, n488, n489 );
nand U2167 ( new_g9357_, n256, n257 );
nor U2168 ( n257, n258, n259 );
nor U2169 ( n256, n269, n270 );
nand U2170 ( n258, n265, n266 );
nand U2171 ( n274, n275, n276 );
nor U2172 ( n275, n284, n285 );
nor U2173 ( n276, n277, n278 );
nand U2174 ( n285, n286, n287 );
nor U2175 ( n358, n360, n328 );
nor U2176 ( n360, n361, n362 );
nand U2177 ( n361, n381, n382 );
nand U2178 ( n362, n363, n364 );
nand U2179 ( new_g9355_, n333, n334 );
and U2180 ( n334, n335, n336 );
nor U2181 ( n333, n352, n353 );
nor U2182 ( n335, n346, n347 );
nand U2183 ( n363, n321, n365 );
nand U2184 ( n365, n366, n367 );
nor U2185 ( n366, n374, n375 );
nor U2186 ( n367, n368, n369 );
nand U2187 ( new_g9356_, n294, n295 );
nor U2188 ( n295, n296, n297 );
nor U2189 ( n294, n306, n307 );
nand U2190 ( n296, n302, n303 );
nand U2191 ( n311, n312, n313 );
nor U2192 ( n312, n322, n323 );
nor U2193 ( n313, n314, n315 );
nand U2194 ( n323, n324, n325 );
nand U2195 ( n228, n106, n229 );
nand U2196 ( n229, n23, n230 );
nand U2197 ( n230, n231, n232 );
nor U2198 ( n231, n241, n242 );
nand U2199 ( new_g9358_, n209, n210 );
nor U2200 ( n210, n211, n212 );
nor U2201 ( n209, n227, n228 );
nand U2202 ( n211, n220, n221 );
or U2203 ( g9297, n1724, new_g9338_ );
or U2204 ( g9280, n1724, new_g9337_ );
not U2205 ( n106, n359 );
or U2206 ( g9299, n1724, new_g9339_ );
or U2207 ( g9305, n1724, new_g9354_ );
or U2208 ( g9308, n1724, new_g9355_ );
or U2209 ( g9312, n1724, new_g9357_ );
or U2210 ( g9310, n1724, new_g9356_ );
or U2211 ( g9314, n1724, new_g9358_ );
nand U2212 ( n648, n1180, n616 );
nand U2213 ( n645, n1180, n614 );
and U2214 ( n1180, n659, n1717 );
not U2215 ( n116, n616 );
nand U2216 ( n655, n893, n659 );
nor U2217 ( n893, n116, n1717 );
not U2218 ( n119, n631 );
not U2219 ( n66, n785 );
nor U2220 ( n935, g6850, n856 );
nor U2221 ( n849, new_g6664_, n66 );
nor U2222 ( n590, n1716, n1693 );
nand U2223 ( n219, n615, n631 );
and U2224 ( n615, n776, n1715 );
and U2225 ( n776, n818, n1717 );
nand U2226 ( n677, n614, n632 );
nor U2227 ( n321, n1792, n1793 );
or U2228 ( n1792, n678, n679 );
nand U2229 ( n1793, n676, n677 );
and U2230 ( n632, n698, n1715 );
and U2231 ( n226, n616, n617 );
and U2232 ( n225, n590, n617 );
and U2233 ( n380, n1180, n631 );
nand U2234 ( n587, n695, n1715 );
and U2235 ( n252, n616, n632 );
not U2236 ( n58, g9132 );
and U2237 ( n255, n626, n616 );
and U2238 ( n264, n615, n616 );
and U2239 ( n341, n614, n615 );
and U2240 ( n392, n626, n614 );
and U2241 ( n391, n626, n631 );
and U2242 ( n620, n617, n631 );
and U2243 ( n621, n614, n617 );
nand U2244 ( n472, n631, n632 );
and U2245 ( n245, n679, n590 );
nand U2246 ( n630, n626, n590 );
and U2247 ( n249, n678, n616 );
and U2248 ( n246, n679, n616 );
nand U2249 ( n505, n678, n590 );
nor U2250 ( g7514, new_g6664_, n1725 );
not U2251 ( g7298, n901 );
nand U2252 ( n936, n856, n189 );
nand U2253 ( g7474, n192, n987 );
nand U2254 ( n987, n1724, n1699 );
not U2255 ( n127, n1279 );
nor U2256 ( n971, n969, n1698 );
not U2257 ( n79, n1680 );
nand U2258 ( n828, n189, n184 );
nor U2259 ( new_g7209_, n1725, n1027 );
nand U2260 ( n1027, n58, n1697 );
not U2261 ( n5, n904 );
nand U2262 ( g4655, n5, n1621 );
not U2263 ( n190, n892 );
nor U2264 ( g4657, n1654, n1655 );
nand U2265 ( n1654, n1660, n1661 );
nand U2266 ( n1655, n1656, n1657 );
and U2267 ( n1661, n1662, n1663 );
nor U2268 ( n967, n1698, n1723 );
nand U2269 ( new_g5440_, n1448, n1449 );
nor U2270 ( n1448, n1462, n1463 );
nor U2271 ( n1449, n1450, n1451 );
nand U2272 ( n1462, n1468, n1469 );
nor U2273 ( new_g7827_, g6850, n901 );
nand U2274 ( n702, n781, n782 );
nand U2275 ( n782, n8, n783 );
not U2276 ( n8, n780 );
nor U2277 ( new_g7537_, g6850, n936 );
nand U2278 ( n1263, g5164, n1279 );
nand U2279 ( new_g6458_, n1278, n1263 );
nor U2280 ( n1278, n1280, n1281 );
nor U2281 ( n1280, n1752, n1286 );
nor U2282 ( n1281, n1282, n60 );
not U2283 ( n84, n1676 );
not U2284 ( n44, n961 );
nand U2285 ( n1683, n1670, n44 );
xnor U2286 ( n1670, n964, n1742 );
nor U2287 ( new_g7312_, n961, n977 );
nand U2288 ( n977, n978, n45 );
nand U2289 ( n978, n979, n1756 );
not U2290 ( n45, n976 );
nand U2291 ( n834, n781, n860 );
nand U2292 ( n860, n799, n783 );
not U2293 ( n7, n801 );
nor U2294 ( n926, n1748, n1123 );
nor U2295 ( n1130, n1735, n1436 );
not U2296 ( n18, n924 );
nor U2297 ( n923, n924, n1753 );
nand U2298 ( n931, n781, n959 );
nand U2299 ( n959, n875, n783 );
not U2300 ( n6, n877 );
nor U2301 ( n1114, n1755, n1235 );
nor U2302 ( n1433, n1702, n1732 );
nand U2303 ( n1245, n1310, n1311 );
nor U2304 ( n1311, n1312, n1313 );
or U2305 ( n1235, n1707, n1236 );
nor U2306 ( new_g6577_, n1241, n1242 );
nand U2307 ( n1242, n1243, n69 );
nand U2308 ( n1243, n1755, n1235 );
not U2309 ( n69, n1114 );
nor U2310 ( n1055, n1751, n1066 );
not U2311 ( n96, n1053 );
nor U2312 ( n1105, n1111, n1746 );
nor U2313 ( new_g7008_, n1759, n1120 );
nand U2314 ( n1120, n1121, n17 );
nand U2315 ( n1121, n1748, n1123 );
not U2316 ( n17, n926 );
nor U2317 ( n1310, n1734, n1704 );
nand U2318 ( new_g6590_, n1766, n1233 );
nand U2319 ( n1233, n1234, n1235 );
nand U2320 ( n1234, n1707, n1236 );
not U2321 ( n48, n1111 );
nand U2322 ( n1074, n781, n1136 );
nand U2323 ( n1136, n783, n1033 );
nand U2324 ( n1034, n1035, n1036 );
nand U2325 ( n1036, n783, n1730 );
not U2326 ( n16, n1127 );
not U2327 ( n141, n783 );
nor U2328 ( n1084, n1700, n140 );
nor U2329 ( n1318, n1425, n1733 );
or U2330 ( n1425, n1419, n1744 );
nor U2331 ( n870, n1750, n918 );
nand U2332 ( new_g6115_, n1766, n1316 );
nand U2333 ( n1316, n1317, n1315 );
nand U2334 ( n1317, n1703, n82 );
nor U2335 ( n1069, n1852, n1055 );
nand U2336 ( n934, n864, n1749 );
nor U2337 ( n881, n934, n1760 );
nand U2338 ( new_g5545_, n1766, n1423 );
nand U2339 ( n1423, n1424, n82 );
nand U2340 ( n1424, n1733, n1425 );
nor U2341 ( n1209, n1208, n1745 );
nor U2342 ( n1203, n1214, n1762 );
not U2343 ( n68, n1240 );
nand U2344 ( n986, n1002, n1003 );
nor U2345 ( n1002, n865, n1757 );
nor U2346 ( n1003, n992, n1004 );
nand U2347 ( n1004, n1005, n985 );
nor U2348 ( new_g8584_, n862, n837 );
xnor U2349 ( n862, n839, n1757 );
nor U2350 ( new_g7449_, n946, n837 );
xnor U2351 ( n946, n934, n1760 );
nor U2352 ( new_g7238_, n993, n837 );
xnor U2353 ( n993, n992, n1739 );
nor U2354 ( new_g7232_, n997, n837 );
xnor U2355 ( n997, n996, n1767 );
nor U2356 ( n976, n1756, n979 );
nor U2357 ( n1672, n964, n1742 );
nor U2358 ( n1217, n1850, n1203 );
not U2359 ( n167, n1059 );
not U2360 ( n128, n1270 );
nand U2361 ( n781, n783, n167 );
nand U2362 ( n1086, n781, n1099 );
nand U2363 ( n1099, n783, n1729 );
and U2364 ( n1062, n1770, n1066 );
nor U2365 ( n990, n992, n1739 );
nor U2366 ( new_g5513_, n1759, n1434 );
nand U2367 ( n1434, n1435, n15 );
nand U2368 ( n1435, n1735, n1436 );
not U2369 ( n15, n1130 );
nand U2370 ( new_g5537_, n1766, n1431 );
nand U2371 ( n1431, n1432, n1425 );
nand U2372 ( n1432, n1744, n1419 );
and U2373 ( n1212, n1770, n1214 );
nor U2374 ( n1013, n1750, n1026 );
not U2375 ( n87, n885 );
not U2376 ( n60, n1283 );
not U2377 ( n80, n1313 );
nor U2378 ( new_g4837_, n1704, n1590 );
nand U2379 ( n1590, n80, n1734 );
nor U2380 ( new_g4819_, n1734, n1594 );
nand U2381 ( n1594, n80, n1704 );
nand U2382 ( new_g5576_, n1397, n1398 );
nor U2383 ( n1397, n1409, n1410 );
nor U2384 ( n1398, n1399, n1400 );
nand U2385 ( n1410, n1411, n1412 );
or U2386 ( n1064, n1740, n1065 );
nor U2387 ( n1206, n1851, n1209 );
nand U2388 ( new_g5672_, n1377, n1378 );
nor U2389 ( n1377, n1387, n1388 );
nor U2390 ( n1378, n1379, n1380 );
nand U2391 ( n1388, n1389, n1390 );
not U2392 ( n89, n1342 );
not U2393 ( n1, n1347 );
not U2394 ( n121, n1359 );
not U2395 ( n108, n1352 );
nor U2396 ( new_g4317_, n1787, n1275 );
not U2397 ( n156, n1474 );
nor U2398 ( new_g4878_, n1313, n1584 );
nand U2399 ( n1584, n1704, n1734 );
and U2400 ( n1221, n1770, n1208 );
nand U2401 ( new_g5698_, n1362, n1363 );
nor U2402 ( n1362, n1370, n1371 );
nor U2403 ( n1363, n1364, n1365 );
nand U2404 ( n1370, n1375, n1376 );
nor U2405 ( n1440, n1701, n1759 );
nand U2406 ( n1634, n1733, n1703 );
nand U2407 ( new_g4280_, n1629, n1630 );
nor U2408 ( n1630, n1631, n1632 );
nor U2409 ( n1629, n1633, n1634 );
nand U2410 ( n1631, n1755, n1708 );
nand U2411 ( n1632, n1765, n1707 );
nor U2412 ( new_g3515_, n1643, n1644 );
nand U2413 ( n1643, n1649, n1650 );
nand U2414 ( n1644, n1645, n1646 );
and U2415 ( n1650, n1651, n1652 );
nand U2416 ( n1628, n1638, n1711 );
not U2417 ( n59, n1592 );
not U2418 ( n56, n1588 );
nor U2419 ( new_g3237_, n1754, n1667 );
nand U2420 ( n1667, n1779, n1709 );
nor U2421 ( new_g4354_, n1712, n1620 );
nand U2422 ( n1620, n1786, n1713 );
nand U2423 ( new_g3339_, n1713, n1666 );
nand U2424 ( n1666, n1712, n1786 );
nand U2425 ( n359, n1046, n892 );
nor U2426 ( n1046, g55, n945 );
nand U2427 ( n945, g44, n192 );
nand U2428 ( n549, n553, n554 );
nand U2429 ( n554, g647, n32 );
nor U2430 ( n553, n31, n555 );
and U2431 ( n555, n41, g524 );
nand U2432 ( n535, n536, n537 );
nor U2433 ( n537, n538, n539 );
nor U2434 ( n536, n540, n359 );
and U2435 ( n538, n27, g225 );
nand U2436 ( new_g9387_, n200, n201 );
nand U2437 ( n200, new_g7480_, n193 );
nand U2438 ( n201, n202, g44 );
not U2439 ( n193, g44 );
not U2440 ( n192, g45 );
nand U2441 ( g9378, g62, n3 );
nand U2442 ( n600, n601, n602 );
nor U2443 ( n602, n603, n604 );
nor U2444 ( n601, n605, n359 );
and U2445 ( n603, n27, g228 );
nand U2446 ( n640, n646, n647 );
nand U2447 ( n647, g648, n32 );
nor U2448 ( n646, n31, n649 );
and U2449 ( n649, n41, g527 );
nor U2450 ( n892, g42, g41 );
nand U2451 ( n428, n432, n373 );
nand U2452 ( n432, g510, n41 );
nand U2453 ( n414, n415, n416 );
nor U2454 ( n416, n417, n418 );
nor U2455 ( n415, n419, n359 );
and U2456 ( n417, n27, g219 );
nand U2457 ( n474, n475, n476 );
nor U2458 ( n476, n477, n478 );
nor U2459 ( n475, n479, n359 );
and U2460 ( n477, n27, g222 );
nand U2461 ( n488, n492, n373 );
nand U2462 ( n492, g513, n41 );
nand U2463 ( n270, n271, n106 );
and U2464 ( n271, n272, n273 );
nand U2465 ( n273, g626, n252 );
nand U2466 ( n272, n23, n274 );
nand U2467 ( n277, n281, n282 );
nand U2468 ( n282, g633, n32 );
nor U2469 ( n281, n239, n283 );
and U2470 ( n283, n41, g501 );
nand U2471 ( n368, n372, n373 );
nand U2472 ( n372, g507, n41 );
nand U2473 ( n353, n354, n355 );
nor U2474 ( n355, n356, n357 );
nor U2475 ( n354, n358, n359 );
and U2476 ( n356, n27, g216 );
nand U2477 ( n307, n308, n106 );
and U2478 ( n308, n309, n310 );
nand U2479 ( n310, g627, n252 );
nand U2480 ( n309, n23, n311 );
nand U2481 ( n314, n318, n319 );
nand U2482 ( n319, g634, n32 );
nor U2483 ( n318, n239, n320 );
and U2484 ( n320, n41, g504 );
nor U2485 ( n232, n233, n234 );
nand U2486 ( n234, n235, n236 );
nand U2487 ( n233, n237, n238 );
nand U2488 ( n236, g706, n34 );
nor U2489 ( n237, n239, n240 );
and U2490 ( n240, n41, g498 );
nand U2491 ( n557, n558, n559 );
nand U2492 ( n558, g468, n40 );
nand U2493 ( n559, g757, n39 );
nand U2494 ( n666, n667, n668 );
nand U2495 ( n667, g471, n40 );
nand U2496 ( n668, g49, n39 );
nand U2497 ( n494, n495, n496 );
nand U2498 ( n495, g465, n40 );
nand U2499 ( n496, g756, n39 );
nand U2500 ( n434, n435, n436 );
nand U2501 ( n435, g462, n40 );
nand U2502 ( n436, g753, n39 );
nand U2503 ( n375, n376, n377 );
nand U2504 ( n376, g459, n40 );
nand U2505 ( n377, g752, n39 );
nand U2506 ( n278, n279, n280 );
nand U2507 ( n280, g661, n34 );
nand U2508 ( n279, g755, n39 );
nand U2509 ( n315, n316, n317 );
nand U2510 ( n317, g665, n34 );
nand U2511 ( n316, g754, n39 );
nand U2512 ( n235, g751, n39 );
and U2513 ( n478, n29, g384 );
and U2514 ( n604, n29, g390 );
and U2515 ( n418, n29, g381 );
and U2516 ( n539, n29, g387 );
and U2517 ( n357, n29, g378 );
nand U2518 ( n473, n506, n507 );
nor U2519 ( n507, n508, n509 );
nor U2520 ( n506, n512, n513 );
and U2521 ( n508, n392, g611 );
and U2522 ( n513, n28, g303 );
nand U2523 ( n599, n688, n689 );
nor U2524 ( n689, n690, n691 );
nor U2525 ( n688, n696, n697 );
and U2526 ( n690, n392, g613 );
and U2527 ( n697, n28, g309 );
nand U2528 ( n413, n443, n444 );
nor U2529 ( n444, n445, n446 );
nor U2530 ( n443, n449, n451 );
and U2531 ( n445, n392, g610 );
and U2532 ( n451, n28, g300 );
nand U2533 ( n534, n568, n569 );
nor U2534 ( n569, n570, n571 );
nor U2535 ( n568, n574, n575 );
and U2536 ( n570, n392, g612 );
and U2537 ( n575, n28, g306 );
nand U2538 ( n352, n385, n386 );
nor U2539 ( n386, n387, n388 );
nor U2540 ( n385, n393, n394 );
and U2541 ( n387, n392, g609 );
and U2542 ( n394, n28, g297 );
nand U2543 ( n429, n430, n431 );
nand U2544 ( n430, g673, n34 );
nand U2545 ( n431, g645, n32 );
nand U2546 ( n556, n560, n561 );
nand U2547 ( n560, g741, n38 );
nand U2548 ( n561, g698, n380 );
nand U2549 ( n665, n672, n673 );
nand U2550 ( n672, g746, n38 );
nand U2551 ( n673, g694, n380 );
nand U2552 ( n433, n437, n438 );
nand U2553 ( n438, g734, n36 );
nand U2554 ( n437, g722, n380 );
nand U2555 ( n493, n497, n498 );
nand U2556 ( n498, g718, n36 );
nand U2557 ( n497, g702, n380 );
nand U2558 ( n369, n370, n371 );
nand U2559 ( n370, g669, n34 );
nand U2560 ( n371, g635, n32 );
nand U2561 ( n374, n378, n379 );
nand U2562 ( n379, g730, n36 );
nand U2563 ( n378, g723, n380 );
nand U2564 ( n197, n198, n199 );
nor U2565 ( n199, g45, g44 );
nor U2566 ( n198, n3, n190 );
nand U2567 ( n196, n1783, n197 );
nand U2568 ( n238, g690, n32 );
nand U2569 ( n662, n755, g77 );
nor U2570 ( n755, n756, n1714 );
nand U2571 ( n756, n1177, n1692 );
nor U2572 ( n1177, g86, g83 );
nand U2573 ( n671, n1252, n1253 );
and U2574 ( n1252, g83, g86 );
nor U2575 ( n1253, n1714, n1692 );
nor U2576 ( n659, n671, g74 );
nand U2577 ( n785, n935, g973 );
and U2578 ( n842, n853, n854 );
nor U2579 ( n854, new_g7406_, n855 );
nor U2580 ( n853, n856, n47 );
or U2581 ( n855, g6425, g979 );
nand U2582 ( n856, n1192, n1193 );
and U2583 ( n1193, n1194, n1195 );
nor U2584 ( n1192, g962, n1196 );
nor U2585 ( n1194, g972, g971 );
nor U2586 ( g1015, n844, n845 );
nand U2587 ( n844, g1, g162 );
nand U2588 ( n845, g1013, n842 );
nor U2589 ( g1006, n851, n852 );
nand U2590 ( n851, g43, n184 );
nand U2591 ( n852, n842, g162 );
not U2592 ( g6850, g43 );
nor U2593 ( n614, n1716, g68 );
and U2594 ( new_g6664_, n1226, g984 );
nor U2595 ( n1226, g979, g6850 );
nand U2596 ( n550, n551, n552 );
nand U2597 ( n551, g714, n36 );
nand U2598 ( n552, g681, n34 );
nand U2599 ( n641, n642, n643 );
nand U2600 ( n642, g710, n36 );
nand U2601 ( n643, g685, n34 );
nand U2602 ( n489, n490, n491 );
nand U2603 ( n490, g677, n34 );
nand U2604 ( n491, g652, n32 );
nor U2605 ( n818, n756, g80 );
nand U2606 ( g8872, g1, n843 );
or U2607 ( n843, n47, g1030 );
and U2608 ( n698, n1045, g80 );
nor U2609 ( n1045, g77, n756 );
and U2610 ( new_g7406_, n935, g976 );
and U2611 ( n617, g74, n776 );
and U2612 ( n695, g77, n818 );
nand U2613 ( g9132, n1251, g1033 );
nor U2614 ( n1251, g1017, g6850 );
nand U2615 ( g8958, g1, n847 );
nand U2616 ( n847, n848, n849 );
nor U2617 ( n848, g1030, n850 );
nor U2618 ( n850, n58, g10 );
and U2619 ( n626, n695, g74 );
nor U2620 ( n679, n662, g74 );
and U2621 ( n678, g74, n698 );
and U2622 ( n544, n1794, n1795 );
nand U2623 ( n1794, n24, g765 );
nand U2624 ( n1795, n249, g773 );
and U2625 ( n483, n1796, n1797 );
nand U2626 ( n1796, n24, g764 );
nand U2627 ( n1797, n249, g772 );
and U2628 ( n635, n1798, n1799 );
nand U2629 ( n1798, n24, g766 );
nand U2630 ( n1799, n249, g774 );
and U2631 ( n439, n1800, n1801 );
nand U2632 ( n1800, n24, g763 );
nand U2633 ( n1801, n249, g771 );
nor U2634 ( n564, n566, n567 );
nor U2635 ( n566, n505, n1694 );
and U2636 ( n567, n245, g849 );
nor U2637 ( n683, n684, n685 );
nor U2638 ( n684, n505, n1695 );
and U2639 ( n685, n245, g852 );
and U2640 ( n381, n1802, n1803 );
nand U2641 ( n1802, n24, g762 );
nand U2642 ( n1803, n249, g770 );
nor U2643 ( n501, n503, n504 );
nor U2644 ( n503, n505, n1696 );
and U2645 ( n504, n245, g846 );
nor U2646 ( n682, n686, n687 );
nor U2647 ( n687, n677, n1718 );
and U2648 ( n686, n246, g48 );
xor U2649 ( new_g7480_, n937, n938 );
xor U2650 ( n938, n939, n940 );
nand U2651 ( n937, g47, n945 );
xor U2652 ( n939, n943, n944 );
nand U2653 ( n284, n288, n289 );
nand U2654 ( n288, g768, n249 );
nand U2655 ( n289, g760, n24 );
nand U2656 ( n322, n326, n327 );
nand U2657 ( n326, g769, n249 );
nand U2658 ( n327, g761, n24 );
nand U2659 ( n424, g4, n246 );
nand U2660 ( n565, g3, n246 );
nand U2661 ( n287, g834, n245 );
nand U2662 ( n286, g7, n246 );
nand U2663 ( n440, g843, n245 );
nand U2664 ( n502, g2, n246 );
nand U2665 ( n325, g837, n245 );
nand U2666 ( n324, g6, n246 );
nand U2667 ( n241, n247, n248 );
nand U2668 ( n247, g767, n249 );
nand U2669 ( n248, g759, n24 );
nand U2670 ( n364, g5, n246 );
nand U2671 ( n382, g840, n245 );
nand U2672 ( n242, n243, n244 );
nand U2673 ( n243, g8, n246 );
nand U2674 ( n244, g831, n245 );
nand U2675 ( n521, n522, n523 );
nand U2676 ( n522, g182, n264 );
nand U2677 ( n523, g162, n26 );
nand U2678 ( n517, n518, n519 );
nor U2679 ( n518, n524, n525 );
nor U2680 ( n519, n520, n521 );
and U2681 ( n525, n255, g607 );
nand U2682 ( n583, n584, n586 );
nand U2683 ( n584, g185, n264 );
nand U2684 ( n586, g168, n26 );
nand U2685 ( n579, n580, n581 );
nor U2686 ( n580, n588, n589 );
nor U2687 ( n581, n582, n583 );
and U2688 ( n589, n255, g608 );
nand U2689 ( n459, n460, n461 );
nand U2690 ( n460, g181, n264 );
nand U2691 ( n461, n26, g158 );
nand U2692 ( n455, n456, n457 );
nor U2693 ( n456, n462, n463 );
nor U2694 ( n457, n458, n459 );
and U2695 ( n463, n255, g606 );
nand U2696 ( n571, n572, n573 );
nand U2697 ( n572, g599, n391 );
nand U2698 ( n573, g620, n30 );
nand U2699 ( n509, n510, n511 );
nand U2700 ( n510, g598, n391 );
nand U2701 ( n511, g619, n30 );
nand U2702 ( n691, n692, n693 );
nand U2703 ( n692, g600, n391 );
nand U2704 ( n693, g621, n30 );
nand U2705 ( n446, n447, n448 );
nand U2706 ( n447, g597, n391 );
nand U2707 ( n448, g618, n30 );
nand U2708 ( n526, n530, n531 );
nand U2709 ( n531, g362, n225 );
nor U2710 ( n530, n532, n533 );
nor U2711 ( n532, n472, n1719 );
and U2712 ( n533, n226, g281 );
nand U2713 ( n591, n595, n596 );
nand U2714 ( n596, g365, n225 );
nor U2715 ( n595, n597, n598 );
nor U2716 ( n597, n472, n1720 );
and U2717 ( n598, n226, g284 );
nor U2718 ( n398, n399, n400 );
nand U2719 ( n400, n401, n402 );
nand U2720 ( n399, n403, n404 );
nand U2721 ( n402, g95, n341 );
and U2722 ( n403, n1804, n1805 );
nand U2723 ( n1804, n226, g267 );
nand U2724 ( n1805, n225, g348 );
nand U2725 ( n388, n389, n390 );
nand U2726 ( n389, g596, n391 );
nand U2727 ( n390, g617, n30 );
nand U2728 ( n464, n468, n469 );
nand U2729 ( n469, g351, n225 );
nor U2730 ( n468, n470, n471 );
nor U2731 ( n470, n472, n1721 );
and U2732 ( n471, n226, g270 );
nand U2733 ( n259, n260, n261 );
nand U2734 ( n261, g420, n218 );
nor U2735 ( n260, n262, n263 );
and U2736 ( n263, g183, n264 );
and U2737 ( n262, n26, g6207 );
nand U2738 ( n901, g1, n856 );
nand U2739 ( n297, n298, n299 );
nand U2740 ( n299, g423, n218 );
nor U2741 ( n298, n300, n301 );
and U2742 ( n301, g184, n264 );
and U2743 ( n520, n218, g443 );
and U2744 ( n300, n26, g150 );
nand U2745 ( n212, n213, n214 );
nand U2746 ( n214, g563, n215 );
nor U2747 ( n213, n216, n217 );
nor U2748 ( n216, n219, n1697 );
and U2749 ( n217, n218, g417 );
nor U2750 ( n336, n337, n338 );
nand U2751 ( n338, n339, n340 );
nand U2752 ( n337, n342, n343 );
nand U2753 ( n340, g89, n341 );
and U2754 ( n342, n1806, n1807 );
nand U2755 ( n1806, n226, g264 );
nand U2756 ( n1807, n225, g345 );
nand U2757 ( n227, n250, n251 );
nand U2758 ( n251, g625, n252 );
nor U2759 ( n250, n253, n254 );
and U2760 ( n253, n255, g601 );
and U2761 ( n254, n30, g614 );
and U2762 ( n458, n218, g432 );
and U2763 ( n524, n215, g550 );
and U2764 ( n582, n218, g446 );
and U2765 ( n462, n215, g547 );
and U2766 ( n588, n215, g553 );
nand U2767 ( n401, g154, n26 );
nand U2768 ( n269, n290, n291 );
nand U2769 ( n291, g615, n30 );
nor U2770 ( n290, n292, n293 );
and U2771 ( n293, n255, g602 );
and U2772 ( n292, n215, g570 );
nand U2773 ( n306, n329, n330 );
nand U2774 ( n330, g616, n30 );
nor U2775 ( n329, n331, n332 );
and U2776 ( n332, n255, g603 );
and U2777 ( n331, n215, g588 );
nand U2778 ( n408, n409, n410 );
nand U2779 ( n409, g605, n255 );
nand U2780 ( n410, g573, n215 );
nand U2781 ( n339, g174, n26 );
nand U2782 ( n407, n411, n412 );
nand U2783 ( n412, g180, n264 );
nand U2784 ( n411, g429, n218 );
and U2785 ( n265, n1808, n1809 );
nand U2786 ( n1808, n226, g258 );
nand U2787 ( n1809, n225, g339 );
and U2788 ( n220, n1810, n1811 );
nand U2789 ( n1810, n226, g255 );
nand U2790 ( n1811, n225, g336 );
nand U2791 ( n527, n528, n529 );
nand U2792 ( n528, g105, n341 );
nand U2793 ( n529, g138, n222 );
nand U2794 ( n347, n348, n349 );
nand U2795 ( n348, g604, n255 );
nand U2796 ( n349, g591, n215 );
and U2797 ( n302, n1812, n1813 );
nand U2798 ( n1812, n226, g261 );
nand U2799 ( n1813, n225, g342 );
and U2800 ( n512, n252, g630 );
and U2801 ( n696, n252, g632 );
and U2802 ( n449, n252, g629 );
and U2803 ( n574, n252, g631 );
nand U2804 ( n346, n350, n351 );
nand U2805 ( n351, g179, n264 );
nand U2806 ( n350, g426, n218 );
nand U2807 ( n592, n593, n594 );
nand U2808 ( n593, g110, n341 );
nand U2809 ( n594, g142, n222 );
not U2810 ( n189, g1 );
nor U2811 ( n968, g786, n969 );
nand U2812 ( n465, n466, n467 );
nand U2813 ( n466, g100, n341 );
nand U2814 ( n467, g134, n222 );
nand U2815 ( g7763, n965, n966 );
nand U2816 ( n965, g786, n970 );
nand U2817 ( n966, n967, n968 );
nand U2818 ( n970, n971, g828 );
nand U2819 ( n404, g130, n222 );
and U2820 ( n393, n252, g628 );
not U2821 ( n184, g1000 );
nand U2822 ( n343, g126, n222 );
nand U2823 ( g9128, n1142, n1143 );
nand U2824 ( n1143, g32, g30 );
nand U2825 ( n1142, g31, n191 );
not U2826 ( n191, g32 );
nand U2827 ( n266, g118, n222 );
nand U2828 ( n221, g114, n222 );
nand U2829 ( n303, g122, n222 );
not U2830 ( g3856, g929 );
not U2831 ( g3857, g955 );
not U2832 ( g3854, g795 );
nor U2833 ( n1195, g1870, g1871 );
nand U2834 ( n1196, n1814, n1815 );
nand U2835 ( new_g8893_, n815, n816 );
nand U2836 ( n816, g547, n710 );
nand U2837 ( n815, g536, n29 );
nand U2838 ( new_g8894_, n813, n814 );
nand U2839 ( n814, g550, n710 );
nand U2840 ( n813, g540, n29 );
nand U2841 ( new_g8895_, n811, n812 );
nand U2842 ( n812, g553, n710 );
nand U2843 ( n811, g544, n29 );
nand U2844 ( new_g8896_, n809, n810 );
nand U2845 ( n810, g588, n710 );
nand U2846 ( n809, g580, n29 );
nand U2847 ( new_g8897_, n807, n808 );
nand U2848 ( n808, g591, n710 );
nand U2849 ( n807, g584, n29 );
nand U2850 ( new_g8900_, n803, n804 );
nand U2851 ( n804, g573, n710 );
nand U2852 ( n803, g560, n29 );
nand U2853 ( new_g8902_, n791, n792 );
nand U2854 ( n792, g570, n710 );
nand U2855 ( n791, g567, n29 );
nand U2856 ( new_g8984_, n764, n765 );
nand U2857 ( n765, g417, n710 );
nand U2858 ( n764, g399, n29 );
nand U2859 ( new_g8987_, n757, n758 );
nand U2860 ( n758, g420, n710 );
nand U2861 ( n757, g402, n29 );
nand U2862 ( new_g8991_, n746, n747 );
nand U2863 ( n747, g423, n710 );
nand U2864 ( n746, g405, n29 );
nand U2865 ( new_g8995_, n738, n739 );
nand U2866 ( n739, g426, n710 );
nand U2867 ( n738, g408, n29 );
nand U2868 ( new_g8998_, n731, n732 );
nand U2869 ( n732, g429, n710 );
nand U2870 ( n731, g411, n29 );
nand U2871 ( new_g9000_, n727, n728 );
nand U2872 ( n728, g432, n710 );
nand U2873 ( n727, g414, n29 );
nand U2874 ( new_g9007_, n711, n712 );
nand U2875 ( n712, g443, n710 );
nand U2876 ( n711, g437, n29 );
nand U2877 ( new_g9008_, n707, n708 );
nand U2878 ( n708, g446, n710 );
nand U2879 ( n707, g440, n29 );
nand U2880 ( new_g8899_, n805, n806 );
nand U2881 ( n806, g563, n710 );
nand U2882 ( n805, g557, n29 );
nand U2883 ( new_g8988_, n752, n753 );
nand U2884 ( n753, g498, n664 );
nand U2885 ( n752, g480, n40 );
nand U2886 ( new_g8992_, n744, n745 );
nand U2887 ( n745, g501, n664 );
nand U2888 ( n744, g483, n40 );
nand U2889 ( new_g8996_, n736, n737 );
nand U2890 ( n737, g504, n664 );
nand U2891 ( n736, g486, n40 );
nand U2892 ( new_g8999_, n729, n730 );
nand U2893 ( n730, g507, n664 );
nand U2894 ( n729, g489, n40 );
nand U2895 ( new_g9001_, n725, n726 );
nand U2896 ( n726, g510, n664 );
nand U2897 ( n725, g492, n40 );
nand U2898 ( new_g9003_, n721, n722 );
nand U2899 ( n722, g513, n664 );
nand U2900 ( n721, g495, n40 );
nand U2901 ( new_g9009_, n705, n706 );
nand U2902 ( n706, g524, n664 );
nand U2903 ( n705, g518, n40 );
nand U2904 ( new_g9010_, n703, n704 );
nand U2905 ( n704, g527, n664 );
nand U2906 ( n703, g521, n40 );
nor U2907 ( new_g8629_, n828, n846 );
nand U2908 ( n846, n842, g998 );
nand U2909 ( new_g8979_, n774, n775 );
nand U2910 ( n775, g255, n720 );
nand U2911 ( n774, g237, n27 );
nand U2912 ( new_g8980_, n772, n773 );
nand U2913 ( n773, g258, n720 );
nand U2914 ( n772, g240, n27 );
nand U2915 ( new_g8982_, n768, n769 );
nand U2916 ( n769, g261, n720 );
nand U2917 ( n768, g243, n27 );
nand U2918 ( new_g8985_, n762, n763 );
nand U2919 ( n763, g264, n720 );
nand U2920 ( n762, g246, n27 );
nand U2921 ( new_g8989_, n750, n751 );
nand U2922 ( n751, g267, n720 );
nand U2923 ( n750, g249, n27 );
nand U2924 ( new_g8993_, n742, n743 );
nand U2925 ( n743, g270, n720 );
nand U2926 ( n742, g252, n27 );
nand U2927 ( new_g9002_, n723, n724 );
nand U2928 ( n724, g281, n720 );
nand U2929 ( n723, g275, n27 );
nand U2930 ( new_g9004_, n718, n719 );
nand U2931 ( n719, g284, n720 );
nand U2932 ( n718, g278, n27 );
nand U2933 ( new_g8981_, n770, n771 );
nand U2934 ( n771, g336, n715 );
nand U2935 ( n770, g318, n28 );
nand U2936 ( new_g8983_, n766, n767 );
nand U2937 ( n767, g339, n715 );
nand U2938 ( n766, g321, n28 );
nand U2939 ( new_g8986_, n760, n761 );
nand U2940 ( n761, g342, n715 );
nand U2941 ( n760, g324, n28 );
nand U2942 ( new_g8990_, n748, n749 );
nand U2943 ( n749, g345, n715 );
nand U2944 ( n748, g327, n28 );
nand U2945 ( new_g8994_, n740, n741 );
nand U2946 ( n741, g348, n715 );
nand U2947 ( n740, g330, n28 );
nand U2948 ( new_g8997_, n733, n735 );
nand U2949 ( n735, g351, n715 );
nand U2950 ( n733, g333, n28 );
nand U2951 ( new_g9005_, n716, n717 );
nand U2952 ( n717, g362, n715 );
nand U2953 ( n716, g356, n28 );
nand U2954 ( new_g9006_, n713, n714 );
nand U2955 ( n714, g365, n715 );
nand U2956 ( n713, g359, n28 );
nor U2957 ( new_g8641_, n840, n841 );
nand U2958 ( n841, g1013, new_g6643_ );
nand U2959 ( n840, n825, n842 );
xor U2960 ( n940, n941, n942 );
xor U2961 ( n942, g3, g2 );
xor U2962 ( n941, g48, g4 );
xor U2963 ( n944, g6, g5 );
xor U2964 ( n943, g8, g7 );
nand U2965 ( n1279, n1668, g933 );
and U2966 ( n1668, g929, g871 );
nor U2967 ( n1269, n1271, g889 );
nor U2968 ( n1271, n127, n1272 );
nor U2969 ( n1272, n1273, g866 );
nor U2970 ( n1266, n1267, n1268 );
nor U2971 ( n1267, n1274, n1275 );
nor U2972 ( n1268, n1269, n128 );
or U2973 ( n1274, g866, g875 );
nand U2974 ( new_g6459_, n1262, n1263 );
nor U2975 ( n1262, n1264, n1265 );
nor U2976 ( n1264, n1276, n1277 );
nor U2977 ( n1265, g926, n1266 );
nor U2978 ( n1290, n1291, n1292 );
nor U2979 ( n1291, n1303, n1763 );
nand U2980 ( n1292, n1293, n1747 );
nand U2981 ( n1293, n1294, n1295 );
nor U2982 ( n1294, n1273, n1752 );
nor U2983 ( n1295, g889, n127 );
nand U2984 ( new_g6457_, n1287, n1288 );
nand U2985 ( n1288, g887, n1279 );
nor U2986 ( n1287, n1283, n1289 );
nor U2987 ( n1289, g785, n1290 );
nand U2988 ( n787, n821, n822 );
or U2989 ( n822, n823, n824 );
nor U2990 ( n821, n66, n827 );
nand U2991 ( n823, n826, g43 );
nor U2992 ( new_g8801_, n819, n820 );
nor U2993 ( n820, g6425, n787 );
nor U2994 ( new_g8911_, new_g7406_, n786 );
nor U2995 ( n786, n787, n788 );
nand U2996 ( n788, n789, g9132 );
nand U2997 ( n789, n790, g1018 );
nand U2998 ( n886, n898, n899 );
or U2999 ( n899, n87, g1025 );
and U3000 ( n898, n900, g43 );
nand U3001 ( n900, g9132, n1725 );
nand U3002 ( new_g7837_, n882, n883 );
nand U3003 ( n883, n884, g1025 );
nor U3004 ( n884, n885, n886 );
nor U3005 ( n1303, g889, n1279 );
nand U3006 ( new_g7832_, n882, n897 );
or U3007 ( n897, n886, g1018 );
nor U3008 ( new_g7833_, n886, n894 );
nand U3009 ( n894, n895, n1782 );
nand U3010 ( n895, n87, n896 );
nand U3011 ( n969, g822, n79 );
nand U3012 ( n1680, g819, g815 );
nor U3013 ( n827, n828, n829 );
nand U3014 ( n829, g999, g998 );
xnor U3015 ( n1331, g831, g1783 );
nor U3016 ( n1327, n1328, n1329 );
nand U3017 ( n1328, n1332, n1333 );
nand U3018 ( n1329, n1330, n1331 );
xnor U3019 ( n1332, g834, g1829 );
nor U3020 ( g6849, n1323, n1324 );
or U3021 ( n1323, g778, g889 );
nand U3022 ( n1324, n1270, n1325 );
nand U3023 ( n1325, n1326, n1327 );
nand U3024 ( n882, g1017, n898 );
xnor U3025 ( n1330, g843, g1810 );
xnor U3026 ( n1337, g849, g1798 );
nor U3027 ( n825, n189, n188 );
not U3028 ( n188, g10 );
nor U3029 ( n1326, n1334, n1335 );
nand U3030 ( n1334, n1338, n1339 );
nand U3031 ( n1335, n1336, n1337 );
xnor U3032 ( n1338, g852, g883 );
nand U3033 ( n824, n825, g1007 );
xnor U3034 ( n1336, g837, g1824 );
xnor U3035 ( n1333, g846, g1804 );
xnor U3036 ( n1339, g840, g1817 );
nor U3037 ( n826, g1016, g1008 );
nor U3038 ( n904, n1722, g940 );
nand U3039 ( n890, n891, g55 );
nor U3040 ( n891, g45, n190 );
nand U3041 ( n889, n1784, n890 );
nor U3042 ( new_g8976_, g979, n785 );
nor U3043 ( n1270, g887, g785 );
nor U3044 ( n1657, g1366, n1658 );
or U3045 ( n1658, g1368, g1367 );
nor U3046 ( new_g6643_, g6850, g162 );
nor U3047 ( g5164, n1816, n1817 );
nand U3048 ( n1816, g887, g889 );
nor U3049 ( n1656, g1363, n1659 );
or U3050 ( n1659, g1365, g1364 );
nor U3051 ( n1660, g1369, n1664 );
or U3052 ( n1664, g1371, g1370 );
nor U3053 ( n1663, g1375, g1374 );
nand U3054 ( n1451, n1452, n1453 );
nand U3055 ( n1453, g677, g652 );
nor U3056 ( n1452, n1454, n1455 );
and U3057 ( n1454, g647, g681 );
and U3058 ( n1455, g648, g685 );
nand U3059 ( n1463, n1464, n1465 );
nand U3060 ( n1465, g723, g730 );
nor U3061 ( n1464, n1466, n1467 );
and U3062 ( n1466, g718, g702 );
and U3063 ( n1467, g734, g722 );
nor U3064 ( n1662, g1373, g1372 );
nand U3065 ( n1450, n1456, n1457 );
nor U3066 ( n1456, n1460, n1461 );
nor U3067 ( n1457, n1458, n1459 );
and U3068 ( n1460, g635, g669 );
and U3069 ( n1459, g634, g665 );
and U3070 ( n1461, g645, g673 );
and U3071 ( n1468, n1818, n1819 );
nand U3072 ( n1818, g690, g706 );
nand U3073 ( n1819, g710, g694 );
and U3074 ( n1458, g633, g661 );
or U3075 ( n1033, n1820, n1078 );
or U3076 ( n799, n1821, n861 );
nand U3077 ( n784, n798, g1061 );
nor U3078 ( n798, n799, n1743 );
nand U3079 ( n960, n1032, g1149 );
nor U3080 ( n1032, n1033, n1730 );
nand U3081 ( n861, n874, g1049 );
nor U3082 ( n874, n875, n1736 );
nand U3083 ( n1078, n1137, g1134 );
nor U3084 ( n1137, n1729, n1700 );
nor U3085 ( n780, n1758, n784 );
or U3086 ( n875, n1823, n960 );
nand U3087 ( new_g9080_, n699, n700 );
nand U3088 ( n700, n701, g1069 );
nand U3089 ( n699, g4267, n702 );
nor U3090 ( n701, n140, n8 );
nand U3091 ( new_g8978_, n777, n778 );
nand U3092 ( n778, n779, n780 );
nand U3093 ( n777, g1069, n702 );
nor U3094 ( n779, g1069, n140 );
nor U3095 ( new_g4728_, n1601, n1788 );
nor U3096 ( n1601, g207, n1602 );
xor U3097 ( n1602, g210, g1206 );
nor U3098 ( new_g4705_, n1607, n1788 );
nor U3099 ( n1607, g202, n1608 );
xor U3100 ( n1608, g205, g1202 );
nor U3101 ( new_g4711_, n1605, n1788 );
nor U3102 ( n1605, g196, n1606 );
xor U3103 ( n1606, g195, g1194 );
nor U3104 ( new_g4720_, n1603, n1788 );
nor U3105 ( n1603, g187, n1604 );
xor U3106 ( n1604, g186, g1198 );
nand U3107 ( n1621, g940, n1722 );
nor U3108 ( new_g4676_, n1612, n4 );
nor U3109 ( n1612, n1781, n1613 );
nand U3110 ( n1613, g945, g955 );
nand U3111 ( n1676, n967, g786 );
nand U3112 ( n1685, n1673, n1674 );
nand U3113 ( n1674, g825, n969 );
nor U3114 ( n1673, n84, n1675 );
nor U3115 ( n1675, g825, n969 );
nand U3116 ( n1469, g698, g714 );
nand U3117 ( n1686, n1677, n1678 );
nand U3118 ( n1677, g822, n1680 );
nand U3119 ( n1678, n79, n1679 );
nand U3120 ( n1679, g822, n1676 );
nand U3121 ( n961, g781, n1100 );
nand U3122 ( n1684, n1671, n44 );
xnor U3123 ( n1671, g809, n1672 );
nor U3124 ( new_g7314_, n975, n961 );
nor U3125 ( n975, g775, n976 );
nor U3126 ( new_g7321_, g799, n961 );
and U3127 ( g4664, n1824, g1400 );
and U3128 ( g4663, n1825, g1397 );
and U3129 ( g4661, n1826, g1394 );
and U3130 ( g4660, n1827, g1392 );
nor U3131 ( new_g7324_, n961, n962 );
nand U3132 ( n962, n963, n964 );
or U3133 ( n963, g799, g803 );
nand U3134 ( g7048, g944, n1695 );
nor U3135 ( new_g6949_, n819, n1145 );
or U3136 ( n1145, g43, g985 );
nand U3137 ( g7731, n1828, n1829 );
xnor U3138 ( n1687, g945, n1681 );
nand U3139 ( n1681, g959, g955 );
xnor U3140 ( n1689, g871, n1682 );
nand U3141 ( n1682, g933, g929 );
nand U3142 ( g7063, g1412, g1405 );
xnor U3143 ( n1690, g933, g3856 );
nor U3144 ( n801, n834, n835 );
nor U3145 ( n835, n141, g1057 );
nand U3146 ( n800, n801, n802 );
or U3147 ( n802, n141, g1061 );
nand U3148 ( new_g8901_, n793, n795 );
nand U3149 ( n795, n796, n797 );
nand U3150 ( n793, g1065, n800 );
nor U3151 ( n796, g1065, n784 );
nand U3152 ( new_g8793_, n830, n831 );
nand U3153 ( n831, n832, n833 );
nand U3154 ( n830, g1061, n7 );
nor U3155 ( n832, n1743, n140 );
nor U3156 ( new_g6951_, g43, n1144 );
xnor U3157 ( n1144, g990, g985 );
nor U3158 ( new_g6954_, g43, n1140 );
xor U3159 ( n1140, n1141, g995 );
nand U3160 ( n1141, g990, g985 );
xnor U3161 ( n1688, n1781, g955 );
nand U3162 ( new_g6445_, n1304, n1305 );
nand U3163 ( n1304, g12, g859 );
nand U3164 ( n1305, g11, n1694 );
nand U3165 ( new_g4747_, n1599, n1600 );
or U3166 ( n1599, n1776, g1176 );
nand U3167 ( n1600, g1080, n1776 );
nand U3168 ( new_g8607_, n857, n858 );
nand U3169 ( n858, n859, n797 );
nand U3170 ( n857, g1057, n834 );
nor U3171 ( n859, g1057, n799 );
nor U3172 ( n833, g1061, n799 );
nand U3173 ( n1123, n1126, g1348 );
nor U3174 ( n1126, n1127, n1738 );
nand U3175 ( n1436, n1437, g1336 );
nor U3176 ( n1437, n1731, n1701 );
nand U3177 ( n1127, g1342, n1130 );
nand U3178 ( n924, g1354, n926 );
nand U3179 ( n922, g1357, n18 );
nor U3180 ( new_g7679_, n1759, n919 );
nand U3181 ( n919, n920, n921 );
nand U3182 ( n920, n923, g1360 );
nand U3183 ( n921, n1771, n922 );
nor U3184 ( n877, n931, n932 );
nor U3185 ( n932, n141, g1045 );
nand U3186 ( n876, n877, n878 );
or U3187 ( n878, n141, g1049 );
nand U3188 ( new_g8068_, n871, n872 );
nand U3189 ( n872, n873, n797 );
nand U3190 ( n871, g1053, n876 );
nor U3191 ( n873, g1053, n861 );
nand U3192 ( new_g7605_, n927, n928 );
nand U3193 ( n928, n929, n930 );
nand U3194 ( n927, g1049, n6 );
nor U3195 ( n929, n1736, n140 );
nor U3196 ( new_g7677_, n925, n1759 );
xnor U3197 ( n925, g1357, n18 );
nand U3198 ( n1313, n1433, g1220 );
nand U3199 ( n1236, n1244, g1227 );
nor U3200 ( n1244, n1245, n1737 );
nand U3201 ( new_g7020_, n1766, n1112 );
nand U3202 ( n1112, g2662, n1113 );
xnor U3203 ( n1113, n1708, n1114 );
nand U3204 ( n1312, n1429, g1225 );
nor U3205 ( n1429, n1733, n1703 );
nand U3206 ( n1065, n1256, n1257 );
nor U3207 ( n1256, n1260, n1261 );
nor U3208 ( n1257, n1258, n1259 );
nand U3209 ( n1261, g1323, g1322 );
nand U3210 ( n1066, n1255, g1325 );
nor U3211 ( n1255, n1065, n1740 );
nand U3212 ( n1259, g1319, g1318 );
nand U3213 ( n1053, g1327, n1055 );
nand U3214 ( n1186, g1328, n96 );
nor U3215 ( new_g6460_, n1851, n1254 );
nor U3216 ( n1254, n95, g5669 );
not U3217 ( n95, n1186 );
nor U3218 ( n1187, n96, g1328 );
nand U3219 ( n1258, g1317, g1313 );
nand U3220 ( new_g6912_, n1183, n1184 );
nand U3221 ( n1183, g93, n1851 );
nand U3222 ( n1184, n1185, n1186 );
nor U3223 ( n1185, n1852, n1187 );
nand U3224 ( new_g7415_, n956, n957 );
nand U3225 ( n957, n958, n797 );
nand U3226 ( n956, g1045, n931 );
nor U3227 ( n958, g1045, n875 );
nand U3228 ( new_g7220_, n1014, n1015 );
nand U3229 ( n1015, g1288, n1710 );
nor U3230 ( n1014, g1304, n1016 );
nor U3231 ( n1016, n1017, n1710 );
nand U3232 ( n1111, g1288, n1020 );
nor U3233 ( n1017, n1018, new_g4681_ );
nor U3234 ( n1018, n48, n1019 );
nor U3235 ( n1019, n1020, g1288 );
and U3236 ( n1020, g1284, n1119 );
and U3237 ( n1094, n1105, g1300 );
and U3238 ( new_g4681_, g1296, n1094 );
nor U3239 ( n1119, n1830, n1831 );
nand U3240 ( n1830, g1272, g1276 );
nor U3241 ( new_g7197_, n1028, n1759 );
xnor U3242 ( n1028, n926, g1354 );
nor U3243 ( n930, g1049, n875 );
nand U3244 ( n1260, g1321, g1320 );
and U3245 ( n1273, n1296, n1297 );
nor U3246 ( n1296, n1301, n1302 );
nor U3247 ( n1297, n1298, n1299 );
or U3248 ( n1301, g1783, g1798 );
or U3249 ( n1299, g1829, g1810 );
or U3250 ( n1302, g883, g1817 );
or U3251 ( n1298, g1804, g1824 );
nand U3252 ( new_g7031_, n1088, n1089 );
nand U3253 ( n1088, n1095, g1296 );
nand U3254 ( n1089, n1090, n1091 );
nor U3255 ( n1090, new_g4681_, n1093 );
nor U3256 ( n1093, n1094, g1296 );
nor U3257 ( n1054, n1055, g1327 );
nand U3258 ( new_g7089_, n1050, n1051 );
nand U3259 ( n1050, g98, n1850 );
nand U3260 ( n1051, n1052, n1053 );
nor U3261 ( n1052, n1850, n1054 );
nor U3262 ( n1035, n1074, n1135 );
nor U3263 ( n1135, n141, g1149 );
nand U3264 ( new_g7177_, n1029, n1030 );
nand U3265 ( n1030, n1031, n797 );
nand U3266 ( n1029, g1041, n1034 );
nor U3267 ( n1031, g1041, n960 );
nor U3268 ( new_g7007_, n1759, n1124 );
nand U3269 ( n1124, n1125, n1123 );
nand U3270 ( n1125, n1772, n1128 );
nand U3271 ( n1128, g1345, n16 );
nand U3272 ( n783, g4267, g1158 );
nand U3273 ( new_g7033_, n1082, n1083 );
nand U3274 ( n1082, g1134, n12 );
nand U3275 ( n1083, n1084, n1085 );
not U3276 ( n12, n1080 );
nand U3277 ( n1315, n1318, g1224 );
nand U3278 ( new_g6120_, n1314, n1766 );
xor U3279 ( n1314, n1315, g1225 );
nand U3280 ( n918, n1024, n1025 );
and U3281 ( n1024, g1114, g1118 );
nor U3282 ( n1025, n1026, n1741 );
or U3283 ( n1026, n1832, n1833 );
nand U3284 ( n1832, g1102, g1106 );
nand U3285 ( n1833, g1087, g1098 );
nor U3286 ( new_g8076_, g1097, n868 );
xor U3287 ( n868, n869, g1142 );
nand U3288 ( n869, n867, g1126 );
and U3289 ( n867, g1122, n870 );
nand U3290 ( new_g6966_, n1131, n1132 );
nand U3291 ( n1132, n1133, n1134 );
or U3292 ( n1131, n1730, n1035 );
nor U3293 ( n1134, g1037, n1033 );
nand U3294 ( new_g6585_, n1766, n1237 );
nand U3295 ( n1237, n1238, n1236 );
nand U3296 ( n1238, n1765, n1239 );
nand U3297 ( n1239, g1226, n81 );
nand U3298 ( new_g7080_, n1067, n1068 );
nand U3299 ( n1067, g103, n1852 );
nand U3300 ( n1068, n1069, n1070 );
nand U3301 ( n1070, n1751, n1066 );
nand U3302 ( new_g7027_, n1101, n1102 );
nand U3303 ( n1101, n1095, g1300 );
nand U3304 ( n1102, n1103, n1091 );
nor U3305 ( n1103, n1094, n1104 );
nor U3306 ( n1104, n1105, g1300 );
nor U3307 ( new_g7002_, n1129, n1759 );
xnor U3308 ( n1129, g1345, n16 );
or U3309 ( n949, n1834, n1835 );
nand U3310 ( n1834, g1494, g1499 );
nand U3311 ( n1835, g1481, g1489 );
nor U3312 ( new_g8059_, n879, n837 );
xor U3313 ( n879, n880, g1467 );
nand U3314 ( n880, n881, g1462 );
nor U3315 ( n864, n1836, n1837 );
nand U3316 ( n1836, g1514, g1509 );
or U3317 ( n1837, n949, n1739 );
nand U3318 ( n1240, g1247, n1319 );
nand U3319 ( n1319, n1320, n1321 );
or U3320 ( n1321, g1257, g1263 );
and U3321 ( n1320, n1426, n1427 );
nor U3322 ( n1426, n1708, n1430 );
nor U3323 ( n1427, n1737, n1428 );
nand U3324 ( n1430, g1228, g1227 );
or U3325 ( n1428, n1312, g1229 );
nand U3326 ( new_g6579_, g1253, n1240 );
nand U3327 ( n1275, g785, n1283 );
nor U3328 ( n1283, n1747, g889 );
nand U3329 ( n1214, n1209, g1321 );
nand U3330 ( n1208, n1225, n1224 );
and U3331 ( n1225, g1318, g1319 );
and U3332 ( n1224, g1317, g1313 );
nand U3333 ( new_g6739_, n1200, n1201 );
nand U3334 ( n1200, g117, n1850 );
nand U3335 ( n1201, n1202, n1770 );
xor U3336 ( n1202, g1323, n1203 );
nand U3337 ( n837, n986, n1000 );
nand U3338 ( n1000, n101, n1001 );
xor U3339 ( n1001, g1911, g1513 );
not U3340 ( n101, n985 );
nand U3341 ( n985, g150, n1725 );
nor U3342 ( new_g8779_, n836, n837 );
xnor U3343 ( n836, g1477, n838 );
nor U3344 ( n838, n1757, n839 );
nor U3345 ( new_g7596_, n933, n837 );
xnor U3346 ( n933, g1462, n881 );
nor U3347 ( new_g7242_, n988, n837 );
xor U3348 ( n988, n989, g1514 );
nand U3349 ( n989, n990, g1509 );
nor U3350 ( new_g7240_, n991, n837 );
xnor U3351 ( n991, g1509, n990 );
nor U3352 ( new_g7235_, n994, n837 );
xnor U3353 ( n994, g1499, n995 );
nor U3354 ( n995, n1767, n996 );
nor U3355 ( new_g7228_, n999, n837 );
xnor U3356 ( n999, n998, g1489 );
nand U3357 ( new_g6123_, n1309, n1766 );
xnor U3358 ( n1309, g1226, n81 );
nor U3359 ( new_g7271_, n837, n980 );
xnor U3360 ( n980, g1481, n1749 );
nand U3361 ( n964, g803, g799 );
nand U3362 ( n979, n1672, g809 );
nand U3363 ( n1100, g775, n976 );
nand U3364 ( new_g6686_, n1215, n1216 );
nand U3365 ( n1215, g121, n1851 );
nand U3366 ( n1216, n1217, n1218 );
nand U3367 ( n1218, n1762, n1214 );
nor U3368 ( n1059, n1705, g8216 );
nand U3369 ( n839, n863, n864 );
nor U3370 ( n863, g8216, n865 );
or U3371 ( n992, n949, g8216 );
nand U3372 ( n1005, n1006, n1007 );
nand U3373 ( n1006, g1514, n1706 );
nand U3374 ( n1007, n1008, g1504 );
and U3375 ( n1008, g174, g1477 );
nor U3376 ( new_g7021_, g1304, n1109 );
xnor U3377 ( n1109, n1110, n1746 );
nand U3378 ( n1110, g1307, n48 );
nor U3379 ( n1080, n1086, n1087 );
nor U3380 ( n1087, n141, g1130 );
nand U3381 ( n1079, n1080, n1081 );
or U3382 ( n1081, n141, g1134 );
nand U3383 ( new_g7036_, n1075, n1076 );
nand U3384 ( n1076, n1077, n797 );
nand U3385 ( n1075, g1138, n1079 );
nor U3386 ( n1077, g1138, n1078 );
nand U3387 ( new_g8155_, n866, n1778 );
xnor U3388 ( n866, g1126, n867 );
nand U3389 ( new_g7041_, n1071, n1072 );
nand U3390 ( n1072, n1073, n797 );
nand U3391 ( n1071, g1149, n1074 );
nor U3392 ( n1073, g1149, n1033 );
nand U3393 ( new_g7254_, n981, n982 );
or U3394 ( n981, n985, g1911 );
nand U3395 ( n982, n984, n985 );
xnor U3396 ( n984, g1486, n986 );
and U3397 ( n1133, g1149, n797 );
nand U3398 ( new_g5686_, g1263, n1320 );
nand U3399 ( new_g5559_, g1257, n1320 );
nand U3400 ( new_g5538_, g1266, n1320 );
nand U3401 ( new_g7426_, n953, n954 );
nor U3402 ( n954, g7425, n955 );
nor U3403 ( n953, g1166, new_g7217_ );
or U3404 ( n955, g7424, g7423 );
and U3405 ( new_g7217_, n1021, n1022 );
and U3406 ( n1021, g1126, g1142 );
nor U3407 ( n1022, n918, n1769 );
nand U3408 ( n865, n1011, g1519 );
and U3409 ( n1011, g1462, g1467 );
nand U3410 ( new_g7086_, n1060, n1061 );
nand U3411 ( n1060, g108, n1851 );
nand U3412 ( n1061, n1062, n1063 );
nand U3413 ( n1063, n1777, n1064 );
nor U3414 ( new_g6091_, n1322, n1759 );
xnor U3415 ( n1322, n1130, g1342 );
nand U3416 ( new_g7030_, n1096, n1097 );
nand U3417 ( n1096, g1130, n1086 );
nand U3418 ( n1097, n1098, n797 );
nor U3419 ( n1098, g1130, n1729 );
nand U3420 ( new_g7697_, n917, n1778 );
xnor U3421 ( n917, n870, g1122 );
nand U3422 ( new_g6718_, n1210, n1211 );
nand U3423 ( n1210, g125, n1852 );
nand U3424 ( n1211, n1212, n1213 );
or U3425 ( n1213, g1321, n1209 );
xnor U3426 ( new_g7029_, g778, n1100 );
or U3427 ( new_g5657_, n1395, n904 );
nor U3428 ( n1395, g943, n4 );
nand U3429 ( new_g7443_, n950, n1778 );
xor U3430 ( n950, n951, g1118 );
nand U3431 ( n951, n952, g1114 );
and U3432 ( n952, n1013, g1110 );
nand U3433 ( n996, n998, g1489 );
and U3434 ( n998, g1481, n1749 );
nor U3435 ( n1282, n1284, n1285 );
nor U3436 ( n1285, g4316, g785 );
nor U3437 ( n1284, g875, n1817 );
nor U3438 ( n885, g1021, g1018 );
xnor U3439 ( n1403, g632, n1731 );
nand U3440 ( n1400, n1401, n1402 );
xnor U3441 ( n1402, g630, g1336 );
nor U3442 ( n1401, n1403, n1404 );
xnor U3443 ( n1404, n1720, g1354 );
nand U3444 ( new_g7227_, n1012, n1778 );
xnor U3445 ( n1012, g1114, n952 );
nand U3446 ( new_g6735_, n1204, n1205 );
nand U3447 ( n1204, g129, n1852 );
nand U3448 ( n1205, n1206, n1207 );
nand U3449 ( n1207, n1745, n1208 );
xnor U3450 ( n1384, g759, n1753 );
nand U3451 ( n1380, n1381, n1382 );
xnor U3452 ( n1382, g761, g1351 );
nor U3453 ( n1381, n1383, n1384 );
xor U3454 ( n1383, g760, g1354 );
xnor U3455 ( n1416, g631, n1701 );
nand U3456 ( n1409, n1413, n1414 );
xnor U3457 ( n1414, g626, g1348 );
nor U3458 ( n1413, n1415, n1416 );
xnor U3459 ( n1415, g627, n1738 );
nand U3460 ( new_g5566_, n1766, n1417 );
nand U3461 ( n1417, n1418, n1419 );
nand U3462 ( n1418, n1732, n1420 );
nand U3463 ( n1420, n1310, g1214 );
nand U3464 ( new_g7017_, n1115, n1116 );
nand U3465 ( n1115, n1095, g1284 );
nand U3466 ( n1116, n1117, n1091 );
nor U3467 ( n1117, n1020, n1118 );
and U3468 ( n1342, g533, n1838 );
and U3469 ( n1347, g452, n1839 );
and U3470 ( n1359, g290, n1840 );
and U3471 ( n1352, g371, n1841 );
nand U3472 ( new_g5231_, n1513, n1514 );
nand U3473 ( n1514, g455, n1342 );
nand U3474 ( n1513, g462, n89 );
nand U3475 ( new_g5254_, n1485, n1486 );
nand U3476 ( n1486, g435, n1347 );
nand U3477 ( n1485, g437, n1 );
nand U3478 ( new_g5219_, n1532, n1533 );
nand U3479 ( n1533, g374, n1347 );
nand U3480 ( n1532, g381, n1 );
nand U3481 ( new_g5221_, n1528, n1529 );
nand U3482 ( n1529, g454, n1342 );
nand U3483 ( n1528, g459, n89 );
nand U3484 ( new_g5229_, n1518, n1519 );
nand U3485 ( n1519, g375, n1347 );
nand U3486 ( n1518, g384, n1 );
nand U3487 ( new_g5235_, n1505, n1506 );
nand U3488 ( n1506, g397, n1347 );
nand U3489 ( n1505, g411, n1 );
nand U3490 ( new_g5707_, n1355, n1356 );
nand U3491 ( n1356, g295, n1352 );
nand U3492 ( n1355, g306, n108 );
nand U3493 ( new_g5243_, n1493, n1494 );
nand U3494 ( n1494, g398, n1347 );
nand U3495 ( n1493, g414, n1 );
nand U3496 ( new_g5203_, n1560, n1561 );
nand U3497 ( n1561, g313, n1352 );
nand U3498 ( n1560, g321, n108 );
nand U3499 ( new_g5211_, n1548, n1549 );
nand U3500 ( n1549, g314, n1352 );
nand U3501 ( n1548, g324, n108 );
nand U3502 ( new_g5711_, n1348, n1349 );
nand U3503 ( n1349, g376, n1347 );
nand U3504 ( n1348, g387, n1 );
nand U3505 ( new_g5210_, n1550, n1551 );
nand U3506 ( n1551, g293, n1352 );
nand U3507 ( n1550, g300, n108 );
nand U3508 ( new_g5264_, n1475, n1476 );
nand U3509 ( n1476, g517, n1342 );
nand U3510 ( n1475, g521, n89 );
nand U3511 ( new_g5227_, n1522, n1523 );
nand U3512 ( n1523, g236, n1359 );
nand U3513 ( n1522, g252, n121 );
nand U3514 ( new_g5193_, n1575, n1576 );
nand U3515 ( n1576, g211, n1359 );
nand U3516 ( n1575, g216, n121 );
nand U3517 ( new_g5220_, n1530, n1531 );
nand U3518 ( n1531, g395, n1347 );
nand U3519 ( n1530, g405, n1 );
nand U3520 ( new_g5212_, n1546, n1547 );
nand U3521 ( n1547, g373, n1347 );
nand U3522 ( n1546, g378, n1 );
nand U3523 ( new_g5202_, n1562, n1563 );
nand U3524 ( n1563, g292, n1352 );
nand U3525 ( n1562, g297, n108 );
nand U3526 ( new_g5200_, n1567, n1568 );
nand U3527 ( n1568, g212, n1359 );
nand U3528 ( n1567, g219, n121 );
nand U3529 ( new_g5208_, n1554, n1555 );
nand U3530 ( n1555, g213, n1359 );
nand U3531 ( n1554, g222, n121 );
nand U3532 ( new_g5236_, n1503, n1504 );
nand U3533 ( n1504, g456, n1342 );
nand U3534 ( n1503, g465, n89 );
nand U3535 ( new_g5217_, n1536, n1537 );
nand U3536 ( n1537, g294, n1352 );
nand U3537 ( n1536, g303, n108 );
nand U3538 ( new_g5704_, n1360, n1361 );
nand U3539 ( n1361, g214, n1359 );
nand U3540 ( n1360, g225, n121 );
nand U3541 ( new_g5716_, n1343, n1344 );
nand U3542 ( n1344, g457, n1342 );
nand U3543 ( n1343, g468, n89 );
nand U3544 ( new_g5706_, n1357, n1358 );
nand U3545 ( n1358, g215, n1359 );
nand U3546 ( n1357, g228, n121 );
nand U3547 ( new_g5710_, n1350, n1351 );
nand U3548 ( n1351, g296, n1352 );
nand U3549 ( n1350, g309, n108 );
nand U3550 ( new_g5715_, n1345, n1346 );
nand U3551 ( n1346, g377, n1347 );
nand U3552 ( n1345, g390, n1 );
nand U3553 ( new_g5722_, n1340, n1341 );
nand U3554 ( n1341, g458, n1342 );
nand U3555 ( n1340, g471, n89 );
nand U3556 ( new_g5222_, n1526, n1527 );
nand U3557 ( n1527, g475, n1342 );
nand U3558 ( n1526, g483, n89 );
nand U3559 ( new_g5194_, n1573, n1574 );
nand U3560 ( n1574, g232, n1359 );
nand U3561 ( n1573, g240, n121 );
nand U3562 ( new_g5213_, n1544, n1545 );
nand U3563 ( n1545, g394, n1347 );
nand U3564 ( n1544, g402, n1 );
nand U3565 ( new_g5214_, n1542, n1543 );
nand U3566 ( n1543, g474, n1342 );
nand U3567 ( n1542, g480, n89 );
nand U3568 ( new_g5188_, n1577, n1578 );
nand U3569 ( n1578, g231, n1359 );
nand U3570 ( n1577, g237, n121 );
nand U3571 ( new_g5204_, n1558, n1559 );
nand U3572 ( n1559, g393, n1347 );
nand U3573 ( n1558, g399, n1 );
nand U3574 ( new_g5195_, n1571, n1572 );
nand U3575 ( n1572, g312, n1352 );
nand U3576 ( n1571, g318, n108 );
nand U3577 ( new_g5230_, n1515, n1517 );
nand U3578 ( n1517, g396, n1347 );
nand U3579 ( n1515, g408, n1 );
nand U3580 ( new_g5209_, n1552, n1553 );
nand U3581 ( n1553, g234, n1359 );
nand U3582 ( n1552, g246, n121 );
nand U3583 ( new_g5237_, n1501, n1502 );
nand U3584 ( n1502, g477, n1342 );
nand U3585 ( n1501, g489, n89 );
nand U3586 ( new_g5218_, n1534, n1535 );
nand U3587 ( n1535, g315, n1352 );
nand U3588 ( n1534, g327, n108 );
nand U3589 ( new_g5216_, n1538, n1539 );
nand U3590 ( n1539, g235, n1359 );
nand U3591 ( n1538, g249, n121 );
nand U3592 ( new_g5228_, n1520, n1521 );
nand U3593 ( n1521, g316, n1352 );
nand U3594 ( n1520, g330, n108 );
nand U3595 ( new_g5244_, n1491, n1492 );
nand U3596 ( n1492, g478, n1342 );
nand U3597 ( n1491, g492, n89 );
nand U3598 ( new_g5255_, n1483, n1484 );
nand U3599 ( n1484, g479, n1342 );
nand U3600 ( n1483, g495, n89 );
nand U3601 ( new_g5234_, n1507, n1508 );
nand U3602 ( n1508, g317, n1352 );
nand U3603 ( n1507, g333, n108 );
nand U3604 ( new_g5201_, n1564, n1565 );
nand U3605 ( n1565, g233, n1359 );
nand U3606 ( n1564, g243, n121 );
nand U3607 ( new_g5232_, n1511, n1512 );
nand U3608 ( n1512, g476, n1342 );
nand U3609 ( n1511, g486, n89 );
nand U3610 ( new_g5260_, n1477, n1478 );
nand U3611 ( n1478, g516, n1342 );
nand U3612 ( n1477, g518, n89 );
nand U3613 ( new_g5242_, n1495, n1496 );
nand U3614 ( n1496, g354, n1352 );
nand U3615 ( n1495, g356, n108 );
nand U3616 ( new_g5233_, n1509, n1510 );
nand U3617 ( n1510, g273, n1359 );
nand U3618 ( n1509, g275, n121 );
nand U3619 ( new_g5259_, n1479, n1480 );
nand U3620 ( n1480, g436, n1347 );
nand U3621 ( n1479, g440, n1 );
nand U3622 ( new_g5241_, n1497, n1498 );
nand U3623 ( n1498, g274, n1359 );
nand U3624 ( n1497, g278, n121 );
nand U3625 ( new_g5253_, n1487, n1488 );
nand U3626 ( n1488, g355, n1352 );
nand U3627 ( n1487, g359, n108 );
nand U3628 ( new_g6740_, n1197, n1198 );
nand U3629 ( n1197, g113, n1850 );
nand U3630 ( n1198, n1199, n1770 );
xnor U3631 ( n1199, g1324, n1065 );
nor U3632 ( n1625, g1459, n1640 );
nor U3633 ( n1640, n1754, n1709 );
nand U3634 ( new_g4256_, g1444, n1625 );
nand U3635 ( new_g4299_, n1623, n1624 );
nand U3636 ( n1624, n1625, g1454 );
or U3637 ( n1623, n1754, new_g4256_ );
nand U3638 ( n1286, n1270, g889 );
nor U3639 ( n1597, n1638, g7507 );
nand U3640 ( n1638, g1439, g1432 );
nor U3641 ( new_g4868_, n1586, n1241 );
xnor U3642 ( n1586, n1310, g1214 );
nand U3643 ( new_g4812_, n1595, n1596 );
nand U3644 ( n1596, n1597, n1773 );
nor U3645 ( n1595, g1443, n1598 );
nor U3646 ( n1598, n1597, n1773 );
nor U3647 ( n1118, n1119, g1284 );
nand U3648 ( new_g7318_, n972, n973 );
nand U3649 ( n973, n974, g825 );
or U3650 ( n972, n1723, n971 );
nor U3651 ( n974, g828, n969 );
xnor U3652 ( n1393, g763, n1738 );
nand U3653 ( n1387, n1391, n1392 );
xnor U3654 ( n1392, g762, g1348 );
nor U3655 ( n1391, n1393, n1394 );
xor U3656 ( n1394, g766, g1336 );
nor U3657 ( new_g5475_, n1759, g1330 );
or U3658 ( n1442, new_g5475_, n1842 );
and U3659 ( n1842, g1247, n1701 );
nand U3660 ( new_g5489_, n1438, n1439 );
nand U3661 ( n1439, n1440, n1441 );
nand U3662 ( n1438, g1336, n1442 );
nor U3663 ( n1441, g1336, n1731 );
xnor U3664 ( n1407, g625, n1748 );
nand U3665 ( n1399, n1405, n1406 );
xnor U3666 ( n1406, g623, g1357 );
nor U3667 ( n1405, n1407, n1408 );
xnor U3668 ( n1408, n1721, g1360 );
nand U3669 ( n1229, g1307, g1272 );
nor U3670 ( new_g6611_, g1304, n1227 );
xnor U3671 ( n1227, g1280, n1228 );
nor U3672 ( n1228, n1764, n1229 );
nand U3673 ( n1276, g874, n1817 );
nor U3674 ( n1250, n1705, n1761 );
nor U3675 ( n1248, g1077, n1249 );
and U3676 ( n1249, n1250, g1179 );
nand U3677 ( new_g6571_, n1246, n1247 );
nand U3678 ( n1246, n1249, n1780 );
nand U3679 ( n1247, n1248, g2888 );
nand U3680 ( n1277, g889, g887 );
nand U3681 ( new_g7025_, n1106, n1778 );
xnor U3682 ( n1106, n1013, g1110 );
nor U3683 ( new_g7087_, n141, n1058 );
xnor U3684 ( n1058, n1059, g1092 );
nand U3685 ( new_g7788_, n909, n910 );
nand U3686 ( n909, n904, g48 );
nand U3687 ( n910, g954, n5 );
nand U3688 ( new_g7783_, n913, n914 );
nand U3689 ( n913, n904, g3 );
nand U3690 ( n914, g953, n5 );
nand U3691 ( new_g7826_, n902, n903 );
nand U3692 ( n902, n904, g2 );
nand U3693 ( n903, g952, n5 );
nand U3694 ( new_g7810_, n905, n906 );
nand U3695 ( n905, n904, g4 );
nand U3696 ( n906, g951, n5 );
nand U3697 ( new_g7791_, n907, n908 );
nand U3698 ( n907, n904, g5 );
nand U3699 ( n908, g950, n5 );
nand U3700 ( new_g7787_, n911, n912 );
nand U3701 ( n911, n904, g6 );
nand U3702 ( n912, g949, n5 );
nand U3703 ( new_g7782_, n915, n916 );
nand U3704 ( n915, n904, g7 );
nand U3705 ( n916, g948, n5 );
and U3706 ( new_g4272_, n1843, n1625 );
xor U3707 ( n1843, g1444, g1450 );
and U3708 ( n1474, g595, n1844 );
nand U3709 ( new_g5265_, n1472, n1473 );
nand U3710 ( n1473, g556, n1474 );
nand U3711 ( n1472, g557, n156 );
nand U3712 ( new_g5205_, n1556, n1557 );
nand U3713 ( n1557, g583, n1474 );
nand U3714 ( n1556, g584, n156 );
nand U3715 ( new_g5223_, n1524, n1525 );
nand U3716 ( n1525, g566, n1474 );
nand U3717 ( n1524, g567, n156 );
nand U3718 ( new_g5196_, n1569, n1570 );
nand U3719 ( n1570, g579, n1474 );
nand U3720 ( n1569, g580, n156 );
nand U3721 ( new_g5215_, n1540, n1541 );
nand U3722 ( n1541, g587, n1474 );
nand U3723 ( n1540, g560, n156 );
nand U3724 ( new_g5238_, n1499, n1500 );
nand U3725 ( n1500, g535, n1474 );
nand U3726 ( n1499, g536, n156 );
nand U3727 ( new_g5245_, n1489, n1490 );
nand U3728 ( n1490, g539, n1474 );
nand U3729 ( n1489, g540, n156 );
nand U3730 ( new_g5256_, n1481, n1482 );
nand U3731 ( n1482, g543, n1474 );
nand U3732 ( n1481, g544, n156 );
nor U3733 ( n790, g1025, g1021 );
or U3734 ( new_g7825_, n5, g8 );
nand U3735 ( new_g6602_, n1230, n1778 );
xor U3736 ( n1230, n1231, g1106 );
nand U3737 ( n1231, n1232, g1102 );
and U3738 ( n1232, n1446, g1098 );
and U3739 ( n1446, g1148, g1087 );
nand U3740 ( new_g6685_, n1219, n1220 );
nand U3741 ( n1219, g133, n1850 );
nand U3742 ( n1220, n1221, n1222 );
nand U3743 ( n1222, n1775, n1223 );
nor U3744 ( n1091, n1710, g1304 );
nand U3745 ( n1365, n1366, n1367 );
xnor U3746 ( n1366, g768, g1300 );
xnor U3747 ( n1367, g767, g1296 );
nor U3748 ( new_g5452_, g1097, n1445 );
xnor U3749 ( n1445, g1102, n1232 );
nand U3750 ( n1371, n1372, n1373 );
xnor U3751 ( n1372, g1280, g772 );
xnor U3752 ( n1373, g771, g1284 );
nand U3753 ( new_g4264_, n1636, n1637 );
nand U3754 ( n1637, g7507, n1638 );
nor U3755 ( n1636, g1443, n1597 );
nor U3756 ( n1095, g1304, g1307 );
nand U3757 ( n1364, n1368, n1369 );
xnor U3758 ( n1368, g769, g1292 );
xnor U3759 ( n1369, g770, g1288 );
xnor U3760 ( n1411, g628, g1342 );
xnor U3761 ( n1389, g764, g1342 );
xnor U3762 ( n1376, g774, g1272 );
nand U3763 ( n1379, n1385, n1386 );
nor U3764 ( n1385, g1333, g1330 );
xnor U3765 ( n1386, g758, g1360 );
nand U3766 ( new_g6262_, n1306, n1307 );
nand U3767 ( n1306, g137, n1851 );
nand U3768 ( n1307, n1308, n1770 );
xor U3769 ( n1308, g1318, n1224 );
xnor U3770 ( n1412, g629, g1339 );
xnor U3771 ( n1390, g765, g1339 );
buf U3772 ( n1850, g1329 );
buf U3773 ( n1851, g1329 );
nand U3774 ( n1223, n1224, g1318 );
buf U3775 ( n1852, g1329 );
nor U3776 ( new_g5563_, g1304, n1421 );
xnor U3777 ( n1421, n1229, n1764 );
xnor U3778 ( n1375, g773, g1276 );
nand U3779 ( new_g4879_, n1582, n1583 );
nor U3780 ( n1583, g1220, g1217 );
nor U3781 ( n1582, n1702, n1734 );
nor U3782 ( n1646, g1379, n1647 );
or U3783 ( n1647, g1381, g1380 );
and U3784 ( new_g4232_, g154, n1725 );
or U3785 ( new_g5572_, new_g4232_, g5571 );
nand U3786 ( n896, g1021, g1018 );
nor U3787 ( n1645, g1376, n1648 );
or U3788 ( n1648, g1378, g1377 );
nand U3789 ( n1241, g2662, n1766 );
nor U3790 ( new_g5441_, g1097, n1447 );
xnor U3791 ( n1447, n1446, g1098 );
and U3792 ( n819, n1146, g995 );
nor U3793 ( n1146, g990, g985 );
nor U3794 ( n1085, g1134, n1729 );
nor U3795 ( new_g4284_, n1627, n1628 );
xnor U3796 ( n1627, g1435, g1439 );
nor U3797 ( new_g4236_, n1641, n1628 );
nor U3798 ( n1641, g1432, n1642 );
and U3799 ( n1642, g1439, g1435 );
nor U3800 ( n1649, g1382, n1653 );
or U3801 ( n1653, g1384, g1383 );
nor U3802 ( n1652, g1388, g1387 );
nor U3803 ( new_g5560_, g1304, n1422 );
xnor U3804 ( n1422, g1272, g1307 );
nor U3805 ( n1651, g1386, g1385 );
nand U3806 ( new_g4688_, n1609, n1610 );
nand U3807 ( n1609, g145, n1851 );
or U3808 ( n1610, g1313, n1850 );
xnor U3809 ( new_g6280_, g600, n1737 );
xnor U3810 ( new_g6283_, g613, n1737 );
nand U3811 ( new_g5708_, n1353, n1354 );
nand U3812 ( n1353, g1077, g2888 );
nand U3813 ( n1354, n1250, g1176 );
xnor U3814 ( new_g6169_, g608, n1704 );
xnor U3815 ( new_g6181_, g621, n1704 );
or U3816 ( n1633, g1225, g1226 );
xnor U3817 ( new_g6170_, g620, n1734 );
xnor U3818 ( new_g6164_, g607, n1734 );
nor U3819 ( new_g5479_, n1444, n1759 );
xnor U3820 ( n1444, g1330, g1333 );
nand U3821 ( new_g5052_, n1579, n1580 );
nand U3822 ( n1579, g141, n1852 );
nand U3823 ( n1580, n1581, n1770 );
xor U3824 ( n1581, g1317, g1313 );
xnor U3825 ( new_g6159_, g606, n1702 );
xnor U3826 ( new_g6165_, g619, n1702 );
xnor U3827 ( new_g5747_, g604, n1744 );
xnor U3828 ( new_g5752_, g617, n1744 );
nor U3829 ( n1592, n1593, g1405 );
nor U3830 ( n1588, n1589, g1412 );
nand U3831 ( n1593, n1845, n1846 );
nand U3832 ( n1589, n1847, n1848 );
or U3833 ( new_g4825_, n1591, n1592 );
nor U3834 ( n1591, g1408, n1593 );
or U3835 ( new_g4840_, n1587, n1588 );
nor U3836 ( n1587, g1415, n1589 );
nand U3837 ( new_g4263_, n1639, g1435 );
and U3838 ( n1639, n1711, n1638 );
xnor U3839 ( new_g6281_, g612, n1765 );
xnor U3840 ( new_g6276_, g599, n1765 );
xnor U3841 ( new_g5753_, g618, n1732 );
xnor U3842 ( new_g5751_, g605, n1732 );
nor U3843 ( new_g3429_, n1779, n1665 );
nand U3844 ( n1665, g1454, n1754 );
or U3845 ( n1616, g4370, g4373 );
nand U3846 ( new_g4374_, n1614, n1615 );
nor U3847 ( n1614, n1617, g4267 );
nor U3848 ( n1615, g4371, n1616 );
or U3849 ( n1617, g4372, g1179 );
xnor U3850 ( new_g6287_, g615, n1703 );
xnor U3851 ( new_g6284_, g602, n1703 );
xnor U3852 ( new_g6275_, g610, n1755 );
xnor U3853 ( new_g6273_, g597, n1755 );
nor U3854 ( new_g5624_, g1097, n1396 );
xnor U3855 ( n1396, g1087, g1148 );
xnor U3856 ( new_g6277_, g611, n1707 );
xnor U3857 ( new_g6274_, g598, n1707 );
xnor U3858 ( new_g5748_, g616, n1733 );
xnor U3859 ( new_g6286_, g603, n1733 );
nand U3860 ( new_g4297_, n1626, n1766 );
xnor U3861 ( n1626, g1207, g1211 );
xnor U3862 ( new_g6188_, g609, n1708 );
xnor U3863 ( new_g6180_, g596, n1708 );
xor U3864 ( new_g6282_, g601, g1225 );
xor U3865 ( new_g6285_, g614, g1225 );
nand U3866 ( new_g4364_, n1618, n1619 );
nand U3867 ( n1618, g1416, g1724 );
nand U3868 ( n1619, g7063, n1712 );
nand U3869 ( new_g4249_, g1207, n1766 );
and U3870 ( new_g4349_, g942, n1621 );
and U3871 ( new_g4327_, n1787, g874 );
xnor U3872 ( new_g7328_, g819, n1785 );
and U3873 ( new_g7128_, n1849, g154 );
nor U3874 ( new_g3259_, g1269, g1268 );
endmodule

